

module top
(
  clk_i,
  reset_i,
  v_i,
  len_i,
  data_i,
  ready_o,
  v_o,
  len_v_o,
  data_o,
  yumi_i
);

  input [5:0] len_i;
  input [1599:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output len_v_o;

  bsg_parallel_in_serial_out_dynamic
  wrapper
  (
    .len_i(len_i),
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .ready_o(ready_o),
    .v_o(v_o),
    .len_v_o(len_v_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p6_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [5:0] w_data_i;
  input [0:0] r_addr_i;
  output [5:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [5:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [11:0] \nz.mem ;
  reg \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [11] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [10] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [9] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [8] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [7] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [6] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_11_sv2v_reg  <= w_data_i[5];
      \nz.mem_10_sv2v_reg  <= w_data_i[4];
      \nz.mem_9_sv2v_reg  <= w_data_i[3];
      \nz.mem_8_sv2v_reg  <= w_data_i[2];
      \nz.mem_7_sv2v_reg  <= w_data_i[1];
      \nz.mem_6_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p6_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [5:0] w_data_i;
  input [0:0] r_addr_i;
  output [5:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [5:0] r_data_o;

  bsg_mem_1r1w_synth_width_p6_els_p2_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p6
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [5:0] data_i;
  output [5:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [5:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p6_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p1600_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [1599:0] w_data_i;
  input [0:0] r_addr_i;
  output [1599:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [1599:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38;
  wire [3199:0] \nz.mem ;
  reg \nz.mem_3199_sv2v_reg ,\nz.mem_3198_sv2v_reg ,\nz.mem_3197_sv2v_reg ,
  \nz.mem_3196_sv2v_reg ,\nz.mem_3195_sv2v_reg ,\nz.mem_3194_sv2v_reg ,
  \nz.mem_3193_sv2v_reg ,\nz.mem_3192_sv2v_reg ,\nz.mem_3191_sv2v_reg ,\nz.mem_3190_sv2v_reg ,
  \nz.mem_3189_sv2v_reg ,\nz.mem_3188_sv2v_reg ,\nz.mem_3187_sv2v_reg ,
  \nz.mem_3186_sv2v_reg ,\nz.mem_3185_sv2v_reg ,\nz.mem_3184_sv2v_reg ,\nz.mem_3183_sv2v_reg ,
  \nz.mem_3182_sv2v_reg ,\nz.mem_3181_sv2v_reg ,\nz.mem_3180_sv2v_reg ,
  \nz.mem_3179_sv2v_reg ,\nz.mem_3178_sv2v_reg ,\nz.mem_3177_sv2v_reg ,\nz.mem_3176_sv2v_reg ,
  \nz.mem_3175_sv2v_reg ,\nz.mem_3174_sv2v_reg ,\nz.mem_3173_sv2v_reg ,
  \nz.mem_3172_sv2v_reg ,\nz.mem_3171_sv2v_reg ,\nz.mem_3170_sv2v_reg ,\nz.mem_3169_sv2v_reg ,
  \nz.mem_3168_sv2v_reg ,\nz.mem_3167_sv2v_reg ,\nz.mem_3166_sv2v_reg ,
  \nz.mem_3165_sv2v_reg ,\nz.mem_3164_sv2v_reg ,\nz.mem_3163_sv2v_reg ,\nz.mem_3162_sv2v_reg ,
  \nz.mem_3161_sv2v_reg ,\nz.mem_3160_sv2v_reg ,\nz.mem_3159_sv2v_reg ,
  \nz.mem_3158_sv2v_reg ,\nz.mem_3157_sv2v_reg ,\nz.mem_3156_sv2v_reg ,\nz.mem_3155_sv2v_reg ,
  \nz.mem_3154_sv2v_reg ,\nz.mem_3153_sv2v_reg ,\nz.mem_3152_sv2v_reg ,
  \nz.mem_3151_sv2v_reg ,\nz.mem_3150_sv2v_reg ,\nz.mem_3149_sv2v_reg ,\nz.mem_3148_sv2v_reg ,
  \nz.mem_3147_sv2v_reg ,\nz.mem_3146_sv2v_reg ,\nz.mem_3145_sv2v_reg ,
  \nz.mem_3144_sv2v_reg ,\nz.mem_3143_sv2v_reg ,\nz.mem_3142_sv2v_reg ,\nz.mem_3141_sv2v_reg ,
  \nz.mem_3140_sv2v_reg ,\nz.mem_3139_sv2v_reg ,\nz.mem_3138_sv2v_reg ,
  \nz.mem_3137_sv2v_reg ,\nz.mem_3136_sv2v_reg ,\nz.mem_3135_sv2v_reg ,\nz.mem_3134_sv2v_reg ,
  \nz.mem_3133_sv2v_reg ,\nz.mem_3132_sv2v_reg ,\nz.mem_3131_sv2v_reg ,
  \nz.mem_3130_sv2v_reg ,\nz.mem_3129_sv2v_reg ,\nz.mem_3128_sv2v_reg ,\nz.mem_3127_sv2v_reg ,
  \nz.mem_3126_sv2v_reg ,\nz.mem_3125_sv2v_reg ,\nz.mem_3124_sv2v_reg ,
  \nz.mem_3123_sv2v_reg ,\nz.mem_3122_sv2v_reg ,\nz.mem_3121_sv2v_reg ,\nz.mem_3120_sv2v_reg ,
  \nz.mem_3119_sv2v_reg ,\nz.mem_3118_sv2v_reg ,\nz.mem_3117_sv2v_reg ,
  \nz.mem_3116_sv2v_reg ,\nz.mem_3115_sv2v_reg ,\nz.mem_3114_sv2v_reg ,
  \nz.mem_3113_sv2v_reg ,\nz.mem_3112_sv2v_reg ,\nz.mem_3111_sv2v_reg ,\nz.mem_3110_sv2v_reg ,
  \nz.mem_3109_sv2v_reg ,\nz.mem_3108_sv2v_reg ,\nz.mem_3107_sv2v_reg ,
  \nz.mem_3106_sv2v_reg ,\nz.mem_3105_sv2v_reg ,\nz.mem_3104_sv2v_reg ,\nz.mem_3103_sv2v_reg ,
  \nz.mem_3102_sv2v_reg ,\nz.mem_3101_sv2v_reg ,\nz.mem_3100_sv2v_reg ,
  \nz.mem_3099_sv2v_reg ,\nz.mem_3098_sv2v_reg ,\nz.mem_3097_sv2v_reg ,\nz.mem_3096_sv2v_reg ,
  \nz.mem_3095_sv2v_reg ,\nz.mem_3094_sv2v_reg ,\nz.mem_3093_sv2v_reg ,
  \nz.mem_3092_sv2v_reg ,\nz.mem_3091_sv2v_reg ,\nz.mem_3090_sv2v_reg ,\nz.mem_3089_sv2v_reg ,
  \nz.mem_3088_sv2v_reg ,\nz.mem_3087_sv2v_reg ,\nz.mem_3086_sv2v_reg ,
  \nz.mem_3085_sv2v_reg ,\nz.mem_3084_sv2v_reg ,\nz.mem_3083_sv2v_reg ,\nz.mem_3082_sv2v_reg ,
  \nz.mem_3081_sv2v_reg ,\nz.mem_3080_sv2v_reg ,\nz.mem_3079_sv2v_reg ,
  \nz.mem_3078_sv2v_reg ,\nz.mem_3077_sv2v_reg ,\nz.mem_3076_sv2v_reg ,\nz.mem_3075_sv2v_reg ,
  \nz.mem_3074_sv2v_reg ,\nz.mem_3073_sv2v_reg ,\nz.mem_3072_sv2v_reg ,
  \nz.mem_3071_sv2v_reg ,\nz.mem_3070_sv2v_reg ,\nz.mem_3069_sv2v_reg ,\nz.mem_3068_sv2v_reg ,
  \nz.mem_3067_sv2v_reg ,\nz.mem_3066_sv2v_reg ,\nz.mem_3065_sv2v_reg ,
  \nz.mem_3064_sv2v_reg ,\nz.mem_3063_sv2v_reg ,\nz.mem_3062_sv2v_reg ,\nz.mem_3061_sv2v_reg ,
  \nz.mem_3060_sv2v_reg ,\nz.mem_3059_sv2v_reg ,\nz.mem_3058_sv2v_reg ,
  \nz.mem_3057_sv2v_reg ,\nz.mem_3056_sv2v_reg ,\nz.mem_3055_sv2v_reg ,\nz.mem_3054_sv2v_reg ,
  \nz.mem_3053_sv2v_reg ,\nz.mem_3052_sv2v_reg ,\nz.mem_3051_sv2v_reg ,
  \nz.mem_3050_sv2v_reg ,\nz.mem_3049_sv2v_reg ,\nz.mem_3048_sv2v_reg ,\nz.mem_3047_sv2v_reg ,
  \nz.mem_3046_sv2v_reg ,\nz.mem_3045_sv2v_reg ,\nz.mem_3044_sv2v_reg ,
  \nz.mem_3043_sv2v_reg ,\nz.mem_3042_sv2v_reg ,\nz.mem_3041_sv2v_reg ,\nz.mem_3040_sv2v_reg ,
  \nz.mem_3039_sv2v_reg ,\nz.mem_3038_sv2v_reg ,\nz.mem_3037_sv2v_reg ,
  \nz.mem_3036_sv2v_reg ,\nz.mem_3035_sv2v_reg ,\nz.mem_3034_sv2v_reg ,
  \nz.mem_3033_sv2v_reg ,\nz.mem_3032_sv2v_reg ,\nz.mem_3031_sv2v_reg ,\nz.mem_3030_sv2v_reg ,
  \nz.mem_3029_sv2v_reg ,\nz.mem_3028_sv2v_reg ,\nz.mem_3027_sv2v_reg ,
  \nz.mem_3026_sv2v_reg ,\nz.mem_3025_sv2v_reg ,\nz.mem_3024_sv2v_reg ,\nz.mem_3023_sv2v_reg ,
  \nz.mem_3022_sv2v_reg ,\nz.mem_3021_sv2v_reg ,\nz.mem_3020_sv2v_reg ,
  \nz.mem_3019_sv2v_reg ,\nz.mem_3018_sv2v_reg ,\nz.mem_3017_sv2v_reg ,\nz.mem_3016_sv2v_reg ,
  \nz.mem_3015_sv2v_reg ,\nz.mem_3014_sv2v_reg ,\nz.mem_3013_sv2v_reg ,
  \nz.mem_3012_sv2v_reg ,\nz.mem_3011_sv2v_reg ,\nz.mem_3010_sv2v_reg ,\nz.mem_3009_sv2v_reg ,
  \nz.mem_3008_sv2v_reg ,\nz.mem_3007_sv2v_reg ,\nz.mem_3006_sv2v_reg ,
  \nz.mem_3005_sv2v_reg ,\nz.mem_3004_sv2v_reg ,\nz.mem_3003_sv2v_reg ,\nz.mem_3002_sv2v_reg ,
  \nz.mem_3001_sv2v_reg ,\nz.mem_3000_sv2v_reg ,\nz.mem_2999_sv2v_reg ,
  \nz.mem_2998_sv2v_reg ,\nz.mem_2997_sv2v_reg ,\nz.mem_2996_sv2v_reg ,\nz.mem_2995_sv2v_reg ,
  \nz.mem_2994_sv2v_reg ,\nz.mem_2993_sv2v_reg ,\nz.mem_2992_sv2v_reg ,
  \nz.mem_2991_sv2v_reg ,\nz.mem_2990_sv2v_reg ,\nz.mem_2989_sv2v_reg ,\nz.mem_2988_sv2v_reg ,
  \nz.mem_2987_sv2v_reg ,\nz.mem_2986_sv2v_reg ,\nz.mem_2985_sv2v_reg ,
  \nz.mem_2984_sv2v_reg ,\nz.mem_2983_sv2v_reg ,\nz.mem_2982_sv2v_reg ,\nz.mem_2981_sv2v_reg ,
  \nz.mem_2980_sv2v_reg ,\nz.mem_2979_sv2v_reg ,\nz.mem_2978_sv2v_reg ,
  \nz.mem_2977_sv2v_reg ,\nz.mem_2976_sv2v_reg ,\nz.mem_2975_sv2v_reg ,\nz.mem_2974_sv2v_reg ,
  \nz.mem_2973_sv2v_reg ,\nz.mem_2972_sv2v_reg ,\nz.mem_2971_sv2v_reg ,
  \nz.mem_2970_sv2v_reg ,\nz.mem_2969_sv2v_reg ,\nz.mem_2968_sv2v_reg ,\nz.mem_2967_sv2v_reg ,
  \nz.mem_2966_sv2v_reg ,\nz.mem_2965_sv2v_reg ,\nz.mem_2964_sv2v_reg ,
  \nz.mem_2963_sv2v_reg ,\nz.mem_2962_sv2v_reg ,\nz.mem_2961_sv2v_reg ,\nz.mem_2960_sv2v_reg ,
  \nz.mem_2959_sv2v_reg ,\nz.mem_2958_sv2v_reg ,\nz.mem_2957_sv2v_reg ,
  \nz.mem_2956_sv2v_reg ,\nz.mem_2955_sv2v_reg ,\nz.mem_2954_sv2v_reg ,
  \nz.mem_2953_sv2v_reg ,\nz.mem_2952_sv2v_reg ,\nz.mem_2951_sv2v_reg ,\nz.mem_2950_sv2v_reg ,
  \nz.mem_2949_sv2v_reg ,\nz.mem_2948_sv2v_reg ,\nz.mem_2947_sv2v_reg ,
  \nz.mem_2946_sv2v_reg ,\nz.mem_2945_sv2v_reg ,\nz.mem_2944_sv2v_reg ,\nz.mem_2943_sv2v_reg ,
  \nz.mem_2942_sv2v_reg ,\nz.mem_2941_sv2v_reg ,\nz.mem_2940_sv2v_reg ,
  \nz.mem_2939_sv2v_reg ,\nz.mem_2938_sv2v_reg ,\nz.mem_2937_sv2v_reg ,\nz.mem_2936_sv2v_reg ,
  \nz.mem_2935_sv2v_reg ,\nz.mem_2934_sv2v_reg ,\nz.mem_2933_sv2v_reg ,
  \nz.mem_2932_sv2v_reg ,\nz.mem_2931_sv2v_reg ,\nz.mem_2930_sv2v_reg ,\nz.mem_2929_sv2v_reg ,
  \nz.mem_2928_sv2v_reg ,\nz.mem_2927_sv2v_reg ,\nz.mem_2926_sv2v_reg ,
  \nz.mem_2925_sv2v_reg ,\nz.mem_2924_sv2v_reg ,\nz.mem_2923_sv2v_reg ,\nz.mem_2922_sv2v_reg ,
  \nz.mem_2921_sv2v_reg ,\nz.mem_2920_sv2v_reg ,\nz.mem_2919_sv2v_reg ,
  \nz.mem_2918_sv2v_reg ,\nz.mem_2917_sv2v_reg ,\nz.mem_2916_sv2v_reg ,\nz.mem_2915_sv2v_reg ,
  \nz.mem_2914_sv2v_reg ,\nz.mem_2913_sv2v_reg ,\nz.mem_2912_sv2v_reg ,
  \nz.mem_2911_sv2v_reg ,\nz.mem_2910_sv2v_reg ,\nz.mem_2909_sv2v_reg ,\nz.mem_2908_sv2v_reg ,
  \nz.mem_2907_sv2v_reg ,\nz.mem_2906_sv2v_reg ,\nz.mem_2905_sv2v_reg ,
  \nz.mem_2904_sv2v_reg ,\nz.mem_2903_sv2v_reg ,\nz.mem_2902_sv2v_reg ,\nz.mem_2901_sv2v_reg ,
  \nz.mem_2900_sv2v_reg ,\nz.mem_2899_sv2v_reg ,\nz.mem_2898_sv2v_reg ,
  \nz.mem_2897_sv2v_reg ,\nz.mem_2896_sv2v_reg ,\nz.mem_2895_sv2v_reg ,\nz.mem_2894_sv2v_reg ,
  \nz.mem_2893_sv2v_reg ,\nz.mem_2892_sv2v_reg ,\nz.mem_2891_sv2v_reg ,
  \nz.mem_2890_sv2v_reg ,\nz.mem_2889_sv2v_reg ,\nz.mem_2888_sv2v_reg ,\nz.mem_2887_sv2v_reg ,
  \nz.mem_2886_sv2v_reg ,\nz.mem_2885_sv2v_reg ,\nz.mem_2884_sv2v_reg ,
  \nz.mem_2883_sv2v_reg ,\nz.mem_2882_sv2v_reg ,\nz.mem_2881_sv2v_reg ,\nz.mem_2880_sv2v_reg ,
  \nz.mem_2879_sv2v_reg ,\nz.mem_2878_sv2v_reg ,\nz.mem_2877_sv2v_reg ,
  \nz.mem_2876_sv2v_reg ,\nz.mem_2875_sv2v_reg ,\nz.mem_2874_sv2v_reg ,
  \nz.mem_2873_sv2v_reg ,\nz.mem_2872_sv2v_reg ,\nz.mem_2871_sv2v_reg ,\nz.mem_2870_sv2v_reg ,
  \nz.mem_2869_sv2v_reg ,\nz.mem_2868_sv2v_reg ,\nz.mem_2867_sv2v_reg ,
  \nz.mem_2866_sv2v_reg ,\nz.mem_2865_sv2v_reg ,\nz.mem_2864_sv2v_reg ,\nz.mem_2863_sv2v_reg ,
  \nz.mem_2862_sv2v_reg ,\nz.mem_2861_sv2v_reg ,\nz.mem_2860_sv2v_reg ,
  \nz.mem_2859_sv2v_reg ,\nz.mem_2858_sv2v_reg ,\nz.mem_2857_sv2v_reg ,\nz.mem_2856_sv2v_reg ,
  \nz.mem_2855_sv2v_reg ,\nz.mem_2854_sv2v_reg ,\nz.mem_2853_sv2v_reg ,
  \nz.mem_2852_sv2v_reg ,\nz.mem_2851_sv2v_reg ,\nz.mem_2850_sv2v_reg ,\nz.mem_2849_sv2v_reg ,
  \nz.mem_2848_sv2v_reg ,\nz.mem_2847_sv2v_reg ,\nz.mem_2846_sv2v_reg ,
  \nz.mem_2845_sv2v_reg ,\nz.mem_2844_sv2v_reg ,\nz.mem_2843_sv2v_reg ,\nz.mem_2842_sv2v_reg ,
  \nz.mem_2841_sv2v_reg ,\nz.mem_2840_sv2v_reg ,\nz.mem_2839_sv2v_reg ,
  \nz.mem_2838_sv2v_reg ,\nz.mem_2837_sv2v_reg ,\nz.mem_2836_sv2v_reg ,\nz.mem_2835_sv2v_reg ,
  \nz.mem_2834_sv2v_reg ,\nz.mem_2833_sv2v_reg ,\nz.mem_2832_sv2v_reg ,
  \nz.mem_2831_sv2v_reg ,\nz.mem_2830_sv2v_reg ,\nz.mem_2829_sv2v_reg ,\nz.mem_2828_sv2v_reg ,
  \nz.mem_2827_sv2v_reg ,\nz.mem_2826_sv2v_reg ,\nz.mem_2825_sv2v_reg ,
  \nz.mem_2824_sv2v_reg ,\nz.mem_2823_sv2v_reg ,\nz.mem_2822_sv2v_reg ,\nz.mem_2821_sv2v_reg ,
  \nz.mem_2820_sv2v_reg ,\nz.mem_2819_sv2v_reg ,\nz.mem_2818_sv2v_reg ,
  \nz.mem_2817_sv2v_reg ,\nz.mem_2816_sv2v_reg ,\nz.mem_2815_sv2v_reg ,\nz.mem_2814_sv2v_reg ,
  \nz.mem_2813_sv2v_reg ,\nz.mem_2812_sv2v_reg ,\nz.mem_2811_sv2v_reg ,
  \nz.mem_2810_sv2v_reg ,\nz.mem_2809_sv2v_reg ,\nz.mem_2808_sv2v_reg ,\nz.mem_2807_sv2v_reg ,
  \nz.mem_2806_sv2v_reg ,\nz.mem_2805_sv2v_reg ,\nz.mem_2804_sv2v_reg ,
  \nz.mem_2803_sv2v_reg ,\nz.mem_2802_sv2v_reg ,\nz.mem_2801_sv2v_reg ,\nz.mem_2800_sv2v_reg ,
  \nz.mem_2799_sv2v_reg ,\nz.mem_2798_sv2v_reg ,\nz.mem_2797_sv2v_reg ,
  \nz.mem_2796_sv2v_reg ,\nz.mem_2795_sv2v_reg ,\nz.mem_2794_sv2v_reg ,
  \nz.mem_2793_sv2v_reg ,\nz.mem_2792_sv2v_reg ,\nz.mem_2791_sv2v_reg ,\nz.mem_2790_sv2v_reg ,
  \nz.mem_2789_sv2v_reg ,\nz.mem_2788_sv2v_reg ,\nz.mem_2787_sv2v_reg ,
  \nz.mem_2786_sv2v_reg ,\nz.mem_2785_sv2v_reg ,\nz.mem_2784_sv2v_reg ,\nz.mem_2783_sv2v_reg ,
  \nz.mem_2782_sv2v_reg ,\nz.mem_2781_sv2v_reg ,\nz.mem_2780_sv2v_reg ,
  \nz.mem_2779_sv2v_reg ,\nz.mem_2778_sv2v_reg ,\nz.mem_2777_sv2v_reg ,\nz.mem_2776_sv2v_reg ,
  \nz.mem_2775_sv2v_reg ,\nz.mem_2774_sv2v_reg ,\nz.mem_2773_sv2v_reg ,
  \nz.mem_2772_sv2v_reg ,\nz.mem_2771_sv2v_reg ,\nz.mem_2770_sv2v_reg ,\nz.mem_2769_sv2v_reg ,
  \nz.mem_2768_sv2v_reg ,\nz.mem_2767_sv2v_reg ,\nz.mem_2766_sv2v_reg ,
  \nz.mem_2765_sv2v_reg ,\nz.mem_2764_sv2v_reg ,\nz.mem_2763_sv2v_reg ,\nz.mem_2762_sv2v_reg ,
  \nz.mem_2761_sv2v_reg ,\nz.mem_2760_sv2v_reg ,\nz.mem_2759_sv2v_reg ,
  \nz.mem_2758_sv2v_reg ,\nz.mem_2757_sv2v_reg ,\nz.mem_2756_sv2v_reg ,\nz.mem_2755_sv2v_reg ,
  \nz.mem_2754_sv2v_reg ,\nz.mem_2753_sv2v_reg ,\nz.mem_2752_sv2v_reg ,
  \nz.mem_2751_sv2v_reg ,\nz.mem_2750_sv2v_reg ,\nz.mem_2749_sv2v_reg ,\nz.mem_2748_sv2v_reg ,
  \nz.mem_2747_sv2v_reg ,\nz.mem_2746_sv2v_reg ,\nz.mem_2745_sv2v_reg ,
  \nz.mem_2744_sv2v_reg ,\nz.mem_2743_sv2v_reg ,\nz.mem_2742_sv2v_reg ,\nz.mem_2741_sv2v_reg ,
  \nz.mem_2740_sv2v_reg ,\nz.mem_2739_sv2v_reg ,\nz.mem_2738_sv2v_reg ,
  \nz.mem_2737_sv2v_reg ,\nz.mem_2736_sv2v_reg ,\nz.mem_2735_sv2v_reg ,\nz.mem_2734_sv2v_reg ,
  \nz.mem_2733_sv2v_reg ,\nz.mem_2732_sv2v_reg ,\nz.mem_2731_sv2v_reg ,
  \nz.mem_2730_sv2v_reg ,\nz.mem_2729_sv2v_reg ,\nz.mem_2728_sv2v_reg ,\nz.mem_2727_sv2v_reg ,
  \nz.mem_2726_sv2v_reg ,\nz.mem_2725_sv2v_reg ,\nz.mem_2724_sv2v_reg ,
  \nz.mem_2723_sv2v_reg ,\nz.mem_2722_sv2v_reg ,\nz.mem_2721_sv2v_reg ,\nz.mem_2720_sv2v_reg ,
  \nz.mem_2719_sv2v_reg ,\nz.mem_2718_sv2v_reg ,\nz.mem_2717_sv2v_reg ,
  \nz.mem_2716_sv2v_reg ,\nz.mem_2715_sv2v_reg ,\nz.mem_2714_sv2v_reg ,
  \nz.mem_2713_sv2v_reg ,\nz.mem_2712_sv2v_reg ,\nz.mem_2711_sv2v_reg ,\nz.mem_2710_sv2v_reg ,
  \nz.mem_2709_sv2v_reg ,\nz.mem_2708_sv2v_reg ,\nz.mem_2707_sv2v_reg ,
  \nz.mem_2706_sv2v_reg ,\nz.mem_2705_sv2v_reg ,\nz.mem_2704_sv2v_reg ,\nz.mem_2703_sv2v_reg ,
  \nz.mem_2702_sv2v_reg ,\nz.mem_2701_sv2v_reg ,\nz.mem_2700_sv2v_reg ,
  \nz.mem_2699_sv2v_reg ,\nz.mem_2698_sv2v_reg ,\nz.mem_2697_sv2v_reg ,\nz.mem_2696_sv2v_reg ,
  \nz.mem_2695_sv2v_reg ,\nz.mem_2694_sv2v_reg ,\nz.mem_2693_sv2v_reg ,
  \nz.mem_2692_sv2v_reg ,\nz.mem_2691_sv2v_reg ,\nz.mem_2690_sv2v_reg ,\nz.mem_2689_sv2v_reg ,
  \nz.mem_2688_sv2v_reg ,\nz.mem_2687_sv2v_reg ,\nz.mem_2686_sv2v_reg ,
  \nz.mem_2685_sv2v_reg ,\nz.mem_2684_sv2v_reg ,\nz.mem_2683_sv2v_reg ,\nz.mem_2682_sv2v_reg ,
  \nz.mem_2681_sv2v_reg ,\nz.mem_2680_sv2v_reg ,\nz.mem_2679_sv2v_reg ,
  \nz.mem_2678_sv2v_reg ,\nz.mem_2677_sv2v_reg ,\nz.mem_2676_sv2v_reg ,\nz.mem_2675_sv2v_reg ,
  \nz.mem_2674_sv2v_reg ,\nz.mem_2673_sv2v_reg ,\nz.mem_2672_sv2v_reg ,
  \nz.mem_2671_sv2v_reg ,\nz.mem_2670_sv2v_reg ,\nz.mem_2669_sv2v_reg ,\nz.mem_2668_sv2v_reg ,
  \nz.mem_2667_sv2v_reg ,\nz.mem_2666_sv2v_reg ,\nz.mem_2665_sv2v_reg ,
  \nz.mem_2664_sv2v_reg ,\nz.mem_2663_sv2v_reg ,\nz.mem_2662_sv2v_reg ,\nz.mem_2661_sv2v_reg ,
  \nz.mem_2660_sv2v_reg ,\nz.mem_2659_sv2v_reg ,\nz.mem_2658_sv2v_reg ,
  \nz.mem_2657_sv2v_reg ,\nz.mem_2656_sv2v_reg ,\nz.mem_2655_sv2v_reg ,\nz.mem_2654_sv2v_reg ,
  \nz.mem_2653_sv2v_reg ,\nz.mem_2652_sv2v_reg ,\nz.mem_2651_sv2v_reg ,
  \nz.mem_2650_sv2v_reg ,\nz.mem_2649_sv2v_reg ,\nz.mem_2648_sv2v_reg ,\nz.mem_2647_sv2v_reg ,
  \nz.mem_2646_sv2v_reg ,\nz.mem_2645_sv2v_reg ,\nz.mem_2644_sv2v_reg ,
  \nz.mem_2643_sv2v_reg ,\nz.mem_2642_sv2v_reg ,\nz.mem_2641_sv2v_reg ,\nz.mem_2640_sv2v_reg ,
  \nz.mem_2639_sv2v_reg ,\nz.mem_2638_sv2v_reg ,\nz.mem_2637_sv2v_reg ,
  \nz.mem_2636_sv2v_reg ,\nz.mem_2635_sv2v_reg ,\nz.mem_2634_sv2v_reg ,
  \nz.mem_2633_sv2v_reg ,\nz.mem_2632_sv2v_reg ,\nz.mem_2631_sv2v_reg ,\nz.mem_2630_sv2v_reg ,
  \nz.mem_2629_sv2v_reg ,\nz.mem_2628_sv2v_reg ,\nz.mem_2627_sv2v_reg ,
  \nz.mem_2626_sv2v_reg ,\nz.mem_2625_sv2v_reg ,\nz.mem_2624_sv2v_reg ,\nz.mem_2623_sv2v_reg ,
  \nz.mem_2622_sv2v_reg ,\nz.mem_2621_sv2v_reg ,\nz.mem_2620_sv2v_reg ,
  \nz.mem_2619_sv2v_reg ,\nz.mem_2618_sv2v_reg ,\nz.mem_2617_sv2v_reg ,\nz.mem_2616_sv2v_reg ,
  \nz.mem_2615_sv2v_reg ,\nz.mem_2614_sv2v_reg ,\nz.mem_2613_sv2v_reg ,
  \nz.mem_2612_sv2v_reg ,\nz.mem_2611_sv2v_reg ,\nz.mem_2610_sv2v_reg ,\nz.mem_2609_sv2v_reg ,
  \nz.mem_2608_sv2v_reg ,\nz.mem_2607_sv2v_reg ,\nz.mem_2606_sv2v_reg ,
  \nz.mem_2605_sv2v_reg ,\nz.mem_2604_sv2v_reg ,\nz.mem_2603_sv2v_reg ,\nz.mem_2602_sv2v_reg ,
  \nz.mem_2601_sv2v_reg ,\nz.mem_2600_sv2v_reg ,\nz.mem_2599_sv2v_reg ,
  \nz.mem_2598_sv2v_reg ,\nz.mem_2597_sv2v_reg ,\nz.mem_2596_sv2v_reg ,\nz.mem_2595_sv2v_reg ,
  \nz.mem_2594_sv2v_reg ,\nz.mem_2593_sv2v_reg ,\nz.mem_2592_sv2v_reg ,
  \nz.mem_2591_sv2v_reg ,\nz.mem_2590_sv2v_reg ,\nz.mem_2589_sv2v_reg ,\nz.mem_2588_sv2v_reg ,
  \nz.mem_2587_sv2v_reg ,\nz.mem_2586_sv2v_reg ,\nz.mem_2585_sv2v_reg ,
  \nz.mem_2584_sv2v_reg ,\nz.mem_2583_sv2v_reg ,\nz.mem_2582_sv2v_reg ,\nz.mem_2581_sv2v_reg ,
  \nz.mem_2580_sv2v_reg ,\nz.mem_2579_sv2v_reg ,\nz.mem_2578_sv2v_reg ,
  \nz.mem_2577_sv2v_reg ,\nz.mem_2576_sv2v_reg ,\nz.mem_2575_sv2v_reg ,\nz.mem_2574_sv2v_reg ,
  \nz.mem_2573_sv2v_reg ,\nz.mem_2572_sv2v_reg ,\nz.mem_2571_sv2v_reg ,
  \nz.mem_2570_sv2v_reg ,\nz.mem_2569_sv2v_reg ,\nz.mem_2568_sv2v_reg ,\nz.mem_2567_sv2v_reg ,
  \nz.mem_2566_sv2v_reg ,\nz.mem_2565_sv2v_reg ,\nz.mem_2564_sv2v_reg ,
  \nz.mem_2563_sv2v_reg ,\nz.mem_2562_sv2v_reg ,\nz.mem_2561_sv2v_reg ,\nz.mem_2560_sv2v_reg ,
  \nz.mem_2559_sv2v_reg ,\nz.mem_2558_sv2v_reg ,\nz.mem_2557_sv2v_reg ,
  \nz.mem_2556_sv2v_reg ,\nz.mem_2555_sv2v_reg ,\nz.mem_2554_sv2v_reg ,
  \nz.mem_2553_sv2v_reg ,\nz.mem_2552_sv2v_reg ,\nz.mem_2551_sv2v_reg ,\nz.mem_2550_sv2v_reg ,
  \nz.mem_2549_sv2v_reg ,\nz.mem_2548_sv2v_reg ,\nz.mem_2547_sv2v_reg ,
  \nz.mem_2546_sv2v_reg ,\nz.mem_2545_sv2v_reg ,\nz.mem_2544_sv2v_reg ,\nz.mem_2543_sv2v_reg ,
  \nz.mem_2542_sv2v_reg ,\nz.mem_2541_sv2v_reg ,\nz.mem_2540_sv2v_reg ,
  \nz.mem_2539_sv2v_reg ,\nz.mem_2538_sv2v_reg ,\nz.mem_2537_sv2v_reg ,\nz.mem_2536_sv2v_reg ,
  \nz.mem_2535_sv2v_reg ,\nz.mem_2534_sv2v_reg ,\nz.mem_2533_sv2v_reg ,
  \nz.mem_2532_sv2v_reg ,\nz.mem_2531_sv2v_reg ,\nz.mem_2530_sv2v_reg ,\nz.mem_2529_sv2v_reg ,
  \nz.mem_2528_sv2v_reg ,\nz.mem_2527_sv2v_reg ,\nz.mem_2526_sv2v_reg ,
  \nz.mem_2525_sv2v_reg ,\nz.mem_2524_sv2v_reg ,\nz.mem_2523_sv2v_reg ,\nz.mem_2522_sv2v_reg ,
  \nz.mem_2521_sv2v_reg ,\nz.mem_2520_sv2v_reg ,\nz.mem_2519_sv2v_reg ,
  \nz.mem_2518_sv2v_reg ,\nz.mem_2517_sv2v_reg ,\nz.mem_2516_sv2v_reg ,\nz.mem_2515_sv2v_reg ,
  \nz.mem_2514_sv2v_reg ,\nz.mem_2513_sv2v_reg ,\nz.mem_2512_sv2v_reg ,
  \nz.mem_2511_sv2v_reg ,\nz.mem_2510_sv2v_reg ,\nz.mem_2509_sv2v_reg ,\nz.mem_2508_sv2v_reg ,
  \nz.mem_2507_sv2v_reg ,\nz.mem_2506_sv2v_reg ,\nz.mem_2505_sv2v_reg ,
  \nz.mem_2504_sv2v_reg ,\nz.mem_2503_sv2v_reg ,\nz.mem_2502_sv2v_reg ,\nz.mem_2501_sv2v_reg ,
  \nz.mem_2500_sv2v_reg ,\nz.mem_2499_sv2v_reg ,\nz.mem_2498_sv2v_reg ,
  \nz.mem_2497_sv2v_reg ,\nz.mem_2496_sv2v_reg ,\nz.mem_2495_sv2v_reg ,\nz.mem_2494_sv2v_reg ,
  \nz.mem_2493_sv2v_reg ,\nz.mem_2492_sv2v_reg ,\nz.mem_2491_sv2v_reg ,
  \nz.mem_2490_sv2v_reg ,\nz.mem_2489_sv2v_reg ,\nz.mem_2488_sv2v_reg ,\nz.mem_2487_sv2v_reg ,
  \nz.mem_2486_sv2v_reg ,\nz.mem_2485_sv2v_reg ,\nz.mem_2484_sv2v_reg ,
  \nz.mem_2483_sv2v_reg ,\nz.mem_2482_sv2v_reg ,\nz.mem_2481_sv2v_reg ,\nz.mem_2480_sv2v_reg ,
  \nz.mem_2479_sv2v_reg ,\nz.mem_2478_sv2v_reg ,\nz.mem_2477_sv2v_reg ,
  \nz.mem_2476_sv2v_reg ,\nz.mem_2475_sv2v_reg ,\nz.mem_2474_sv2v_reg ,
  \nz.mem_2473_sv2v_reg ,\nz.mem_2472_sv2v_reg ,\nz.mem_2471_sv2v_reg ,\nz.mem_2470_sv2v_reg ,
  \nz.mem_2469_sv2v_reg ,\nz.mem_2468_sv2v_reg ,\nz.mem_2467_sv2v_reg ,
  \nz.mem_2466_sv2v_reg ,\nz.mem_2465_sv2v_reg ,\nz.mem_2464_sv2v_reg ,\nz.mem_2463_sv2v_reg ,
  \nz.mem_2462_sv2v_reg ,\nz.mem_2461_sv2v_reg ,\nz.mem_2460_sv2v_reg ,
  \nz.mem_2459_sv2v_reg ,\nz.mem_2458_sv2v_reg ,\nz.mem_2457_sv2v_reg ,\nz.mem_2456_sv2v_reg ,
  \nz.mem_2455_sv2v_reg ,\nz.mem_2454_sv2v_reg ,\nz.mem_2453_sv2v_reg ,
  \nz.mem_2452_sv2v_reg ,\nz.mem_2451_sv2v_reg ,\nz.mem_2450_sv2v_reg ,\nz.mem_2449_sv2v_reg ,
  \nz.mem_2448_sv2v_reg ,\nz.mem_2447_sv2v_reg ,\nz.mem_2446_sv2v_reg ,
  \nz.mem_2445_sv2v_reg ,\nz.mem_2444_sv2v_reg ,\nz.mem_2443_sv2v_reg ,\nz.mem_2442_sv2v_reg ,
  \nz.mem_2441_sv2v_reg ,\nz.mem_2440_sv2v_reg ,\nz.mem_2439_sv2v_reg ,
  \nz.mem_2438_sv2v_reg ,\nz.mem_2437_sv2v_reg ,\nz.mem_2436_sv2v_reg ,\nz.mem_2435_sv2v_reg ,
  \nz.mem_2434_sv2v_reg ,\nz.mem_2433_sv2v_reg ,\nz.mem_2432_sv2v_reg ,
  \nz.mem_2431_sv2v_reg ,\nz.mem_2430_sv2v_reg ,\nz.mem_2429_sv2v_reg ,\nz.mem_2428_sv2v_reg ,
  \nz.mem_2427_sv2v_reg ,\nz.mem_2426_sv2v_reg ,\nz.mem_2425_sv2v_reg ,
  \nz.mem_2424_sv2v_reg ,\nz.mem_2423_sv2v_reg ,\nz.mem_2422_sv2v_reg ,\nz.mem_2421_sv2v_reg ,
  \nz.mem_2420_sv2v_reg ,\nz.mem_2419_sv2v_reg ,\nz.mem_2418_sv2v_reg ,
  \nz.mem_2417_sv2v_reg ,\nz.mem_2416_sv2v_reg ,\nz.mem_2415_sv2v_reg ,\nz.mem_2414_sv2v_reg ,
  \nz.mem_2413_sv2v_reg ,\nz.mem_2412_sv2v_reg ,\nz.mem_2411_sv2v_reg ,
  \nz.mem_2410_sv2v_reg ,\nz.mem_2409_sv2v_reg ,\nz.mem_2408_sv2v_reg ,\nz.mem_2407_sv2v_reg ,
  \nz.mem_2406_sv2v_reg ,\nz.mem_2405_sv2v_reg ,\nz.mem_2404_sv2v_reg ,
  \nz.mem_2403_sv2v_reg ,\nz.mem_2402_sv2v_reg ,\nz.mem_2401_sv2v_reg ,\nz.mem_2400_sv2v_reg ,
  \nz.mem_2399_sv2v_reg ,\nz.mem_2398_sv2v_reg ,\nz.mem_2397_sv2v_reg ,
  \nz.mem_2396_sv2v_reg ,\nz.mem_2395_sv2v_reg ,\nz.mem_2394_sv2v_reg ,
  \nz.mem_2393_sv2v_reg ,\nz.mem_2392_sv2v_reg ,\nz.mem_2391_sv2v_reg ,\nz.mem_2390_sv2v_reg ,
  \nz.mem_2389_sv2v_reg ,\nz.mem_2388_sv2v_reg ,\nz.mem_2387_sv2v_reg ,
  \nz.mem_2386_sv2v_reg ,\nz.mem_2385_sv2v_reg ,\nz.mem_2384_sv2v_reg ,\nz.mem_2383_sv2v_reg ,
  \nz.mem_2382_sv2v_reg ,\nz.mem_2381_sv2v_reg ,\nz.mem_2380_sv2v_reg ,
  \nz.mem_2379_sv2v_reg ,\nz.mem_2378_sv2v_reg ,\nz.mem_2377_sv2v_reg ,\nz.mem_2376_sv2v_reg ,
  \nz.mem_2375_sv2v_reg ,\nz.mem_2374_sv2v_reg ,\nz.mem_2373_sv2v_reg ,
  \nz.mem_2372_sv2v_reg ,\nz.mem_2371_sv2v_reg ,\nz.mem_2370_sv2v_reg ,\nz.mem_2369_sv2v_reg ,
  \nz.mem_2368_sv2v_reg ,\nz.mem_2367_sv2v_reg ,\nz.mem_2366_sv2v_reg ,
  \nz.mem_2365_sv2v_reg ,\nz.mem_2364_sv2v_reg ,\nz.mem_2363_sv2v_reg ,\nz.mem_2362_sv2v_reg ,
  \nz.mem_2361_sv2v_reg ,\nz.mem_2360_sv2v_reg ,\nz.mem_2359_sv2v_reg ,
  \nz.mem_2358_sv2v_reg ,\nz.mem_2357_sv2v_reg ,\nz.mem_2356_sv2v_reg ,\nz.mem_2355_sv2v_reg ,
  \nz.mem_2354_sv2v_reg ,\nz.mem_2353_sv2v_reg ,\nz.mem_2352_sv2v_reg ,
  \nz.mem_2351_sv2v_reg ,\nz.mem_2350_sv2v_reg ,\nz.mem_2349_sv2v_reg ,\nz.mem_2348_sv2v_reg ,
  \nz.mem_2347_sv2v_reg ,\nz.mem_2346_sv2v_reg ,\nz.mem_2345_sv2v_reg ,
  \nz.mem_2344_sv2v_reg ,\nz.mem_2343_sv2v_reg ,\nz.mem_2342_sv2v_reg ,\nz.mem_2341_sv2v_reg ,
  \nz.mem_2340_sv2v_reg ,\nz.mem_2339_sv2v_reg ,\nz.mem_2338_sv2v_reg ,
  \nz.mem_2337_sv2v_reg ,\nz.mem_2336_sv2v_reg ,\nz.mem_2335_sv2v_reg ,\nz.mem_2334_sv2v_reg ,
  \nz.mem_2333_sv2v_reg ,\nz.mem_2332_sv2v_reg ,\nz.mem_2331_sv2v_reg ,
  \nz.mem_2330_sv2v_reg ,\nz.mem_2329_sv2v_reg ,\nz.mem_2328_sv2v_reg ,\nz.mem_2327_sv2v_reg ,
  \nz.mem_2326_sv2v_reg ,\nz.mem_2325_sv2v_reg ,\nz.mem_2324_sv2v_reg ,
  \nz.mem_2323_sv2v_reg ,\nz.mem_2322_sv2v_reg ,\nz.mem_2321_sv2v_reg ,\nz.mem_2320_sv2v_reg ,
  \nz.mem_2319_sv2v_reg ,\nz.mem_2318_sv2v_reg ,\nz.mem_2317_sv2v_reg ,
  \nz.mem_2316_sv2v_reg ,\nz.mem_2315_sv2v_reg ,\nz.mem_2314_sv2v_reg ,
  \nz.mem_2313_sv2v_reg ,\nz.mem_2312_sv2v_reg ,\nz.mem_2311_sv2v_reg ,\nz.mem_2310_sv2v_reg ,
  \nz.mem_2309_sv2v_reg ,\nz.mem_2308_sv2v_reg ,\nz.mem_2307_sv2v_reg ,
  \nz.mem_2306_sv2v_reg ,\nz.mem_2305_sv2v_reg ,\nz.mem_2304_sv2v_reg ,\nz.mem_2303_sv2v_reg ,
  \nz.mem_2302_sv2v_reg ,\nz.mem_2301_sv2v_reg ,\nz.mem_2300_sv2v_reg ,
  \nz.mem_2299_sv2v_reg ,\nz.mem_2298_sv2v_reg ,\nz.mem_2297_sv2v_reg ,\nz.mem_2296_sv2v_reg ,
  \nz.mem_2295_sv2v_reg ,\nz.mem_2294_sv2v_reg ,\nz.mem_2293_sv2v_reg ,
  \nz.mem_2292_sv2v_reg ,\nz.mem_2291_sv2v_reg ,\nz.mem_2290_sv2v_reg ,\nz.mem_2289_sv2v_reg ,
  \nz.mem_2288_sv2v_reg ,\nz.mem_2287_sv2v_reg ,\nz.mem_2286_sv2v_reg ,
  \nz.mem_2285_sv2v_reg ,\nz.mem_2284_sv2v_reg ,\nz.mem_2283_sv2v_reg ,\nz.mem_2282_sv2v_reg ,
  \nz.mem_2281_sv2v_reg ,\nz.mem_2280_sv2v_reg ,\nz.mem_2279_sv2v_reg ,
  \nz.mem_2278_sv2v_reg ,\nz.mem_2277_sv2v_reg ,\nz.mem_2276_sv2v_reg ,\nz.mem_2275_sv2v_reg ,
  \nz.mem_2274_sv2v_reg ,\nz.mem_2273_sv2v_reg ,\nz.mem_2272_sv2v_reg ,
  \nz.mem_2271_sv2v_reg ,\nz.mem_2270_sv2v_reg ,\nz.mem_2269_sv2v_reg ,\nz.mem_2268_sv2v_reg ,
  \nz.mem_2267_sv2v_reg ,\nz.mem_2266_sv2v_reg ,\nz.mem_2265_sv2v_reg ,
  \nz.mem_2264_sv2v_reg ,\nz.mem_2263_sv2v_reg ,\nz.mem_2262_sv2v_reg ,\nz.mem_2261_sv2v_reg ,
  \nz.mem_2260_sv2v_reg ,\nz.mem_2259_sv2v_reg ,\nz.mem_2258_sv2v_reg ,
  \nz.mem_2257_sv2v_reg ,\nz.mem_2256_sv2v_reg ,\nz.mem_2255_sv2v_reg ,\nz.mem_2254_sv2v_reg ,
  \nz.mem_2253_sv2v_reg ,\nz.mem_2252_sv2v_reg ,\nz.mem_2251_sv2v_reg ,
  \nz.mem_2250_sv2v_reg ,\nz.mem_2249_sv2v_reg ,\nz.mem_2248_sv2v_reg ,\nz.mem_2247_sv2v_reg ,
  \nz.mem_2246_sv2v_reg ,\nz.mem_2245_sv2v_reg ,\nz.mem_2244_sv2v_reg ,
  \nz.mem_2243_sv2v_reg ,\nz.mem_2242_sv2v_reg ,\nz.mem_2241_sv2v_reg ,\nz.mem_2240_sv2v_reg ,
  \nz.mem_2239_sv2v_reg ,\nz.mem_2238_sv2v_reg ,\nz.mem_2237_sv2v_reg ,
  \nz.mem_2236_sv2v_reg ,\nz.mem_2235_sv2v_reg ,\nz.mem_2234_sv2v_reg ,
  \nz.mem_2233_sv2v_reg ,\nz.mem_2232_sv2v_reg ,\nz.mem_2231_sv2v_reg ,\nz.mem_2230_sv2v_reg ,
  \nz.mem_2229_sv2v_reg ,\nz.mem_2228_sv2v_reg ,\nz.mem_2227_sv2v_reg ,
  \nz.mem_2226_sv2v_reg ,\nz.mem_2225_sv2v_reg ,\nz.mem_2224_sv2v_reg ,\nz.mem_2223_sv2v_reg ,
  \nz.mem_2222_sv2v_reg ,\nz.mem_2221_sv2v_reg ,\nz.mem_2220_sv2v_reg ,
  \nz.mem_2219_sv2v_reg ,\nz.mem_2218_sv2v_reg ,\nz.mem_2217_sv2v_reg ,\nz.mem_2216_sv2v_reg ,
  \nz.mem_2215_sv2v_reg ,\nz.mem_2214_sv2v_reg ,\nz.mem_2213_sv2v_reg ,
  \nz.mem_2212_sv2v_reg ,\nz.mem_2211_sv2v_reg ,\nz.mem_2210_sv2v_reg ,\nz.mem_2209_sv2v_reg ,
  \nz.mem_2208_sv2v_reg ,\nz.mem_2207_sv2v_reg ,\nz.mem_2206_sv2v_reg ,
  \nz.mem_2205_sv2v_reg ,\nz.mem_2204_sv2v_reg ,\nz.mem_2203_sv2v_reg ,\nz.mem_2202_sv2v_reg ,
  \nz.mem_2201_sv2v_reg ,\nz.mem_2200_sv2v_reg ,\nz.mem_2199_sv2v_reg ,
  \nz.mem_2198_sv2v_reg ,\nz.mem_2197_sv2v_reg ,\nz.mem_2196_sv2v_reg ,\nz.mem_2195_sv2v_reg ,
  \nz.mem_2194_sv2v_reg ,\nz.mem_2193_sv2v_reg ,\nz.mem_2192_sv2v_reg ,
  \nz.mem_2191_sv2v_reg ,\nz.mem_2190_sv2v_reg ,\nz.mem_2189_sv2v_reg ,\nz.mem_2188_sv2v_reg ,
  \nz.mem_2187_sv2v_reg ,\nz.mem_2186_sv2v_reg ,\nz.mem_2185_sv2v_reg ,
  \nz.mem_2184_sv2v_reg ,\nz.mem_2183_sv2v_reg ,\nz.mem_2182_sv2v_reg ,\nz.mem_2181_sv2v_reg ,
  \nz.mem_2180_sv2v_reg ,\nz.mem_2179_sv2v_reg ,\nz.mem_2178_sv2v_reg ,
  \nz.mem_2177_sv2v_reg ,\nz.mem_2176_sv2v_reg ,\nz.mem_2175_sv2v_reg ,\nz.mem_2174_sv2v_reg ,
  \nz.mem_2173_sv2v_reg ,\nz.mem_2172_sv2v_reg ,\nz.mem_2171_sv2v_reg ,
  \nz.mem_2170_sv2v_reg ,\nz.mem_2169_sv2v_reg ,\nz.mem_2168_sv2v_reg ,\nz.mem_2167_sv2v_reg ,
  \nz.mem_2166_sv2v_reg ,\nz.mem_2165_sv2v_reg ,\nz.mem_2164_sv2v_reg ,
  \nz.mem_2163_sv2v_reg ,\nz.mem_2162_sv2v_reg ,\nz.mem_2161_sv2v_reg ,\nz.mem_2160_sv2v_reg ,
  \nz.mem_2159_sv2v_reg ,\nz.mem_2158_sv2v_reg ,\nz.mem_2157_sv2v_reg ,
  \nz.mem_2156_sv2v_reg ,\nz.mem_2155_sv2v_reg ,\nz.mem_2154_sv2v_reg ,
  \nz.mem_2153_sv2v_reg ,\nz.mem_2152_sv2v_reg ,\nz.mem_2151_sv2v_reg ,\nz.mem_2150_sv2v_reg ,
  \nz.mem_2149_sv2v_reg ,\nz.mem_2148_sv2v_reg ,\nz.mem_2147_sv2v_reg ,
  \nz.mem_2146_sv2v_reg ,\nz.mem_2145_sv2v_reg ,\nz.mem_2144_sv2v_reg ,\nz.mem_2143_sv2v_reg ,
  \nz.mem_2142_sv2v_reg ,\nz.mem_2141_sv2v_reg ,\nz.mem_2140_sv2v_reg ,
  \nz.mem_2139_sv2v_reg ,\nz.mem_2138_sv2v_reg ,\nz.mem_2137_sv2v_reg ,\nz.mem_2136_sv2v_reg ,
  \nz.mem_2135_sv2v_reg ,\nz.mem_2134_sv2v_reg ,\nz.mem_2133_sv2v_reg ,
  \nz.mem_2132_sv2v_reg ,\nz.mem_2131_sv2v_reg ,\nz.mem_2130_sv2v_reg ,\nz.mem_2129_sv2v_reg ,
  \nz.mem_2128_sv2v_reg ,\nz.mem_2127_sv2v_reg ,\nz.mem_2126_sv2v_reg ,
  \nz.mem_2125_sv2v_reg ,\nz.mem_2124_sv2v_reg ,\nz.mem_2123_sv2v_reg ,\nz.mem_2122_sv2v_reg ,
  \nz.mem_2121_sv2v_reg ,\nz.mem_2120_sv2v_reg ,\nz.mem_2119_sv2v_reg ,
  \nz.mem_2118_sv2v_reg ,\nz.mem_2117_sv2v_reg ,\nz.mem_2116_sv2v_reg ,\nz.mem_2115_sv2v_reg ,
  \nz.mem_2114_sv2v_reg ,\nz.mem_2113_sv2v_reg ,\nz.mem_2112_sv2v_reg ,
  \nz.mem_2111_sv2v_reg ,\nz.mem_2110_sv2v_reg ,\nz.mem_2109_sv2v_reg ,\nz.mem_2108_sv2v_reg ,
  \nz.mem_2107_sv2v_reg ,\nz.mem_2106_sv2v_reg ,\nz.mem_2105_sv2v_reg ,
  \nz.mem_2104_sv2v_reg ,\nz.mem_2103_sv2v_reg ,\nz.mem_2102_sv2v_reg ,\nz.mem_2101_sv2v_reg ,
  \nz.mem_2100_sv2v_reg ,\nz.mem_2099_sv2v_reg ,\nz.mem_2098_sv2v_reg ,
  \nz.mem_2097_sv2v_reg ,\nz.mem_2096_sv2v_reg ,\nz.mem_2095_sv2v_reg ,\nz.mem_2094_sv2v_reg ,
  \nz.mem_2093_sv2v_reg ,\nz.mem_2092_sv2v_reg ,\nz.mem_2091_sv2v_reg ,
  \nz.mem_2090_sv2v_reg ,\nz.mem_2089_sv2v_reg ,\nz.mem_2088_sv2v_reg ,\nz.mem_2087_sv2v_reg ,
  \nz.mem_2086_sv2v_reg ,\nz.mem_2085_sv2v_reg ,\nz.mem_2084_sv2v_reg ,
  \nz.mem_2083_sv2v_reg ,\nz.mem_2082_sv2v_reg ,\nz.mem_2081_sv2v_reg ,\nz.mem_2080_sv2v_reg ,
  \nz.mem_2079_sv2v_reg ,\nz.mem_2078_sv2v_reg ,\nz.mem_2077_sv2v_reg ,
  \nz.mem_2076_sv2v_reg ,\nz.mem_2075_sv2v_reg ,\nz.mem_2074_sv2v_reg ,
  \nz.mem_2073_sv2v_reg ,\nz.mem_2072_sv2v_reg ,\nz.mem_2071_sv2v_reg ,\nz.mem_2070_sv2v_reg ,
  \nz.mem_2069_sv2v_reg ,\nz.mem_2068_sv2v_reg ,\nz.mem_2067_sv2v_reg ,
  \nz.mem_2066_sv2v_reg ,\nz.mem_2065_sv2v_reg ,\nz.mem_2064_sv2v_reg ,\nz.mem_2063_sv2v_reg ,
  \nz.mem_2062_sv2v_reg ,\nz.mem_2061_sv2v_reg ,\nz.mem_2060_sv2v_reg ,
  \nz.mem_2059_sv2v_reg ,\nz.mem_2058_sv2v_reg ,\nz.mem_2057_sv2v_reg ,\nz.mem_2056_sv2v_reg ,
  \nz.mem_2055_sv2v_reg ,\nz.mem_2054_sv2v_reg ,\nz.mem_2053_sv2v_reg ,
  \nz.mem_2052_sv2v_reg ,\nz.mem_2051_sv2v_reg ,\nz.mem_2050_sv2v_reg ,\nz.mem_2049_sv2v_reg ,
  \nz.mem_2048_sv2v_reg ,\nz.mem_2047_sv2v_reg ,\nz.mem_2046_sv2v_reg ,
  \nz.mem_2045_sv2v_reg ,\nz.mem_2044_sv2v_reg ,\nz.mem_2043_sv2v_reg ,\nz.mem_2042_sv2v_reg ,
  \nz.mem_2041_sv2v_reg ,\nz.mem_2040_sv2v_reg ,\nz.mem_2039_sv2v_reg ,
  \nz.mem_2038_sv2v_reg ,\nz.mem_2037_sv2v_reg ,\nz.mem_2036_sv2v_reg ,\nz.mem_2035_sv2v_reg ,
  \nz.mem_2034_sv2v_reg ,\nz.mem_2033_sv2v_reg ,\nz.mem_2032_sv2v_reg ,
  \nz.mem_2031_sv2v_reg ,\nz.mem_2030_sv2v_reg ,\nz.mem_2029_sv2v_reg ,\nz.mem_2028_sv2v_reg ,
  \nz.mem_2027_sv2v_reg ,\nz.mem_2026_sv2v_reg ,\nz.mem_2025_sv2v_reg ,
  \nz.mem_2024_sv2v_reg ,\nz.mem_2023_sv2v_reg ,\nz.mem_2022_sv2v_reg ,\nz.mem_2021_sv2v_reg ,
  \nz.mem_2020_sv2v_reg ,\nz.mem_2019_sv2v_reg ,\nz.mem_2018_sv2v_reg ,
  \nz.mem_2017_sv2v_reg ,\nz.mem_2016_sv2v_reg ,\nz.mem_2015_sv2v_reg ,\nz.mem_2014_sv2v_reg ,
  \nz.mem_2013_sv2v_reg ,\nz.mem_2012_sv2v_reg ,\nz.mem_2011_sv2v_reg ,
  \nz.mem_2010_sv2v_reg ,\nz.mem_2009_sv2v_reg ,\nz.mem_2008_sv2v_reg ,\nz.mem_2007_sv2v_reg ,
  \nz.mem_2006_sv2v_reg ,\nz.mem_2005_sv2v_reg ,\nz.mem_2004_sv2v_reg ,
  \nz.mem_2003_sv2v_reg ,\nz.mem_2002_sv2v_reg ,\nz.mem_2001_sv2v_reg ,\nz.mem_2000_sv2v_reg ,
  \nz.mem_1999_sv2v_reg ,\nz.mem_1998_sv2v_reg ,\nz.mem_1997_sv2v_reg ,
  \nz.mem_1996_sv2v_reg ,\nz.mem_1995_sv2v_reg ,\nz.mem_1994_sv2v_reg ,
  \nz.mem_1993_sv2v_reg ,\nz.mem_1992_sv2v_reg ,\nz.mem_1991_sv2v_reg ,\nz.mem_1990_sv2v_reg ,
  \nz.mem_1989_sv2v_reg ,\nz.mem_1988_sv2v_reg ,\nz.mem_1987_sv2v_reg ,
  \nz.mem_1986_sv2v_reg ,\nz.mem_1985_sv2v_reg ,\nz.mem_1984_sv2v_reg ,\nz.mem_1983_sv2v_reg ,
  \nz.mem_1982_sv2v_reg ,\nz.mem_1981_sv2v_reg ,\nz.mem_1980_sv2v_reg ,
  \nz.mem_1979_sv2v_reg ,\nz.mem_1978_sv2v_reg ,\nz.mem_1977_sv2v_reg ,\nz.mem_1976_sv2v_reg ,
  \nz.mem_1975_sv2v_reg ,\nz.mem_1974_sv2v_reg ,\nz.mem_1973_sv2v_reg ,
  \nz.mem_1972_sv2v_reg ,\nz.mem_1971_sv2v_reg ,\nz.mem_1970_sv2v_reg ,\nz.mem_1969_sv2v_reg ,
  \nz.mem_1968_sv2v_reg ,\nz.mem_1967_sv2v_reg ,\nz.mem_1966_sv2v_reg ,
  \nz.mem_1965_sv2v_reg ,\nz.mem_1964_sv2v_reg ,\nz.mem_1963_sv2v_reg ,\nz.mem_1962_sv2v_reg ,
  \nz.mem_1961_sv2v_reg ,\nz.mem_1960_sv2v_reg ,\nz.mem_1959_sv2v_reg ,
  \nz.mem_1958_sv2v_reg ,\nz.mem_1957_sv2v_reg ,\nz.mem_1956_sv2v_reg ,\nz.mem_1955_sv2v_reg ,
  \nz.mem_1954_sv2v_reg ,\nz.mem_1953_sv2v_reg ,\nz.mem_1952_sv2v_reg ,
  \nz.mem_1951_sv2v_reg ,\nz.mem_1950_sv2v_reg ,\nz.mem_1949_sv2v_reg ,\nz.mem_1948_sv2v_reg ,
  \nz.mem_1947_sv2v_reg ,\nz.mem_1946_sv2v_reg ,\nz.mem_1945_sv2v_reg ,
  \nz.mem_1944_sv2v_reg ,\nz.mem_1943_sv2v_reg ,\nz.mem_1942_sv2v_reg ,\nz.mem_1941_sv2v_reg ,
  \nz.mem_1940_sv2v_reg ,\nz.mem_1939_sv2v_reg ,\nz.mem_1938_sv2v_reg ,
  \nz.mem_1937_sv2v_reg ,\nz.mem_1936_sv2v_reg ,\nz.mem_1935_sv2v_reg ,\nz.mem_1934_sv2v_reg ,
  \nz.mem_1933_sv2v_reg ,\nz.mem_1932_sv2v_reg ,\nz.mem_1931_sv2v_reg ,
  \nz.mem_1930_sv2v_reg ,\nz.mem_1929_sv2v_reg ,\nz.mem_1928_sv2v_reg ,\nz.mem_1927_sv2v_reg ,
  \nz.mem_1926_sv2v_reg ,\nz.mem_1925_sv2v_reg ,\nz.mem_1924_sv2v_reg ,
  \nz.mem_1923_sv2v_reg ,\nz.mem_1922_sv2v_reg ,\nz.mem_1921_sv2v_reg ,\nz.mem_1920_sv2v_reg ,
  \nz.mem_1919_sv2v_reg ,\nz.mem_1918_sv2v_reg ,\nz.mem_1917_sv2v_reg ,
  \nz.mem_1916_sv2v_reg ,\nz.mem_1915_sv2v_reg ,\nz.mem_1914_sv2v_reg ,
  \nz.mem_1913_sv2v_reg ,\nz.mem_1912_sv2v_reg ,\nz.mem_1911_sv2v_reg ,\nz.mem_1910_sv2v_reg ,
  \nz.mem_1909_sv2v_reg ,\nz.mem_1908_sv2v_reg ,\nz.mem_1907_sv2v_reg ,
  \nz.mem_1906_sv2v_reg ,\nz.mem_1905_sv2v_reg ,\nz.mem_1904_sv2v_reg ,\nz.mem_1903_sv2v_reg ,
  \nz.mem_1902_sv2v_reg ,\nz.mem_1901_sv2v_reg ,\nz.mem_1900_sv2v_reg ,
  \nz.mem_1899_sv2v_reg ,\nz.mem_1898_sv2v_reg ,\nz.mem_1897_sv2v_reg ,\nz.mem_1896_sv2v_reg ,
  \nz.mem_1895_sv2v_reg ,\nz.mem_1894_sv2v_reg ,\nz.mem_1893_sv2v_reg ,
  \nz.mem_1892_sv2v_reg ,\nz.mem_1891_sv2v_reg ,\nz.mem_1890_sv2v_reg ,\nz.mem_1889_sv2v_reg ,
  \nz.mem_1888_sv2v_reg ,\nz.mem_1887_sv2v_reg ,\nz.mem_1886_sv2v_reg ,
  \nz.mem_1885_sv2v_reg ,\nz.mem_1884_sv2v_reg ,\nz.mem_1883_sv2v_reg ,\nz.mem_1882_sv2v_reg ,
  \nz.mem_1881_sv2v_reg ,\nz.mem_1880_sv2v_reg ,\nz.mem_1879_sv2v_reg ,
  \nz.mem_1878_sv2v_reg ,\nz.mem_1877_sv2v_reg ,\nz.mem_1876_sv2v_reg ,\nz.mem_1875_sv2v_reg ,
  \nz.mem_1874_sv2v_reg ,\nz.mem_1873_sv2v_reg ,\nz.mem_1872_sv2v_reg ,
  \nz.mem_1871_sv2v_reg ,\nz.mem_1870_sv2v_reg ,\nz.mem_1869_sv2v_reg ,\nz.mem_1868_sv2v_reg ,
  \nz.mem_1867_sv2v_reg ,\nz.mem_1866_sv2v_reg ,\nz.mem_1865_sv2v_reg ,
  \nz.mem_1864_sv2v_reg ,\nz.mem_1863_sv2v_reg ,\nz.mem_1862_sv2v_reg ,\nz.mem_1861_sv2v_reg ,
  \nz.mem_1860_sv2v_reg ,\nz.mem_1859_sv2v_reg ,\nz.mem_1858_sv2v_reg ,
  \nz.mem_1857_sv2v_reg ,\nz.mem_1856_sv2v_reg ,\nz.mem_1855_sv2v_reg ,\nz.mem_1854_sv2v_reg ,
  \nz.mem_1853_sv2v_reg ,\nz.mem_1852_sv2v_reg ,\nz.mem_1851_sv2v_reg ,
  \nz.mem_1850_sv2v_reg ,\nz.mem_1849_sv2v_reg ,\nz.mem_1848_sv2v_reg ,\nz.mem_1847_sv2v_reg ,
  \nz.mem_1846_sv2v_reg ,\nz.mem_1845_sv2v_reg ,\nz.mem_1844_sv2v_reg ,
  \nz.mem_1843_sv2v_reg ,\nz.mem_1842_sv2v_reg ,\nz.mem_1841_sv2v_reg ,\nz.mem_1840_sv2v_reg ,
  \nz.mem_1839_sv2v_reg ,\nz.mem_1838_sv2v_reg ,\nz.mem_1837_sv2v_reg ,
  \nz.mem_1836_sv2v_reg ,\nz.mem_1835_sv2v_reg ,\nz.mem_1834_sv2v_reg ,
  \nz.mem_1833_sv2v_reg ,\nz.mem_1832_sv2v_reg ,\nz.mem_1831_sv2v_reg ,\nz.mem_1830_sv2v_reg ,
  \nz.mem_1829_sv2v_reg ,\nz.mem_1828_sv2v_reg ,\nz.mem_1827_sv2v_reg ,
  \nz.mem_1826_sv2v_reg ,\nz.mem_1825_sv2v_reg ,\nz.mem_1824_sv2v_reg ,\nz.mem_1823_sv2v_reg ,
  \nz.mem_1822_sv2v_reg ,\nz.mem_1821_sv2v_reg ,\nz.mem_1820_sv2v_reg ,
  \nz.mem_1819_sv2v_reg ,\nz.mem_1818_sv2v_reg ,\nz.mem_1817_sv2v_reg ,\nz.mem_1816_sv2v_reg ,
  \nz.mem_1815_sv2v_reg ,\nz.mem_1814_sv2v_reg ,\nz.mem_1813_sv2v_reg ,
  \nz.mem_1812_sv2v_reg ,\nz.mem_1811_sv2v_reg ,\nz.mem_1810_sv2v_reg ,\nz.mem_1809_sv2v_reg ,
  \nz.mem_1808_sv2v_reg ,\nz.mem_1807_sv2v_reg ,\nz.mem_1806_sv2v_reg ,
  \nz.mem_1805_sv2v_reg ,\nz.mem_1804_sv2v_reg ,\nz.mem_1803_sv2v_reg ,\nz.mem_1802_sv2v_reg ,
  \nz.mem_1801_sv2v_reg ,\nz.mem_1800_sv2v_reg ,\nz.mem_1799_sv2v_reg ,
  \nz.mem_1798_sv2v_reg ,\nz.mem_1797_sv2v_reg ,\nz.mem_1796_sv2v_reg ,\nz.mem_1795_sv2v_reg ,
  \nz.mem_1794_sv2v_reg ,\nz.mem_1793_sv2v_reg ,\nz.mem_1792_sv2v_reg ,
  \nz.mem_1791_sv2v_reg ,\nz.mem_1790_sv2v_reg ,\nz.mem_1789_sv2v_reg ,\nz.mem_1788_sv2v_reg ,
  \nz.mem_1787_sv2v_reg ,\nz.mem_1786_sv2v_reg ,\nz.mem_1785_sv2v_reg ,
  \nz.mem_1784_sv2v_reg ,\nz.mem_1783_sv2v_reg ,\nz.mem_1782_sv2v_reg ,\nz.mem_1781_sv2v_reg ,
  \nz.mem_1780_sv2v_reg ,\nz.mem_1779_sv2v_reg ,\nz.mem_1778_sv2v_reg ,
  \nz.mem_1777_sv2v_reg ,\nz.mem_1776_sv2v_reg ,\nz.mem_1775_sv2v_reg ,\nz.mem_1774_sv2v_reg ,
  \nz.mem_1773_sv2v_reg ,\nz.mem_1772_sv2v_reg ,\nz.mem_1771_sv2v_reg ,
  \nz.mem_1770_sv2v_reg ,\nz.mem_1769_sv2v_reg ,\nz.mem_1768_sv2v_reg ,\nz.mem_1767_sv2v_reg ,
  \nz.mem_1766_sv2v_reg ,\nz.mem_1765_sv2v_reg ,\nz.mem_1764_sv2v_reg ,
  \nz.mem_1763_sv2v_reg ,\nz.mem_1762_sv2v_reg ,\nz.mem_1761_sv2v_reg ,\nz.mem_1760_sv2v_reg ,
  \nz.mem_1759_sv2v_reg ,\nz.mem_1758_sv2v_reg ,\nz.mem_1757_sv2v_reg ,
  \nz.mem_1756_sv2v_reg ,\nz.mem_1755_sv2v_reg ,\nz.mem_1754_sv2v_reg ,
  \nz.mem_1753_sv2v_reg ,\nz.mem_1752_sv2v_reg ,\nz.mem_1751_sv2v_reg ,\nz.mem_1750_sv2v_reg ,
  \nz.mem_1749_sv2v_reg ,\nz.mem_1748_sv2v_reg ,\nz.mem_1747_sv2v_reg ,
  \nz.mem_1746_sv2v_reg ,\nz.mem_1745_sv2v_reg ,\nz.mem_1744_sv2v_reg ,\nz.mem_1743_sv2v_reg ,
  \nz.mem_1742_sv2v_reg ,\nz.mem_1741_sv2v_reg ,\nz.mem_1740_sv2v_reg ,
  \nz.mem_1739_sv2v_reg ,\nz.mem_1738_sv2v_reg ,\nz.mem_1737_sv2v_reg ,\nz.mem_1736_sv2v_reg ,
  \nz.mem_1735_sv2v_reg ,\nz.mem_1734_sv2v_reg ,\nz.mem_1733_sv2v_reg ,
  \nz.mem_1732_sv2v_reg ,\nz.mem_1731_sv2v_reg ,\nz.mem_1730_sv2v_reg ,\nz.mem_1729_sv2v_reg ,
  \nz.mem_1728_sv2v_reg ,\nz.mem_1727_sv2v_reg ,\nz.mem_1726_sv2v_reg ,
  \nz.mem_1725_sv2v_reg ,\nz.mem_1724_sv2v_reg ,\nz.mem_1723_sv2v_reg ,\nz.mem_1722_sv2v_reg ,
  \nz.mem_1721_sv2v_reg ,\nz.mem_1720_sv2v_reg ,\nz.mem_1719_sv2v_reg ,
  \nz.mem_1718_sv2v_reg ,\nz.mem_1717_sv2v_reg ,\nz.mem_1716_sv2v_reg ,\nz.mem_1715_sv2v_reg ,
  \nz.mem_1714_sv2v_reg ,\nz.mem_1713_sv2v_reg ,\nz.mem_1712_sv2v_reg ,
  \nz.mem_1711_sv2v_reg ,\nz.mem_1710_sv2v_reg ,\nz.mem_1709_sv2v_reg ,\nz.mem_1708_sv2v_reg ,
  \nz.mem_1707_sv2v_reg ,\nz.mem_1706_sv2v_reg ,\nz.mem_1705_sv2v_reg ,
  \nz.mem_1704_sv2v_reg ,\nz.mem_1703_sv2v_reg ,\nz.mem_1702_sv2v_reg ,\nz.mem_1701_sv2v_reg ,
  \nz.mem_1700_sv2v_reg ,\nz.mem_1699_sv2v_reg ,\nz.mem_1698_sv2v_reg ,
  \nz.mem_1697_sv2v_reg ,\nz.mem_1696_sv2v_reg ,\nz.mem_1695_sv2v_reg ,\nz.mem_1694_sv2v_reg ,
  \nz.mem_1693_sv2v_reg ,\nz.mem_1692_sv2v_reg ,\nz.mem_1691_sv2v_reg ,
  \nz.mem_1690_sv2v_reg ,\nz.mem_1689_sv2v_reg ,\nz.mem_1688_sv2v_reg ,\nz.mem_1687_sv2v_reg ,
  \nz.mem_1686_sv2v_reg ,\nz.mem_1685_sv2v_reg ,\nz.mem_1684_sv2v_reg ,
  \nz.mem_1683_sv2v_reg ,\nz.mem_1682_sv2v_reg ,\nz.mem_1681_sv2v_reg ,\nz.mem_1680_sv2v_reg ,
  \nz.mem_1679_sv2v_reg ,\nz.mem_1678_sv2v_reg ,\nz.mem_1677_sv2v_reg ,
  \nz.mem_1676_sv2v_reg ,\nz.mem_1675_sv2v_reg ,\nz.mem_1674_sv2v_reg ,
  \nz.mem_1673_sv2v_reg ,\nz.mem_1672_sv2v_reg ,\nz.mem_1671_sv2v_reg ,\nz.mem_1670_sv2v_reg ,
  \nz.mem_1669_sv2v_reg ,\nz.mem_1668_sv2v_reg ,\nz.mem_1667_sv2v_reg ,
  \nz.mem_1666_sv2v_reg ,\nz.mem_1665_sv2v_reg ,\nz.mem_1664_sv2v_reg ,\nz.mem_1663_sv2v_reg ,
  \nz.mem_1662_sv2v_reg ,\nz.mem_1661_sv2v_reg ,\nz.mem_1660_sv2v_reg ,
  \nz.mem_1659_sv2v_reg ,\nz.mem_1658_sv2v_reg ,\nz.mem_1657_sv2v_reg ,\nz.mem_1656_sv2v_reg ,
  \nz.mem_1655_sv2v_reg ,\nz.mem_1654_sv2v_reg ,\nz.mem_1653_sv2v_reg ,
  \nz.mem_1652_sv2v_reg ,\nz.mem_1651_sv2v_reg ,\nz.mem_1650_sv2v_reg ,\nz.mem_1649_sv2v_reg ,
  \nz.mem_1648_sv2v_reg ,\nz.mem_1647_sv2v_reg ,\nz.mem_1646_sv2v_reg ,
  \nz.mem_1645_sv2v_reg ,\nz.mem_1644_sv2v_reg ,\nz.mem_1643_sv2v_reg ,\nz.mem_1642_sv2v_reg ,
  \nz.mem_1641_sv2v_reg ,\nz.mem_1640_sv2v_reg ,\nz.mem_1639_sv2v_reg ,
  \nz.mem_1638_sv2v_reg ,\nz.mem_1637_sv2v_reg ,\nz.mem_1636_sv2v_reg ,\nz.mem_1635_sv2v_reg ,
  \nz.mem_1634_sv2v_reg ,\nz.mem_1633_sv2v_reg ,\nz.mem_1632_sv2v_reg ,
  \nz.mem_1631_sv2v_reg ,\nz.mem_1630_sv2v_reg ,\nz.mem_1629_sv2v_reg ,\nz.mem_1628_sv2v_reg ,
  \nz.mem_1627_sv2v_reg ,\nz.mem_1626_sv2v_reg ,\nz.mem_1625_sv2v_reg ,
  \nz.mem_1624_sv2v_reg ,\nz.mem_1623_sv2v_reg ,\nz.mem_1622_sv2v_reg ,\nz.mem_1621_sv2v_reg ,
  \nz.mem_1620_sv2v_reg ,\nz.mem_1619_sv2v_reg ,\nz.mem_1618_sv2v_reg ,
  \nz.mem_1617_sv2v_reg ,\nz.mem_1616_sv2v_reg ,\nz.mem_1615_sv2v_reg ,\nz.mem_1614_sv2v_reg ,
  \nz.mem_1613_sv2v_reg ,\nz.mem_1612_sv2v_reg ,\nz.mem_1611_sv2v_reg ,
  \nz.mem_1610_sv2v_reg ,\nz.mem_1609_sv2v_reg ,\nz.mem_1608_sv2v_reg ,\nz.mem_1607_sv2v_reg ,
  \nz.mem_1606_sv2v_reg ,\nz.mem_1605_sv2v_reg ,\nz.mem_1604_sv2v_reg ,
  \nz.mem_1603_sv2v_reg ,\nz.mem_1602_sv2v_reg ,\nz.mem_1601_sv2v_reg ,\nz.mem_1600_sv2v_reg ,
  \nz.mem_1599_sv2v_reg ,\nz.mem_1598_sv2v_reg ,\nz.mem_1597_sv2v_reg ,
  \nz.mem_1596_sv2v_reg ,\nz.mem_1595_sv2v_reg ,\nz.mem_1594_sv2v_reg ,
  \nz.mem_1593_sv2v_reg ,\nz.mem_1592_sv2v_reg ,\nz.mem_1591_sv2v_reg ,\nz.mem_1590_sv2v_reg ,
  \nz.mem_1589_sv2v_reg ,\nz.mem_1588_sv2v_reg ,\nz.mem_1587_sv2v_reg ,
  \nz.mem_1586_sv2v_reg ,\nz.mem_1585_sv2v_reg ,\nz.mem_1584_sv2v_reg ,\nz.mem_1583_sv2v_reg ,
  \nz.mem_1582_sv2v_reg ,\nz.mem_1581_sv2v_reg ,\nz.mem_1580_sv2v_reg ,
  \nz.mem_1579_sv2v_reg ,\nz.mem_1578_sv2v_reg ,\nz.mem_1577_sv2v_reg ,\nz.mem_1576_sv2v_reg ,
  \nz.mem_1575_sv2v_reg ,\nz.mem_1574_sv2v_reg ,\nz.mem_1573_sv2v_reg ,
  \nz.mem_1572_sv2v_reg ,\nz.mem_1571_sv2v_reg ,\nz.mem_1570_sv2v_reg ,\nz.mem_1569_sv2v_reg ,
  \nz.mem_1568_sv2v_reg ,\nz.mem_1567_sv2v_reg ,\nz.mem_1566_sv2v_reg ,
  \nz.mem_1565_sv2v_reg ,\nz.mem_1564_sv2v_reg ,\nz.mem_1563_sv2v_reg ,\nz.mem_1562_sv2v_reg ,
  \nz.mem_1561_sv2v_reg ,\nz.mem_1560_sv2v_reg ,\nz.mem_1559_sv2v_reg ,
  \nz.mem_1558_sv2v_reg ,\nz.mem_1557_sv2v_reg ,\nz.mem_1556_sv2v_reg ,\nz.mem_1555_sv2v_reg ,
  \nz.mem_1554_sv2v_reg ,\nz.mem_1553_sv2v_reg ,\nz.mem_1552_sv2v_reg ,
  \nz.mem_1551_sv2v_reg ,\nz.mem_1550_sv2v_reg ,\nz.mem_1549_sv2v_reg ,\nz.mem_1548_sv2v_reg ,
  \nz.mem_1547_sv2v_reg ,\nz.mem_1546_sv2v_reg ,\nz.mem_1545_sv2v_reg ,
  \nz.mem_1544_sv2v_reg ,\nz.mem_1543_sv2v_reg ,\nz.mem_1542_sv2v_reg ,\nz.mem_1541_sv2v_reg ,
  \nz.mem_1540_sv2v_reg ,\nz.mem_1539_sv2v_reg ,\nz.mem_1538_sv2v_reg ,
  \nz.mem_1537_sv2v_reg ,\nz.mem_1536_sv2v_reg ,\nz.mem_1535_sv2v_reg ,\nz.mem_1534_sv2v_reg ,
  \nz.mem_1533_sv2v_reg ,\nz.mem_1532_sv2v_reg ,\nz.mem_1531_sv2v_reg ,
  \nz.mem_1530_sv2v_reg ,\nz.mem_1529_sv2v_reg ,\nz.mem_1528_sv2v_reg ,\nz.mem_1527_sv2v_reg ,
  \nz.mem_1526_sv2v_reg ,\nz.mem_1525_sv2v_reg ,\nz.mem_1524_sv2v_reg ,
  \nz.mem_1523_sv2v_reg ,\nz.mem_1522_sv2v_reg ,\nz.mem_1521_sv2v_reg ,\nz.mem_1520_sv2v_reg ,
  \nz.mem_1519_sv2v_reg ,\nz.mem_1518_sv2v_reg ,\nz.mem_1517_sv2v_reg ,
  \nz.mem_1516_sv2v_reg ,\nz.mem_1515_sv2v_reg ,\nz.mem_1514_sv2v_reg ,
  \nz.mem_1513_sv2v_reg ,\nz.mem_1512_sv2v_reg ,\nz.mem_1511_sv2v_reg ,\nz.mem_1510_sv2v_reg ,
  \nz.mem_1509_sv2v_reg ,\nz.mem_1508_sv2v_reg ,\nz.mem_1507_sv2v_reg ,
  \nz.mem_1506_sv2v_reg ,\nz.mem_1505_sv2v_reg ,\nz.mem_1504_sv2v_reg ,\nz.mem_1503_sv2v_reg ,
  \nz.mem_1502_sv2v_reg ,\nz.mem_1501_sv2v_reg ,\nz.mem_1500_sv2v_reg ,
  \nz.mem_1499_sv2v_reg ,\nz.mem_1498_sv2v_reg ,\nz.mem_1497_sv2v_reg ,\nz.mem_1496_sv2v_reg ,
  \nz.mem_1495_sv2v_reg ,\nz.mem_1494_sv2v_reg ,\nz.mem_1493_sv2v_reg ,
  \nz.mem_1492_sv2v_reg ,\nz.mem_1491_sv2v_reg ,\nz.mem_1490_sv2v_reg ,\nz.mem_1489_sv2v_reg ,
  \nz.mem_1488_sv2v_reg ,\nz.mem_1487_sv2v_reg ,\nz.mem_1486_sv2v_reg ,
  \nz.mem_1485_sv2v_reg ,\nz.mem_1484_sv2v_reg ,\nz.mem_1483_sv2v_reg ,\nz.mem_1482_sv2v_reg ,
  \nz.mem_1481_sv2v_reg ,\nz.mem_1480_sv2v_reg ,\nz.mem_1479_sv2v_reg ,
  \nz.mem_1478_sv2v_reg ,\nz.mem_1477_sv2v_reg ,\nz.mem_1476_sv2v_reg ,\nz.mem_1475_sv2v_reg ,
  \nz.mem_1474_sv2v_reg ,\nz.mem_1473_sv2v_reg ,\nz.mem_1472_sv2v_reg ,
  \nz.mem_1471_sv2v_reg ,\nz.mem_1470_sv2v_reg ,\nz.mem_1469_sv2v_reg ,\nz.mem_1468_sv2v_reg ,
  \nz.mem_1467_sv2v_reg ,\nz.mem_1466_sv2v_reg ,\nz.mem_1465_sv2v_reg ,
  \nz.mem_1464_sv2v_reg ,\nz.mem_1463_sv2v_reg ,\nz.mem_1462_sv2v_reg ,\nz.mem_1461_sv2v_reg ,
  \nz.mem_1460_sv2v_reg ,\nz.mem_1459_sv2v_reg ,\nz.mem_1458_sv2v_reg ,
  \nz.mem_1457_sv2v_reg ,\nz.mem_1456_sv2v_reg ,\nz.mem_1455_sv2v_reg ,\nz.mem_1454_sv2v_reg ,
  \nz.mem_1453_sv2v_reg ,\nz.mem_1452_sv2v_reg ,\nz.mem_1451_sv2v_reg ,
  \nz.mem_1450_sv2v_reg ,\nz.mem_1449_sv2v_reg ,\nz.mem_1448_sv2v_reg ,\nz.mem_1447_sv2v_reg ,
  \nz.mem_1446_sv2v_reg ,\nz.mem_1445_sv2v_reg ,\nz.mem_1444_sv2v_reg ,
  \nz.mem_1443_sv2v_reg ,\nz.mem_1442_sv2v_reg ,\nz.mem_1441_sv2v_reg ,\nz.mem_1440_sv2v_reg ,
  \nz.mem_1439_sv2v_reg ,\nz.mem_1438_sv2v_reg ,\nz.mem_1437_sv2v_reg ,
  \nz.mem_1436_sv2v_reg ,\nz.mem_1435_sv2v_reg ,\nz.mem_1434_sv2v_reg ,
  \nz.mem_1433_sv2v_reg ,\nz.mem_1432_sv2v_reg ,\nz.mem_1431_sv2v_reg ,\nz.mem_1430_sv2v_reg ,
  \nz.mem_1429_sv2v_reg ,\nz.mem_1428_sv2v_reg ,\nz.mem_1427_sv2v_reg ,
  \nz.mem_1426_sv2v_reg ,\nz.mem_1425_sv2v_reg ,\nz.mem_1424_sv2v_reg ,\nz.mem_1423_sv2v_reg ,
  \nz.mem_1422_sv2v_reg ,\nz.mem_1421_sv2v_reg ,\nz.mem_1420_sv2v_reg ,
  \nz.mem_1419_sv2v_reg ,\nz.mem_1418_sv2v_reg ,\nz.mem_1417_sv2v_reg ,\nz.mem_1416_sv2v_reg ,
  \nz.mem_1415_sv2v_reg ,\nz.mem_1414_sv2v_reg ,\nz.mem_1413_sv2v_reg ,
  \nz.mem_1412_sv2v_reg ,\nz.mem_1411_sv2v_reg ,\nz.mem_1410_sv2v_reg ,\nz.mem_1409_sv2v_reg ,
  \nz.mem_1408_sv2v_reg ,\nz.mem_1407_sv2v_reg ,\nz.mem_1406_sv2v_reg ,
  \nz.mem_1405_sv2v_reg ,\nz.mem_1404_sv2v_reg ,\nz.mem_1403_sv2v_reg ,\nz.mem_1402_sv2v_reg ,
  \nz.mem_1401_sv2v_reg ,\nz.mem_1400_sv2v_reg ,\nz.mem_1399_sv2v_reg ,
  \nz.mem_1398_sv2v_reg ,\nz.mem_1397_sv2v_reg ,\nz.mem_1396_sv2v_reg ,\nz.mem_1395_sv2v_reg ,
  \nz.mem_1394_sv2v_reg ,\nz.mem_1393_sv2v_reg ,\nz.mem_1392_sv2v_reg ,
  \nz.mem_1391_sv2v_reg ,\nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,\nz.mem_1388_sv2v_reg ,
  \nz.mem_1387_sv2v_reg ,\nz.mem_1386_sv2v_reg ,\nz.mem_1385_sv2v_reg ,
  \nz.mem_1384_sv2v_reg ,\nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,\nz.mem_1381_sv2v_reg ,
  \nz.mem_1380_sv2v_reg ,\nz.mem_1379_sv2v_reg ,\nz.mem_1378_sv2v_reg ,
  \nz.mem_1377_sv2v_reg ,\nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,\nz.mem_1374_sv2v_reg ,
  \nz.mem_1373_sv2v_reg ,\nz.mem_1372_sv2v_reg ,\nz.mem_1371_sv2v_reg ,
  \nz.mem_1370_sv2v_reg ,\nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,\nz.mem_1367_sv2v_reg ,
  \nz.mem_1366_sv2v_reg ,\nz.mem_1365_sv2v_reg ,\nz.mem_1364_sv2v_reg ,
  \nz.mem_1363_sv2v_reg ,\nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,\nz.mem_1360_sv2v_reg ,
  \nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,\nz.mem_1357_sv2v_reg ,
  \nz.mem_1356_sv2v_reg ,\nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,
  \nz.mem_1353_sv2v_reg ,\nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,\nz.mem_1350_sv2v_reg ,
  \nz.mem_1349_sv2v_reg ,\nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,
  \nz.mem_1346_sv2v_reg ,\nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,\nz.mem_1343_sv2v_reg ,
  \nz.mem_1342_sv2v_reg ,\nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,
  \nz.mem_1339_sv2v_reg ,\nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,\nz.mem_1336_sv2v_reg ,
  \nz.mem_1335_sv2v_reg ,\nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,
  \nz.mem_1332_sv2v_reg ,\nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,\nz.mem_1329_sv2v_reg ,
  \nz.mem_1328_sv2v_reg ,\nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,
  \nz.mem_1325_sv2v_reg ,\nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,\nz.mem_1322_sv2v_reg ,
  \nz.mem_1321_sv2v_reg ,\nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,
  \nz.mem_1318_sv2v_reg ,\nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,\nz.mem_1315_sv2v_reg ,
  \nz.mem_1314_sv2v_reg ,\nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,
  \nz.mem_1311_sv2v_reg ,\nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,\nz.mem_1308_sv2v_reg ,
  \nz.mem_1307_sv2v_reg ,\nz.mem_1306_sv2v_reg ,\nz.mem_1305_sv2v_reg ,
  \nz.mem_1304_sv2v_reg ,\nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,\nz.mem_1301_sv2v_reg ,
  \nz.mem_1300_sv2v_reg ,\nz.mem_1299_sv2v_reg ,\nz.mem_1298_sv2v_reg ,
  \nz.mem_1297_sv2v_reg ,\nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,\nz.mem_1294_sv2v_reg ,
  \nz.mem_1293_sv2v_reg ,\nz.mem_1292_sv2v_reg ,\nz.mem_1291_sv2v_reg ,
  \nz.mem_1290_sv2v_reg ,\nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,\nz.mem_1287_sv2v_reg ,
  \nz.mem_1286_sv2v_reg ,\nz.mem_1285_sv2v_reg ,\nz.mem_1284_sv2v_reg ,
  \nz.mem_1283_sv2v_reg ,\nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,\nz.mem_1280_sv2v_reg ,
  \nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,\nz.mem_1277_sv2v_reg ,
  \nz.mem_1276_sv2v_reg ,\nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,
  \nz.mem_1273_sv2v_reg ,\nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,\nz.mem_1270_sv2v_reg ,
  \nz.mem_1269_sv2v_reg ,\nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,
  \nz.mem_1266_sv2v_reg ,\nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,\nz.mem_1263_sv2v_reg ,
  \nz.mem_1262_sv2v_reg ,\nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,
  \nz.mem_1259_sv2v_reg ,\nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,\nz.mem_1256_sv2v_reg ,
  \nz.mem_1255_sv2v_reg ,\nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,
  \nz.mem_1252_sv2v_reg ,\nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,\nz.mem_1249_sv2v_reg ,
  \nz.mem_1248_sv2v_reg ,\nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,
  \nz.mem_1245_sv2v_reg ,\nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,\nz.mem_1242_sv2v_reg ,
  \nz.mem_1241_sv2v_reg ,\nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,
  \nz.mem_1238_sv2v_reg ,\nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,\nz.mem_1235_sv2v_reg ,
  \nz.mem_1234_sv2v_reg ,\nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,
  \nz.mem_1231_sv2v_reg ,\nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,\nz.mem_1228_sv2v_reg ,
  \nz.mem_1227_sv2v_reg ,\nz.mem_1226_sv2v_reg ,\nz.mem_1225_sv2v_reg ,
  \nz.mem_1224_sv2v_reg ,\nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,\nz.mem_1221_sv2v_reg ,
  \nz.mem_1220_sv2v_reg ,\nz.mem_1219_sv2v_reg ,\nz.mem_1218_sv2v_reg ,
  \nz.mem_1217_sv2v_reg ,\nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,\nz.mem_1214_sv2v_reg ,
  \nz.mem_1213_sv2v_reg ,\nz.mem_1212_sv2v_reg ,\nz.mem_1211_sv2v_reg ,
  \nz.mem_1210_sv2v_reg ,\nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,\nz.mem_1207_sv2v_reg ,
  \nz.mem_1206_sv2v_reg ,\nz.mem_1205_sv2v_reg ,\nz.mem_1204_sv2v_reg ,
  \nz.mem_1203_sv2v_reg ,\nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,\nz.mem_1200_sv2v_reg ,
  \nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,\nz.mem_1197_sv2v_reg ,
  \nz.mem_1196_sv2v_reg ,\nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,
  \nz.mem_1193_sv2v_reg ,\nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,\nz.mem_1190_sv2v_reg ,
  \nz.mem_1189_sv2v_reg ,\nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,
  \nz.mem_1186_sv2v_reg ,\nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,\nz.mem_1183_sv2v_reg ,
  \nz.mem_1182_sv2v_reg ,\nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,
  \nz.mem_1179_sv2v_reg ,\nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,\nz.mem_1176_sv2v_reg ,
  \nz.mem_1175_sv2v_reg ,\nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,
  \nz.mem_1172_sv2v_reg ,\nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,\nz.mem_1169_sv2v_reg ,
  \nz.mem_1168_sv2v_reg ,\nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,
  \nz.mem_1165_sv2v_reg ,\nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,\nz.mem_1162_sv2v_reg ,
  \nz.mem_1161_sv2v_reg ,\nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,
  \nz.mem_1158_sv2v_reg ,\nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,\nz.mem_1155_sv2v_reg ,
  \nz.mem_1154_sv2v_reg ,\nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,
  \nz.mem_1151_sv2v_reg ,\nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,\nz.mem_1148_sv2v_reg ,
  \nz.mem_1147_sv2v_reg ,\nz.mem_1146_sv2v_reg ,\nz.mem_1145_sv2v_reg ,
  \nz.mem_1144_sv2v_reg ,\nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,\nz.mem_1141_sv2v_reg ,
  \nz.mem_1140_sv2v_reg ,\nz.mem_1139_sv2v_reg ,\nz.mem_1138_sv2v_reg ,
  \nz.mem_1137_sv2v_reg ,\nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,\nz.mem_1134_sv2v_reg ,
  \nz.mem_1133_sv2v_reg ,\nz.mem_1132_sv2v_reg ,\nz.mem_1131_sv2v_reg ,
  \nz.mem_1130_sv2v_reg ,\nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,\nz.mem_1127_sv2v_reg ,
  \nz.mem_1126_sv2v_reg ,\nz.mem_1125_sv2v_reg ,\nz.mem_1124_sv2v_reg ,
  \nz.mem_1123_sv2v_reg ,\nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,\nz.mem_1120_sv2v_reg ,
  \nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,\nz.mem_1117_sv2v_reg ,
  \nz.mem_1116_sv2v_reg ,\nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,
  \nz.mem_1113_sv2v_reg ,\nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,\nz.mem_1110_sv2v_reg ,
  \nz.mem_1109_sv2v_reg ,\nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,
  \nz.mem_1106_sv2v_reg ,\nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,\nz.mem_1103_sv2v_reg ,
  \nz.mem_1102_sv2v_reg ,\nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,
  \nz.mem_1099_sv2v_reg ,\nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,\nz.mem_1096_sv2v_reg ,
  \nz.mem_1095_sv2v_reg ,\nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,
  \nz.mem_1092_sv2v_reg ,\nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,\nz.mem_1089_sv2v_reg ,
  \nz.mem_1088_sv2v_reg ,\nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,
  \nz.mem_1085_sv2v_reg ,\nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,\nz.mem_1082_sv2v_reg ,
  \nz.mem_1081_sv2v_reg ,\nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,
  \nz.mem_1078_sv2v_reg ,\nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,\nz.mem_1075_sv2v_reg ,
  \nz.mem_1074_sv2v_reg ,\nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,
  \nz.mem_1071_sv2v_reg ,\nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,\nz.mem_1068_sv2v_reg ,
  \nz.mem_1067_sv2v_reg ,\nz.mem_1066_sv2v_reg ,\nz.mem_1065_sv2v_reg ,
  \nz.mem_1064_sv2v_reg ,\nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,\nz.mem_1061_sv2v_reg ,
  \nz.mem_1060_sv2v_reg ,\nz.mem_1059_sv2v_reg ,\nz.mem_1058_sv2v_reg ,
  \nz.mem_1057_sv2v_reg ,\nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,\nz.mem_1054_sv2v_reg ,
  \nz.mem_1053_sv2v_reg ,\nz.mem_1052_sv2v_reg ,\nz.mem_1051_sv2v_reg ,
  \nz.mem_1050_sv2v_reg ,\nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,\nz.mem_1047_sv2v_reg ,
  \nz.mem_1046_sv2v_reg ,\nz.mem_1045_sv2v_reg ,\nz.mem_1044_sv2v_reg ,
  \nz.mem_1043_sv2v_reg ,\nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,\nz.mem_1040_sv2v_reg ,
  \nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,\nz.mem_1037_sv2v_reg ,
  \nz.mem_1036_sv2v_reg ,\nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,
  \nz.mem_1033_sv2v_reg ,\nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,\nz.mem_1030_sv2v_reg ,
  \nz.mem_1029_sv2v_reg ,\nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,
  \nz.mem_1026_sv2v_reg ,\nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,\nz.mem_1023_sv2v_reg ,
  \nz.mem_1022_sv2v_reg ,\nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,
  \nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,\nz.mem_1016_sv2v_reg ,
  \nz.mem_1015_sv2v_reg ,\nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,
  \nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,\nz.mem_1009_sv2v_reg ,
  \nz.mem_1008_sv2v_reg ,\nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,
  \nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,\nz.mem_1002_sv2v_reg ,
  \nz.mem_1001_sv2v_reg ,\nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,
  \nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,
  \nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,\nz.mem_991_sv2v_reg ,
  \nz.mem_990_sv2v_reg ,\nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,
  \nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,\nz.mem_984_sv2v_reg ,
  \nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,\nz.mem_980_sv2v_reg ,
  \nz.mem_979_sv2v_reg ,\nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,
  \nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,\nz.mem_973_sv2v_reg ,
  \nz.mem_972_sv2v_reg ,\nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,
  \nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,
  \nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,\nz.mem_962_sv2v_reg ,
  \nz.mem_961_sv2v_reg ,\nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,
  \nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,
  \nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,\nz.mem_951_sv2v_reg ,
  \nz.mem_950_sv2v_reg ,\nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,
  \nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,\nz.mem_944_sv2v_reg ,
  \nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,\nz.mem_940_sv2v_reg ,
  \nz.mem_939_sv2v_reg ,\nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,
  \nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,\nz.mem_933_sv2v_reg ,
  \nz.mem_932_sv2v_reg ,\nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,
  \nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,
  \nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,\nz.mem_922_sv2v_reg ,
  \nz.mem_921_sv2v_reg ,\nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,
  \nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,
  \nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,\nz.mem_911_sv2v_reg ,
  \nz.mem_910_sv2v_reg ,\nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,
  \nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,\nz.mem_904_sv2v_reg ,
  \nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,\nz.mem_900_sv2v_reg ,
  \nz.mem_899_sv2v_reg ,\nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,
  \nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,\nz.mem_893_sv2v_reg ,
  \nz.mem_892_sv2v_reg ,\nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,
  \nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,
  \nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,\nz.mem_882_sv2v_reg ,
  \nz.mem_881_sv2v_reg ,\nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,
  \nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,
  \nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,\nz.mem_871_sv2v_reg ,
  \nz.mem_870_sv2v_reg ,\nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,
  \nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,\nz.mem_864_sv2v_reg ,
  \nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,\nz.mem_860_sv2v_reg ,
  \nz.mem_859_sv2v_reg ,\nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,
  \nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,\nz.mem_853_sv2v_reg ,
  \nz.mem_852_sv2v_reg ,\nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,
  \nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,
  \nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,\nz.mem_842_sv2v_reg ,
  \nz.mem_841_sv2v_reg ,\nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,
  \nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,
  \nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,\nz.mem_831_sv2v_reg ,
  \nz.mem_830_sv2v_reg ,\nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,
  \nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,\nz.mem_824_sv2v_reg ,
  \nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,\nz.mem_820_sv2v_reg ,
  \nz.mem_819_sv2v_reg ,\nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,
  \nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,\nz.mem_813_sv2v_reg ,
  \nz.mem_812_sv2v_reg ,\nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,
  \nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,
  \nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,\nz.mem_802_sv2v_reg ,
  \nz.mem_801_sv2v_reg ,\nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,
  \nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,
  \nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,\nz.mem_791_sv2v_reg ,
  \nz.mem_790_sv2v_reg ,\nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,
  \nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,\nz.mem_784_sv2v_reg ,
  \nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,\nz.mem_780_sv2v_reg ,
  \nz.mem_779_sv2v_reg ,\nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,
  \nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,\nz.mem_773_sv2v_reg ,
  \nz.mem_772_sv2v_reg ,\nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,
  \nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,
  \nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,\nz.mem_762_sv2v_reg ,
  \nz.mem_761_sv2v_reg ,\nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,
  \nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,
  \nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,\nz.mem_751_sv2v_reg ,
  \nz.mem_750_sv2v_reg ,\nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,
  \nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,\nz.mem_744_sv2v_reg ,
  \nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,\nz.mem_740_sv2v_reg ,
  \nz.mem_739_sv2v_reg ,\nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,
  \nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,\nz.mem_733_sv2v_reg ,
  \nz.mem_732_sv2v_reg ,\nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,
  \nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,
  \nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,\nz.mem_722_sv2v_reg ,
  \nz.mem_721_sv2v_reg ,\nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,
  \nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,
  \nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,\nz.mem_711_sv2v_reg ,
  \nz.mem_710_sv2v_reg ,\nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,
  \nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,\nz.mem_704_sv2v_reg ,
  \nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,\nz.mem_700_sv2v_reg ,
  \nz.mem_699_sv2v_reg ,\nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,
  \nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,\nz.mem_693_sv2v_reg ,
  \nz.mem_692_sv2v_reg ,\nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,
  \nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,
  \nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,\nz.mem_682_sv2v_reg ,
  \nz.mem_681_sv2v_reg ,\nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,
  \nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,
  \nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,\nz.mem_671_sv2v_reg ,
  \nz.mem_670_sv2v_reg ,\nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,
  \nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,
  \nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,\nz.mem_660_sv2v_reg ,
  \nz.mem_659_sv2v_reg ,\nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,
  \nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,\nz.mem_653_sv2v_reg ,
  \nz.mem_652_sv2v_reg ,\nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,
  \nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,
  \nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,\nz.mem_642_sv2v_reg ,
  \nz.mem_641_sv2v_reg ,\nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,
  \nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,
  \nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,
  \nz.mem_630_sv2v_reg ,\nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,
  \nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,
  \nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,
  \nz.mem_619_sv2v_reg ,\nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,
  \nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,
  \nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,
  \nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,
  \nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,
  \nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,
  \nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,
  \nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,
  \nz.mem_590_sv2v_reg ,\nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,
  \nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,
  \nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,
  \nz.mem_579_sv2v_reg ,\nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,
  \nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,
  \nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,
  \nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,
  \nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,
  \nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,
  \nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,
  \nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,
  \nz.mem_550_sv2v_reg ,\nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,
  \nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,
  \nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,
  \nz.mem_539_sv2v_reg ,\nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,
  \nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,
  \nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,
  \nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,
  \nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,
  \nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,
  \nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,
  \nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,
  \nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,
  \nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,
  \nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,
  \nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,
  \nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,
  \nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,
  \nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,
  \nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,
  \nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,
  \nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,
  \nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,
  \nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,
  \nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,
  \nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,
  \nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,
  \nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,
  \nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,
  \nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,
  \nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,
  \nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,
  \nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,
  \nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,
  \nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,
  \nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,
  \nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,
  \nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,
  \nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,
  \nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,
  \nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,
  \nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,
  \nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,
  \nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,
  \nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,
  \nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,
  \nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,
  \nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,
  \nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,
  \nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,
  \nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,
  \nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,
  \nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,
  \nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,
  \nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,
  \nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,
  \nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,
  \nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,
  \nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,
  \nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,
  \nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,
  \nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,
  \nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,
  \nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,
  \nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,
  \nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,
  \nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,
  \nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,
  \nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,
  \nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,
  \nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,
  \nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,
  \nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,
  \nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,
  \nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,
  \nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,
  \nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,
  \nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,
  \nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,
  \nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,
  \nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,
  \nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,
  \nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,
  \nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,
  \nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,
  \nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,
  \nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,
  \nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,
  \nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,
  \nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,
  \nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,
  \nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,
  \nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,
  \nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,
  \nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,
  \nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,
  \nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,
  \nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,
  \nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,
  \nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,
  \nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.mem [3199] = \nz.mem_3199_sv2v_reg ;
  assign \nz.mem [3198] = \nz.mem_3198_sv2v_reg ;
  assign \nz.mem [3197] = \nz.mem_3197_sv2v_reg ;
  assign \nz.mem [3196] = \nz.mem_3196_sv2v_reg ;
  assign \nz.mem [3195] = \nz.mem_3195_sv2v_reg ;
  assign \nz.mem [3194] = \nz.mem_3194_sv2v_reg ;
  assign \nz.mem [3193] = \nz.mem_3193_sv2v_reg ;
  assign \nz.mem [3192] = \nz.mem_3192_sv2v_reg ;
  assign \nz.mem [3191] = \nz.mem_3191_sv2v_reg ;
  assign \nz.mem [3190] = \nz.mem_3190_sv2v_reg ;
  assign \nz.mem [3189] = \nz.mem_3189_sv2v_reg ;
  assign \nz.mem [3188] = \nz.mem_3188_sv2v_reg ;
  assign \nz.mem [3187] = \nz.mem_3187_sv2v_reg ;
  assign \nz.mem [3186] = \nz.mem_3186_sv2v_reg ;
  assign \nz.mem [3185] = \nz.mem_3185_sv2v_reg ;
  assign \nz.mem [3184] = \nz.mem_3184_sv2v_reg ;
  assign \nz.mem [3183] = \nz.mem_3183_sv2v_reg ;
  assign \nz.mem [3182] = \nz.mem_3182_sv2v_reg ;
  assign \nz.mem [3181] = \nz.mem_3181_sv2v_reg ;
  assign \nz.mem [3180] = \nz.mem_3180_sv2v_reg ;
  assign \nz.mem [3179] = \nz.mem_3179_sv2v_reg ;
  assign \nz.mem [3178] = \nz.mem_3178_sv2v_reg ;
  assign \nz.mem [3177] = \nz.mem_3177_sv2v_reg ;
  assign \nz.mem [3176] = \nz.mem_3176_sv2v_reg ;
  assign \nz.mem [3175] = \nz.mem_3175_sv2v_reg ;
  assign \nz.mem [3174] = \nz.mem_3174_sv2v_reg ;
  assign \nz.mem [3173] = \nz.mem_3173_sv2v_reg ;
  assign \nz.mem [3172] = \nz.mem_3172_sv2v_reg ;
  assign \nz.mem [3171] = \nz.mem_3171_sv2v_reg ;
  assign \nz.mem [3170] = \nz.mem_3170_sv2v_reg ;
  assign \nz.mem [3169] = \nz.mem_3169_sv2v_reg ;
  assign \nz.mem [3168] = \nz.mem_3168_sv2v_reg ;
  assign \nz.mem [3167] = \nz.mem_3167_sv2v_reg ;
  assign \nz.mem [3166] = \nz.mem_3166_sv2v_reg ;
  assign \nz.mem [3165] = \nz.mem_3165_sv2v_reg ;
  assign \nz.mem [3164] = \nz.mem_3164_sv2v_reg ;
  assign \nz.mem [3163] = \nz.mem_3163_sv2v_reg ;
  assign \nz.mem [3162] = \nz.mem_3162_sv2v_reg ;
  assign \nz.mem [3161] = \nz.mem_3161_sv2v_reg ;
  assign \nz.mem [3160] = \nz.mem_3160_sv2v_reg ;
  assign \nz.mem [3159] = \nz.mem_3159_sv2v_reg ;
  assign \nz.mem [3158] = \nz.mem_3158_sv2v_reg ;
  assign \nz.mem [3157] = \nz.mem_3157_sv2v_reg ;
  assign \nz.mem [3156] = \nz.mem_3156_sv2v_reg ;
  assign \nz.mem [3155] = \nz.mem_3155_sv2v_reg ;
  assign \nz.mem [3154] = \nz.mem_3154_sv2v_reg ;
  assign \nz.mem [3153] = \nz.mem_3153_sv2v_reg ;
  assign \nz.mem [3152] = \nz.mem_3152_sv2v_reg ;
  assign \nz.mem [3151] = \nz.mem_3151_sv2v_reg ;
  assign \nz.mem [3150] = \nz.mem_3150_sv2v_reg ;
  assign \nz.mem [3149] = \nz.mem_3149_sv2v_reg ;
  assign \nz.mem [3148] = \nz.mem_3148_sv2v_reg ;
  assign \nz.mem [3147] = \nz.mem_3147_sv2v_reg ;
  assign \nz.mem [3146] = \nz.mem_3146_sv2v_reg ;
  assign \nz.mem [3145] = \nz.mem_3145_sv2v_reg ;
  assign \nz.mem [3144] = \nz.mem_3144_sv2v_reg ;
  assign \nz.mem [3143] = \nz.mem_3143_sv2v_reg ;
  assign \nz.mem [3142] = \nz.mem_3142_sv2v_reg ;
  assign \nz.mem [3141] = \nz.mem_3141_sv2v_reg ;
  assign \nz.mem [3140] = \nz.mem_3140_sv2v_reg ;
  assign \nz.mem [3139] = \nz.mem_3139_sv2v_reg ;
  assign \nz.mem [3138] = \nz.mem_3138_sv2v_reg ;
  assign \nz.mem [3137] = \nz.mem_3137_sv2v_reg ;
  assign \nz.mem [3136] = \nz.mem_3136_sv2v_reg ;
  assign \nz.mem [3135] = \nz.mem_3135_sv2v_reg ;
  assign \nz.mem [3134] = \nz.mem_3134_sv2v_reg ;
  assign \nz.mem [3133] = \nz.mem_3133_sv2v_reg ;
  assign \nz.mem [3132] = \nz.mem_3132_sv2v_reg ;
  assign \nz.mem [3131] = \nz.mem_3131_sv2v_reg ;
  assign \nz.mem [3130] = \nz.mem_3130_sv2v_reg ;
  assign \nz.mem [3129] = \nz.mem_3129_sv2v_reg ;
  assign \nz.mem [3128] = \nz.mem_3128_sv2v_reg ;
  assign \nz.mem [3127] = \nz.mem_3127_sv2v_reg ;
  assign \nz.mem [3126] = \nz.mem_3126_sv2v_reg ;
  assign \nz.mem [3125] = \nz.mem_3125_sv2v_reg ;
  assign \nz.mem [3124] = \nz.mem_3124_sv2v_reg ;
  assign \nz.mem [3123] = \nz.mem_3123_sv2v_reg ;
  assign \nz.mem [3122] = \nz.mem_3122_sv2v_reg ;
  assign \nz.mem [3121] = \nz.mem_3121_sv2v_reg ;
  assign \nz.mem [3120] = \nz.mem_3120_sv2v_reg ;
  assign \nz.mem [3119] = \nz.mem_3119_sv2v_reg ;
  assign \nz.mem [3118] = \nz.mem_3118_sv2v_reg ;
  assign \nz.mem [3117] = \nz.mem_3117_sv2v_reg ;
  assign \nz.mem [3116] = \nz.mem_3116_sv2v_reg ;
  assign \nz.mem [3115] = \nz.mem_3115_sv2v_reg ;
  assign \nz.mem [3114] = \nz.mem_3114_sv2v_reg ;
  assign \nz.mem [3113] = \nz.mem_3113_sv2v_reg ;
  assign \nz.mem [3112] = \nz.mem_3112_sv2v_reg ;
  assign \nz.mem [3111] = \nz.mem_3111_sv2v_reg ;
  assign \nz.mem [3110] = \nz.mem_3110_sv2v_reg ;
  assign \nz.mem [3109] = \nz.mem_3109_sv2v_reg ;
  assign \nz.mem [3108] = \nz.mem_3108_sv2v_reg ;
  assign \nz.mem [3107] = \nz.mem_3107_sv2v_reg ;
  assign \nz.mem [3106] = \nz.mem_3106_sv2v_reg ;
  assign \nz.mem [3105] = \nz.mem_3105_sv2v_reg ;
  assign \nz.mem [3104] = \nz.mem_3104_sv2v_reg ;
  assign \nz.mem [3103] = \nz.mem_3103_sv2v_reg ;
  assign \nz.mem [3102] = \nz.mem_3102_sv2v_reg ;
  assign \nz.mem [3101] = \nz.mem_3101_sv2v_reg ;
  assign \nz.mem [3100] = \nz.mem_3100_sv2v_reg ;
  assign \nz.mem [3099] = \nz.mem_3099_sv2v_reg ;
  assign \nz.mem [3098] = \nz.mem_3098_sv2v_reg ;
  assign \nz.mem [3097] = \nz.mem_3097_sv2v_reg ;
  assign \nz.mem [3096] = \nz.mem_3096_sv2v_reg ;
  assign \nz.mem [3095] = \nz.mem_3095_sv2v_reg ;
  assign \nz.mem [3094] = \nz.mem_3094_sv2v_reg ;
  assign \nz.mem [3093] = \nz.mem_3093_sv2v_reg ;
  assign \nz.mem [3092] = \nz.mem_3092_sv2v_reg ;
  assign \nz.mem [3091] = \nz.mem_3091_sv2v_reg ;
  assign \nz.mem [3090] = \nz.mem_3090_sv2v_reg ;
  assign \nz.mem [3089] = \nz.mem_3089_sv2v_reg ;
  assign \nz.mem [3088] = \nz.mem_3088_sv2v_reg ;
  assign \nz.mem [3087] = \nz.mem_3087_sv2v_reg ;
  assign \nz.mem [3086] = \nz.mem_3086_sv2v_reg ;
  assign \nz.mem [3085] = \nz.mem_3085_sv2v_reg ;
  assign \nz.mem [3084] = \nz.mem_3084_sv2v_reg ;
  assign \nz.mem [3083] = \nz.mem_3083_sv2v_reg ;
  assign \nz.mem [3082] = \nz.mem_3082_sv2v_reg ;
  assign \nz.mem [3081] = \nz.mem_3081_sv2v_reg ;
  assign \nz.mem [3080] = \nz.mem_3080_sv2v_reg ;
  assign \nz.mem [3079] = \nz.mem_3079_sv2v_reg ;
  assign \nz.mem [3078] = \nz.mem_3078_sv2v_reg ;
  assign \nz.mem [3077] = \nz.mem_3077_sv2v_reg ;
  assign \nz.mem [3076] = \nz.mem_3076_sv2v_reg ;
  assign \nz.mem [3075] = \nz.mem_3075_sv2v_reg ;
  assign \nz.mem [3074] = \nz.mem_3074_sv2v_reg ;
  assign \nz.mem [3073] = \nz.mem_3073_sv2v_reg ;
  assign \nz.mem [3072] = \nz.mem_3072_sv2v_reg ;
  assign \nz.mem [3071] = \nz.mem_3071_sv2v_reg ;
  assign \nz.mem [3070] = \nz.mem_3070_sv2v_reg ;
  assign \nz.mem [3069] = \nz.mem_3069_sv2v_reg ;
  assign \nz.mem [3068] = \nz.mem_3068_sv2v_reg ;
  assign \nz.mem [3067] = \nz.mem_3067_sv2v_reg ;
  assign \nz.mem [3066] = \nz.mem_3066_sv2v_reg ;
  assign \nz.mem [3065] = \nz.mem_3065_sv2v_reg ;
  assign \nz.mem [3064] = \nz.mem_3064_sv2v_reg ;
  assign \nz.mem [3063] = \nz.mem_3063_sv2v_reg ;
  assign \nz.mem [3062] = \nz.mem_3062_sv2v_reg ;
  assign \nz.mem [3061] = \nz.mem_3061_sv2v_reg ;
  assign \nz.mem [3060] = \nz.mem_3060_sv2v_reg ;
  assign \nz.mem [3059] = \nz.mem_3059_sv2v_reg ;
  assign \nz.mem [3058] = \nz.mem_3058_sv2v_reg ;
  assign \nz.mem [3057] = \nz.mem_3057_sv2v_reg ;
  assign \nz.mem [3056] = \nz.mem_3056_sv2v_reg ;
  assign \nz.mem [3055] = \nz.mem_3055_sv2v_reg ;
  assign \nz.mem [3054] = \nz.mem_3054_sv2v_reg ;
  assign \nz.mem [3053] = \nz.mem_3053_sv2v_reg ;
  assign \nz.mem [3052] = \nz.mem_3052_sv2v_reg ;
  assign \nz.mem [3051] = \nz.mem_3051_sv2v_reg ;
  assign \nz.mem [3050] = \nz.mem_3050_sv2v_reg ;
  assign \nz.mem [3049] = \nz.mem_3049_sv2v_reg ;
  assign \nz.mem [3048] = \nz.mem_3048_sv2v_reg ;
  assign \nz.mem [3047] = \nz.mem_3047_sv2v_reg ;
  assign \nz.mem [3046] = \nz.mem_3046_sv2v_reg ;
  assign \nz.mem [3045] = \nz.mem_3045_sv2v_reg ;
  assign \nz.mem [3044] = \nz.mem_3044_sv2v_reg ;
  assign \nz.mem [3043] = \nz.mem_3043_sv2v_reg ;
  assign \nz.mem [3042] = \nz.mem_3042_sv2v_reg ;
  assign \nz.mem [3041] = \nz.mem_3041_sv2v_reg ;
  assign \nz.mem [3040] = \nz.mem_3040_sv2v_reg ;
  assign \nz.mem [3039] = \nz.mem_3039_sv2v_reg ;
  assign \nz.mem [3038] = \nz.mem_3038_sv2v_reg ;
  assign \nz.mem [3037] = \nz.mem_3037_sv2v_reg ;
  assign \nz.mem [3036] = \nz.mem_3036_sv2v_reg ;
  assign \nz.mem [3035] = \nz.mem_3035_sv2v_reg ;
  assign \nz.mem [3034] = \nz.mem_3034_sv2v_reg ;
  assign \nz.mem [3033] = \nz.mem_3033_sv2v_reg ;
  assign \nz.mem [3032] = \nz.mem_3032_sv2v_reg ;
  assign \nz.mem [3031] = \nz.mem_3031_sv2v_reg ;
  assign \nz.mem [3030] = \nz.mem_3030_sv2v_reg ;
  assign \nz.mem [3029] = \nz.mem_3029_sv2v_reg ;
  assign \nz.mem [3028] = \nz.mem_3028_sv2v_reg ;
  assign \nz.mem [3027] = \nz.mem_3027_sv2v_reg ;
  assign \nz.mem [3026] = \nz.mem_3026_sv2v_reg ;
  assign \nz.mem [3025] = \nz.mem_3025_sv2v_reg ;
  assign \nz.mem [3024] = \nz.mem_3024_sv2v_reg ;
  assign \nz.mem [3023] = \nz.mem_3023_sv2v_reg ;
  assign \nz.mem [3022] = \nz.mem_3022_sv2v_reg ;
  assign \nz.mem [3021] = \nz.mem_3021_sv2v_reg ;
  assign \nz.mem [3020] = \nz.mem_3020_sv2v_reg ;
  assign \nz.mem [3019] = \nz.mem_3019_sv2v_reg ;
  assign \nz.mem [3018] = \nz.mem_3018_sv2v_reg ;
  assign \nz.mem [3017] = \nz.mem_3017_sv2v_reg ;
  assign \nz.mem [3016] = \nz.mem_3016_sv2v_reg ;
  assign \nz.mem [3015] = \nz.mem_3015_sv2v_reg ;
  assign \nz.mem [3014] = \nz.mem_3014_sv2v_reg ;
  assign \nz.mem [3013] = \nz.mem_3013_sv2v_reg ;
  assign \nz.mem [3012] = \nz.mem_3012_sv2v_reg ;
  assign \nz.mem [3011] = \nz.mem_3011_sv2v_reg ;
  assign \nz.mem [3010] = \nz.mem_3010_sv2v_reg ;
  assign \nz.mem [3009] = \nz.mem_3009_sv2v_reg ;
  assign \nz.mem [3008] = \nz.mem_3008_sv2v_reg ;
  assign \nz.mem [3007] = \nz.mem_3007_sv2v_reg ;
  assign \nz.mem [3006] = \nz.mem_3006_sv2v_reg ;
  assign \nz.mem [3005] = \nz.mem_3005_sv2v_reg ;
  assign \nz.mem [3004] = \nz.mem_3004_sv2v_reg ;
  assign \nz.mem [3003] = \nz.mem_3003_sv2v_reg ;
  assign \nz.mem [3002] = \nz.mem_3002_sv2v_reg ;
  assign \nz.mem [3001] = \nz.mem_3001_sv2v_reg ;
  assign \nz.mem [3000] = \nz.mem_3000_sv2v_reg ;
  assign \nz.mem [2999] = \nz.mem_2999_sv2v_reg ;
  assign \nz.mem [2998] = \nz.mem_2998_sv2v_reg ;
  assign \nz.mem [2997] = \nz.mem_2997_sv2v_reg ;
  assign \nz.mem [2996] = \nz.mem_2996_sv2v_reg ;
  assign \nz.mem [2995] = \nz.mem_2995_sv2v_reg ;
  assign \nz.mem [2994] = \nz.mem_2994_sv2v_reg ;
  assign \nz.mem [2993] = \nz.mem_2993_sv2v_reg ;
  assign \nz.mem [2992] = \nz.mem_2992_sv2v_reg ;
  assign \nz.mem [2991] = \nz.mem_2991_sv2v_reg ;
  assign \nz.mem [2990] = \nz.mem_2990_sv2v_reg ;
  assign \nz.mem [2989] = \nz.mem_2989_sv2v_reg ;
  assign \nz.mem [2988] = \nz.mem_2988_sv2v_reg ;
  assign \nz.mem [2987] = \nz.mem_2987_sv2v_reg ;
  assign \nz.mem [2986] = \nz.mem_2986_sv2v_reg ;
  assign \nz.mem [2985] = \nz.mem_2985_sv2v_reg ;
  assign \nz.mem [2984] = \nz.mem_2984_sv2v_reg ;
  assign \nz.mem [2983] = \nz.mem_2983_sv2v_reg ;
  assign \nz.mem [2982] = \nz.mem_2982_sv2v_reg ;
  assign \nz.mem [2981] = \nz.mem_2981_sv2v_reg ;
  assign \nz.mem [2980] = \nz.mem_2980_sv2v_reg ;
  assign \nz.mem [2979] = \nz.mem_2979_sv2v_reg ;
  assign \nz.mem [2978] = \nz.mem_2978_sv2v_reg ;
  assign \nz.mem [2977] = \nz.mem_2977_sv2v_reg ;
  assign \nz.mem [2976] = \nz.mem_2976_sv2v_reg ;
  assign \nz.mem [2975] = \nz.mem_2975_sv2v_reg ;
  assign \nz.mem [2974] = \nz.mem_2974_sv2v_reg ;
  assign \nz.mem [2973] = \nz.mem_2973_sv2v_reg ;
  assign \nz.mem [2972] = \nz.mem_2972_sv2v_reg ;
  assign \nz.mem [2971] = \nz.mem_2971_sv2v_reg ;
  assign \nz.mem [2970] = \nz.mem_2970_sv2v_reg ;
  assign \nz.mem [2969] = \nz.mem_2969_sv2v_reg ;
  assign \nz.mem [2968] = \nz.mem_2968_sv2v_reg ;
  assign \nz.mem [2967] = \nz.mem_2967_sv2v_reg ;
  assign \nz.mem [2966] = \nz.mem_2966_sv2v_reg ;
  assign \nz.mem [2965] = \nz.mem_2965_sv2v_reg ;
  assign \nz.mem [2964] = \nz.mem_2964_sv2v_reg ;
  assign \nz.mem [2963] = \nz.mem_2963_sv2v_reg ;
  assign \nz.mem [2962] = \nz.mem_2962_sv2v_reg ;
  assign \nz.mem [2961] = \nz.mem_2961_sv2v_reg ;
  assign \nz.mem [2960] = \nz.mem_2960_sv2v_reg ;
  assign \nz.mem [2959] = \nz.mem_2959_sv2v_reg ;
  assign \nz.mem [2958] = \nz.mem_2958_sv2v_reg ;
  assign \nz.mem [2957] = \nz.mem_2957_sv2v_reg ;
  assign \nz.mem [2956] = \nz.mem_2956_sv2v_reg ;
  assign \nz.mem [2955] = \nz.mem_2955_sv2v_reg ;
  assign \nz.mem [2954] = \nz.mem_2954_sv2v_reg ;
  assign \nz.mem [2953] = \nz.mem_2953_sv2v_reg ;
  assign \nz.mem [2952] = \nz.mem_2952_sv2v_reg ;
  assign \nz.mem [2951] = \nz.mem_2951_sv2v_reg ;
  assign \nz.mem [2950] = \nz.mem_2950_sv2v_reg ;
  assign \nz.mem [2949] = \nz.mem_2949_sv2v_reg ;
  assign \nz.mem [2948] = \nz.mem_2948_sv2v_reg ;
  assign \nz.mem [2947] = \nz.mem_2947_sv2v_reg ;
  assign \nz.mem [2946] = \nz.mem_2946_sv2v_reg ;
  assign \nz.mem [2945] = \nz.mem_2945_sv2v_reg ;
  assign \nz.mem [2944] = \nz.mem_2944_sv2v_reg ;
  assign \nz.mem [2943] = \nz.mem_2943_sv2v_reg ;
  assign \nz.mem [2942] = \nz.mem_2942_sv2v_reg ;
  assign \nz.mem [2941] = \nz.mem_2941_sv2v_reg ;
  assign \nz.mem [2940] = \nz.mem_2940_sv2v_reg ;
  assign \nz.mem [2939] = \nz.mem_2939_sv2v_reg ;
  assign \nz.mem [2938] = \nz.mem_2938_sv2v_reg ;
  assign \nz.mem [2937] = \nz.mem_2937_sv2v_reg ;
  assign \nz.mem [2936] = \nz.mem_2936_sv2v_reg ;
  assign \nz.mem [2935] = \nz.mem_2935_sv2v_reg ;
  assign \nz.mem [2934] = \nz.mem_2934_sv2v_reg ;
  assign \nz.mem [2933] = \nz.mem_2933_sv2v_reg ;
  assign \nz.mem [2932] = \nz.mem_2932_sv2v_reg ;
  assign \nz.mem [2931] = \nz.mem_2931_sv2v_reg ;
  assign \nz.mem [2930] = \nz.mem_2930_sv2v_reg ;
  assign \nz.mem [2929] = \nz.mem_2929_sv2v_reg ;
  assign \nz.mem [2928] = \nz.mem_2928_sv2v_reg ;
  assign \nz.mem [2927] = \nz.mem_2927_sv2v_reg ;
  assign \nz.mem [2926] = \nz.mem_2926_sv2v_reg ;
  assign \nz.mem [2925] = \nz.mem_2925_sv2v_reg ;
  assign \nz.mem [2924] = \nz.mem_2924_sv2v_reg ;
  assign \nz.mem [2923] = \nz.mem_2923_sv2v_reg ;
  assign \nz.mem [2922] = \nz.mem_2922_sv2v_reg ;
  assign \nz.mem [2921] = \nz.mem_2921_sv2v_reg ;
  assign \nz.mem [2920] = \nz.mem_2920_sv2v_reg ;
  assign \nz.mem [2919] = \nz.mem_2919_sv2v_reg ;
  assign \nz.mem [2918] = \nz.mem_2918_sv2v_reg ;
  assign \nz.mem [2917] = \nz.mem_2917_sv2v_reg ;
  assign \nz.mem [2916] = \nz.mem_2916_sv2v_reg ;
  assign \nz.mem [2915] = \nz.mem_2915_sv2v_reg ;
  assign \nz.mem [2914] = \nz.mem_2914_sv2v_reg ;
  assign \nz.mem [2913] = \nz.mem_2913_sv2v_reg ;
  assign \nz.mem [2912] = \nz.mem_2912_sv2v_reg ;
  assign \nz.mem [2911] = \nz.mem_2911_sv2v_reg ;
  assign \nz.mem [2910] = \nz.mem_2910_sv2v_reg ;
  assign \nz.mem [2909] = \nz.mem_2909_sv2v_reg ;
  assign \nz.mem [2908] = \nz.mem_2908_sv2v_reg ;
  assign \nz.mem [2907] = \nz.mem_2907_sv2v_reg ;
  assign \nz.mem [2906] = \nz.mem_2906_sv2v_reg ;
  assign \nz.mem [2905] = \nz.mem_2905_sv2v_reg ;
  assign \nz.mem [2904] = \nz.mem_2904_sv2v_reg ;
  assign \nz.mem [2903] = \nz.mem_2903_sv2v_reg ;
  assign \nz.mem [2902] = \nz.mem_2902_sv2v_reg ;
  assign \nz.mem [2901] = \nz.mem_2901_sv2v_reg ;
  assign \nz.mem [2900] = \nz.mem_2900_sv2v_reg ;
  assign \nz.mem [2899] = \nz.mem_2899_sv2v_reg ;
  assign \nz.mem [2898] = \nz.mem_2898_sv2v_reg ;
  assign \nz.mem [2897] = \nz.mem_2897_sv2v_reg ;
  assign \nz.mem [2896] = \nz.mem_2896_sv2v_reg ;
  assign \nz.mem [2895] = \nz.mem_2895_sv2v_reg ;
  assign \nz.mem [2894] = \nz.mem_2894_sv2v_reg ;
  assign \nz.mem [2893] = \nz.mem_2893_sv2v_reg ;
  assign \nz.mem [2892] = \nz.mem_2892_sv2v_reg ;
  assign \nz.mem [2891] = \nz.mem_2891_sv2v_reg ;
  assign \nz.mem [2890] = \nz.mem_2890_sv2v_reg ;
  assign \nz.mem [2889] = \nz.mem_2889_sv2v_reg ;
  assign \nz.mem [2888] = \nz.mem_2888_sv2v_reg ;
  assign \nz.mem [2887] = \nz.mem_2887_sv2v_reg ;
  assign \nz.mem [2886] = \nz.mem_2886_sv2v_reg ;
  assign \nz.mem [2885] = \nz.mem_2885_sv2v_reg ;
  assign \nz.mem [2884] = \nz.mem_2884_sv2v_reg ;
  assign \nz.mem [2883] = \nz.mem_2883_sv2v_reg ;
  assign \nz.mem [2882] = \nz.mem_2882_sv2v_reg ;
  assign \nz.mem [2881] = \nz.mem_2881_sv2v_reg ;
  assign \nz.mem [2880] = \nz.mem_2880_sv2v_reg ;
  assign \nz.mem [2879] = \nz.mem_2879_sv2v_reg ;
  assign \nz.mem [2878] = \nz.mem_2878_sv2v_reg ;
  assign \nz.mem [2877] = \nz.mem_2877_sv2v_reg ;
  assign \nz.mem [2876] = \nz.mem_2876_sv2v_reg ;
  assign \nz.mem [2875] = \nz.mem_2875_sv2v_reg ;
  assign \nz.mem [2874] = \nz.mem_2874_sv2v_reg ;
  assign \nz.mem [2873] = \nz.mem_2873_sv2v_reg ;
  assign \nz.mem [2872] = \nz.mem_2872_sv2v_reg ;
  assign \nz.mem [2871] = \nz.mem_2871_sv2v_reg ;
  assign \nz.mem [2870] = \nz.mem_2870_sv2v_reg ;
  assign \nz.mem [2869] = \nz.mem_2869_sv2v_reg ;
  assign \nz.mem [2868] = \nz.mem_2868_sv2v_reg ;
  assign \nz.mem [2867] = \nz.mem_2867_sv2v_reg ;
  assign \nz.mem [2866] = \nz.mem_2866_sv2v_reg ;
  assign \nz.mem [2865] = \nz.mem_2865_sv2v_reg ;
  assign \nz.mem [2864] = \nz.mem_2864_sv2v_reg ;
  assign \nz.mem [2863] = \nz.mem_2863_sv2v_reg ;
  assign \nz.mem [2862] = \nz.mem_2862_sv2v_reg ;
  assign \nz.mem [2861] = \nz.mem_2861_sv2v_reg ;
  assign \nz.mem [2860] = \nz.mem_2860_sv2v_reg ;
  assign \nz.mem [2859] = \nz.mem_2859_sv2v_reg ;
  assign \nz.mem [2858] = \nz.mem_2858_sv2v_reg ;
  assign \nz.mem [2857] = \nz.mem_2857_sv2v_reg ;
  assign \nz.mem [2856] = \nz.mem_2856_sv2v_reg ;
  assign \nz.mem [2855] = \nz.mem_2855_sv2v_reg ;
  assign \nz.mem [2854] = \nz.mem_2854_sv2v_reg ;
  assign \nz.mem [2853] = \nz.mem_2853_sv2v_reg ;
  assign \nz.mem [2852] = \nz.mem_2852_sv2v_reg ;
  assign \nz.mem [2851] = \nz.mem_2851_sv2v_reg ;
  assign \nz.mem [2850] = \nz.mem_2850_sv2v_reg ;
  assign \nz.mem [2849] = \nz.mem_2849_sv2v_reg ;
  assign \nz.mem [2848] = \nz.mem_2848_sv2v_reg ;
  assign \nz.mem [2847] = \nz.mem_2847_sv2v_reg ;
  assign \nz.mem [2846] = \nz.mem_2846_sv2v_reg ;
  assign \nz.mem [2845] = \nz.mem_2845_sv2v_reg ;
  assign \nz.mem [2844] = \nz.mem_2844_sv2v_reg ;
  assign \nz.mem [2843] = \nz.mem_2843_sv2v_reg ;
  assign \nz.mem [2842] = \nz.mem_2842_sv2v_reg ;
  assign \nz.mem [2841] = \nz.mem_2841_sv2v_reg ;
  assign \nz.mem [2840] = \nz.mem_2840_sv2v_reg ;
  assign \nz.mem [2839] = \nz.mem_2839_sv2v_reg ;
  assign \nz.mem [2838] = \nz.mem_2838_sv2v_reg ;
  assign \nz.mem [2837] = \nz.mem_2837_sv2v_reg ;
  assign \nz.mem [2836] = \nz.mem_2836_sv2v_reg ;
  assign \nz.mem [2835] = \nz.mem_2835_sv2v_reg ;
  assign \nz.mem [2834] = \nz.mem_2834_sv2v_reg ;
  assign \nz.mem [2833] = \nz.mem_2833_sv2v_reg ;
  assign \nz.mem [2832] = \nz.mem_2832_sv2v_reg ;
  assign \nz.mem [2831] = \nz.mem_2831_sv2v_reg ;
  assign \nz.mem [2830] = \nz.mem_2830_sv2v_reg ;
  assign \nz.mem [2829] = \nz.mem_2829_sv2v_reg ;
  assign \nz.mem [2828] = \nz.mem_2828_sv2v_reg ;
  assign \nz.mem [2827] = \nz.mem_2827_sv2v_reg ;
  assign \nz.mem [2826] = \nz.mem_2826_sv2v_reg ;
  assign \nz.mem [2825] = \nz.mem_2825_sv2v_reg ;
  assign \nz.mem [2824] = \nz.mem_2824_sv2v_reg ;
  assign \nz.mem [2823] = \nz.mem_2823_sv2v_reg ;
  assign \nz.mem [2822] = \nz.mem_2822_sv2v_reg ;
  assign \nz.mem [2821] = \nz.mem_2821_sv2v_reg ;
  assign \nz.mem [2820] = \nz.mem_2820_sv2v_reg ;
  assign \nz.mem [2819] = \nz.mem_2819_sv2v_reg ;
  assign \nz.mem [2818] = \nz.mem_2818_sv2v_reg ;
  assign \nz.mem [2817] = \nz.mem_2817_sv2v_reg ;
  assign \nz.mem [2816] = \nz.mem_2816_sv2v_reg ;
  assign \nz.mem [2815] = \nz.mem_2815_sv2v_reg ;
  assign \nz.mem [2814] = \nz.mem_2814_sv2v_reg ;
  assign \nz.mem [2813] = \nz.mem_2813_sv2v_reg ;
  assign \nz.mem [2812] = \nz.mem_2812_sv2v_reg ;
  assign \nz.mem [2811] = \nz.mem_2811_sv2v_reg ;
  assign \nz.mem [2810] = \nz.mem_2810_sv2v_reg ;
  assign \nz.mem [2809] = \nz.mem_2809_sv2v_reg ;
  assign \nz.mem [2808] = \nz.mem_2808_sv2v_reg ;
  assign \nz.mem [2807] = \nz.mem_2807_sv2v_reg ;
  assign \nz.mem [2806] = \nz.mem_2806_sv2v_reg ;
  assign \nz.mem [2805] = \nz.mem_2805_sv2v_reg ;
  assign \nz.mem [2804] = \nz.mem_2804_sv2v_reg ;
  assign \nz.mem [2803] = \nz.mem_2803_sv2v_reg ;
  assign \nz.mem [2802] = \nz.mem_2802_sv2v_reg ;
  assign \nz.mem [2801] = \nz.mem_2801_sv2v_reg ;
  assign \nz.mem [2800] = \nz.mem_2800_sv2v_reg ;
  assign \nz.mem [2799] = \nz.mem_2799_sv2v_reg ;
  assign \nz.mem [2798] = \nz.mem_2798_sv2v_reg ;
  assign \nz.mem [2797] = \nz.mem_2797_sv2v_reg ;
  assign \nz.mem [2796] = \nz.mem_2796_sv2v_reg ;
  assign \nz.mem [2795] = \nz.mem_2795_sv2v_reg ;
  assign \nz.mem [2794] = \nz.mem_2794_sv2v_reg ;
  assign \nz.mem [2793] = \nz.mem_2793_sv2v_reg ;
  assign \nz.mem [2792] = \nz.mem_2792_sv2v_reg ;
  assign \nz.mem [2791] = \nz.mem_2791_sv2v_reg ;
  assign \nz.mem [2790] = \nz.mem_2790_sv2v_reg ;
  assign \nz.mem [2789] = \nz.mem_2789_sv2v_reg ;
  assign \nz.mem [2788] = \nz.mem_2788_sv2v_reg ;
  assign \nz.mem [2787] = \nz.mem_2787_sv2v_reg ;
  assign \nz.mem [2786] = \nz.mem_2786_sv2v_reg ;
  assign \nz.mem [2785] = \nz.mem_2785_sv2v_reg ;
  assign \nz.mem [2784] = \nz.mem_2784_sv2v_reg ;
  assign \nz.mem [2783] = \nz.mem_2783_sv2v_reg ;
  assign \nz.mem [2782] = \nz.mem_2782_sv2v_reg ;
  assign \nz.mem [2781] = \nz.mem_2781_sv2v_reg ;
  assign \nz.mem [2780] = \nz.mem_2780_sv2v_reg ;
  assign \nz.mem [2779] = \nz.mem_2779_sv2v_reg ;
  assign \nz.mem [2778] = \nz.mem_2778_sv2v_reg ;
  assign \nz.mem [2777] = \nz.mem_2777_sv2v_reg ;
  assign \nz.mem [2776] = \nz.mem_2776_sv2v_reg ;
  assign \nz.mem [2775] = \nz.mem_2775_sv2v_reg ;
  assign \nz.mem [2774] = \nz.mem_2774_sv2v_reg ;
  assign \nz.mem [2773] = \nz.mem_2773_sv2v_reg ;
  assign \nz.mem [2772] = \nz.mem_2772_sv2v_reg ;
  assign \nz.mem [2771] = \nz.mem_2771_sv2v_reg ;
  assign \nz.mem [2770] = \nz.mem_2770_sv2v_reg ;
  assign \nz.mem [2769] = \nz.mem_2769_sv2v_reg ;
  assign \nz.mem [2768] = \nz.mem_2768_sv2v_reg ;
  assign \nz.mem [2767] = \nz.mem_2767_sv2v_reg ;
  assign \nz.mem [2766] = \nz.mem_2766_sv2v_reg ;
  assign \nz.mem [2765] = \nz.mem_2765_sv2v_reg ;
  assign \nz.mem [2764] = \nz.mem_2764_sv2v_reg ;
  assign \nz.mem [2763] = \nz.mem_2763_sv2v_reg ;
  assign \nz.mem [2762] = \nz.mem_2762_sv2v_reg ;
  assign \nz.mem [2761] = \nz.mem_2761_sv2v_reg ;
  assign \nz.mem [2760] = \nz.mem_2760_sv2v_reg ;
  assign \nz.mem [2759] = \nz.mem_2759_sv2v_reg ;
  assign \nz.mem [2758] = \nz.mem_2758_sv2v_reg ;
  assign \nz.mem [2757] = \nz.mem_2757_sv2v_reg ;
  assign \nz.mem [2756] = \nz.mem_2756_sv2v_reg ;
  assign \nz.mem [2755] = \nz.mem_2755_sv2v_reg ;
  assign \nz.mem [2754] = \nz.mem_2754_sv2v_reg ;
  assign \nz.mem [2753] = \nz.mem_2753_sv2v_reg ;
  assign \nz.mem [2752] = \nz.mem_2752_sv2v_reg ;
  assign \nz.mem [2751] = \nz.mem_2751_sv2v_reg ;
  assign \nz.mem [2750] = \nz.mem_2750_sv2v_reg ;
  assign \nz.mem [2749] = \nz.mem_2749_sv2v_reg ;
  assign \nz.mem [2748] = \nz.mem_2748_sv2v_reg ;
  assign \nz.mem [2747] = \nz.mem_2747_sv2v_reg ;
  assign \nz.mem [2746] = \nz.mem_2746_sv2v_reg ;
  assign \nz.mem [2745] = \nz.mem_2745_sv2v_reg ;
  assign \nz.mem [2744] = \nz.mem_2744_sv2v_reg ;
  assign \nz.mem [2743] = \nz.mem_2743_sv2v_reg ;
  assign \nz.mem [2742] = \nz.mem_2742_sv2v_reg ;
  assign \nz.mem [2741] = \nz.mem_2741_sv2v_reg ;
  assign \nz.mem [2740] = \nz.mem_2740_sv2v_reg ;
  assign \nz.mem [2739] = \nz.mem_2739_sv2v_reg ;
  assign \nz.mem [2738] = \nz.mem_2738_sv2v_reg ;
  assign \nz.mem [2737] = \nz.mem_2737_sv2v_reg ;
  assign \nz.mem [2736] = \nz.mem_2736_sv2v_reg ;
  assign \nz.mem [2735] = \nz.mem_2735_sv2v_reg ;
  assign \nz.mem [2734] = \nz.mem_2734_sv2v_reg ;
  assign \nz.mem [2733] = \nz.mem_2733_sv2v_reg ;
  assign \nz.mem [2732] = \nz.mem_2732_sv2v_reg ;
  assign \nz.mem [2731] = \nz.mem_2731_sv2v_reg ;
  assign \nz.mem [2730] = \nz.mem_2730_sv2v_reg ;
  assign \nz.mem [2729] = \nz.mem_2729_sv2v_reg ;
  assign \nz.mem [2728] = \nz.mem_2728_sv2v_reg ;
  assign \nz.mem [2727] = \nz.mem_2727_sv2v_reg ;
  assign \nz.mem [2726] = \nz.mem_2726_sv2v_reg ;
  assign \nz.mem [2725] = \nz.mem_2725_sv2v_reg ;
  assign \nz.mem [2724] = \nz.mem_2724_sv2v_reg ;
  assign \nz.mem [2723] = \nz.mem_2723_sv2v_reg ;
  assign \nz.mem [2722] = \nz.mem_2722_sv2v_reg ;
  assign \nz.mem [2721] = \nz.mem_2721_sv2v_reg ;
  assign \nz.mem [2720] = \nz.mem_2720_sv2v_reg ;
  assign \nz.mem [2719] = \nz.mem_2719_sv2v_reg ;
  assign \nz.mem [2718] = \nz.mem_2718_sv2v_reg ;
  assign \nz.mem [2717] = \nz.mem_2717_sv2v_reg ;
  assign \nz.mem [2716] = \nz.mem_2716_sv2v_reg ;
  assign \nz.mem [2715] = \nz.mem_2715_sv2v_reg ;
  assign \nz.mem [2714] = \nz.mem_2714_sv2v_reg ;
  assign \nz.mem [2713] = \nz.mem_2713_sv2v_reg ;
  assign \nz.mem [2712] = \nz.mem_2712_sv2v_reg ;
  assign \nz.mem [2711] = \nz.mem_2711_sv2v_reg ;
  assign \nz.mem [2710] = \nz.mem_2710_sv2v_reg ;
  assign \nz.mem [2709] = \nz.mem_2709_sv2v_reg ;
  assign \nz.mem [2708] = \nz.mem_2708_sv2v_reg ;
  assign \nz.mem [2707] = \nz.mem_2707_sv2v_reg ;
  assign \nz.mem [2706] = \nz.mem_2706_sv2v_reg ;
  assign \nz.mem [2705] = \nz.mem_2705_sv2v_reg ;
  assign \nz.mem [2704] = \nz.mem_2704_sv2v_reg ;
  assign \nz.mem [2703] = \nz.mem_2703_sv2v_reg ;
  assign \nz.mem [2702] = \nz.mem_2702_sv2v_reg ;
  assign \nz.mem [2701] = \nz.mem_2701_sv2v_reg ;
  assign \nz.mem [2700] = \nz.mem_2700_sv2v_reg ;
  assign \nz.mem [2699] = \nz.mem_2699_sv2v_reg ;
  assign \nz.mem [2698] = \nz.mem_2698_sv2v_reg ;
  assign \nz.mem [2697] = \nz.mem_2697_sv2v_reg ;
  assign \nz.mem [2696] = \nz.mem_2696_sv2v_reg ;
  assign \nz.mem [2695] = \nz.mem_2695_sv2v_reg ;
  assign \nz.mem [2694] = \nz.mem_2694_sv2v_reg ;
  assign \nz.mem [2693] = \nz.mem_2693_sv2v_reg ;
  assign \nz.mem [2692] = \nz.mem_2692_sv2v_reg ;
  assign \nz.mem [2691] = \nz.mem_2691_sv2v_reg ;
  assign \nz.mem [2690] = \nz.mem_2690_sv2v_reg ;
  assign \nz.mem [2689] = \nz.mem_2689_sv2v_reg ;
  assign \nz.mem [2688] = \nz.mem_2688_sv2v_reg ;
  assign \nz.mem [2687] = \nz.mem_2687_sv2v_reg ;
  assign \nz.mem [2686] = \nz.mem_2686_sv2v_reg ;
  assign \nz.mem [2685] = \nz.mem_2685_sv2v_reg ;
  assign \nz.mem [2684] = \nz.mem_2684_sv2v_reg ;
  assign \nz.mem [2683] = \nz.mem_2683_sv2v_reg ;
  assign \nz.mem [2682] = \nz.mem_2682_sv2v_reg ;
  assign \nz.mem [2681] = \nz.mem_2681_sv2v_reg ;
  assign \nz.mem [2680] = \nz.mem_2680_sv2v_reg ;
  assign \nz.mem [2679] = \nz.mem_2679_sv2v_reg ;
  assign \nz.mem [2678] = \nz.mem_2678_sv2v_reg ;
  assign \nz.mem [2677] = \nz.mem_2677_sv2v_reg ;
  assign \nz.mem [2676] = \nz.mem_2676_sv2v_reg ;
  assign \nz.mem [2675] = \nz.mem_2675_sv2v_reg ;
  assign \nz.mem [2674] = \nz.mem_2674_sv2v_reg ;
  assign \nz.mem [2673] = \nz.mem_2673_sv2v_reg ;
  assign \nz.mem [2672] = \nz.mem_2672_sv2v_reg ;
  assign \nz.mem [2671] = \nz.mem_2671_sv2v_reg ;
  assign \nz.mem [2670] = \nz.mem_2670_sv2v_reg ;
  assign \nz.mem [2669] = \nz.mem_2669_sv2v_reg ;
  assign \nz.mem [2668] = \nz.mem_2668_sv2v_reg ;
  assign \nz.mem [2667] = \nz.mem_2667_sv2v_reg ;
  assign \nz.mem [2666] = \nz.mem_2666_sv2v_reg ;
  assign \nz.mem [2665] = \nz.mem_2665_sv2v_reg ;
  assign \nz.mem [2664] = \nz.mem_2664_sv2v_reg ;
  assign \nz.mem [2663] = \nz.mem_2663_sv2v_reg ;
  assign \nz.mem [2662] = \nz.mem_2662_sv2v_reg ;
  assign \nz.mem [2661] = \nz.mem_2661_sv2v_reg ;
  assign \nz.mem [2660] = \nz.mem_2660_sv2v_reg ;
  assign \nz.mem [2659] = \nz.mem_2659_sv2v_reg ;
  assign \nz.mem [2658] = \nz.mem_2658_sv2v_reg ;
  assign \nz.mem [2657] = \nz.mem_2657_sv2v_reg ;
  assign \nz.mem [2656] = \nz.mem_2656_sv2v_reg ;
  assign \nz.mem [2655] = \nz.mem_2655_sv2v_reg ;
  assign \nz.mem [2654] = \nz.mem_2654_sv2v_reg ;
  assign \nz.mem [2653] = \nz.mem_2653_sv2v_reg ;
  assign \nz.mem [2652] = \nz.mem_2652_sv2v_reg ;
  assign \nz.mem [2651] = \nz.mem_2651_sv2v_reg ;
  assign \nz.mem [2650] = \nz.mem_2650_sv2v_reg ;
  assign \nz.mem [2649] = \nz.mem_2649_sv2v_reg ;
  assign \nz.mem [2648] = \nz.mem_2648_sv2v_reg ;
  assign \nz.mem [2647] = \nz.mem_2647_sv2v_reg ;
  assign \nz.mem [2646] = \nz.mem_2646_sv2v_reg ;
  assign \nz.mem [2645] = \nz.mem_2645_sv2v_reg ;
  assign \nz.mem [2644] = \nz.mem_2644_sv2v_reg ;
  assign \nz.mem [2643] = \nz.mem_2643_sv2v_reg ;
  assign \nz.mem [2642] = \nz.mem_2642_sv2v_reg ;
  assign \nz.mem [2641] = \nz.mem_2641_sv2v_reg ;
  assign \nz.mem [2640] = \nz.mem_2640_sv2v_reg ;
  assign \nz.mem [2639] = \nz.mem_2639_sv2v_reg ;
  assign \nz.mem [2638] = \nz.mem_2638_sv2v_reg ;
  assign \nz.mem [2637] = \nz.mem_2637_sv2v_reg ;
  assign \nz.mem [2636] = \nz.mem_2636_sv2v_reg ;
  assign \nz.mem [2635] = \nz.mem_2635_sv2v_reg ;
  assign \nz.mem [2634] = \nz.mem_2634_sv2v_reg ;
  assign \nz.mem [2633] = \nz.mem_2633_sv2v_reg ;
  assign \nz.mem [2632] = \nz.mem_2632_sv2v_reg ;
  assign \nz.mem [2631] = \nz.mem_2631_sv2v_reg ;
  assign \nz.mem [2630] = \nz.mem_2630_sv2v_reg ;
  assign \nz.mem [2629] = \nz.mem_2629_sv2v_reg ;
  assign \nz.mem [2628] = \nz.mem_2628_sv2v_reg ;
  assign \nz.mem [2627] = \nz.mem_2627_sv2v_reg ;
  assign \nz.mem [2626] = \nz.mem_2626_sv2v_reg ;
  assign \nz.mem [2625] = \nz.mem_2625_sv2v_reg ;
  assign \nz.mem [2624] = \nz.mem_2624_sv2v_reg ;
  assign \nz.mem [2623] = \nz.mem_2623_sv2v_reg ;
  assign \nz.mem [2622] = \nz.mem_2622_sv2v_reg ;
  assign \nz.mem [2621] = \nz.mem_2621_sv2v_reg ;
  assign \nz.mem [2620] = \nz.mem_2620_sv2v_reg ;
  assign \nz.mem [2619] = \nz.mem_2619_sv2v_reg ;
  assign \nz.mem [2618] = \nz.mem_2618_sv2v_reg ;
  assign \nz.mem [2617] = \nz.mem_2617_sv2v_reg ;
  assign \nz.mem [2616] = \nz.mem_2616_sv2v_reg ;
  assign \nz.mem [2615] = \nz.mem_2615_sv2v_reg ;
  assign \nz.mem [2614] = \nz.mem_2614_sv2v_reg ;
  assign \nz.mem [2613] = \nz.mem_2613_sv2v_reg ;
  assign \nz.mem [2612] = \nz.mem_2612_sv2v_reg ;
  assign \nz.mem [2611] = \nz.mem_2611_sv2v_reg ;
  assign \nz.mem [2610] = \nz.mem_2610_sv2v_reg ;
  assign \nz.mem [2609] = \nz.mem_2609_sv2v_reg ;
  assign \nz.mem [2608] = \nz.mem_2608_sv2v_reg ;
  assign \nz.mem [2607] = \nz.mem_2607_sv2v_reg ;
  assign \nz.mem [2606] = \nz.mem_2606_sv2v_reg ;
  assign \nz.mem [2605] = \nz.mem_2605_sv2v_reg ;
  assign \nz.mem [2604] = \nz.mem_2604_sv2v_reg ;
  assign \nz.mem [2603] = \nz.mem_2603_sv2v_reg ;
  assign \nz.mem [2602] = \nz.mem_2602_sv2v_reg ;
  assign \nz.mem [2601] = \nz.mem_2601_sv2v_reg ;
  assign \nz.mem [2600] = \nz.mem_2600_sv2v_reg ;
  assign \nz.mem [2599] = \nz.mem_2599_sv2v_reg ;
  assign \nz.mem [2598] = \nz.mem_2598_sv2v_reg ;
  assign \nz.mem [2597] = \nz.mem_2597_sv2v_reg ;
  assign \nz.mem [2596] = \nz.mem_2596_sv2v_reg ;
  assign \nz.mem [2595] = \nz.mem_2595_sv2v_reg ;
  assign \nz.mem [2594] = \nz.mem_2594_sv2v_reg ;
  assign \nz.mem [2593] = \nz.mem_2593_sv2v_reg ;
  assign \nz.mem [2592] = \nz.mem_2592_sv2v_reg ;
  assign \nz.mem [2591] = \nz.mem_2591_sv2v_reg ;
  assign \nz.mem [2590] = \nz.mem_2590_sv2v_reg ;
  assign \nz.mem [2589] = \nz.mem_2589_sv2v_reg ;
  assign \nz.mem [2588] = \nz.mem_2588_sv2v_reg ;
  assign \nz.mem [2587] = \nz.mem_2587_sv2v_reg ;
  assign \nz.mem [2586] = \nz.mem_2586_sv2v_reg ;
  assign \nz.mem [2585] = \nz.mem_2585_sv2v_reg ;
  assign \nz.mem [2584] = \nz.mem_2584_sv2v_reg ;
  assign \nz.mem [2583] = \nz.mem_2583_sv2v_reg ;
  assign \nz.mem [2582] = \nz.mem_2582_sv2v_reg ;
  assign \nz.mem [2581] = \nz.mem_2581_sv2v_reg ;
  assign \nz.mem [2580] = \nz.mem_2580_sv2v_reg ;
  assign \nz.mem [2579] = \nz.mem_2579_sv2v_reg ;
  assign \nz.mem [2578] = \nz.mem_2578_sv2v_reg ;
  assign \nz.mem [2577] = \nz.mem_2577_sv2v_reg ;
  assign \nz.mem [2576] = \nz.mem_2576_sv2v_reg ;
  assign \nz.mem [2575] = \nz.mem_2575_sv2v_reg ;
  assign \nz.mem [2574] = \nz.mem_2574_sv2v_reg ;
  assign \nz.mem [2573] = \nz.mem_2573_sv2v_reg ;
  assign \nz.mem [2572] = \nz.mem_2572_sv2v_reg ;
  assign \nz.mem [2571] = \nz.mem_2571_sv2v_reg ;
  assign \nz.mem [2570] = \nz.mem_2570_sv2v_reg ;
  assign \nz.mem [2569] = \nz.mem_2569_sv2v_reg ;
  assign \nz.mem [2568] = \nz.mem_2568_sv2v_reg ;
  assign \nz.mem [2567] = \nz.mem_2567_sv2v_reg ;
  assign \nz.mem [2566] = \nz.mem_2566_sv2v_reg ;
  assign \nz.mem [2565] = \nz.mem_2565_sv2v_reg ;
  assign \nz.mem [2564] = \nz.mem_2564_sv2v_reg ;
  assign \nz.mem [2563] = \nz.mem_2563_sv2v_reg ;
  assign \nz.mem [2562] = \nz.mem_2562_sv2v_reg ;
  assign \nz.mem [2561] = \nz.mem_2561_sv2v_reg ;
  assign \nz.mem [2560] = \nz.mem_2560_sv2v_reg ;
  assign \nz.mem [2559] = \nz.mem_2559_sv2v_reg ;
  assign \nz.mem [2558] = \nz.mem_2558_sv2v_reg ;
  assign \nz.mem [2557] = \nz.mem_2557_sv2v_reg ;
  assign \nz.mem [2556] = \nz.mem_2556_sv2v_reg ;
  assign \nz.mem [2555] = \nz.mem_2555_sv2v_reg ;
  assign \nz.mem [2554] = \nz.mem_2554_sv2v_reg ;
  assign \nz.mem [2553] = \nz.mem_2553_sv2v_reg ;
  assign \nz.mem [2552] = \nz.mem_2552_sv2v_reg ;
  assign \nz.mem [2551] = \nz.mem_2551_sv2v_reg ;
  assign \nz.mem [2550] = \nz.mem_2550_sv2v_reg ;
  assign \nz.mem [2549] = \nz.mem_2549_sv2v_reg ;
  assign \nz.mem [2548] = \nz.mem_2548_sv2v_reg ;
  assign \nz.mem [2547] = \nz.mem_2547_sv2v_reg ;
  assign \nz.mem [2546] = \nz.mem_2546_sv2v_reg ;
  assign \nz.mem [2545] = \nz.mem_2545_sv2v_reg ;
  assign \nz.mem [2544] = \nz.mem_2544_sv2v_reg ;
  assign \nz.mem [2543] = \nz.mem_2543_sv2v_reg ;
  assign \nz.mem [2542] = \nz.mem_2542_sv2v_reg ;
  assign \nz.mem [2541] = \nz.mem_2541_sv2v_reg ;
  assign \nz.mem [2540] = \nz.mem_2540_sv2v_reg ;
  assign \nz.mem [2539] = \nz.mem_2539_sv2v_reg ;
  assign \nz.mem [2538] = \nz.mem_2538_sv2v_reg ;
  assign \nz.mem [2537] = \nz.mem_2537_sv2v_reg ;
  assign \nz.mem [2536] = \nz.mem_2536_sv2v_reg ;
  assign \nz.mem [2535] = \nz.mem_2535_sv2v_reg ;
  assign \nz.mem [2534] = \nz.mem_2534_sv2v_reg ;
  assign \nz.mem [2533] = \nz.mem_2533_sv2v_reg ;
  assign \nz.mem [2532] = \nz.mem_2532_sv2v_reg ;
  assign \nz.mem [2531] = \nz.mem_2531_sv2v_reg ;
  assign \nz.mem [2530] = \nz.mem_2530_sv2v_reg ;
  assign \nz.mem [2529] = \nz.mem_2529_sv2v_reg ;
  assign \nz.mem [2528] = \nz.mem_2528_sv2v_reg ;
  assign \nz.mem [2527] = \nz.mem_2527_sv2v_reg ;
  assign \nz.mem [2526] = \nz.mem_2526_sv2v_reg ;
  assign \nz.mem [2525] = \nz.mem_2525_sv2v_reg ;
  assign \nz.mem [2524] = \nz.mem_2524_sv2v_reg ;
  assign \nz.mem [2523] = \nz.mem_2523_sv2v_reg ;
  assign \nz.mem [2522] = \nz.mem_2522_sv2v_reg ;
  assign \nz.mem [2521] = \nz.mem_2521_sv2v_reg ;
  assign \nz.mem [2520] = \nz.mem_2520_sv2v_reg ;
  assign \nz.mem [2519] = \nz.mem_2519_sv2v_reg ;
  assign \nz.mem [2518] = \nz.mem_2518_sv2v_reg ;
  assign \nz.mem [2517] = \nz.mem_2517_sv2v_reg ;
  assign \nz.mem [2516] = \nz.mem_2516_sv2v_reg ;
  assign \nz.mem [2515] = \nz.mem_2515_sv2v_reg ;
  assign \nz.mem [2514] = \nz.mem_2514_sv2v_reg ;
  assign \nz.mem [2513] = \nz.mem_2513_sv2v_reg ;
  assign \nz.mem [2512] = \nz.mem_2512_sv2v_reg ;
  assign \nz.mem [2511] = \nz.mem_2511_sv2v_reg ;
  assign \nz.mem [2510] = \nz.mem_2510_sv2v_reg ;
  assign \nz.mem [2509] = \nz.mem_2509_sv2v_reg ;
  assign \nz.mem [2508] = \nz.mem_2508_sv2v_reg ;
  assign \nz.mem [2507] = \nz.mem_2507_sv2v_reg ;
  assign \nz.mem [2506] = \nz.mem_2506_sv2v_reg ;
  assign \nz.mem [2505] = \nz.mem_2505_sv2v_reg ;
  assign \nz.mem [2504] = \nz.mem_2504_sv2v_reg ;
  assign \nz.mem [2503] = \nz.mem_2503_sv2v_reg ;
  assign \nz.mem [2502] = \nz.mem_2502_sv2v_reg ;
  assign \nz.mem [2501] = \nz.mem_2501_sv2v_reg ;
  assign \nz.mem [2500] = \nz.mem_2500_sv2v_reg ;
  assign \nz.mem [2499] = \nz.mem_2499_sv2v_reg ;
  assign \nz.mem [2498] = \nz.mem_2498_sv2v_reg ;
  assign \nz.mem [2497] = \nz.mem_2497_sv2v_reg ;
  assign \nz.mem [2496] = \nz.mem_2496_sv2v_reg ;
  assign \nz.mem [2495] = \nz.mem_2495_sv2v_reg ;
  assign \nz.mem [2494] = \nz.mem_2494_sv2v_reg ;
  assign \nz.mem [2493] = \nz.mem_2493_sv2v_reg ;
  assign \nz.mem [2492] = \nz.mem_2492_sv2v_reg ;
  assign \nz.mem [2491] = \nz.mem_2491_sv2v_reg ;
  assign \nz.mem [2490] = \nz.mem_2490_sv2v_reg ;
  assign \nz.mem [2489] = \nz.mem_2489_sv2v_reg ;
  assign \nz.mem [2488] = \nz.mem_2488_sv2v_reg ;
  assign \nz.mem [2487] = \nz.mem_2487_sv2v_reg ;
  assign \nz.mem [2486] = \nz.mem_2486_sv2v_reg ;
  assign \nz.mem [2485] = \nz.mem_2485_sv2v_reg ;
  assign \nz.mem [2484] = \nz.mem_2484_sv2v_reg ;
  assign \nz.mem [2483] = \nz.mem_2483_sv2v_reg ;
  assign \nz.mem [2482] = \nz.mem_2482_sv2v_reg ;
  assign \nz.mem [2481] = \nz.mem_2481_sv2v_reg ;
  assign \nz.mem [2480] = \nz.mem_2480_sv2v_reg ;
  assign \nz.mem [2479] = \nz.mem_2479_sv2v_reg ;
  assign \nz.mem [2478] = \nz.mem_2478_sv2v_reg ;
  assign \nz.mem [2477] = \nz.mem_2477_sv2v_reg ;
  assign \nz.mem [2476] = \nz.mem_2476_sv2v_reg ;
  assign \nz.mem [2475] = \nz.mem_2475_sv2v_reg ;
  assign \nz.mem [2474] = \nz.mem_2474_sv2v_reg ;
  assign \nz.mem [2473] = \nz.mem_2473_sv2v_reg ;
  assign \nz.mem [2472] = \nz.mem_2472_sv2v_reg ;
  assign \nz.mem [2471] = \nz.mem_2471_sv2v_reg ;
  assign \nz.mem [2470] = \nz.mem_2470_sv2v_reg ;
  assign \nz.mem [2469] = \nz.mem_2469_sv2v_reg ;
  assign \nz.mem [2468] = \nz.mem_2468_sv2v_reg ;
  assign \nz.mem [2467] = \nz.mem_2467_sv2v_reg ;
  assign \nz.mem [2466] = \nz.mem_2466_sv2v_reg ;
  assign \nz.mem [2465] = \nz.mem_2465_sv2v_reg ;
  assign \nz.mem [2464] = \nz.mem_2464_sv2v_reg ;
  assign \nz.mem [2463] = \nz.mem_2463_sv2v_reg ;
  assign \nz.mem [2462] = \nz.mem_2462_sv2v_reg ;
  assign \nz.mem [2461] = \nz.mem_2461_sv2v_reg ;
  assign \nz.mem [2460] = \nz.mem_2460_sv2v_reg ;
  assign \nz.mem [2459] = \nz.mem_2459_sv2v_reg ;
  assign \nz.mem [2458] = \nz.mem_2458_sv2v_reg ;
  assign \nz.mem [2457] = \nz.mem_2457_sv2v_reg ;
  assign \nz.mem [2456] = \nz.mem_2456_sv2v_reg ;
  assign \nz.mem [2455] = \nz.mem_2455_sv2v_reg ;
  assign \nz.mem [2454] = \nz.mem_2454_sv2v_reg ;
  assign \nz.mem [2453] = \nz.mem_2453_sv2v_reg ;
  assign \nz.mem [2452] = \nz.mem_2452_sv2v_reg ;
  assign \nz.mem [2451] = \nz.mem_2451_sv2v_reg ;
  assign \nz.mem [2450] = \nz.mem_2450_sv2v_reg ;
  assign \nz.mem [2449] = \nz.mem_2449_sv2v_reg ;
  assign \nz.mem [2448] = \nz.mem_2448_sv2v_reg ;
  assign \nz.mem [2447] = \nz.mem_2447_sv2v_reg ;
  assign \nz.mem [2446] = \nz.mem_2446_sv2v_reg ;
  assign \nz.mem [2445] = \nz.mem_2445_sv2v_reg ;
  assign \nz.mem [2444] = \nz.mem_2444_sv2v_reg ;
  assign \nz.mem [2443] = \nz.mem_2443_sv2v_reg ;
  assign \nz.mem [2442] = \nz.mem_2442_sv2v_reg ;
  assign \nz.mem [2441] = \nz.mem_2441_sv2v_reg ;
  assign \nz.mem [2440] = \nz.mem_2440_sv2v_reg ;
  assign \nz.mem [2439] = \nz.mem_2439_sv2v_reg ;
  assign \nz.mem [2438] = \nz.mem_2438_sv2v_reg ;
  assign \nz.mem [2437] = \nz.mem_2437_sv2v_reg ;
  assign \nz.mem [2436] = \nz.mem_2436_sv2v_reg ;
  assign \nz.mem [2435] = \nz.mem_2435_sv2v_reg ;
  assign \nz.mem [2434] = \nz.mem_2434_sv2v_reg ;
  assign \nz.mem [2433] = \nz.mem_2433_sv2v_reg ;
  assign \nz.mem [2432] = \nz.mem_2432_sv2v_reg ;
  assign \nz.mem [2431] = \nz.mem_2431_sv2v_reg ;
  assign \nz.mem [2430] = \nz.mem_2430_sv2v_reg ;
  assign \nz.mem [2429] = \nz.mem_2429_sv2v_reg ;
  assign \nz.mem [2428] = \nz.mem_2428_sv2v_reg ;
  assign \nz.mem [2427] = \nz.mem_2427_sv2v_reg ;
  assign \nz.mem [2426] = \nz.mem_2426_sv2v_reg ;
  assign \nz.mem [2425] = \nz.mem_2425_sv2v_reg ;
  assign \nz.mem [2424] = \nz.mem_2424_sv2v_reg ;
  assign \nz.mem [2423] = \nz.mem_2423_sv2v_reg ;
  assign \nz.mem [2422] = \nz.mem_2422_sv2v_reg ;
  assign \nz.mem [2421] = \nz.mem_2421_sv2v_reg ;
  assign \nz.mem [2420] = \nz.mem_2420_sv2v_reg ;
  assign \nz.mem [2419] = \nz.mem_2419_sv2v_reg ;
  assign \nz.mem [2418] = \nz.mem_2418_sv2v_reg ;
  assign \nz.mem [2417] = \nz.mem_2417_sv2v_reg ;
  assign \nz.mem [2416] = \nz.mem_2416_sv2v_reg ;
  assign \nz.mem [2415] = \nz.mem_2415_sv2v_reg ;
  assign \nz.mem [2414] = \nz.mem_2414_sv2v_reg ;
  assign \nz.mem [2413] = \nz.mem_2413_sv2v_reg ;
  assign \nz.mem [2412] = \nz.mem_2412_sv2v_reg ;
  assign \nz.mem [2411] = \nz.mem_2411_sv2v_reg ;
  assign \nz.mem [2410] = \nz.mem_2410_sv2v_reg ;
  assign \nz.mem [2409] = \nz.mem_2409_sv2v_reg ;
  assign \nz.mem [2408] = \nz.mem_2408_sv2v_reg ;
  assign \nz.mem [2407] = \nz.mem_2407_sv2v_reg ;
  assign \nz.mem [2406] = \nz.mem_2406_sv2v_reg ;
  assign \nz.mem [2405] = \nz.mem_2405_sv2v_reg ;
  assign \nz.mem [2404] = \nz.mem_2404_sv2v_reg ;
  assign \nz.mem [2403] = \nz.mem_2403_sv2v_reg ;
  assign \nz.mem [2402] = \nz.mem_2402_sv2v_reg ;
  assign \nz.mem [2401] = \nz.mem_2401_sv2v_reg ;
  assign \nz.mem [2400] = \nz.mem_2400_sv2v_reg ;
  assign \nz.mem [2399] = \nz.mem_2399_sv2v_reg ;
  assign \nz.mem [2398] = \nz.mem_2398_sv2v_reg ;
  assign \nz.mem [2397] = \nz.mem_2397_sv2v_reg ;
  assign \nz.mem [2396] = \nz.mem_2396_sv2v_reg ;
  assign \nz.mem [2395] = \nz.mem_2395_sv2v_reg ;
  assign \nz.mem [2394] = \nz.mem_2394_sv2v_reg ;
  assign \nz.mem [2393] = \nz.mem_2393_sv2v_reg ;
  assign \nz.mem [2392] = \nz.mem_2392_sv2v_reg ;
  assign \nz.mem [2391] = \nz.mem_2391_sv2v_reg ;
  assign \nz.mem [2390] = \nz.mem_2390_sv2v_reg ;
  assign \nz.mem [2389] = \nz.mem_2389_sv2v_reg ;
  assign \nz.mem [2388] = \nz.mem_2388_sv2v_reg ;
  assign \nz.mem [2387] = \nz.mem_2387_sv2v_reg ;
  assign \nz.mem [2386] = \nz.mem_2386_sv2v_reg ;
  assign \nz.mem [2385] = \nz.mem_2385_sv2v_reg ;
  assign \nz.mem [2384] = \nz.mem_2384_sv2v_reg ;
  assign \nz.mem [2383] = \nz.mem_2383_sv2v_reg ;
  assign \nz.mem [2382] = \nz.mem_2382_sv2v_reg ;
  assign \nz.mem [2381] = \nz.mem_2381_sv2v_reg ;
  assign \nz.mem [2380] = \nz.mem_2380_sv2v_reg ;
  assign \nz.mem [2379] = \nz.mem_2379_sv2v_reg ;
  assign \nz.mem [2378] = \nz.mem_2378_sv2v_reg ;
  assign \nz.mem [2377] = \nz.mem_2377_sv2v_reg ;
  assign \nz.mem [2376] = \nz.mem_2376_sv2v_reg ;
  assign \nz.mem [2375] = \nz.mem_2375_sv2v_reg ;
  assign \nz.mem [2374] = \nz.mem_2374_sv2v_reg ;
  assign \nz.mem [2373] = \nz.mem_2373_sv2v_reg ;
  assign \nz.mem [2372] = \nz.mem_2372_sv2v_reg ;
  assign \nz.mem [2371] = \nz.mem_2371_sv2v_reg ;
  assign \nz.mem [2370] = \nz.mem_2370_sv2v_reg ;
  assign \nz.mem [2369] = \nz.mem_2369_sv2v_reg ;
  assign \nz.mem [2368] = \nz.mem_2368_sv2v_reg ;
  assign \nz.mem [2367] = \nz.mem_2367_sv2v_reg ;
  assign \nz.mem [2366] = \nz.mem_2366_sv2v_reg ;
  assign \nz.mem [2365] = \nz.mem_2365_sv2v_reg ;
  assign \nz.mem [2364] = \nz.mem_2364_sv2v_reg ;
  assign \nz.mem [2363] = \nz.mem_2363_sv2v_reg ;
  assign \nz.mem [2362] = \nz.mem_2362_sv2v_reg ;
  assign \nz.mem [2361] = \nz.mem_2361_sv2v_reg ;
  assign \nz.mem [2360] = \nz.mem_2360_sv2v_reg ;
  assign \nz.mem [2359] = \nz.mem_2359_sv2v_reg ;
  assign \nz.mem [2358] = \nz.mem_2358_sv2v_reg ;
  assign \nz.mem [2357] = \nz.mem_2357_sv2v_reg ;
  assign \nz.mem [2356] = \nz.mem_2356_sv2v_reg ;
  assign \nz.mem [2355] = \nz.mem_2355_sv2v_reg ;
  assign \nz.mem [2354] = \nz.mem_2354_sv2v_reg ;
  assign \nz.mem [2353] = \nz.mem_2353_sv2v_reg ;
  assign \nz.mem [2352] = \nz.mem_2352_sv2v_reg ;
  assign \nz.mem [2351] = \nz.mem_2351_sv2v_reg ;
  assign \nz.mem [2350] = \nz.mem_2350_sv2v_reg ;
  assign \nz.mem [2349] = \nz.mem_2349_sv2v_reg ;
  assign \nz.mem [2348] = \nz.mem_2348_sv2v_reg ;
  assign \nz.mem [2347] = \nz.mem_2347_sv2v_reg ;
  assign \nz.mem [2346] = \nz.mem_2346_sv2v_reg ;
  assign \nz.mem [2345] = \nz.mem_2345_sv2v_reg ;
  assign \nz.mem [2344] = \nz.mem_2344_sv2v_reg ;
  assign \nz.mem [2343] = \nz.mem_2343_sv2v_reg ;
  assign \nz.mem [2342] = \nz.mem_2342_sv2v_reg ;
  assign \nz.mem [2341] = \nz.mem_2341_sv2v_reg ;
  assign \nz.mem [2340] = \nz.mem_2340_sv2v_reg ;
  assign \nz.mem [2339] = \nz.mem_2339_sv2v_reg ;
  assign \nz.mem [2338] = \nz.mem_2338_sv2v_reg ;
  assign \nz.mem [2337] = \nz.mem_2337_sv2v_reg ;
  assign \nz.mem [2336] = \nz.mem_2336_sv2v_reg ;
  assign \nz.mem [2335] = \nz.mem_2335_sv2v_reg ;
  assign \nz.mem [2334] = \nz.mem_2334_sv2v_reg ;
  assign \nz.mem [2333] = \nz.mem_2333_sv2v_reg ;
  assign \nz.mem [2332] = \nz.mem_2332_sv2v_reg ;
  assign \nz.mem [2331] = \nz.mem_2331_sv2v_reg ;
  assign \nz.mem [2330] = \nz.mem_2330_sv2v_reg ;
  assign \nz.mem [2329] = \nz.mem_2329_sv2v_reg ;
  assign \nz.mem [2328] = \nz.mem_2328_sv2v_reg ;
  assign \nz.mem [2327] = \nz.mem_2327_sv2v_reg ;
  assign \nz.mem [2326] = \nz.mem_2326_sv2v_reg ;
  assign \nz.mem [2325] = \nz.mem_2325_sv2v_reg ;
  assign \nz.mem [2324] = \nz.mem_2324_sv2v_reg ;
  assign \nz.mem [2323] = \nz.mem_2323_sv2v_reg ;
  assign \nz.mem [2322] = \nz.mem_2322_sv2v_reg ;
  assign \nz.mem [2321] = \nz.mem_2321_sv2v_reg ;
  assign \nz.mem [2320] = \nz.mem_2320_sv2v_reg ;
  assign \nz.mem [2319] = \nz.mem_2319_sv2v_reg ;
  assign \nz.mem [2318] = \nz.mem_2318_sv2v_reg ;
  assign \nz.mem [2317] = \nz.mem_2317_sv2v_reg ;
  assign \nz.mem [2316] = \nz.mem_2316_sv2v_reg ;
  assign \nz.mem [2315] = \nz.mem_2315_sv2v_reg ;
  assign \nz.mem [2314] = \nz.mem_2314_sv2v_reg ;
  assign \nz.mem [2313] = \nz.mem_2313_sv2v_reg ;
  assign \nz.mem [2312] = \nz.mem_2312_sv2v_reg ;
  assign \nz.mem [2311] = \nz.mem_2311_sv2v_reg ;
  assign \nz.mem [2310] = \nz.mem_2310_sv2v_reg ;
  assign \nz.mem [2309] = \nz.mem_2309_sv2v_reg ;
  assign \nz.mem [2308] = \nz.mem_2308_sv2v_reg ;
  assign \nz.mem [2307] = \nz.mem_2307_sv2v_reg ;
  assign \nz.mem [2306] = \nz.mem_2306_sv2v_reg ;
  assign \nz.mem [2305] = \nz.mem_2305_sv2v_reg ;
  assign \nz.mem [2304] = \nz.mem_2304_sv2v_reg ;
  assign \nz.mem [2303] = \nz.mem_2303_sv2v_reg ;
  assign \nz.mem [2302] = \nz.mem_2302_sv2v_reg ;
  assign \nz.mem [2301] = \nz.mem_2301_sv2v_reg ;
  assign \nz.mem [2300] = \nz.mem_2300_sv2v_reg ;
  assign \nz.mem [2299] = \nz.mem_2299_sv2v_reg ;
  assign \nz.mem [2298] = \nz.mem_2298_sv2v_reg ;
  assign \nz.mem [2297] = \nz.mem_2297_sv2v_reg ;
  assign \nz.mem [2296] = \nz.mem_2296_sv2v_reg ;
  assign \nz.mem [2295] = \nz.mem_2295_sv2v_reg ;
  assign \nz.mem [2294] = \nz.mem_2294_sv2v_reg ;
  assign \nz.mem [2293] = \nz.mem_2293_sv2v_reg ;
  assign \nz.mem [2292] = \nz.mem_2292_sv2v_reg ;
  assign \nz.mem [2291] = \nz.mem_2291_sv2v_reg ;
  assign \nz.mem [2290] = \nz.mem_2290_sv2v_reg ;
  assign \nz.mem [2289] = \nz.mem_2289_sv2v_reg ;
  assign \nz.mem [2288] = \nz.mem_2288_sv2v_reg ;
  assign \nz.mem [2287] = \nz.mem_2287_sv2v_reg ;
  assign \nz.mem [2286] = \nz.mem_2286_sv2v_reg ;
  assign \nz.mem [2285] = \nz.mem_2285_sv2v_reg ;
  assign \nz.mem [2284] = \nz.mem_2284_sv2v_reg ;
  assign \nz.mem [2283] = \nz.mem_2283_sv2v_reg ;
  assign \nz.mem [2282] = \nz.mem_2282_sv2v_reg ;
  assign \nz.mem [2281] = \nz.mem_2281_sv2v_reg ;
  assign \nz.mem [2280] = \nz.mem_2280_sv2v_reg ;
  assign \nz.mem [2279] = \nz.mem_2279_sv2v_reg ;
  assign \nz.mem [2278] = \nz.mem_2278_sv2v_reg ;
  assign \nz.mem [2277] = \nz.mem_2277_sv2v_reg ;
  assign \nz.mem [2276] = \nz.mem_2276_sv2v_reg ;
  assign \nz.mem [2275] = \nz.mem_2275_sv2v_reg ;
  assign \nz.mem [2274] = \nz.mem_2274_sv2v_reg ;
  assign \nz.mem [2273] = \nz.mem_2273_sv2v_reg ;
  assign \nz.mem [2272] = \nz.mem_2272_sv2v_reg ;
  assign \nz.mem [2271] = \nz.mem_2271_sv2v_reg ;
  assign \nz.mem [2270] = \nz.mem_2270_sv2v_reg ;
  assign \nz.mem [2269] = \nz.mem_2269_sv2v_reg ;
  assign \nz.mem [2268] = \nz.mem_2268_sv2v_reg ;
  assign \nz.mem [2267] = \nz.mem_2267_sv2v_reg ;
  assign \nz.mem [2266] = \nz.mem_2266_sv2v_reg ;
  assign \nz.mem [2265] = \nz.mem_2265_sv2v_reg ;
  assign \nz.mem [2264] = \nz.mem_2264_sv2v_reg ;
  assign \nz.mem [2263] = \nz.mem_2263_sv2v_reg ;
  assign \nz.mem [2262] = \nz.mem_2262_sv2v_reg ;
  assign \nz.mem [2261] = \nz.mem_2261_sv2v_reg ;
  assign \nz.mem [2260] = \nz.mem_2260_sv2v_reg ;
  assign \nz.mem [2259] = \nz.mem_2259_sv2v_reg ;
  assign \nz.mem [2258] = \nz.mem_2258_sv2v_reg ;
  assign \nz.mem [2257] = \nz.mem_2257_sv2v_reg ;
  assign \nz.mem [2256] = \nz.mem_2256_sv2v_reg ;
  assign \nz.mem [2255] = \nz.mem_2255_sv2v_reg ;
  assign \nz.mem [2254] = \nz.mem_2254_sv2v_reg ;
  assign \nz.mem [2253] = \nz.mem_2253_sv2v_reg ;
  assign \nz.mem [2252] = \nz.mem_2252_sv2v_reg ;
  assign \nz.mem [2251] = \nz.mem_2251_sv2v_reg ;
  assign \nz.mem [2250] = \nz.mem_2250_sv2v_reg ;
  assign \nz.mem [2249] = \nz.mem_2249_sv2v_reg ;
  assign \nz.mem [2248] = \nz.mem_2248_sv2v_reg ;
  assign \nz.mem [2247] = \nz.mem_2247_sv2v_reg ;
  assign \nz.mem [2246] = \nz.mem_2246_sv2v_reg ;
  assign \nz.mem [2245] = \nz.mem_2245_sv2v_reg ;
  assign \nz.mem [2244] = \nz.mem_2244_sv2v_reg ;
  assign \nz.mem [2243] = \nz.mem_2243_sv2v_reg ;
  assign \nz.mem [2242] = \nz.mem_2242_sv2v_reg ;
  assign \nz.mem [2241] = \nz.mem_2241_sv2v_reg ;
  assign \nz.mem [2240] = \nz.mem_2240_sv2v_reg ;
  assign \nz.mem [2239] = \nz.mem_2239_sv2v_reg ;
  assign \nz.mem [2238] = \nz.mem_2238_sv2v_reg ;
  assign \nz.mem [2237] = \nz.mem_2237_sv2v_reg ;
  assign \nz.mem [2236] = \nz.mem_2236_sv2v_reg ;
  assign \nz.mem [2235] = \nz.mem_2235_sv2v_reg ;
  assign \nz.mem [2234] = \nz.mem_2234_sv2v_reg ;
  assign \nz.mem [2233] = \nz.mem_2233_sv2v_reg ;
  assign \nz.mem [2232] = \nz.mem_2232_sv2v_reg ;
  assign \nz.mem [2231] = \nz.mem_2231_sv2v_reg ;
  assign \nz.mem [2230] = \nz.mem_2230_sv2v_reg ;
  assign \nz.mem [2229] = \nz.mem_2229_sv2v_reg ;
  assign \nz.mem [2228] = \nz.mem_2228_sv2v_reg ;
  assign \nz.mem [2227] = \nz.mem_2227_sv2v_reg ;
  assign \nz.mem [2226] = \nz.mem_2226_sv2v_reg ;
  assign \nz.mem [2225] = \nz.mem_2225_sv2v_reg ;
  assign \nz.mem [2224] = \nz.mem_2224_sv2v_reg ;
  assign \nz.mem [2223] = \nz.mem_2223_sv2v_reg ;
  assign \nz.mem [2222] = \nz.mem_2222_sv2v_reg ;
  assign \nz.mem [2221] = \nz.mem_2221_sv2v_reg ;
  assign \nz.mem [2220] = \nz.mem_2220_sv2v_reg ;
  assign \nz.mem [2219] = \nz.mem_2219_sv2v_reg ;
  assign \nz.mem [2218] = \nz.mem_2218_sv2v_reg ;
  assign \nz.mem [2217] = \nz.mem_2217_sv2v_reg ;
  assign \nz.mem [2216] = \nz.mem_2216_sv2v_reg ;
  assign \nz.mem [2215] = \nz.mem_2215_sv2v_reg ;
  assign \nz.mem [2214] = \nz.mem_2214_sv2v_reg ;
  assign \nz.mem [2213] = \nz.mem_2213_sv2v_reg ;
  assign \nz.mem [2212] = \nz.mem_2212_sv2v_reg ;
  assign \nz.mem [2211] = \nz.mem_2211_sv2v_reg ;
  assign \nz.mem [2210] = \nz.mem_2210_sv2v_reg ;
  assign \nz.mem [2209] = \nz.mem_2209_sv2v_reg ;
  assign \nz.mem [2208] = \nz.mem_2208_sv2v_reg ;
  assign \nz.mem [2207] = \nz.mem_2207_sv2v_reg ;
  assign \nz.mem [2206] = \nz.mem_2206_sv2v_reg ;
  assign \nz.mem [2205] = \nz.mem_2205_sv2v_reg ;
  assign \nz.mem [2204] = \nz.mem_2204_sv2v_reg ;
  assign \nz.mem [2203] = \nz.mem_2203_sv2v_reg ;
  assign \nz.mem [2202] = \nz.mem_2202_sv2v_reg ;
  assign \nz.mem [2201] = \nz.mem_2201_sv2v_reg ;
  assign \nz.mem [2200] = \nz.mem_2200_sv2v_reg ;
  assign \nz.mem [2199] = \nz.mem_2199_sv2v_reg ;
  assign \nz.mem [2198] = \nz.mem_2198_sv2v_reg ;
  assign \nz.mem [2197] = \nz.mem_2197_sv2v_reg ;
  assign \nz.mem [2196] = \nz.mem_2196_sv2v_reg ;
  assign \nz.mem [2195] = \nz.mem_2195_sv2v_reg ;
  assign \nz.mem [2194] = \nz.mem_2194_sv2v_reg ;
  assign \nz.mem [2193] = \nz.mem_2193_sv2v_reg ;
  assign \nz.mem [2192] = \nz.mem_2192_sv2v_reg ;
  assign \nz.mem [2191] = \nz.mem_2191_sv2v_reg ;
  assign \nz.mem [2190] = \nz.mem_2190_sv2v_reg ;
  assign \nz.mem [2189] = \nz.mem_2189_sv2v_reg ;
  assign \nz.mem [2188] = \nz.mem_2188_sv2v_reg ;
  assign \nz.mem [2187] = \nz.mem_2187_sv2v_reg ;
  assign \nz.mem [2186] = \nz.mem_2186_sv2v_reg ;
  assign \nz.mem [2185] = \nz.mem_2185_sv2v_reg ;
  assign \nz.mem [2184] = \nz.mem_2184_sv2v_reg ;
  assign \nz.mem [2183] = \nz.mem_2183_sv2v_reg ;
  assign \nz.mem [2182] = \nz.mem_2182_sv2v_reg ;
  assign \nz.mem [2181] = \nz.mem_2181_sv2v_reg ;
  assign \nz.mem [2180] = \nz.mem_2180_sv2v_reg ;
  assign \nz.mem [2179] = \nz.mem_2179_sv2v_reg ;
  assign \nz.mem [2178] = \nz.mem_2178_sv2v_reg ;
  assign \nz.mem [2177] = \nz.mem_2177_sv2v_reg ;
  assign \nz.mem [2176] = \nz.mem_2176_sv2v_reg ;
  assign \nz.mem [2175] = \nz.mem_2175_sv2v_reg ;
  assign \nz.mem [2174] = \nz.mem_2174_sv2v_reg ;
  assign \nz.mem [2173] = \nz.mem_2173_sv2v_reg ;
  assign \nz.mem [2172] = \nz.mem_2172_sv2v_reg ;
  assign \nz.mem [2171] = \nz.mem_2171_sv2v_reg ;
  assign \nz.mem [2170] = \nz.mem_2170_sv2v_reg ;
  assign \nz.mem [2169] = \nz.mem_2169_sv2v_reg ;
  assign \nz.mem [2168] = \nz.mem_2168_sv2v_reg ;
  assign \nz.mem [2167] = \nz.mem_2167_sv2v_reg ;
  assign \nz.mem [2166] = \nz.mem_2166_sv2v_reg ;
  assign \nz.mem [2165] = \nz.mem_2165_sv2v_reg ;
  assign \nz.mem [2164] = \nz.mem_2164_sv2v_reg ;
  assign \nz.mem [2163] = \nz.mem_2163_sv2v_reg ;
  assign \nz.mem [2162] = \nz.mem_2162_sv2v_reg ;
  assign \nz.mem [2161] = \nz.mem_2161_sv2v_reg ;
  assign \nz.mem [2160] = \nz.mem_2160_sv2v_reg ;
  assign \nz.mem [2159] = \nz.mem_2159_sv2v_reg ;
  assign \nz.mem [2158] = \nz.mem_2158_sv2v_reg ;
  assign \nz.mem [2157] = \nz.mem_2157_sv2v_reg ;
  assign \nz.mem [2156] = \nz.mem_2156_sv2v_reg ;
  assign \nz.mem [2155] = \nz.mem_2155_sv2v_reg ;
  assign \nz.mem [2154] = \nz.mem_2154_sv2v_reg ;
  assign \nz.mem [2153] = \nz.mem_2153_sv2v_reg ;
  assign \nz.mem [2152] = \nz.mem_2152_sv2v_reg ;
  assign \nz.mem [2151] = \nz.mem_2151_sv2v_reg ;
  assign \nz.mem [2150] = \nz.mem_2150_sv2v_reg ;
  assign \nz.mem [2149] = \nz.mem_2149_sv2v_reg ;
  assign \nz.mem [2148] = \nz.mem_2148_sv2v_reg ;
  assign \nz.mem [2147] = \nz.mem_2147_sv2v_reg ;
  assign \nz.mem [2146] = \nz.mem_2146_sv2v_reg ;
  assign \nz.mem [2145] = \nz.mem_2145_sv2v_reg ;
  assign \nz.mem [2144] = \nz.mem_2144_sv2v_reg ;
  assign \nz.mem [2143] = \nz.mem_2143_sv2v_reg ;
  assign \nz.mem [2142] = \nz.mem_2142_sv2v_reg ;
  assign \nz.mem [2141] = \nz.mem_2141_sv2v_reg ;
  assign \nz.mem [2140] = \nz.mem_2140_sv2v_reg ;
  assign \nz.mem [2139] = \nz.mem_2139_sv2v_reg ;
  assign \nz.mem [2138] = \nz.mem_2138_sv2v_reg ;
  assign \nz.mem [2137] = \nz.mem_2137_sv2v_reg ;
  assign \nz.mem [2136] = \nz.mem_2136_sv2v_reg ;
  assign \nz.mem [2135] = \nz.mem_2135_sv2v_reg ;
  assign \nz.mem [2134] = \nz.mem_2134_sv2v_reg ;
  assign \nz.mem [2133] = \nz.mem_2133_sv2v_reg ;
  assign \nz.mem [2132] = \nz.mem_2132_sv2v_reg ;
  assign \nz.mem [2131] = \nz.mem_2131_sv2v_reg ;
  assign \nz.mem [2130] = \nz.mem_2130_sv2v_reg ;
  assign \nz.mem [2129] = \nz.mem_2129_sv2v_reg ;
  assign \nz.mem [2128] = \nz.mem_2128_sv2v_reg ;
  assign \nz.mem [2127] = \nz.mem_2127_sv2v_reg ;
  assign \nz.mem [2126] = \nz.mem_2126_sv2v_reg ;
  assign \nz.mem [2125] = \nz.mem_2125_sv2v_reg ;
  assign \nz.mem [2124] = \nz.mem_2124_sv2v_reg ;
  assign \nz.mem [2123] = \nz.mem_2123_sv2v_reg ;
  assign \nz.mem [2122] = \nz.mem_2122_sv2v_reg ;
  assign \nz.mem [2121] = \nz.mem_2121_sv2v_reg ;
  assign \nz.mem [2120] = \nz.mem_2120_sv2v_reg ;
  assign \nz.mem [2119] = \nz.mem_2119_sv2v_reg ;
  assign \nz.mem [2118] = \nz.mem_2118_sv2v_reg ;
  assign \nz.mem [2117] = \nz.mem_2117_sv2v_reg ;
  assign \nz.mem [2116] = \nz.mem_2116_sv2v_reg ;
  assign \nz.mem [2115] = \nz.mem_2115_sv2v_reg ;
  assign \nz.mem [2114] = \nz.mem_2114_sv2v_reg ;
  assign \nz.mem [2113] = \nz.mem_2113_sv2v_reg ;
  assign \nz.mem [2112] = \nz.mem_2112_sv2v_reg ;
  assign \nz.mem [2111] = \nz.mem_2111_sv2v_reg ;
  assign \nz.mem [2110] = \nz.mem_2110_sv2v_reg ;
  assign \nz.mem [2109] = \nz.mem_2109_sv2v_reg ;
  assign \nz.mem [2108] = \nz.mem_2108_sv2v_reg ;
  assign \nz.mem [2107] = \nz.mem_2107_sv2v_reg ;
  assign \nz.mem [2106] = \nz.mem_2106_sv2v_reg ;
  assign \nz.mem [2105] = \nz.mem_2105_sv2v_reg ;
  assign \nz.mem [2104] = \nz.mem_2104_sv2v_reg ;
  assign \nz.mem [2103] = \nz.mem_2103_sv2v_reg ;
  assign \nz.mem [2102] = \nz.mem_2102_sv2v_reg ;
  assign \nz.mem [2101] = \nz.mem_2101_sv2v_reg ;
  assign \nz.mem [2100] = \nz.mem_2100_sv2v_reg ;
  assign \nz.mem [2099] = \nz.mem_2099_sv2v_reg ;
  assign \nz.mem [2098] = \nz.mem_2098_sv2v_reg ;
  assign \nz.mem [2097] = \nz.mem_2097_sv2v_reg ;
  assign \nz.mem [2096] = \nz.mem_2096_sv2v_reg ;
  assign \nz.mem [2095] = \nz.mem_2095_sv2v_reg ;
  assign \nz.mem [2094] = \nz.mem_2094_sv2v_reg ;
  assign \nz.mem [2093] = \nz.mem_2093_sv2v_reg ;
  assign \nz.mem [2092] = \nz.mem_2092_sv2v_reg ;
  assign \nz.mem [2091] = \nz.mem_2091_sv2v_reg ;
  assign \nz.mem [2090] = \nz.mem_2090_sv2v_reg ;
  assign \nz.mem [2089] = \nz.mem_2089_sv2v_reg ;
  assign \nz.mem [2088] = \nz.mem_2088_sv2v_reg ;
  assign \nz.mem [2087] = \nz.mem_2087_sv2v_reg ;
  assign \nz.mem [2086] = \nz.mem_2086_sv2v_reg ;
  assign \nz.mem [2085] = \nz.mem_2085_sv2v_reg ;
  assign \nz.mem [2084] = \nz.mem_2084_sv2v_reg ;
  assign \nz.mem [2083] = \nz.mem_2083_sv2v_reg ;
  assign \nz.mem [2082] = \nz.mem_2082_sv2v_reg ;
  assign \nz.mem [2081] = \nz.mem_2081_sv2v_reg ;
  assign \nz.mem [2080] = \nz.mem_2080_sv2v_reg ;
  assign \nz.mem [2079] = \nz.mem_2079_sv2v_reg ;
  assign \nz.mem [2078] = \nz.mem_2078_sv2v_reg ;
  assign \nz.mem [2077] = \nz.mem_2077_sv2v_reg ;
  assign \nz.mem [2076] = \nz.mem_2076_sv2v_reg ;
  assign \nz.mem [2075] = \nz.mem_2075_sv2v_reg ;
  assign \nz.mem [2074] = \nz.mem_2074_sv2v_reg ;
  assign \nz.mem [2073] = \nz.mem_2073_sv2v_reg ;
  assign \nz.mem [2072] = \nz.mem_2072_sv2v_reg ;
  assign \nz.mem [2071] = \nz.mem_2071_sv2v_reg ;
  assign \nz.mem [2070] = \nz.mem_2070_sv2v_reg ;
  assign \nz.mem [2069] = \nz.mem_2069_sv2v_reg ;
  assign \nz.mem [2068] = \nz.mem_2068_sv2v_reg ;
  assign \nz.mem [2067] = \nz.mem_2067_sv2v_reg ;
  assign \nz.mem [2066] = \nz.mem_2066_sv2v_reg ;
  assign \nz.mem [2065] = \nz.mem_2065_sv2v_reg ;
  assign \nz.mem [2064] = \nz.mem_2064_sv2v_reg ;
  assign \nz.mem [2063] = \nz.mem_2063_sv2v_reg ;
  assign \nz.mem [2062] = \nz.mem_2062_sv2v_reg ;
  assign \nz.mem [2061] = \nz.mem_2061_sv2v_reg ;
  assign \nz.mem [2060] = \nz.mem_2060_sv2v_reg ;
  assign \nz.mem [2059] = \nz.mem_2059_sv2v_reg ;
  assign \nz.mem [2058] = \nz.mem_2058_sv2v_reg ;
  assign \nz.mem [2057] = \nz.mem_2057_sv2v_reg ;
  assign \nz.mem [2056] = \nz.mem_2056_sv2v_reg ;
  assign \nz.mem [2055] = \nz.mem_2055_sv2v_reg ;
  assign \nz.mem [2054] = \nz.mem_2054_sv2v_reg ;
  assign \nz.mem [2053] = \nz.mem_2053_sv2v_reg ;
  assign \nz.mem [2052] = \nz.mem_2052_sv2v_reg ;
  assign \nz.mem [2051] = \nz.mem_2051_sv2v_reg ;
  assign \nz.mem [2050] = \nz.mem_2050_sv2v_reg ;
  assign \nz.mem [2049] = \nz.mem_2049_sv2v_reg ;
  assign \nz.mem [2048] = \nz.mem_2048_sv2v_reg ;
  assign \nz.mem [2047] = \nz.mem_2047_sv2v_reg ;
  assign \nz.mem [2046] = \nz.mem_2046_sv2v_reg ;
  assign \nz.mem [2045] = \nz.mem_2045_sv2v_reg ;
  assign \nz.mem [2044] = \nz.mem_2044_sv2v_reg ;
  assign \nz.mem [2043] = \nz.mem_2043_sv2v_reg ;
  assign \nz.mem [2042] = \nz.mem_2042_sv2v_reg ;
  assign \nz.mem [2041] = \nz.mem_2041_sv2v_reg ;
  assign \nz.mem [2040] = \nz.mem_2040_sv2v_reg ;
  assign \nz.mem [2039] = \nz.mem_2039_sv2v_reg ;
  assign \nz.mem [2038] = \nz.mem_2038_sv2v_reg ;
  assign \nz.mem [2037] = \nz.mem_2037_sv2v_reg ;
  assign \nz.mem [2036] = \nz.mem_2036_sv2v_reg ;
  assign \nz.mem [2035] = \nz.mem_2035_sv2v_reg ;
  assign \nz.mem [2034] = \nz.mem_2034_sv2v_reg ;
  assign \nz.mem [2033] = \nz.mem_2033_sv2v_reg ;
  assign \nz.mem [2032] = \nz.mem_2032_sv2v_reg ;
  assign \nz.mem [2031] = \nz.mem_2031_sv2v_reg ;
  assign \nz.mem [2030] = \nz.mem_2030_sv2v_reg ;
  assign \nz.mem [2029] = \nz.mem_2029_sv2v_reg ;
  assign \nz.mem [2028] = \nz.mem_2028_sv2v_reg ;
  assign \nz.mem [2027] = \nz.mem_2027_sv2v_reg ;
  assign \nz.mem [2026] = \nz.mem_2026_sv2v_reg ;
  assign \nz.mem [2025] = \nz.mem_2025_sv2v_reg ;
  assign \nz.mem [2024] = \nz.mem_2024_sv2v_reg ;
  assign \nz.mem [2023] = \nz.mem_2023_sv2v_reg ;
  assign \nz.mem [2022] = \nz.mem_2022_sv2v_reg ;
  assign \nz.mem [2021] = \nz.mem_2021_sv2v_reg ;
  assign \nz.mem [2020] = \nz.mem_2020_sv2v_reg ;
  assign \nz.mem [2019] = \nz.mem_2019_sv2v_reg ;
  assign \nz.mem [2018] = \nz.mem_2018_sv2v_reg ;
  assign \nz.mem [2017] = \nz.mem_2017_sv2v_reg ;
  assign \nz.mem [2016] = \nz.mem_2016_sv2v_reg ;
  assign \nz.mem [2015] = \nz.mem_2015_sv2v_reg ;
  assign \nz.mem [2014] = \nz.mem_2014_sv2v_reg ;
  assign \nz.mem [2013] = \nz.mem_2013_sv2v_reg ;
  assign \nz.mem [2012] = \nz.mem_2012_sv2v_reg ;
  assign \nz.mem [2011] = \nz.mem_2011_sv2v_reg ;
  assign \nz.mem [2010] = \nz.mem_2010_sv2v_reg ;
  assign \nz.mem [2009] = \nz.mem_2009_sv2v_reg ;
  assign \nz.mem [2008] = \nz.mem_2008_sv2v_reg ;
  assign \nz.mem [2007] = \nz.mem_2007_sv2v_reg ;
  assign \nz.mem [2006] = \nz.mem_2006_sv2v_reg ;
  assign \nz.mem [2005] = \nz.mem_2005_sv2v_reg ;
  assign \nz.mem [2004] = \nz.mem_2004_sv2v_reg ;
  assign \nz.mem [2003] = \nz.mem_2003_sv2v_reg ;
  assign \nz.mem [2002] = \nz.mem_2002_sv2v_reg ;
  assign \nz.mem [2001] = \nz.mem_2001_sv2v_reg ;
  assign \nz.mem [2000] = \nz.mem_2000_sv2v_reg ;
  assign \nz.mem [1999] = \nz.mem_1999_sv2v_reg ;
  assign \nz.mem [1998] = \nz.mem_1998_sv2v_reg ;
  assign \nz.mem [1997] = \nz.mem_1997_sv2v_reg ;
  assign \nz.mem [1996] = \nz.mem_1996_sv2v_reg ;
  assign \nz.mem [1995] = \nz.mem_1995_sv2v_reg ;
  assign \nz.mem [1994] = \nz.mem_1994_sv2v_reg ;
  assign \nz.mem [1993] = \nz.mem_1993_sv2v_reg ;
  assign \nz.mem [1992] = \nz.mem_1992_sv2v_reg ;
  assign \nz.mem [1991] = \nz.mem_1991_sv2v_reg ;
  assign \nz.mem [1990] = \nz.mem_1990_sv2v_reg ;
  assign \nz.mem [1989] = \nz.mem_1989_sv2v_reg ;
  assign \nz.mem [1988] = \nz.mem_1988_sv2v_reg ;
  assign \nz.mem [1987] = \nz.mem_1987_sv2v_reg ;
  assign \nz.mem [1986] = \nz.mem_1986_sv2v_reg ;
  assign \nz.mem [1985] = \nz.mem_1985_sv2v_reg ;
  assign \nz.mem [1984] = \nz.mem_1984_sv2v_reg ;
  assign \nz.mem [1983] = \nz.mem_1983_sv2v_reg ;
  assign \nz.mem [1982] = \nz.mem_1982_sv2v_reg ;
  assign \nz.mem [1981] = \nz.mem_1981_sv2v_reg ;
  assign \nz.mem [1980] = \nz.mem_1980_sv2v_reg ;
  assign \nz.mem [1979] = \nz.mem_1979_sv2v_reg ;
  assign \nz.mem [1978] = \nz.mem_1978_sv2v_reg ;
  assign \nz.mem [1977] = \nz.mem_1977_sv2v_reg ;
  assign \nz.mem [1976] = \nz.mem_1976_sv2v_reg ;
  assign \nz.mem [1975] = \nz.mem_1975_sv2v_reg ;
  assign \nz.mem [1974] = \nz.mem_1974_sv2v_reg ;
  assign \nz.mem [1973] = \nz.mem_1973_sv2v_reg ;
  assign \nz.mem [1972] = \nz.mem_1972_sv2v_reg ;
  assign \nz.mem [1971] = \nz.mem_1971_sv2v_reg ;
  assign \nz.mem [1970] = \nz.mem_1970_sv2v_reg ;
  assign \nz.mem [1969] = \nz.mem_1969_sv2v_reg ;
  assign \nz.mem [1968] = \nz.mem_1968_sv2v_reg ;
  assign \nz.mem [1967] = \nz.mem_1967_sv2v_reg ;
  assign \nz.mem [1966] = \nz.mem_1966_sv2v_reg ;
  assign \nz.mem [1965] = \nz.mem_1965_sv2v_reg ;
  assign \nz.mem [1964] = \nz.mem_1964_sv2v_reg ;
  assign \nz.mem [1963] = \nz.mem_1963_sv2v_reg ;
  assign \nz.mem [1962] = \nz.mem_1962_sv2v_reg ;
  assign \nz.mem [1961] = \nz.mem_1961_sv2v_reg ;
  assign \nz.mem [1960] = \nz.mem_1960_sv2v_reg ;
  assign \nz.mem [1959] = \nz.mem_1959_sv2v_reg ;
  assign \nz.mem [1958] = \nz.mem_1958_sv2v_reg ;
  assign \nz.mem [1957] = \nz.mem_1957_sv2v_reg ;
  assign \nz.mem [1956] = \nz.mem_1956_sv2v_reg ;
  assign \nz.mem [1955] = \nz.mem_1955_sv2v_reg ;
  assign \nz.mem [1954] = \nz.mem_1954_sv2v_reg ;
  assign \nz.mem [1953] = \nz.mem_1953_sv2v_reg ;
  assign \nz.mem [1952] = \nz.mem_1952_sv2v_reg ;
  assign \nz.mem [1951] = \nz.mem_1951_sv2v_reg ;
  assign \nz.mem [1950] = \nz.mem_1950_sv2v_reg ;
  assign \nz.mem [1949] = \nz.mem_1949_sv2v_reg ;
  assign \nz.mem [1948] = \nz.mem_1948_sv2v_reg ;
  assign \nz.mem [1947] = \nz.mem_1947_sv2v_reg ;
  assign \nz.mem [1946] = \nz.mem_1946_sv2v_reg ;
  assign \nz.mem [1945] = \nz.mem_1945_sv2v_reg ;
  assign \nz.mem [1944] = \nz.mem_1944_sv2v_reg ;
  assign \nz.mem [1943] = \nz.mem_1943_sv2v_reg ;
  assign \nz.mem [1942] = \nz.mem_1942_sv2v_reg ;
  assign \nz.mem [1941] = \nz.mem_1941_sv2v_reg ;
  assign \nz.mem [1940] = \nz.mem_1940_sv2v_reg ;
  assign \nz.mem [1939] = \nz.mem_1939_sv2v_reg ;
  assign \nz.mem [1938] = \nz.mem_1938_sv2v_reg ;
  assign \nz.mem [1937] = \nz.mem_1937_sv2v_reg ;
  assign \nz.mem [1936] = \nz.mem_1936_sv2v_reg ;
  assign \nz.mem [1935] = \nz.mem_1935_sv2v_reg ;
  assign \nz.mem [1934] = \nz.mem_1934_sv2v_reg ;
  assign \nz.mem [1933] = \nz.mem_1933_sv2v_reg ;
  assign \nz.mem [1932] = \nz.mem_1932_sv2v_reg ;
  assign \nz.mem [1931] = \nz.mem_1931_sv2v_reg ;
  assign \nz.mem [1930] = \nz.mem_1930_sv2v_reg ;
  assign \nz.mem [1929] = \nz.mem_1929_sv2v_reg ;
  assign \nz.mem [1928] = \nz.mem_1928_sv2v_reg ;
  assign \nz.mem [1927] = \nz.mem_1927_sv2v_reg ;
  assign \nz.mem [1926] = \nz.mem_1926_sv2v_reg ;
  assign \nz.mem [1925] = \nz.mem_1925_sv2v_reg ;
  assign \nz.mem [1924] = \nz.mem_1924_sv2v_reg ;
  assign \nz.mem [1923] = \nz.mem_1923_sv2v_reg ;
  assign \nz.mem [1922] = \nz.mem_1922_sv2v_reg ;
  assign \nz.mem [1921] = \nz.mem_1921_sv2v_reg ;
  assign \nz.mem [1920] = \nz.mem_1920_sv2v_reg ;
  assign \nz.mem [1919] = \nz.mem_1919_sv2v_reg ;
  assign \nz.mem [1918] = \nz.mem_1918_sv2v_reg ;
  assign \nz.mem [1917] = \nz.mem_1917_sv2v_reg ;
  assign \nz.mem [1916] = \nz.mem_1916_sv2v_reg ;
  assign \nz.mem [1915] = \nz.mem_1915_sv2v_reg ;
  assign \nz.mem [1914] = \nz.mem_1914_sv2v_reg ;
  assign \nz.mem [1913] = \nz.mem_1913_sv2v_reg ;
  assign \nz.mem [1912] = \nz.mem_1912_sv2v_reg ;
  assign \nz.mem [1911] = \nz.mem_1911_sv2v_reg ;
  assign \nz.mem [1910] = \nz.mem_1910_sv2v_reg ;
  assign \nz.mem [1909] = \nz.mem_1909_sv2v_reg ;
  assign \nz.mem [1908] = \nz.mem_1908_sv2v_reg ;
  assign \nz.mem [1907] = \nz.mem_1907_sv2v_reg ;
  assign \nz.mem [1906] = \nz.mem_1906_sv2v_reg ;
  assign \nz.mem [1905] = \nz.mem_1905_sv2v_reg ;
  assign \nz.mem [1904] = \nz.mem_1904_sv2v_reg ;
  assign \nz.mem [1903] = \nz.mem_1903_sv2v_reg ;
  assign \nz.mem [1902] = \nz.mem_1902_sv2v_reg ;
  assign \nz.mem [1901] = \nz.mem_1901_sv2v_reg ;
  assign \nz.mem [1900] = \nz.mem_1900_sv2v_reg ;
  assign \nz.mem [1899] = \nz.mem_1899_sv2v_reg ;
  assign \nz.mem [1898] = \nz.mem_1898_sv2v_reg ;
  assign \nz.mem [1897] = \nz.mem_1897_sv2v_reg ;
  assign \nz.mem [1896] = \nz.mem_1896_sv2v_reg ;
  assign \nz.mem [1895] = \nz.mem_1895_sv2v_reg ;
  assign \nz.mem [1894] = \nz.mem_1894_sv2v_reg ;
  assign \nz.mem [1893] = \nz.mem_1893_sv2v_reg ;
  assign \nz.mem [1892] = \nz.mem_1892_sv2v_reg ;
  assign \nz.mem [1891] = \nz.mem_1891_sv2v_reg ;
  assign \nz.mem [1890] = \nz.mem_1890_sv2v_reg ;
  assign \nz.mem [1889] = \nz.mem_1889_sv2v_reg ;
  assign \nz.mem [1888] = \nz.mem_1888_sv2v_reg ;
  assign \nz.mem [1887] = \nz.mem_1887_sv2v_reg ;
  assign \nz.mem [1886] = \nz.mem_1886_sv2v_reg ;
  assign \nz.mem [1885] = \nz.mem_1885_sv2v_reg ;
  assign \nz.mem [1884] = \nz.mem_1884_sv2v_reg ;
  assign \nz.mem [1883] = \nz.mem_1883_sv2v_reg ;
  assign \nz.mem [1882] = \nz.mem_1882_sv2v_reg ;
  assign \nz.mem [1881] = \nz.mem_1881_sv2v_reg ;
  assign \nz.mem [1880] = \nz.mem_1880_sv2v_reg ;
  assign \nz.mem [1879] = \nz.mem_1879_sv2v_reg ;
  assign \nz.mem [1878] = \nz.mem_1878_sv2v_reg ;
  assign \nz.mem [1877] = \nz.mem_1877_sv2v_reg ;
  assign \nz.mem [1876] = \nz.mem_1876_sv2v_reg ;
  assign \nz.mem [1875] = \nz.mem_1875_sv2v_reg ;
  assign \nz.mem [1874] = \nz.mem_1874_sv2v_reg ;
  assign \nz.mem [1873] = \nz.mem_1873_sv2v_reg ;
  assign \nz.mem [1872] = \nz.mem_1872_sv2v_reg ;
  assign \nz.mem [1871] = \nz.mem_1871_sv2v_reg ;
  assign \nz.mem [1870] = \nz.mem_1870_sv2v_reg ;
  assign \nz.mem [1869] = \nz.mem_1869_sv2v_reg ;
  assign \nz.mem [1868] = \nz.mem_1868_sv2v_reg ;
  assign \nz.mem [1867] = \nz.mem_1867_sv2v_reg ;
  assign \nz.mem [1866] = \nz.mem_1866_sv2v_reg ;
  assign \nz.mem [1865] = \nz.mem_1865_sv2v_reg ;
  assign \nz.mem [1864] = \nz.mem_1864_sv2v_reg ;
  assign \nz.mem [1863] = \nz.mem_1863_sv2v_reg ;
  assign \nz.mem [1862] = \nz.mem_1862_sv2v_reg ;
  assign \nz.mem [1861] = \nz.mem_1861_sv2v_reg ;
  assign \nz.mem [1860] = \nz.mem_1860_sv2v_reg ;
  assign \nz.mem [1859] = \nz.mem_1859_sv2v_reg ;
  assign \nz.mem [1858] = \nz.mem_1858_sv2v_reg ;
  assign \nz.mem [1857] = \nz.mem_1857_sv2v_reg ;
  assign \nz.mem [1856] = \nz.mem_1856_sv2v_reg ;
  assign \nz.mem [1855] = \nz.mem_1855_sv2v_reg ;
  assign \nz.mem [1854] = \nz.mem_1854_sv2v_reg ;
  assign \nz.mem [1853] = \nz.mem_1853_sv2v_reg ;
  assign \nz.mem [1852] = \nz.mem_1852_sv2v_reg ;
  assign \nz.mem [1851] = \nz.mem_1851_sv2v_reg ;
  assign \nz.mem [1850] = \nz.mem_1850_sv2v_reg ;
  assign \nz.mem [1849] = \nz.mem_1849_sv2v_reg ;
  assign \nz.mem [1848] = \nz.mem_1848_sv2v_reg ;
  assign \nz.mem [1847] = \nz.mem_1847_sv2v_reg ;
  assign \nz.mem [1846] = \nz.mem_1846_sv2v_reg ;
  assign \nz.mem [1845] = \nz.mem_1845_sv2v_reg ;
  assign \nz.mem [1844] = \nz.mem_1844_sv2v_reg ;
  assign \nz.mem [1843] = \nz.mem_1843_sv2v_reg ;
  assign \nz.mem [1842] = \nz.mem_1842_sv2v_reg ;
  assign \nz.mem [1841] = \nz.mem_1841_sv2v_reg ;
  assign \nz.mem [1840] = \nz.mem_1840_sv2v_reg ;
  assign \nz.mem [1839] = \nz.mem_1839_sv2v_reg ;
  assign \nz.mem [1838] = \nz.mem_1838_sv2v_reg ;
  assign \nz.mem [1837] = \nz.mem_1837_sv2v_reg ;
  assign \nz.mem [1836] = \nz.mem_1836_sv2v_reg ;
  assign \nz.mem [1835] = \nz.mem_1835_sv2v_reg ;
  assign \nz.mem [1834] = \nz.mem_1834_sv2v_reg ;
  assign \nz.mem [1833] = \nz.mem_1833_sv2v_reg ;
  assign \nz.mem [1832] = \nz.mem_1832_sv2v_reg ;
  assign \nz.mem [1831] = \nz.mem_1831_sv2v_reg ;
  assign \nz.mem [1830] = \nz.mem_1830_sv2v_reg ;
  assign \nz.mem [1829] = \nz.mem_1829_sv2v_reg ;
  assign \nz.mem [1828] = \nz.mem_1828_sv2v_reg ;
  assign \nz.mem [1827] = \nz.mem_1827_sv2v_reg ;
  assign \nz.mem [1826] = \nz.mem_1826_sv2v_reg ;
  assign \nz.mem [1825] = \nz.mem_1825_sv2v_reg ;
  assign \nz.mem [1824] = \nz.mem_1824_sv2v_reg ;
  assign \nz.mem [1823] = \nz.mem_1823_sv2v_reg ;
  assign \nz.mem [1822] = \nz.mem_1822_sv2v_reg ;
  assign \nz.mem [1821] = \nz.mem_1821_sv2v_reg ;
  assign \nz.mem [1820] = \nz.mem_1820_sv2v_reg ;
  assign \nz.mem [1819] = \nz.mem_1819_sv2v_reg ;
  assign \nz.mem [1818] = \nz.mem_1818_sv2v_reg ;
  assign \nz.mem [1817] = \nz.mem_1817_sv2v_reg ;
  assign \nz.mem [1816] = \nz.mem_1816_sv2v_reg ;
  assign \nz.mem [1815] = \nz.mem_1815_sv2v_reg ;
  assign \nz.mem [1814] = \nz.mem_1814_sv2v_reg ;
  assign \nz.mem [1813] = \nz.mem_1813_sv2v_reg ;
  assign \nz.mem [1812] = \nz.mem_1812_sv2v_reg ;
  assign \nz.mem [1811] = \nz.mem_1811_sv2v_reg ;
  assign \nz.mem [1810] = \nz.mem_1810_sv2v_reg ;
  assign \nz.mem [1809] = \nz.mem_1809_sv2v_reg ;
  assign \nz.mem [1808] = \nz.mem_1808_sv2v_reg ;
  assign \nz.mem [1807] = \nz.mem_1807_sv2v_reg ;
  assign \nz.mem [1806] = \nz.mem_1806_sv2v_reg ;
  assign \nz.mem [1805] = \nz.mem_1805_sv2v_reg ;
  assign \nz.mem [1804] = \nz.mem_1804_sv2v_reg ;
  assign \nz.mem [1803] = \nz.mem_1803_sv2v_reg ;
  assign \nz.mem [1802] = \nz.mem_1802_sv2v_reg ;
  assign \nz.mem [1801] = \nz.mem_1801_sv2v_reg ;
  assign \nz.mem [1800] = \nz.mem_1800_sv2v_reg ;
  assign \nz.mem [1799] = \nz.mem_1799_sv2v_reg ;
  assign \nz.mem [1798] = \nz.mem_1798_sv2v_reg ;
  assign \nz.mem [1797] = \nz.mem_1797_sv2v_reg ;
  assign \nz.mem [1796] = \nz.mem_1796_sv2v_reg ;
  assign \nz.mem [1795] = \nz.mem_1795_sv2v_reg ;
  assign \nz.mem [1794] = \nz.mem_1794_sv2v_reg ;
  assign \nz.mem [1793] = \nz.mem_1793_sv2v_reg ;
  assign \nz.mem [1792] = \nz.mem_1792_sv2v_reg ;
  assign \nz.mem [1791] = \nz.mem_1791_sv2v_reg ;
  assign \nz.mem [1790] = \nz.mem_1790_sv2v_reg ;
  assign \nz.mem [1789] = \nz.mem_1789_sv2v_reg ;
  assign \nz.mem [1788] = \nz.mem_1788_sv2v_reg ;
  assign \nz.mem [1787] = \nz.mem_1787_sv2v_reg ;
  assign \nz.mem [1786] = \nz.mem_1786_sv2v_reg ;
  assign \nz.mem [1785] = \nz.mem_1785_sv2v_reg ;
  assign \nz.mem [1784] = \nz.mem_1784_sv2v_reg ;
  assign \nz.mem [1783] = \nz.mem_1783_sv2v_reg ;
  assign \nz.mem [1782] = \nz.mem_1782_sv2v_reg ;
  assign \nz.mem [1781] = \nz.mem_1781_sv2v_reg ;
  assign \nz.mem [1780] = \nz.mem_1780_sv2v_reg ;
  assign \nz.mem [1779] = \nz.mem_1779_sv2v_reg ;
  assign \nz.mem [1778] = \nz.mem_1778_sv2v_reg ;
  assign \nz.mem [1777] = \nz.mem_1777_sv2v_reg ;
  assign \nz.mem [1776] = \nz.mem_1776_sv2v_reg ;
  assign \nz.mem [1775] = \nz.mem_1775_sv2v_reg ;
  assign \nz.mem [1774] = \nz.mem_1774_sv2v_reg ;
  assign \nz.mem [1773] = \nz.mem_1773_sv2v_reg ;
  assign \nz.mem [1772] = \nz.mem_1772_sv2v_reg ;
  assign \nz.mem [1771] = \nz.mem_1771_sv2v_reg ;
  assign \nz.mem [1770] = \nz.mem_1770_sv2v_reg ;
  assign \nz.mem [1769] = \nz.mem_1769_sv2v_reg ;
  assign \nz.mem [1768] = \nz.mem_1768_sv2v_reg ;
  assign \nz.mem [1767] = \nz.mem_1767_sv2v_reg ;
  assign \nz.mem [1766] = \nz.mem_1766_sv2v_reg ;
  assign \nz.mem [1765] = \nz.mem_1765_sv2v_reg ;
  assign \nz.mem [1764] = \nz.mem_1764_sv2v_reg ;
  assign \nz.mem [1763] = \nz.mem_1763_sv2v_reg ;
  assign \nz.mem [1762] = \nz.mem_1762_sv2v_reg ;
  assign \nz.mem [1761] = \nz.mem_1761_sv2v_reg ;
  assign \nz.mem [1760] = \nz.mem_1760_sv2v_reg ;
  assign \nz.mem [1759] = \nz.mem_1759_sv2v_reg ;
  assign \nz.mem [1758] = \nz.mem_1758_sv2v_reg ;
  assign \nz.mem [1757] = \nz.mem_1757_sv2v_reg ;
  assign \nz.mem [1756] = \nz.mem_1756_sv2v_reg ;
  assign \nz.mem [1755] = \nz.mem_1755_sv2v_reg ;
  assign \nz.mem [1754] = \nz.mem_1754_sv2v_reg ;
  assign \nz.mem [1753] = \nz.mem_1753_sv2v_reg ;
  assign \nz.mem [1752] = \nz.mem_1752_sv2v_reg ;
  assign \nz.mem [1751] = \nz.mem_1751_sv2v_reg ;
  assign \nz.mem [1750] = \nz.mem_1750_sv2v_reg ;
  assign \nz.mem [1749] = \nz.mem_1749_sv2v_reg ;
  assign \nz.mem [1748] = \nz.mem_1748_sv2v_reg ;
  assign \nz.mem [1747] = \nz.mem_1747_sv2v_reg ;
  assign \nz.mem [1746] = \nz.mem_1746_sv2v_reg ;
  assign \nz.mem [1745] = \nz.mem_1745_sv2v_reg ;
  assign \nz.mem [1744] = \nz.mem_1744_sv2v_reg ;
  assign \nz.mem [1743] = \nz.mem_1743_sv2v_reg ;
  assign \nz.mem [1742] = \nz.mem_1742_sv2v_reg ;
  assign \nz.mem [1741] = \nz.mem_1741_sv2v_reg ;
  assign \nz.mem [1740] = \nz.mem_1740_sv2v_reg ;
  assign \nz.mem [1739] = \nz.mem_1739_sv2v_reg ;
  assign \nz.mem [1738] = \nz.mem_1738_sv2v_reg ;
  assign \nz.mem [1737] = \nz.mem_1737_sv2v_reg ;
  assign \nz.mem [1736] = \nz.mem_1736_sv2v_reg ;
  assign \nz.mem [1735] = \nz.mem_1735_sv2v_reg ;
  assign \nz.mem [1734] = \nz.mem_1734_sv2v_reg ;
  assign \nz.mem [1733] = \nz.mem_1733_sv2v_reg ;
  assign \nz.mem [1732] = \nz.mem_1732_sv2v_reg ;
  assign \nz.mem [1731] = \nz.mem_1731_sv2v_reg ;
  assign \nz.mem [1730] = \nz.mem_1730_sv2v_reg ;
  assign \nz.mem [1729] = \nz.mem_1729_sv2v_reg ;
  assign \nz.mem [1728] = \nz.mem_1728_sv2v_reg ;
  assign \nz.mem [1727] = \nz.mem_1727_sv2v_reg ;
  assign \nz.mem [1726] = \nz.mem_1726_sv2v_reg ;
  assign \nz.mem [1725] = \nz.mem_1725_sv2v_reg ;
  assign \nz.mem [1724] = \nz.mem_1724_sv2v_reg ;
  assign \nz.mem [1723] = \nz.mem_1723_sv2v_reg ;
  assign \nz.mem [1722] = \nz.mem_1722_sv2v_reg ;
  assign \nz.mem [1721] = \nz.mem_1721_sv2v_reg ;
  assign \nz.mem [1720] = \nz.mem_1720_sv2v_reg ;
  assign \nz.mem [1719] = \nz.mem_1719_sv2v_reg ;
  assign \nz.mem [1718] = \nz.mem_1718_sv2v_reg ;
  assign \nz.mem [1717] = \nz.mem_1717_sv2v_reg ;
  assign \nz.mem [1716] = \nz.mem_1716_sv2v_reg ;
  assign \nz.mem [1715] = \nz.mem_1715_sv2v_reg ;
  assign \nz.mem [1714] = \nz.mem_1714_sv2v_reg ;
  assign \nz.mem [1713] = \nz.mem_1713_sv2v_reg ;
  assign \nz.mem [1712] = \nz.mem_1712_sv2v_reg ;
  assign \nz.mem [1711] = \nz.mem_1711_sv2v_reg ;
  assign \nz.mem [1710] = \nz.mem_1710_sv2v_reg ;
  assign \nz.mem [1709] = \nz.mem_1709_sv2v_reg ;
  assign \nz.mem [1708] = \nz.mem_1708_sv2v_reg ;
  assign \nz.mem [1707] = \nz.mem_1707_sv2v_reg ;
  assign \nz.mem [1706] = \nz.mem_1706_sv2v_reg ;
  assign \nz.mem [1705] = \nz.mem_1705_sv2v_reg ;
  assign \nz.mem [1704] = \nz.mem_1704_sv2v_reg ;
  assign \nz.mem [1703] = \nz.mem_1703_sv2v_reg ;
  assign \nz.mem [1702] = \nz.mem_1702_sv2v_reg ;
  assign \nz.mem [1701] = \nz.mem_1701_sv2v_reg ;
  assign \nz.mem [1700] = \nz.mem_1700_sv2v_reg ;
  assign \nz.mem [1699] = \nz.mem_1699_sv2v_reg ;
  assign \nz.mem [1698] = \nz.mem_1698_sv2v_reg ;
  assign \nz.mem [1697] = \nz.mem_1697_sv2v_reg ;
  assign \nz.mem [1696] = \nz.mem_1696_sv2v_reg ;
  assign \nz.mem [1695] = \nz.mem_1695_sv2v_reg ;
  assign \nz.mem [1694] = \nz.mem_1694_sv2v_reg ;
  assign \nz.mem [1693] = \nz.mem_1693_sv2v_reg ;
  assign \nz.mem [1692] = \nz.mem_1692_sv2v_reg ;
  assign \nz.mem [1691] = \nz.mem_1691_sv2v_reg ;
  assign \nz.mem [1690] = \nz.mem_1690_sv2v_reg ;
  assign \nz.mem [1689] = \nz.mem_1689_sv2v_reg ;
  assign \nz.mem [1688] = \nz.mem_1688_sv2v_reg ;
  assign \nz.mem [1687] = \nz.mem_1687_sv2v_reg ;
  assign \nz.mem [1686] = \nz.mem_1686_sv2v_reg ;
  assign \nz.mem [1685] = \nz.mem_1685_sv2v_reg ;
  assign \nz.mem [1684] = \nz.mem_1684_sv2v_reg ;
  assign \nz.mem [1683] = \nz.mem_1683_sv2v_reg ;
  assign \nz.mem [1682] = \nz.mem_1682_sv2v_reg ;
  assign \nz.mem [1681] = \nz.mem_1681_sv2v_reg ;
  assign \nz.mem [1680] = \nz.mem_1680_sv2v_reg ;
  assign \nz.mem [1679] = \nz.mem_1679_sv2v_reg ;
  assign \nz.mem [1678] = \nz.mem_1678_sv2v_reg ;
  assign \nz.mem [1677] = \nz.mem_1677_sv2v_reg ;
  assign \nz.mem [1676] = \nz.mem_1676_sv2v_reg ;
  assign \nz.mem [1675] = \nz.mem_1675_sv2v_reg ;
  assign \nz.mem [1674] = \nz.mem_1674_sv2v_reg ;
  assign \nz.mem [1673] = \nz.mem_1673_sv2v_reg ;
  assign \nz.mem [1672] = \nz.mem_1672_sv2v_reg ;
  assign \nz.mem [1671] = \nz.mem_1671_sv2v_reg ;
  assign \nz.mem [1670] = \nz.mem_1670_sv2v_reg ;
  assign \nz.mem [1669] = \nz.mem_1669_sv2v_reg ;
  assign \nz.mem [1668] = \nz.mem_1668_sv2v_reg ;
  assign \nz.mem [1667] = \nz.mem_1667_sv2v_reg ;
  assign \nz.mem [1666] = \nz.mem_1666_sv2v_reg ;
  assign \nz.mem [1665] = \nz.mem_1665_sv2v_reg ;
  assign \nz.mem [1664] = \nz.mem_1664_sv2v_reg ;
  assign \nz.mem [1663] = \nz.mem_1663_sv2v_reg ;
  assign \nz.mem [1662] = \nz.mem_1662_sv2v_reg ;
  assign \nz.mem [1661] = \nz.mem_1661_sv2v_reg ;
  assign \nz.mem [1660] = \nz.mem_1660_sv2v_reg ;
  assign \nz.mem [1659] = \nz.mem_1659_sv2v_reg ;
  assign \nz.mem [1658] = \nz.mem_1658_sv2v_reg ;
  assign \nz.mem [1657] = \nz.mem_1657_sv2v_reg ;
  assign \nz.mem [1656] = \nz.mem_1656_sv2v_reg ;
  assign \nz.mem [1655] = \nz.mem_1655_sv2v_reg ;
  assign \nz.mem [1654] = \nz.mem_1654_sv2v_reg ;
  assign \nz.mem [1653] = \nz.mem_1653_sv2v_reg ;
  assign \nz.mem [1652] = \nz.mem_1652_sv2v_reg ;
  assign \nz.mem [1651] = \nz.mem_1651_sv2v_reg ;
  assign \nz.mem [1650] = \nz.mem_1650_sv2v_reg ;
  assign \nz.mem [1649] = \nz.mem_1649_sv2v_reg ;
  assign \nz.mem [1648] = \nz.mem_1648_sv2v_reg ;
  assign \nz.mem [1647] = \nz.mem_1647_sv2v_reg ;
  assign \nz.mem [1646] = \nz.mem_1646_sv2v_reg ;
  assign \nz.mem [1645] = \nz.mem_1645_sv2v_reg ;
  assign \nz.mem [1644] = \nz.mem_1644_sv2v_reg ;
  assign \nz.mem [1643] = \nz.mem_1643_sv2v_reg ;
  assign \nz.mem [1642] = \nz.mem_1642_sv2v_reg ;
  assign \nz.mem [1641] = \nz.mem_1641_sv2v_reg ;
  assign \nz.mem [1640] = \nz.mem_1640_sv2v_reg ;
  assign \nz.mem [1639] = \nz.mem_1639_sv2v_reg ;
  assign \nz.mem [1638] = \nz.mem_1638_sv2v_reg ;
  assign \nz.mem [1637] = \nz.mem_1637_sv2v_reg ;
  assign \nz.mem [1636] = \nz.mem_1636_sv2v_reg ;
  assign \nz.mem [1635] = \nz.mem_1635_sv2v_reg ;
  assign \nz.mem [1634] = \nz.mem_1634_sv2v_reg ;
  assign \nz.mem [1633] = \nz.mem_1633_sv2v_reg ;
  assign \nz.mem [1632] = \nz.mem_1632_sv2v_reg ;
  assign \nz.mem [1631] = \nz.mem_1631_sv2v_reg ;
  assign \nz.mem [1630] = \nz.mem_1630_sv2v_reg ;
  assign \nz.mem [1629] = \nz.mem_1629_sv2v_reg ;
  assign \nz.mem [1628] = \nz.mem_1628_sv2v_reg ;
  assign \nz.mem [1627] = \nz.mem_1627_sv2v_reg ;
  assign \nz.mem [1626] = \nz.mem_1626_sv2v_reg ;
  assign \nz.mem [1625] = \nz.mem_1625_sv2v_reg ;
  assign \nz.mem [1624] = \nz.mem_1624_sv2v_reg ;
  assign \nz.mem [1623] = \nz.mem_1623_sv2v_reg ;
  assign \nz.mem [1622] = \nz.mem_1622_sv2v_reg ;
  assign \nz.mem [1621] = \nz.mem_1621_sv2v_reg ;
  assign \nz.mem [1620] = \nz.mem_1620_sv2v_reg ;
  assign \nz.mem [1619] = \nz.mem_1619_sv2v_reg ;
  assign \nz.mem [1618] = \nz.mem_1618_sv2v_reg ;
  assign \nz.mem [1617] = \nz.mem_1617_sv2v_reg ;
  assign \nz.mem [1616] = \nz.mem_1616_sv2v_reg ;
  assign \nz.mem [1615] = \nz.mem_1615_sv2v_reg ;
  assign \nz.mem [1614] = \nz.mem_1614_sv2v_reg ;
  assign \nz.mem [1613] = \nz.mem_1613_sv2v_reg ;
  assign \nz.mem [1612] = \nz.mem_1612_sv2v_reg ;
  assign \nz.mem [1611] = \nz.mem_1611_sv2v_reg ;
  assign \nz.mem [1610] = \nz.mem_1610_sv2v_reg ;
  assign \nz.mem [1609] = \nz.mem_1609_sv2v_reg ;
  assign \nz.mem [1608] = \nz.mem_1608_sv2v_reg ;
  assign \nz.mem [1607] = \nz.mem_1607_sv2v_reg ;
  assign \nz.mem [1606] = \nz.mem_1606_sv2v_reg ;
  assign \nz.mem [1605] = \nz.mem_1605_sv2v_reg ;
  assign \nz.mem [1604] = \nz.mem_1604_sv2v_reg ;
  assign \nz.mem [1603] = \nz.mem_1603_sv2v_reg ;
  assign \nz.mem [1602] = \nz.mem_1602_sv2v_reg ;
  assign \nz.mem [1601] = \nz.mem_1601_sv2v_reg ;
  assign \nz.mem [1600] = \nz.mem_1600_sv2v_reg ;
  assign \nz.mem [1599] = \nz.mem_1599_sv2v_reg ;
  assign \nz.mem [1598] = \nz.mem_1598_sv2v_reg ;
  assign \nz.mem [1597] = \nz.mem_1597_sv2v_reg ;
  assign \nz.mem [1596] = \nz.mem_1596_sv2v_reg ;
  assign \nz.mem [1595] = \nz.mem_1595_sv2v_reg ;
  assign \nz.mem [1594] = \nz.mem_1594_sv2v_reg ;
  assign \nz.mem [1593] = \nz.mem_1593_sv2v_reg ;
  assign \nz.mem [1592] = \nz.mem_1592_sv2v_reg ;
  assign \nz.mem [1591] = \nz.mem_1591_sv2v_reg ;
  assign \nz.mem [1590] = \nz.mem_1590_sv2v_reg ;
  assign \nz.mem [1589] = \nz.mem_1589_sv2v_reg ;
  assign \nz.mem [1588] = \nz.mem_1588_sv2v_reg ;
  assign \nz.mem [1587] = \nz.mem_1587_sv2v_reg ;
  assign \nz.mem [1586] = \nz.mem_1586_sv2v_reg ;
  assign \nz.mem [1585] = \nz.mem_1585_sv2v_reg ;
  assign \nz.mem [1584] = \nz.mem_1584_sv2v_reg ;
  assign \nz.mem [1583] = \nz.mem_1583_sv2v_reg ;
  assign \nz.mem [1582] = \nz.mem_1582_sv2v_reg ;
  assign \nz.mem [1581] = \nz.mem_1581_sv2v_reg ;
  assign \nz.mem [1580] = \nz.mem_1580_sv2v_reg ;
  assign \nz.mem [1579] = \nz.mem_1579_sv2v_reg ;
  assign \nz.mem [1578] = \nz.mem_1578_sv2v_reg ;
  assign \nz.mem [1577] = \nz.mem_1577_sv2v_reg ;
  assign \nz.mem [1576] = \nz.mem_1576_sv2v_reg ;
  assign \nz.mem [1575] = \nz.mem_1575_sv2v_reg ;
  assign \nz.mem [1574] = \nz.mem_1574_sv2v_reg ;
  assign \nz.mem [1573] = \nz.mem_1573_sv2v_reg ;
  assign \nz.mem [1572] = \nz.mem_1572_sv2v_reg ;
  assign \nz.mem [1571] = \nz.mem_1571_sv2v_reg ;
  assign \nz.mem [1570] = \nz.mem_1570_sv2v_reg ;
  assign \nz.mem [1569] = \nz.mem_1569_sv2v_reg ;
  assign \nz.mem [1568] = \nz.mem_1568_sv2v_reg ;
  assign \nz.mem [1567] = \nz.mem_1567_sv2v_reg ;
  assign \nz.mem [1566] = \nz.mem_1566_sv2v_reg ;
  assign \nz.mem [1565] = \nz.mem_1565_sv2v_reg ;
  assign \nz.mem [1564] = \nz.mem_1564_sv2v_reg ;
  assign \nz.mem [1563] = \nz.mem_1563_sv2v_reg ;
  assign \nz.mem [1562] = \nz.mem_1562_sv2v_reg ;
  assign \nz.mem [1561] = \nz.mem_1561_sv2v_reg ;
  assign \nz.mem [1560] = \nz.mem_1560_sv2v_reg ;
  assign \nz.mem [1559] = \nz.mem_1559_sv2v_reg ;
  assign \nz.mem [1558] = \nz.mem_1558_sv2v_reg ;
  assign \nz.mem [1557] = \nz.mem_1557_sv2v_reg ;
  assign \nz.mem [1556] = \nz.mem_1556_sv2v_reg ;
  assign \nz.mem [1555] = \nz.mem_1555_sv2v_reg ;
  assign \nz.mem [1554] = \nz.mem_1554_sv2v_reg ;
  assign \nz.mem [1553] = \nz.mem_1553_sv2v_reg ;
  assign \nz.mem [1552] = \nz.mem_1552_sv2v_reg ;
  assign \nz.mem [1551] = \nz.mem_1551_sv2v_reg ;
  assign \nz.mem [1550] = \nz.mem_1550_sv2v_reg ;
  assign \nz.mem [1549] = \nz.mem_1549_sv2v_reg ;
  assign \nz.mem [1548] = \nz.mem_1548_sv2v_reg ;
  assign \nz.mem [1547] = \nz.mem_1547_sv2v_reg ;
  assign \nz.mem [1546] = \nz.mem_1546_sv2v_reg ;
  assign \nz.mem [1545] = \nz.mem_1545_sv2v_reg ;
  assign \nz.mem [1544] = \nz.mem_1544_sv2v_reg ;
  assign \nz.mem [1543] = \nz.mem_1543_sv2v_reg ;
  assign \nz.mem [1542] = \nz.mem_1542_sv2v_reg ;
  assign \nz.mem [1541] = \nz.mem_1541_sv2v_reg ;
  assign \nz.mem [1540] = \nz.mem_1540_sv2v_reg ;
  assign \nz.mem [1539] = \nz.mem_1539_sv2v_reg ;
  assign \nz.mem [1538] = \nz.mem_1538_sv2v_reg ;
  assign \nz.mem [1537] = \nz.mem_1537_sv2v_reg ;
  assign \nz.mem [1536] = \nz.mem_1536_sv2v_reg ;
  assign \nz.mem [1535] = \nz.mem_1535_sv2v_reg ;
  assign \nz.mem [1534] = \nz.mem_1534_sv2v_reg ;
  assign \nz.mem [1533] = \nz.mem_1533_sv2v_reg ;
  assign \nz.mem [1532] = \nz.mem_1532_sv2v_reg ;
  assign \nz.mem [1531] = \nz.mem_1531_sv2v_reg ;
  assign \nz.mem [1530] = \nz.mem_1530_sv2v_reg ;
  assign \nz.mem [1529] = \nz.mem_1529_sv2v_reg ;
  assign \nz.mem [1528] = \nz.mem_1528_sv2v_reg ;
  assign \nz.mem [1527] = \nz.mem_1527_sv2v_reg ;
  assign \nz.mem [1526] = \nz.mem_1526_sv2v_reg ;
  assign \nz.mem [1525] = \nz.mem_1525_sv2v_reg ;
  assign \nz.mem [1524] = \nz.mem_1524_sv2v_reg ;
  assign \nz.mem [1523] = \nz.mem_1523_sv2v_reg ;
  assign \nz.mem [1522] = \nz.mem_1522_sv2v_reg ;
  assign \nz.mem [1521] = \nz.mem_1521_sv2v_reg ;
  assign \nz.mem [1520] = \nz.mem_1520_sv2v_reg ;
  assign \nz.mem [1519] = \nz.mem_1519_sv2v_reg ;
  assign \nz.mem [1518] = \nz.mem_1518_sv2v_reg ;
  assign \nz.mem [1517] = \nz.mem_1517_sv2v_reg ;
  assign \nz.mem [1516] = \nz.mem_1516_sv2v_reg ;
  assign \nz.mem [1515] = \nz.mem_1515_sv2v_reg ;
  assign \nz.mem [1514] = \nz.mem_1514_sv2v_reg ;
  assign \nz.mem [1513] = \nz.mem_1513_sv2v_reg ;
  assign \nz.mem [1512] = \nz.mem_1512_sv2v_reg ;
  assign \nz.mem [1511] = \nz.mem_1511_sv2v_reg ;
  assign \nz.mem [1510] = \nz.mem_1510_sv2v_reg ;
  assign \nz.mem [1509] = \nz.mem_1509_sv2v_reg ;
  assign \nz.mem [1508] = \nz.mem_1508_sv2v_reg ;
  assign \nz.mem [1507] = \nz.mem_1507_sv2v_reg ;
  assign \nz.mem [1506] = \nz.mem_1506_sv2v_reg ;
  assign \nz.mem [1505] = \nz.mem_1505_sv2v_reg ;
  assign \nz.mem [1504] = \nz.mem_1504_sv2v_reg ;
  assign \nz.mem [1503] = \nz.mem_1503_sv2v_reg ;
  assign \nz.mem [1502] = \nz.mem_1502_sv2v_reg ;
  assign \nz.mem [1501] = \nz.mem_1501_sv2v_reg ;
  assign \nz.mem [1500] = \nz.mem_1500_sv2v_reg ;
  assign \nz.mem [1499] = \nz.mem_1499_sv2v_reg ;
  assign \nz.mem [1498] = \nz.mem_1498_sv2v_reg ;
  assign \nz.mem [1497] = \nz.mem_1497_sv2v_reg ;
  assign \nz.mem [1496] = \nz.mem_1496_sv2v_reg ;
  assign \nz.mem [1495] = \nz.mem_1495_sv2v_reg ;
  assign \nz.mem [1494] = \nz.mem_1494_sv2v_reg ;
  assign \nz.mem [1493] = \nz.mem_1493_sv2v_reg ;
  assign \nz.mem [1492] = \nz.mem_1492_sv2v_reg ;
  assign \nz.mem [1491] = \nz.mem_1491_sv2v_reg ;
  assign \nz.mem [1490] = \nz.mem_1490_sv2v_reg ;
  assign \nz.mem [1489] = \nz.mem_1489_sv2v_reg ;
  assign \nz.mem [1488] = \nz.mem_1488_sv2v_reg ;
  assign \nz.mem [1487] = \nz.mem_1487_sv2v_reg ;
  assign \nz.mem [1486] = \nz.mem_1486_sv2v_reg ;
  assign \nz.mem [1485] = \nz.mem_1485_sv2v_reg ;
  assign \nz.mem [1484] = \nz.mem_1484_sv2v_reg ;
  assign \nz.mem [1483] = \nz.mem_1483_sv2v_reg ;
  assign \nz.mem [1482] = \nz.mem_1482_sv2v_reg ;
  assign \nz.mem [1481] = \nz.mem_1481_sv2v_reg ;
  assign \nz.mem [1480] = \nz.mem_1480_sv2v_reg ;
  assign \nz.mem [1479] = \nz.mem_1479_sv2v_reg ;
  assign \nz.mem [1478] = \nz.mem_1478_sv2v_reg ;
  assign \nz.mem [1477] = \nz.mem_1477_sv2v_reg ;
  assign \nz.mem [1476] = \nz.mem_1476_sv2v_reg ;
  assign \nz.mem [1475] = \nz.mem_1475_sv2v_reg ;
  assign \nz.mem [1474] = \nz.mem_1474_sv2v_reg ;
  assign \nz.mem [1473] = \nz.mem_1473_sv2v_reg ;
  assign \nz.mem [1472] = \nz.mem_1472_sv2v_reg ;
  assign \nz.mem [1471] = \nz.mem_1471_sv2v_reg ;
  assign \nz.mem [1470] = \nz.mem_1470_sv2v_reg ;
  assign \nz.mem [1469] = \nz.mem_1469_sv2v_reg ;
  assign \nz.mem [1468] = \nz.mem_1468_sv2v_reg ;
  assign \nz.mem [1467] = \nz.mem_1467_sv2v_reg ;
  assign \nz.mem [1466] = \nz.mem_1466_sv2v_reg ;
  assign \nz.mem [1465] = \nz.mem_1465_sv2v_reg ;
  assign \nz.mem [1464] = \nz.mem_1464_sv2v_reg ;
  assign \nz.mem [1463] = \nz.mem_1463_sv2v_reg ;
  assign \nz.mem [1462] = \nz.mem_1462_sv2v_reg ;
  assign \nz.mem [1461] = \nz.mem_1461_sv2v_reg ;
  assign \nz.mem [1460] = \nz.mem_1460_sv2v_reg ;
  assign \nz.mem [1459] = \nz.mem_1459_sv2v_reg ;
  assign \nz.mem [1458] = \nz.mem_1458_sv2v_reg ;
  assign \nz.mem [1457] = \nz.mem_1457_sv2v_reg ;
  assign \nz.mem [1456] = \nz.mem_1456_sv2v_reg ;
  assign \nz.mem [1455] = \nz.mem_1455_sv2v_reg ;
  assign \nz.mem [1454] = \nz.mem_1454_sv2v_reg ;
  assign \nz.mem [1453] = \nz.mem_1453_sv2v_reg ;
  assign \nz.mem [1452] = \nz.mem_1452_sv2v_reg ;
  assign \nz.mem [1451] = \nz.mem_1451_sv2v_reg ;
  assign \nz.mem [1450] = \nz.mem_1450_sv2v_reg ;
  assign \nz.mem [1449] = \nz.mem_1449_sv2v_reg ;
  assign \nz.mem [1448] = \nz.mem_1448_sv2v_reg ;
  assign \nz.mem [1447] = \nz.mem_1447_sv2v_reg ;
  assign \nz.mem [1446] = \nz.mem_1446_sv2v_reg ;
  assign \nz.mem [1445] = \nz.mem_1445_sv2v_reg ;
  assign \nz.mem [1444] = \nz.mem_1444_sv2v_reg ;
  assign \nz.mem [1443] = \nz.mem_1443_sv2v_reg ;
  assign \nz.mem [1442] = \nz.mem_1442_sv2v_reg ;
  assign \nz.mem [1441] = \nz.mem_1441_sv2v_reg ;
  assign \nz.mem [1440] = \nz.mem_1440_sv2v_reg ;
  assign \nz.mem [1439] = \nz.mem_1439_sv2v_reg ;
  assign \nz.mem [1438] = \nz.mem_1438_sv2v_reg ;
  assign \nz.mem [1437] = \nz.mem_1437_sv2v_reg ;
  assign \nz.mem [1436] = \nz.mem_1436_sv2v_reg ;
  assign \nz.mem [1435] = \nz.mem_1435_sv2v_reg ;
  assign \nz.mem [1434] = \nz.mem_1434_sv2v_reg ;
  assign \nz.mem [1433] = \nz.mem_1433_sv2v_reg ;
  assign \nz.mem [1432] = \nz.mem_1432_sv2v_reg ;
  assign \nz.mem [1431] = \nz.mem_1431_sv2v_reg ;
  assign \nz.mem [1430] = \nz.mem_1430_sv2v_reg ;
  assign \nz.mem [1429] = \nz.mem_1429_sv2v_reg ;
  assign \nz.mem [1428] = \nz.mem_1428_sv2v_reg ;
  assign \nz.mem [1427] = \nz.mem_1427_sv2v_reg ;
  assign \nz.mem [1426] = \nz.mem_1426_sv2v_reg ;
  assign \nz.mem [1425] = \nz.mem_1425_sv2v_reg ;
  assign \nz.mem [1424] = \nz.mem_1424_sv2v_reg ;
  assign \nz.mem [1423] = \nz.mem_1423_sv2v_reg ;
  assign \nz.mem [1422] = \nz.mem_1422_sv2v_reg ;
  assign \nz.mem [1421] = \nz.mem_1421_sv2v_reg ;
  assign \nz.mem [1420] = \nz.mem_1420_sv2v_reg ;
  assign \nz.mem [1419] = \nz.mem_1419_sv2v_reg ;
  assign \nz.mem [1418] = \nz.mem_1418_sv2v_reg ;
  assign \nz.mem [1417] = \nz.mem_1417_sv2v_reg ;
  assign \nz.mem [1416] = \nz.mem_1416_sv2v_reg ;
  assign \nz.mem [1415] = \nz.mem_1415_sv2v_reg ;
  assign \nz.mem [1414] = \nz.mem_1414_sv2v_reg ;
  assign \nz.mem [1413] = \nz.mem_1413_sv2v_reg ;
  assign \nz.mem [1412] = \nz.mem_1412_sv2v_reg ;
  assign \nz.mem [1411] = \nz.mem_1411_sv2v_reg ;
  assign \nz.mem [1410] = \nz.mem_1410_sv2v_reg ;
  assign \nz.mem [1409] = \nz.mem_1409_sv2v_reg ;
  assign \nz.mem [1408] = \nz.mem_1408_sv2v_reg ;
  assign \nz.mem [1407] = \nz.mem_1407_sv2v_reg ;
  assign \nz.mem [1406] = \nz.mem_1406_sv2v_reg ;
  assign \nz.mem [1405] = \nz.mem_1405_sv2v_reg ;
  assign \nz.mem [1404] = \nz.mem_1404_sv2v_reg ;
  assign \nz.mem [1403] = \nz.mem_1403_sv2v_reg ;
  assign \nz.mem [1402] = \nz.mem_1402_sv2v_reg ;
  assign \nz.mem [1401] = \nz.mem_1401_sv2v_reg ;
  assign \nz.mem [1400] = \nz.mem_1400_sv2v_reg ;
  assign \nz.mem [1399] = \nz.mem_1399_sv2v_reg ;
  assign \nz.mem [1398] = \nz.mem_1398_sv2v_reg ;
  assign \nz.mem [1397] = \nz.mem_1397_sv2v_reg ;
  assign \nz.mem [1396] = \nz.mem_1396_sv2v_reg ;
  assign \nz.mem [1395] = \nz.mem_1395_sv2v_reg ;
  assign \nz.mem [1394] = \nz.mem_1394_sv2v_reg ;
  assign \nz.mem [1393] = \nz.mem_1393_sv2v_reg ;
  assign \nz.mem [1392] = \nz.mem_1392_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[1599] = (N3)? \nz.mem [1599] : 
                          (N0)? \nz.mem [3199] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[1598] = (N3)? \nz.mem [1598] : 
                          (N0)? \nz.mem [3198] : 1'b0;
  assign r_data_o[1597] = (N3)? \nz.mem [1597] : 
                          (N0)? \nz.mem [3197] : 1'b0;
  assign r_data_o[1596] = (N3)? \nz.mem [1596] : 
                          (N0)? \nz.mem [3196] : 1'b0;
  assign r_data_o[1595] = (N3)? \nz.mem [1595] : 
                          (N0)? \nz.mem [3195] : 1'b0;
  assign r_data_o[1594] = (N3)? \nz.mem [1594] : 
                          (N0)? \nz.mem [3194] : 1'b0;
  assign r_data_o[1593] = (N3)? \nz.mem [1593] : 
                          (N0)? \nz.mem [3193] : 1'b0;
  assign r_data_o[1592] = (N3)? \nz.mem [1592] : 
                          (N0)? \nz.mem [3192] : 1'b0;
  assign r_data_o[1591] = (N3)? \nz.mem [1591] : 
                          (N0)? \nz.mem [3191] : 1'b0;
  assign r_data_o[1590] = (N3)? \nz.mem [1590] : 
                          (N0)? \nz.mem [3190] : 1'b0;
  assign r_data_o[1589] = (N3)? \nz.mem [1589] : 
                          (N0)? \nz.mem [3189] : 1'b0;
  assign r_data_o[1588] = (N3)? \nz.mem [1588] : 
                          (N0)? \nz.mem [3188] : 1'b0;
  assign r_data_o[1587] = (N3)? \nz.mem [1587] : 
                          (N0)? \nz.mem [3187] : 1'b0;
  assign r_data_o[1586] = (N3)? \nz.mem [1586] : 
                          (N0)? \nz.mem [3186] : 1'b0;
  assign r_data_o[1585] = (N3)? \nz.mem [1585] : 
                          (N0)? \nz.mem [3185] : 1'b0;
  assign r_data_o[1584] = (N3)? \nz.mem [1584] : 
                          (N0)? \nz.mem [3184] : 1'b0;
  assign r_data_o[1583] = (N3)? \nz.mem [1583] : 
                          (N0)? \nz.mem [3183] : 1'b0;
  assign r_data_o[1582] = (N3)? \nz.mem [1582] : 
                          (N0)? \nz.mem [3182] : 1'b0;
  assign r_data_o[1581] = (N3)? \nz.mem [1581] : 
                          (N0)? \nz.mem [3181] : 1'b0;
  assign r_data_o[1580] = (N3)? \nz.mem [1580] : 
                          (N0)? \nz.mem [3180] : 1'b0;
  assign r_data_o[1579] = (N3)? \nz.mem [1579] : 
                          (N0)? \nz.mem [3179] : 1'b0;
  assign r_data_o[1578] = (N3)? \nz.mem [1578] : 
                          (N0)? \nz.mem [3178] : 1'b0;
  assign r_data_o[1577] = (N3)? \nz.mem [1577] : 
                          (N0)? \nz.mem [3177] : 1'b0;
  assign r_data_o[1576] = (N3)? \nz.mem [1576] : 
                          (N0)? \nz.mem [3176] : 1'b0;
  assign r_data_o[1575] = (N3)? \nz.mem [1575] : 
                          (N0)? \nz.mem [3175] : 1'b0;
  assign r_data_o[1574] = (N3)? \nz.mem [1574] : 
                          (N0)? \nz.mem [3174] : 1'b0;
  assign r_data_o[1573] = (N3)? \nz.mem [1573] : 
                          (N0)? \nz.mem [3173] : 1'b0;
  assign r_data_o[1572] = (N3)? \nz.mem [1572] : 
                          (N0)? \nz.mem [3172] : 1'b0;
  assign r_data_o[1571] = (N3)? \nz.mem [1571] : 
                          (N0)? \nz.mem [3171] : 1'b0;
  assign r_data_o[1570] = (N3)? \nz.mem [1570] : 
                          (N0)? \nz.mem [3170] : 1'b0;
  assign r_data_o[1569] = (N3)? \nz.mem [1569] : 
                          (N0)? \nz.mem [3169] : 1'b0;
  assign r_data_o[1568] = (N3)? \nz.mem [1568] : 
                          (N0)? \nz.mem [3168] : 1'b0;
  assign r_data_o[1567] = (N3)? \nz.mem [1567] : 
                          (N0)? \nz.mem [3167] : 1'b0;
  assign r_data_o[1566] = (N3)? \nz.mem [1566] : 
                          (N0)? \nz.mem [3166] : 1'b0;
  assign r_data_o[1565] = (N3)? \nz.mem [1565] : 
                          (N0)? \nz.mem [3165] : 1'b0;
  assign r_data_o[1564] = (N3)? \nz.mem [1564] : 
                          (N0)? \nz.mem [3164] : 1'b0;
  assign r_data_o[1563] = (N3)? \nz.mem [1563] : 
                          (N0)? \nz.mem [3163] : 1'b0;
  assign r_data_o[1562] = (N3)? \nz.mem [1562] : 
                          (N0)? \nz.mem [3162] : 1'b0;
  assign r_data_o[1561] = (N3)? \nz.mem [1561] : 
                          (N0)? \nz.mem [3161] : 1'b0;
  assign r_data_o[1560] = (N3)? \nz.mem [1560] : 
                          (N0)? \nz.mem [3160] : 1'b0;
  assign r_data_o[1559] = (N3)? \nz.mem [1559] : 
                          (N0)? \nz.mem [3159] : 1'b0;
  assign r_data_o[1558] = (N3)? \nz.mem [1558] : 
                          (N0)? \nz.mem [3158] : 1'b0;
  assign r_data_o[1557] = (N3)? \nz.mem [1557] : 
                          (N0)? \nz.mem [3157] : 1'b0;
  assign r_data_o[1556] = (N3)? \nz.mem [1556] : 
                          (N0)? \nz.mem [3156] : 1'b0;
  assign r_data_o[1555] = (N3)? \nz.mem [1555] : 
                          (N0)? \nz.mem [3155] : 1'b0;
  assign r_data_o[1554] = (N3)? \nz.mem [1554] : 
                          (N0)? \nz.mem [3154] : 1'b0;
  assign r_data_o[1553] = (N3)? \nz.mem [1553] : 
                          (N0)? \nz.mem [3153] : 1'b0;
  assign r_data_o[1552] = (N3)? \nz.mem [1552] : 
                          (N0)? \nz.mem [3152] : 1'b0;
  assign r_data_o[1551] = (N3)? \nz.mem [1551] : 
                          (N0)? \nz.mem [3151] : 1'b0;
  assign r_data_o[1550] = (N3)? \nz.mem [1550] : 
                          (N0)? \nz.mem [3150] : 1'b0;
  assign r_data_o[1549] = (N3)? \nz.mem [1549] : 
                          (N0)? \nz.mem [3149] : 1'b0;
  assign r_data_o[1548] = (N3)? \nz.mem [1548] : 
                          (N0)? \nz.mem [3148] : 1'b0;
  assign r_data_o[1547] = (N3)? \nz.mem [1547] : 
                          (N0)? \nz.mem [3147] : 1'b0;
  assign r_data_o[1546] = (N3)? \nz.mem [1546] : 
                          (N0)? \nz.mem [3146] : 1'b0;
  assign r_data_o[1545] = (N3)? \nz.mem [1545] : 
                          (N0)? \nz.mem [3145] : 1'b0;
  assign r_data_o[1544] = (N3)? \nz.mem [1544] : 
                          (N0)? \nz.mem [3144] : 1'b0;
  assign r_data_o[1543] = (N3)? \nz.mem [1543] : 
                          (N0)? \nz.mem [3143] : 1'b0;
  assign r_data_o[1542] = (N3)? \nz.mem [1542] : 
                          (N0)? \nz.mem [3142] : 1'b0;
  assign r_data_o[1541] = (N3)? \nz.mem [1541] : 
                          (N0)? \nz.mem [3141] : 1'b0;
  assign r_data_o[1540] = (N3)? \nz.mem [1540] : 
                          (N0)? \nz.mem [3140] : 1'b0;
  assign r_data_o[1539] = (N3)? \nz.mem [1539] : 
                          (N0)? \nz.mem [3139] : 1'b0;
  assign r_data_o[1538] = (N3)? \nz.mem [1538] : 
                          (N0)? \nz.mem [3138] : 1'b0;
  assign r_data_o[1537] = (N3)? \nz.mem [1537] : 
                          (N0)? \nz.mem [3137] : 1'b0;
  assign r_data_o[1536] = (N3)? \nz.mem [1536] : 
                          (N0)? \nz.mem [3136] : 1'b0;
  assign r_data_o[1535] = (N3)? \nz.mem [1535] : 
                          (N0)? \nz.mem [3135] : 1'b0;
  assign r_data_o[1534] = (N3)? \nz.mem [1534] : 
                          (N0)? \nz.mem [3134] : 1'b0;
  assign r_data_o[1533] = (N3)? \nz.mem [1533] : 
                          (N0)? \nz.mem [3133] : 1'b0;
  assign r_data_o[1532] = (N3)? \nz.mem [1532] : 
                          (N0)? \nz.mem [3132] : 1'b0;
  assign r_data_o[1531] = (N3)? \nz.mem [1531] : 
                          (N0)? \nz.mem [3131] : 1'b0;
  assign r_data_o[1530] = (N3)? \nz.mem [1530] : 
                          (N0)? \nz.mem [3130] : 1'b0;
  assign r_data_o[1529] = (N3)? \nz.mem [1529] : 
                          (N0)? \nz.mem [3129] : 1'b0;
  assign r_data_o[1528] = (N3)? \nz.mem [1528] : 
                          (N0)? \nz.mem [3128] : 1'b0;
  assign r_data_o[1527] = (N3)? \nz.mem [1527] : 
                          (N0)? \nz.mem [3127] : 1'b0;
  assign r_data_o[1526] = (N3)? \nz.mem [1526] : 
                          (N0)? \nz.mem [3126] : 1'b0;
  assign r_data_o[1525] = (N3)? \nz.mem [1525] : 
                          (N0)? \nz.mem [3125] : 1'b0;
  assign r_data_o[1524] = (N3)? \nz.mem [1524] : 
                          (N0)? \nz.mem [3124] : 1'b0;
  assign r_data_o[1523] = (N3)? \nz.mem [1523] : 
                          (N0)? \nz.mem [3123] : 1'b0;
  assign r_data_o[1522] = (N3)? \nz.mem [1522] : 
                          (N0)? \nz.mem [3122] : 1'b0;
  assign r_data_o[1521] = (N3)? \nz.mem [1521] : 
                          (N0)? \nz.mem [3121] : 1'b0;
  assign r_data_o[1520] = (N3)? \nz.mem [1520] : 
                          (N0)? \nz.mem [3120] : 1'b0;
  assign r_data_o[1519] = (N3)? \nz.mem [1519] : 
                          (N0)? \nz.mem [3119] : 1'b0;
  assign r_data_o[1518] = (N3)? \nz.mem [1518] : 
                          (N0)? \nz.mem [3118] : 1'b0;
  assign r_data_o[1517] = (N3)? \nz.mem [1517] : 
                          (N0)? \nz.mem [3117] : 1'b0;
  assign r_data_o[1516] = (N3)? \nz.mem [1516] : 
                          (N0)? \nz.mem [3116] : 1'b0;
  assign r_data_o[1515] = (N3)? \nz.mem [1515] : 
                          (N0)? \nz.mem [3115] : 1'b0;
  assign r_data_o[1514] = (N3)? \nz.mem [1514] : 
                          (N0)? \nz.mem [3114] : 1'b0;
  assign r_data_o[1513] = (N3)? \nz.mem [1513] : 
                          (N0)? \nz.mem [3113] : 1'b0;
  assign r_data_o[1512] = (N3)? \nz.mem [1512] : 
                          (N0)? \nz.mem [3112] : 1'b0;
  assign r_data_o[1511] = (N3)? \nz.mem [1511] : 
                          (N0)? \nz.mem [3111] : 1'b0;
  assign r_data_o[1510] = (N3)? \nz.mem [1510] : 
                          (N0)? \nz.mem [3110] : 1'b0;
  assign r_data_o[1509] = (N3)? \nz.mem [1509] : 
                          (N0)? \nz.mem [3109] : 1'b0;
  assign r_data_o[1508] = (N3)? \nz.mem [1508] : 
                          (N0)? \nz.mem [3108] : 1'b0;
  assign r_data_o[1507] = (N3)? \nz.mem [1507] : 
                          (N0)? \nz.mem [3107] : 1'b0;
  assign r_data_o[1506] = (N3)? \nz.mem [1506] : 
                          (N0)? \nz.mem [3106] : 1'b0;
  assign r_data_o[1505] = (N3)? \nz.mem [1505] : 
                          (N0)? \nz.mem [3105] : 1'b0;
  assign r_data_o[1504] = (N3)? \nz.mem [1504] : 
                          (N0)? \nz.mem [3104] : 1'b0;
  assign r_data_o[1503] = (N3)? \nz.mem [1503] : 
                          (N0)? \nz.mem [3103] : 1'b0;
  assign r_data_o[1502] = (N3)? \nz.mem [1502] : 
                          (N0)? \nz.mem [3102] : 1'b0;
  assign r_data_o[1501] = (N3)? \nz.mem [1501] : 
                          (N0)? \nz.mem [3101] : 1'b0;
  assign r_data_o[1500] = (N3)? \nz.mem [1500] : 
                          (N0)? \nz.mem [3100] : 1'b0;
  assign r_data_o[1499] = (N3)? \nz.mem [1499] : 
                          (N0)? \nz.mem [3099] : 1'b0;
  assign r_data_o[1498] = (N3)? \nz.mem [1498] : 
                          (N0)? \nz.mem [3098] : 1'b0;
  assign r_data_o[1497] = (N3)? \nz.mem [1497] : 
                          (N0)? \nz.mem [3097] : 1'b0;
  assign r_data_o[1496] = (N3)? \nz.mem [1496] : 
                          (N0)? \nz.mem [3096] : 1'b0;
  assign r_data_o[1495] = (N3)? \nz.mem [1495] : 
                          (N0)? \nz.mem [3095] : 1'b0;
  assign r_data_o[1494] = (N3)? \nz.mem [1494] : 
                          (N0)? \nz.mem [3094] : 1'b0;
  assign r_data_o[1493] = (N3)? \nz.mem [1493] : 
                          (N0)? \nz.mem [3093] : 1'b0;
  assign r_data_o[1492] = (N3)? \nz.mem [1492] : 
                          (N0)? \nz.mem [3092] : 1'b0;
  assign r_data_o[1491] = (N3)? \nz.mem [1491] : 
                          (N0)? \nz.mem [3091] : 1'b0;
  assign r_data_o[1490] = (N3)? \nz.mem [1490] : 
                          (N0)? \nz.mem [3090] : 1'b0;
  assign r_data_o[1489] = (N3)? \nz.mem [1489] : 
                          (N0)? \nz.mem [3089] : 1'b0;
  assign r_data_o[1488] = (N3)? \nz.mem [1488] : 
                          (N0)? \nz.mem [3088] : 1'b0;
  assign r_data_o[1487] = (N3)? \nz.mem [1487] : 
                          (N0)? \nz.mem [3087] : 1'b0;
  assign r_data_o[1486] = (N3)? \nz.mem [1486] : 
                          (N0)? \nz.mem [3086] : 1'b0;
  assign r_data_o[1485] = (N3)? \nz.mem [1485] : 
                          (N0)? \nz.mem [3085] : 1'b0;
  assign r_data_o[1484] = (N3)? \nz.mem [1484] : 
                          (N0)? \nz.mem [3084] : 1'b0;
  assign r_data_o[1483] = (N3)? \nz.mem [1483] : 
                          (N0)? \nz.mem [3083] : 1'b0;
  assign r_data_o[1482] = (N3)? \nz.mem [1482] : 
                          (N0)? \nz.mem [3082] : 1'b0;
  assign r_data_o[1481] = (N3)? \nz.mem [1481] : 
                          (N0)? \nz.mem [3081] : 1'b0;
  assign r_data_o[1480] = (N3)? \nz.mem [1480] : 
                          (N0)? \nz.mem [3080] : 1'b0;
  assign r_data_o[1479] = (N3)? \nz.mem [1479] : 
                          (N0)? \nz.mem [3079] : 1'b0;
  assign r_data_o[1478] = (N3)? \nz.mem [1478] : 
                          (N0)? \nz.mem [3078] : 1'b0;
  assign r_data_o[1477] = (N3)? \nz.mem [1477] : 
                          (N0)? \nz.mem [3077] : 1'b0;
  assign r_data_o[1476] = (N3)? \nz.mem [1476] : 
                          (N0)? \nz.mem [3076] : 1'b0;
  assign r_data_o[1475] = (N3)? \nz.mem [1475] : 
                          (N0)? \nz.mem [3075] : 1'b0;
  assign r_data_o[1474] = (N3)? \nz.mem [1474] : 
                          (N0)? \nz.mem [3074] : 1'b0;
  assign r_data_o[1473] = (N3)? \nz.mem [1473] : 
                          (N0)? \nz.mem [3073] : 1'b0;
  assign r_data_o[1472] = (N3)? \nz.mem [1472] : 
                          (N0)? \nz.mem [3072] : 1'b0;
  assign r_data_o[1471] = (N3)? \nz.mem [1471] : 
                          (N0)? \nz.mem [3071] : 1'b0;
  assign r_data_o[1470] = (N3)? \nz.mem [1470] : 
                          (N0)? \nz.mem [3070] : 1'b0;
  assign r_data_o[1469] = (N3)? \nz.mem [1469] : 
                          (N0)? \nz.mem [3069] : 1'b0;
  assign r_data_o[1468] = (N3)? \nz.mem [1468] : 
                          (N0)? \nz.mem [3068] : 1'b0;
  assign r_data_o[1467] = (N3)? \nz.mem [1467] : 
                          (N0)? \nz.mem [3067] : 1'b0;
  assign r_data_o[1466] = (N3)? \nz.mem [1466] : 
                          (N0)? \nz.mem [3066] : 1'b0;
  assign r_data_o[1465] = (N3)? \nz.mem [1465] : 
                          (N0)? \nz.mem [3065] : 1'b0;
  assign r_data_o[1464] = (N3)? \nz.mem [1464] : 
                          (N0)? \nz.mem [3064] : 1'b0;
  assign r_data_o[1463] = (N3)? \nz.mem [1463] : 
                          (N0)? \nz.mem [3063] : 1'b0;
  assign r_data_o[1462] = (N3)? \nz.mem [1462] : 
                          (N0)? \nz.mem [3062] : 1'b0;
  assign r_data_o[1461] = (N3)? \nz.mem [1461] : 
                          (N0)? \nz.mem [3061] : 1'b0;
  assign r_data_o[1460] = (N3)? \nz.mem [1460] : 
                          (N0)? \nz.mem [3060] : 1'b0;
  assign r_data_o[1459] = (N3)? \nz.mem [1459] : 
                          (N0)? \nz.mem [3059] : 1'b0;
  assign r_data_o[1458] = (N3)? \nz.mem [1458] : 
                          (N0)? \nz.mem [3058] : 1'b0;
  assign r_data_o[1457] = (N3)? \nz.mem [1457] : 
                          (N0)? \nz.mem [3057] : 1'b0;
  assign r_data_o[1456] = (N3)? \nz.mem [1456] : 
                          (N0)? \nz.mem [3056] : 1'b0;
  assign r_data_o[1455] = (N3)? \nz.mem [1455] : 
                          (N0)? \nz.mem [3055] : 1'b0;
  assign r_data_o[1454] = (N3)? \nz.mem [1454] : 
                          (N0)? \nz.mem [3054] : 1'b0;
  assign r_data_o[1453] = (N3)? \nz.mem [1453] : 
                          (N0)? \nz.mem [3053] : 1'b0;
  assign r_data_o[1452] = (N3)? \nz.mem [1452] : 
                          (N0)? \nz.mem [3052] : 1'b0;
  assign r_data_o[1451] = (N3)? \nz.mem [1451] : 
                          (N0)? \nz.mem [3051] : 1'b0;
  assign r_data_o[1450] = (N3)? \nz.mem [1450] : 
                          (N0)? \nz.mem [3050] : 1'b0;
  assign r_data_o[1449] = (N3)? \nz.mem [1449] : 
                          (N0)? \nz.mem [3049] : 1'b0;
  assign r_data_o[1448] = (N3)? \nz.mem [1448] : 
                          (N0)? \nz.mem [3048] : 1'b0;
  assign r_data_o[1447] = (N3)? \nz.mem [1447] : 
                          (N0)? \nz.mem [3047] : 1'b0;
  assign r_data_o[1446] = (N3)? \nz.mem [1446] : 
                          (N0)? \nz.mem [3046] : 1'b0;
  assign r_data_o[1445] = (N3)? \nz.mem [1445] : 
                          (N0)? \nz.mem [3045] : 1'b0;
  assign r_data_o[1444] = (N3)? \nz.mem [1444] : 
                          (N0)? \nz.mem [3044] : 1'b0;
  assign r_data_o[1443] = (N3)? \nz.mem [1443] : 
                          (N0)? \nz.mem [3043] : 1'b0;
  assign r_data_o[1442] = (N3)? \nz.mem [1442] : 
                          (N0)? \nz.mem [3042] : 1'b0;
  assign r_data_o[1441] = (N3)? \nz.mem [1441] : 
                          (N0)? \nz.mem [3041] : 1'b0;
  assign r_data_o[1440] = (N3)? \nz.mem [1440] : 
                          (N0)? \nz.mem [3040] : 1'b0;
  assign r_data_o[1439] = (N3)? \nz.mem [1439] : 
                          (N0)? \nz.mem [3039] : 1'b0;
  assign r_data_o[1438] = (N3)? \nz.mem [1438] : 
                          (N0)? \nz.mem [3038] : 1'b0;
  assign r_data_o[1437] = (N3)? \nz.mem [1437] : 
                          (N0)? \nz.mem [3037] : 1'b0;
  assign r_data_o[1436] = (N3)? \nz.mem [1436] : 
                          (N0)? \nz.mem [3036] : 1'b0;
  assign r_data_o[1435] = (N3)? \nz.mem [1435] : 
                          (N0)? \nz.mem [3035] : 1'b0;
  assign r_data_o[1434] = (N3)? \nz.mem [1434] : 
                          (N0)? \nz.mem [3034] : 1'b0;
  assign r_data_o[1433] = (N3)? \nz.mem [1433] : 
                          (N0)? \nz.mem [3033] : 1'b0;
  assign r_data_o[1432] = (N3)? \nz.mem [1432] : 
                          (N0)? \nz.mem [3032] : 1'b0;
  assign r_data_o[1431] = (N3)? \nz.mem [1431] : 
                          (N0)? \nz.mem [3031] : 1'b0;
  assign r_data_o[1430] = (N3)? \nz.mem [1430] : 
                          (N0)? \nz.mem [3030] : 1'b0;
  assign r_data_o[1429] = (N3)? \nz.mem [1429] : 
                          (N0)? \nz.mem [3029] : 1'b0;
  assign r_data_o[1428] = (N3)? \nz.mem [1428] : 
                          (N0)? \nz.mem [3028] : 1'b0;
  assign r_data_o[1427] = (N3)? \nz.mem [1427] : 
                          (N0)? \nz.mem [3027] : 1'b0;
  assign r_data_o[1426] = (N3)? \nz.mem [1426] : 
                          (N0)? \nz.mem [3026] : 1'b0;
  assign r_data_o[1425] = (N3)? \nz.mem [1425] : 
                          (N0)? \nz.mem [3025] : 1'b0;
  assign r_data_o[1424] = (N3)? \nz.mem [1424] : 
                          (N0)? \nz.mem [3024] : 1'b0;
  assign r_data_o[1423] = (N3)? \nz.mem [1423] : 
                          (N0)? \nz.mem [3023] : 1'b0;
  assign r_data_o[1422] = (N3)? \nz.mem [1422] : 
                          (N0)? \nz.mem [3022] : 1'b0;
  assign r_data_o[1421] = (N3)? \nz.mem [1421] : 
                          (N0)? \nz.mem [3021] : 1'b0;
  assign r_data_o[1420] = (N3)? \nz.mem [1420] : 
                          (N0)? \nz.mem [3020] : 1'b0;
  assign r_data_o[1419] = (N3)? \nz.mem [1419] : 
                          (N0)? \nz.mem [3019] : 1'b0;
  assign r_data_o[1418] = (N3)? \nz.mem [1418] : 
                          (N0)? \nz.mem [3018] : 1'b0;
  assign r_data_o[1417] = (N3)? \nz.mem [1417] : 
                          (N0)? \nz.mem [3017] : 1'b0;
  assign r_data_o[1416] = (N3)? \nz.mem [1416] : 
                          (N0)? \nz.mem [3016] : 1'b0;
  assign r_data_o[1415] = (N3)? \nz.mem [1415] : 
                          (N0)? \nz.mem [3015] : 1'b0;
  assign r_data_o[1414] = (N3)? \nz.mem [1414] : 
                          (N0)? \nz.mem [3014] : 1'b0;
  assign r_data_o[1413] = (N3)? \nz.mem [1413] : 
                          (N0)? \nz.mem [3013] : 1'b0;
  assign r_data_o[1412] = (N3)? \nz.mem [1412] : 
                          (N0)? \nz.mem [3012] : 1'b0;
  assign r_data_o[1411] = (N3)? \nz.mem [1411] : 
                          (N0)? \nz.mem [3011] : 1'b0;
  assign r_data_o[1410] = (N3)? \nz.mem [1410] : 
                          (N0)? \nz.mem [3010] : 1'b0;
  assign r_data_o[1409] = (N3)? \nz.mem [1409] : 
                          (N0)? \nz.mem [3009] : 1'b0;
  assign r_data_o[1408] = (N3)? \nz.mem [1408] : 
                          (N0)? \nz.mem [3008] : 1'b0;
  assign r_data_o[1407] = (N3)? \nz.mem [1407] : 
                          (N0)? \nz.mem [3007] : 1'b0;
  assign r_data_o[1406] = (N3)? \nz.mem [1406] : 
                          (N0)? \nz.mem [3006] : 1'b0;
  assign r_data_o[1405] = (N3)? \nz.mem [1405] : 
                          (N0)? \nz.mem [3005] : 1'b0;
  assign r_data_o[1404] = (N3)? \nz.mem [1404] : 
                          (N0)? \nz.mem [3004] : 1'b0;
  assign r_data_o[1403] = (N3)? \nz.mem [1403] : 
                          (N0)? \nz.mem [3003] : 1'b0;
  assign r_data_o[1402] = (N3)? \nz.mem [1402] : 
                          (N0)? \nz.mem [3002] : 1'b0;
  assign r_data_o[1401] = (N3)? \nz.mem [1401] : 
                          (N0)? \nz.mem [3001] : 1'b0;
  assign r_data_o[1400] = (N3)? \nz.mem [1400] : 
                          (N0)? \nz.mem [3000] : 1'b0;
  assign r_data_o[1399] = (N3)? \nz.mem [1399] : 
                          (N0)? \nz.mem [2999] : 1'b0;
  assign r_data_o[1398] = (N3)? \nz.mem [1398] : 
                          (N0)? \nz.mem [2998] : 1'b0;
  assign r_data_o[1397] = (N3)? \nz.mem [1397] : 
                          (N0)? \nz.mem [2997] : 1'b0;
  assign r_data_o[1396] = (N3)? \nz.mem [1396] : 
                          (N0)? \nz.mem [2996] : 1'b0;
  assign r_data_o[1395] = (N3)? \nz.mem [1395] : 
                          (N0)? \nz.mem [2995] : 1'b0;
  assign r_data_o[1394] = (N3)? \nz.mem [1394] : 
                          (N0)? \nz.mem [2994] : 1'b0;
  assign r_data_o[1393] = (N3)? \nz.mem [1393] : 
                          (N0)? \nz.mem [2993] : 1'b0;
  assign r_data_o[1392] = (N3)? \nz.mem [1392] : 
                          (N0)? \nz.mem [2992] : 1'b0;
  assign r_data_o[1391] = (N3)? \nz.mem [1391] : 
                          (N0)? \nz.mem [2991] : 1'b0;
  assign r_data_o[1390] = (N3)? \nz.mem [1390] : 
                          (N0)? \nz.mem [2990] : 1'b0;
  assign r_data_o[1389] = (N3)? \nz.mem [1389] : 
                          (N0)? \nz.mem [2989] : 1'b0;
  assign r_data_o[1388] = (N3)? \nz.mem [1388] : 
                          (N0)? \nz.mem [2988] : 1'b0;
  assign r_data_o[1387] = (N3)? \nz.mem [1387] : 
                          (N0)? \nz.mem [2987] : 1'b0;
  assign r_data_o[1386] = (N3)? \nz.mem [1386] : 
                          (N0)? \nz.mem [2986] : 1'b0;
  assign r_data_o[1385] = (N3)? \nz.mem [1385] : 
                          (N0)? \nz.mem [2985] : 1'b0;
  assign r_data_o[1384] = (N3)? \nz.mem [1384] : 
                          (N0)? \nz.mem [2984] : 1'b0;
  assign r_data_o[1383] = (N3)? \nz.mem [1383] : 
                          (N0)? \nz.mem [2983] : 1'b0;
  assign r_data_o[1382] = (N3)? \nz.mem [1382] : 
                          (N0)? \nz.mem [2982] : 1'b0;
  assign r_data_o[1381] = (N3)? \nz.mem [1381] : 
                          (N0)? \nz.mem [2981] : 1'b0;
  assign r_data_o[1380] = (N3)? \nz.mem [1380] : 
                          (N0)? \nz.mem [2980] : 1'b0;
  assign r_data_o[1379] = (N3)? \nz.mem [1379] : 
                          (N0)? \nz.mem [2979] : 1'b0;
  assign r_data_o[1378] = (N3)? \nz.mem [1378] : 
                          (N0)? \nz.mem [2978] : 1'b0;
  assign r_data_o[1377] = (N3)? \nz.mem [1377] : 
                          (N0)? \nz.mem [2977] : 1'b0;
  assign r_data_o[1376] = (N3)? \nz.mem [1376] : 
                          (N0)? \nz.mem [2976] : 1'b0;
  assign r_data_o[1375] = (N3)? \nz.mem [1375] : 
                          (N0)? \nz.mem [2975] : 1'b0;
  assign r_data_o[1374] = (N3)? \nz.mem [1374] : 
                          (N0)? \nz.mem [2974] : 1'b0;
  assign r_data_o[1373] = (N3)? \nz.mem [1373] : 
                          (N0)? \nz.mem [2973] : 1'b0;
  assign r_data_o[1372] = (N3)? \nz.mem [1372] : 
                          (N0)? \nz.mem [2972] : 1'b0;
  assign r_data_o[1371] = (N3)? \nz.mem [1371] : 
                          (N0)? \nz.mem [2971] : 1'b0;
  assign r_data_o[1370] = (N3)? \nz.mem [1370] : 
                          (N0)? \nz.mem [2970] : 1'b0;
  assign r_data_o[1369] = (N3)? \nz.mem [1369] : 
                          (N0)? \nz.mem [2969] : 1'b0;
  assign r_data_o[1368] = (N3)? \nz.mem [1368] : 
                          (N0)? \nz.mem [2968] : 1'b0;
  assign r_data_o[1367] = (N3)? \nz.mem [1367] : 
                          (N0)? \nz.mem [2967] : 1'b0;
  assign r_data_o[1366] = (N3)? \nz.mem [1366] : 
                          (N0)? \nz.mem [2966] : 1'b0;
  assign r_data_o[1365] = (N3)? \nz.mem [1365] : 
                          (N0)? \nz.mem [2965] : 1'b0;
  assign r_data_o[1364] = (N3)? \nz.mem [1364] : 
                          (N0)? \nz.mem [2964] : 1'b0;
  assign r_data_o[1363] = (N3)? \nz.mem [1363] : 
                          (N0)? \nz.mem [2963] : 1'b0;
  assign r_data_o[1362] = (N3)? \nz.mem [1362] : 
                          (N0)? \nz.mem [2962] : 1'b0;
  assign r_data_o[1361] = (N3)? \nz.mem [1361] : 
                          (N0)? \nz.mem [2961] : 1'b0;
  assign r_data_o[1360] = (N3)? \nz.mem [1360] : 
                          (N0)? \nz.mem [2960] : 1'b0;
  assign r_data_o[1359] = (N3)? \nz.mem [1359] : 
                          (N0)? \nz.mem [2959] : 1'b0;
  assign r_data_o[1358] = (N3)? \nz.mem [1358] : 
                          (N0)? \nz.mem [2958] : 1'b0;
  assign r_data_o[1357] = (N3)? \nz.mem [1357] : 
                          (N0)? \nz.mem [2957] : 1'b0;
  assign r_data_o[1356] = (N3)? \nz.mem [1356] : 
                          (N0)? \nz.mem [2956] : 1'b0;
  assign r_data_o[1355] = (N3)? \nz.mem [1355] : 
                          (N0)? \nz.mem [2955] : 1'b0;
  assign r_data_o[1354] = (N3)? \nz.mem [1354] : 
                          (N0)? \nz.mem [2954] : 1'b0;
  assign r_data_o[1353] = (N3)? \nz.mem [1353] : 
                          (N0)? \nz.mem [2953] : 1'b0;
  assign r_data_o[1352] = (N3)? \nz.mem [1352] : 
                          (N0)? \nz.mem [2952] : 1'b0;
  assign r_data_o[1351] = (N3)? \nz.mem [1351] : 
                          (N0)? \nz.mem [2951] : 1'b0;
  assign r_data_o[1350] = (N3)? \nz.mem [1350] : 
                          (N0)? \nz.mem [2950] : 1'b0;
  assign r_data_o[1349] = (N3)? \nz.mem [1349] : 
                          (N0)? \nz.mem [2949] : 1'b0;
  assign r_data_o[1348] = (N3)? \nz.mem [1348] : 
                          (N0)? \nz.mem [2948] : 1'b0;
  assign r_data_o[1347] = (N3)? \nz.mem [1347] : 
                          (N0)? \nz.mem [2947] : 1'b0;
  assign r_data_o[1346] = (N3)? \nz.mem [1346] : 
                          (N0)? \nz.mem [2946] : 1'b0;
  assign r_data_o[1345] = (N3)? \nz.mem [1345] : 
                          (N0)? \nz.mem [2945] : 1'b0;
  assign r_data_o[1344] = (N3)? \nz.mem [1344] : 
                          (N0)? \nz.mem [2944] : 1'b0;
  assign r_data_o[1343] = (N3)? \nz.mem [1343] : 
                          (N0)? \nz.mem [2943] : 1'b0;
  assign r_data_o[1342] = (N3)? \nz.mem [1342] : 
                          (N0)? \nz.mem [2942] : 1'b0;
  assign r_data_o[1341] = (N3)? \nz.mem [1341] : 
                          (N0)? \nz.mem [2941] : 1'b0;
  assign r_data_o[1340] = (N3)? \nz.mem [1340] : 
                          (N0)? \nz.mem [2940] : 1'b0;
  assign r_data_o[1339] = (N3)? \nz.mem [1339] : 
                          (N0)? \nz.mem [2939] : 1'b0;
  assign r_data_o[1338] = (N3)? \nz.mem [1338] : 
                          (N0)? \nz.mem [2938] : 1'b0;
  assign r_data_o[1337] = (N3)? \nz.mem [1337] : 
                          (N0)? \nz.mem [2937] : 1'b0;
  assign r_data_o[1336] = (N3)? \nz.mem [1336] : 
                          (N0)? \nz.mem [2936] : 1'b0;
  assign r_data_o[1335] = (N3)? \nz.mem [1335] : 
                          (N0)? \nz.mem [2935] : 1'b0;
  assign r_data_o[1334] = (N3)? \nz.mem [1334] : 
                          (N0)? \nz.mem [2934] : 1'b0;
  assign r_data_o[1333] = (N3)? \nz.mem [1333] : 
                          (N0)? \nz.mem [2933] : 1'b0;
  assign r_data_o[1332] = (N3)? \nz.mem [1332] : 
                          (N0)? \nz.mem [2932] : 1'b0;
  assign r_data_o[1331] = (N3)? \nz.mem [1331] : 
                          (N0)? \nz.mem [2931] : 1'b0;
  assign r_data_o[1330] = (N3)? \nz.mem [1330] : 
                          (N0)? \nz.mem [2930] : 1'b0;
  assign r_data_o[1329] = (N3)? \nz.mem [1329] : 
                          (N0)? \nz.mem [2929] : 1'b0;
  assign r_data_o[1328] = (N3)? \nz.mem [1328] : 
                          (N0)? \nz.mem [2928] : 1'b0;
  assign r_data_o[1327] = (N3)? \nz.mem [1327] : 
                          (N0)? \nz.mem [2927] : 1'b0;
  assign r_data_o[1326] = (N3)? \nz.mem [1326] : 
                          (N0)? \nz.mem [2926] : 1'b0;
  assign r_data_o[1325] = (N3)? \nz.mem [1325] : 
                          (N0)? \nz.mem [2925] : 1'b0;
  assign r_data_o[1324] = (N3)? \nz.mem [1324] : 
                          (N0)? \nz.mem [2924] : 1'b0;
  assign r_data_o[1323] = (N3)? \nz.mem [1323] : 
                          (N0)? \nz.mem [2923] : 1'b0;
  assign r_data_o[1322] = (N3)? \nz.mem [1322] : 
                          (N0)? \nz.mem [2922] : 1'b0;
  assign r_data_o[1321] = (N3)? \nz.mem [1321] : 
                          (N0)? \nz.mem [2921] : 1'b0;
  assign r_data_o[1320] = (N3)? \nz.mem [1320] : 
                          (N0)? \nz.mem [2920] : 1'b0;
  assign r_data_o[1319] = (N3)? \nz.mem [1319] : 
                          (N0)? \nz.mem [2919] : 1'b0;
  assign r_data_o[1318] = (N3)? \nz.mem [1318] : 
                          (N0)? \nz.mem [2918] : 1'b0;
  assign r_data_o[1317] = (N3)? \nz.mem [1317] : 
                          (N0)? \nz.mem [2917] : 1'b0;
  assign r_data_o[1316] = (N3)? \nz.mem [1316] : 
                          (N0)? \nz.mem [2916] : 1'b0;
  assign r_data_o[1315] = (N3)? \nz.mem [1315] : 
                          (N0)? \nz.mem [2915] : 1'b0;
  assign r_data_o[1314] = (N3)? \nz.mem [1314] : 
                          (N0)? \nz.mem [2914] : 1'b0;
  assign r_data_o[1313] = (N3)? \nz.mem [1313] : 
                          (N0)? \nz.mem [2913] : 1'b0;
  assign r_data_o[1312] = (N3)? \nz.mem [1312] : 
                          (N0)? \nz.mem [2912] : 1'b0;
  assign r_data_o[1311] = (N3)? \nz.mem [1311] : 
                          (N0)? \nz.mem [2911] : 1'b0;
  assign r_data_o[1310] = (N3)? \nz.mem [1310] : 
                          (N0)? \nz.mem [2910] : 1'b0;
  assign r_data_o[1309] = (N3)? \nz.mem [1309] : 
                          (N0)? \nz.mem [2909] : 1'b0;
  assign r_data_o[1308] = (N3)? \nz.mem [1308] : 
                          (N0)? \nz.mem [2908] : 1'b0;
  assign r_data_o[1307] = (N3)? \nz.mem [1307] : 
                          (N0)? \nz.mem [2907] : 1'b0;
  assign r_data_o[1306] = (N3)? \nz.mem [1306] : 
                          (N0)? \nz.mem [2906] : 1'b0;
  assign r_data_o[1305] = (N3)? \nz.mem [1305] : 
                          (N0)? \nz.mem [2905] : 1'b0;
  assign r_data_o[1304] = (N3)? \nz.mem [1304] : 
                          (N0)? \nz.mem [2904] : 1'b0;
  assign r_data_o[1303] = (N3)? \nz.mem [1303] : 
                          (N0)? \nz.mem [2903] : 1'b0;
  assign r_data_o[1302] = (N3)? \nz.mem [1302] : 
                          (N0)? \nz.mem [2902] : 1'b0;
  assign r_data_o[1301] = (N3)? \nz.mem [1301] : 
                          (N0)? \nz.mem [2901] : 1'b0;
  assign r_data_o[1300] = (N3)? \nz.mem [1300] : 
                          (N0)? \nz.mem [2900] : 1'b0;
  assign r_data_o[1299] = (N3)? \nz.mem [1299] : 
                          (N0)? \nz.mem [2899] : 1'b0;
  assign r_data_o[1298] = (N3)? \nz.mem [1298] : 
                          (N0)? \nz.mem [2898] : 1'b0;
  assign r_data_o[1297] = (N3)? \nz.mem [1297] : 
                          (N0)? \nz.mem [2897] : 1'b0;
  assign r_data_o[1296] = (N3)? \nz.mem [1296] : 
                          (N0)? \nz.mem [2896] : 1'b0;
  assign r_data_o[1295] = (N3)? \nz.mem [1295] : 
                          (N0)? \nz.mem [2895] : 1'b0;
  assign r_data_o[1294] = (N3)? \nz.mem [1294] : 
                          (N0)? \nz.mem [2894] : 1'b0;
  assign r_data_o[1293] = (N3)? \nz.mem [1293] : 
                          (N0)? \nz.mem [2893] : 1'b0;
  assign r_data_o[1292] = (N3)? \nz.mem [1292] : 
                          (N0)? \nz.mem [2892] : 1'b0;
  assign r_data_o[1291] = (N3)? \nz.mem [1291] : 
                          (N0)? \nz.mem [2891] : 1'b0;
  assign r_data_o[1290] = (N3)? \nz.mem [1290] : 
                          (N0)? \nz.mem [2890] : 1'b0;
  assign r_data_o[1289] = (N3)? \nz.mem [1289] : 
                          (N0)? \nz.mem [2889] : 1'b0;
  assign r_data_o[1288] = (N3)? \nz.mem [1288] : 
                          (N0)? \nz.mem [2888] : 1'b0;
  assign r_data_o[1287] = (N3)? \nz.mem [1287] : 
                          (N0)? \nz.mem [2887] : 1'b0;
  assign r_data_o[1286] = (N3)? \nz.mem [1286] : 
                          (N0)? \nz.mem [2886] : 1'b0;
  assign r_data_o[1285] = (N3)? \nz.mem [1285] : 
                          (N0)? \nz.mem [2885] : 1'b0;
  assign r_data_o[1284] = (N3)? \nz.mem [1284] : 
                          (N0)? \nz.mem [2884] : 1'b0;
  assign r_data_o[1283] = (N3)? \nz.mem [1283] : 
                          (N0)? \nz.mem [2883] : 1'b0;
  assign r_data_o[1282] = (N3)? \nz.mem [1282] : 
                          (N0)? \nz.mem [2882] : 1'b0;
  assign r_data_o[1281] = (N3)? \nz.mem [1281] : 
                          (N0)? \nz.mem [2881] : 1'b0;
  assign r_data_o[1280] = (N3)? \nz.mem [1280] : 
                          (N0)? \nz.mem [2880] : 1'b0;
  assign r_data_o[1279] = (N3)? \nz.mem [1279] : 
                          (N0)? \nz.mem [2879] : 1'b0;
  assign r_data_o[1278] = (N3)? \nz.mem [1278] : 
                          (N0)? \nz.mem [2878] : 1'b0;
  assign r_data_o[1277] = (N3)? \nz.mem [1277] : 
                          (N0)? \nz.mem [2877] : 1'b0;
  assign r_data_o[1276] = (N3)? \nz.mem [1276] : 
                          (N0)? \nz.mem [2876] : 1'b0;
  assign r_data_o[1275] = (N3)? \nz.mem [1275] : 
                          (N0)? \nz.mem [2875] : 1'b0;
  assign r_data_o[1274] = (N3)? \nz.mem [1274] : 
                          (N0)? \nz.mem [2874] : 1'b0;
  assign r_data_o[1273] = (N3)? \nz.mem [1273] : 
                          (N0)? \nz.mem [2873] : 1'b0;
  assign r_data_o[1272] = (N3)? \nz.mem [1272] : 
                          (N0)? \nz.mem [2872] : 1'b0;
  assign r_data_o[1271] = (N3)? \nz.mem [1271] : 
                          (N0)? \nz.mem [2871] : 1'b0;
  assign r_data_o[1270] = (N3)? \nz.mem [1270] : 
                          (N0)? \nz.mem [2870] : 1'b0;
  assign r_data_o[1269] = (N3)? \nz.mem [1269] : 
                          (N0)? \nz.mem [2869] : 1'b0;
  assign r_data_o[1268] = (N3)? \nz.mem [1268] : 
                          (N0)? \nz.mem [2868] : 1'b0;
  assign r_data_o[1267] = (N3)? \nz.mem [1267] : 
                          (N0)? \nz.mem [2867] : 1'b0;
  assign r_data_o[1266] = (N3)? \nz.mem [1266] : 
                          (N0)? \nz.mem [2866] : 1'b0;
  assign r_data_o[1265] = (N3)? \nz.mem [1265] : 
                          (N0)? \nz.mem [2865] : 1'b0;
  assign r_data_o[1264] = (N3)? \nz.mem [1264] : 
                          (N0)? \nz.mem [2864] : 1'b0;
  assign r_data_o[1263] = (N3)? \nz.mem [1263] : 
                          (N0)? \nz.mem [2863] : 1'b0;
  assign r_data_o[1262] = (N3)? \nz.mem [1262] : 
                          (N0)? \nz.mem [2862] : 1'b0;
  assign r_data_o[1261] = (N3)? \nz.mem [1261] : 
                          (N0)? \nz.mem [2861] : 1'b0;
  assign r_data_o[1260] = (N3)? \nz.mem [1260] : 
                          (N0)? \nz.mem [2860] : 1'b0;
  assign r_data_o[1259] = (N3)? \nz.mem [1259] : 
                          (N0)? \nz.mem [2859] : 1'b0;
  assign r_data_o[1258] = (N3)? \nz.mem [1258] : 
                          (N0)? \nz.mem [2858] : 1'b0;
  assign r_data_o[1257] = (N3)? \nz.mem [1257] : 
                          (N0)? \nz.mem [2857] : 1'b0;
  assign r_data_o[1256] = (N3)? \nz.mem [1256] : 
                          (N0)? \nz.mem [2856] : 1'b0;
  assign r_data_o[1255] = (N3)? \nz.mem [1255] : 
                          (N0)? \nz.mem [2855] : 1'b0;
  assign r_data_o[1254] = (N3)? \nz.mem [1254] : 
                          (N0)? \nz.mem [2854] : 1'b0;
  assign r_data_o[1253] = (N3)? \nz.mem [1253] : 
                          (N0)? \nz.mem [2853] : 1'b0;
  assign r_data_o[1252] = (N3)? \nz.mem [1252] : 
                          (N0)? \nz.mem [2852] : 1'b0;
  assign r_data_o[1251] = (N3)? \nz.mem [1251] : 
                          (N0)? \nz.mem [2851] : 1'b0;
  assign r_data_o[1250] = (N3)? \nz.mem [1250] : 
                          (N0)? \nz.mem [2850] : 1'b0;
  assign r_data_o[1249] = (N3)? \nz.mem [1249] : 
                          (N0)? \nz.mem [2849] : 1'b0;
  assign r_data_o[1248] = (N3)? \nz.mem [1248] : 
                          (N0)? \nz.mem [2848] : 1'b0;
  assign r_data_o[1247] = (N3)? \nz.mem [1247] : 
                          (N0)? \nz.mem [2847] : 1'b0;
  assign r_data_o[1246] = (N3)? \nz.mem [1246] : 
                          (N0)? \nz.mem [2846] : 1'b0;
  assign r_data_o[1245] = (N3)? \nz.mem [1245] : 
                          (N0)? \nz.mem [2845] : 1'b0;
  assign r_data_o[1244] = (N3)? \nz.mem [1244] : 
                          (N0)? \nz.mem [2844] : 1'b0;
  assign r_data_o[1243] = (N3)? \nz.mem [1243] : 
                          (N0)? \nz.mem [2843] : 1'b0;
  assign r_data_o[1242] = (N3)? \nz.mem [1242] : 
                          (N0)? \nz.mem [2842] : 1'b0;
  assign r_data_o[1241] = (N3)? \nz.mem [1241] : 
                          (N0)? \nz.mem [2841] : 1'b0;
  assign r_data_o[1240] = (N3)? \nz.mem [1240] : 
                          (N0)? \nz.mem [2840] : 1'b0;
  assign r_data_o[1239] = (N3)? \nz.mem [1239] : 
                          (N0)? \nz.mem [2839] : 1'b0;
  assign r_data_o[1238] = (N3)? \nz.mem [1238] : 
                          (N0)? \nz.mem [2838] : 1'b0;
  assign r_data_o[1237] = (N3)? \nz.mem [1237] : 
                          (N0)? \nz.mem [2837] : 1'b0;
  assign r_data_o[1236] = (N3)? \nz.mem [1236] : 
                          (N0)? \nz.mem [2836] : 1'b0;
  assign r_data_o[1235] = (N3)? \nz.mem [1235] : 
                          (N0)? \nz.mem [2835] : 1'b0;
  assign r_data_o[1234] = (N3)? \nz.mem [1234] : 
                          (N0)? \nz.mem [2834] : 1'b0;
  assign r_data_o[1233] = (N3)? \nz.mem [1233] : 
                          (N0)? \nz.mem [2833] : 1'b0;
  assign r_data_o[1232] = (N3)? \nz.mem [1232] : 
                          (N0)? \nz.mem [2832] : 1'b0;
  assign r_data_o[1231] = (N3)? \nz.mem [1231] : 
                          (N0)? \nz.mem [2831] : 1'b0;
  assign r_data_o[1230] = (N3)? \nz.mem [1230] : 
                          (N0)? \nz.mem [2830] : 1'b0;
  assign r_data_o[1229] = (N3)? \nz.mem [1229] : 
                          (N0)? \nz.mem [2829] : 1'b0;
  assign r_data_o[1228] = (N3)? \nz.mem [1228] : 
                          (N0)? \nz.mem [2828] : 1'b0;
  assign r_data_o[1227] = (N3)? \nz.mem [1227] : 
                          (N0)? \nz.mem [2827] : 1'b0;
  assign r_data_o[1226] = (N3)? \nz.mem [1226] : 
                          (N0)? \nz.mem [2826] : 1'b0;
  assign r_data_o[1225] = (N3)? \nz.mem [1225] : 
                          (N0)? \nz.mem [2825] : 1'b0;
  assign r_data_o[1224] = (N3)? \nz.mem [1224] : 
                          (N0)? \nz.mem [2824] : 1'b0;
  assign r_data_o[1223] = (N3)? \nz.mem [1223] : 
                          (N0)? \nz.mem [2823] : 1'b0;
  assign r_data_o[1222] = (N3)? \nz.mem [1222] : 
                          (N0)? \nz.mem [2822] : 1'b0;
  assign r_data_o[1221] = (N3)? \nz.mem [1221] : 
                          (N0)? \nz.mem [2821] : 1'b0;
  assign r_data_o[1220] = (N3)? \nz.mem [1220] : 
                          (N0)? \nz.mem [2820] : 1'b0;
  assign r_data_o[1219] = (N3)? \nz.mem [1219] : 
                          (N0)? \nz.mem [2819] : 1'b0;
  assign r_data_o[1218] = (N3)? \nz.mem [1218] : 
                          (N0)? \nz.mem [2818] : 1'b0;
  assign r_data_o[1217] = (N3)? \nz.mem [1217] : 
                          (N0)? \nz.mem [2817] : 1'b0;
  assign r_data_o[1216] = (N3)? \nz.mem [1216] : 
                          (N0)? \nz.mem [2816] : 1'b0;
  assign r_data_o[1215] = (N3)? \nz.mem [1215] : 
                          (N0)? \nz.mem [2815] : 1'b0;
  assign r_data_o[1214] = (N3)? \nz.mem [1214] : 
                          (N0)? \nz.mem [2814] : 1'b0;
  assign r_data_o[1213] = (N3)? \nz.mem [1213] : 
                          (N0)? \nz.mem [2813] : 1'b0;
  assign r_data_o[1212] = (N3)? \nz.mem [1212] : 
                          (N0)? \nz.mem [2812] : 1'b0;
  assign r_data_o[1211] = (N3)? \nz.mem [1211] : 
                          (N0)? \nz.mem [2811] : 1'b0;
  assign r_data_o[1210] = (N3)? \nz.mem [1210] : 
                          (N0)? \nz.mem [2810] : 1'b0;
  assign r_data_o[1209] = (N3)? \nz.mem [1209] : 
                          (N0)? \nz.mem [2809] : 1'b0;
  assign r_data_o[1208] = (N3)? \nz.mem [1208] : 
                          (N0)? \nz.mem [2808] : 1'b0;
  assign r_data_o[1207] = (N3)? \nz.mem [1207] : 
                          (N0)? \nz.mem [2807] : 1'b0;
  assign r_data_o[1206] = (N3)? \nz.mem [1206] : 
                          (N0)? \nz.mem [2806] : 1'b0;
  assign r_data_o[1205] = (N3)? \nz.mem [1205] : 
                          (N0)? \nz.mem [2805] : 1'b0;
  assign r_data_o[1204] = (N3)? \nz.mem [1204] : 
                          (N0)? \nz.mem [2804] : 1'b0;
  assign r_data_o[1203] = (N3)? \nz.mem [1203] : 
                          (N0)? \nz.mem [2803] : 1'b0;
  assign r_data_o[1202] = (N3)? \nz.mem [1202] : 
                          (N0)? \nz.mem [2802] : 1'b0;
  assign r_data_o[1201] = (N3)? \nz.mem [1201] : 
                          (N0)? \nz.mem [2801] : 1'b0;
  assign r_data_o[1200] = (N3)? \nz.mem [1200] : 
                          (N0)? \nz.mem [2800] : 1'b0;
  assign r_data_o[1199] = (N3)? \nz.mem [1199] : 
                          (N0)? \nz.mem [2799] : 1'b0;
  assign r_data_o[1198] = (N3)? \nz.mem [1198] : 
                          (N0)? \nz.mem [2798] : 1'b0;
  assign r_data_o[1197] = (N3)? \nz.mem [1197] : 
                          (N0)? \nz.mem [2797] : 1'b0;
  assign r_data_o[1196] = (N3)? \nz.mem [1196] : 
                          (N0)? \nz.mem [2796] : 1'b0;
  assign r_data_o[1195] = (N3)? \nz.mem [1195] : 
                          (N0)? \nz.mem [2795] : 1'b0;
  assign r_data_o[1194] = (N3)? \nz.mem [1194] : 
                          (N0)? \nz.mem [2794] : 1'b0;
  assign r_data_o[1193] = (N3)? \nz.mem [1193] : 
                          (N0)? \nz.mem [2793] : 1'b0;
  assign r_data_o[1192] = (N3)? \nz.mem [1192] : 
                          (N0)? \nz.mem [2792] : 1'b0;
  assign r_data_o[1191] = (N3)? \nz.mem [1191] : 
                          (N0)? \nz.mem [2791] : 1'b0;
  assign r_data_o[1190] = (N3)? \nz.mem [1190] : 
                          (N0)? \nz.mem [2790] : 1'b0;
  assign r_data_o[1189] = (N3)? \nz.mem [1189] : 
                          (N0)? \nz.mem [2789] : 1'b0;
  assign r_data_o[1188] = (N3)? \nz.mem [1188] : 
                          (N0)? \nz.mem [2788] : 1'b0;
  assign r_data_o[1187] = (N3)? \nz.mem [1187] : 
                          (N0)? \nz.mem [2787] : 1'b0;
  assign r_data_o[1186] = (N3)? \nz.mem [1186] : 
                          (N0)? \nz.mem [2786] : 1'b0;
  assign r_data_o[1185] = (N3)? \nz.mem [1185] : 
                          (N0)? \nz.mem [2785] : 1'b0;
  assign r_data_o[1184] = (N3)? \nz.mem [1184] : 
                          (N0)? \nz.mem [2784] : 1'b0;
  assign r_data_o[1183] = (N3)? \nz.mem [1183] : 
                          (N0)? \nz.mem [2783] : 1'b0;
  assign r_data_o[1182] = (N3)? \nz.mem [1182] : 
                          (N0)? \nz.mem [2782] : 1'b0;
  assign r_data_o[1181] = (N3)? \nz.mem [1181] : 
                          (N0)? \nz.mem [2781] : 1'b0;
  assign r_data_o[1180] = (N3)? \nz.mem [1180] : 
                          (N0)? \nz.mem [2780] : 1'b0;
  assign r_data_o[1179] = (N3)? \nz.mem [1179] : 
                          (N0)? \nz.mem [2779] : 1'b0;
  assign r_data_o[1178] = (N3)? \nz.mem [1178] : 
                          (N0)? \nz.mem [2778] : 1'b0;
  assign r_data_o[1177] = (N3)? \nz.mem [1177] : 
                          (N0)? \nz.mem [2777] : 1'b0;
  assign r_data_o[1176] = (N3)? \nz.mem [1176] : 
                          (N0)? \nz.mem [2776] : 1'b0;
  assign r_data_o[1175] = (N3)? \nz.mem [1175] : 
                          (N0)? \nz.mem [2775] : 1'b0;
  assign r_data_o[1174] = (N3)? \nz.mem [1174] : 
                          (N0)? \nz.mem [2774] : 1'b0;
  assign r_data_o[1173] = (N3)? \nz.mem [1173] : 
                          (N0)? \nz.mem [2773] : 1'b0;
  assign r_data_o[1172] = (N3)? \nz.mem [1172] : 
                          (N0)? \nz.mem [2772] : 1'b0;
  assign r_data_o[1171] = (N3)? \nz.mem [1171] : 
                          (N0)? \nz.mem [2771] : 1'b0;
  assign r_data_o[1170] = (N3)? \nz.mem [1170] : 
                          (N0)? \nz.mem [2770] : 1'b0;
  assign r_data_o[1169] = (N3)? \nz.mem [1169] : 
                          (N0)? \nz.mem [2769] : 1'b0;
  assign r_data_o[1168] = (N3)? \nz.mem [1168] : 
                          (N0)? \nz.mem [2768] : 1'b0;
  assign r_data_o[1167] = (N3)? \nz.mem [1167] : 
                          (N0)? \nz.mem [2767] : 1'b0;
  assign r_data_o[1166] = (N3)? \nz.mem [1166] : 
                          (N0)? \nz.mem [2766] : 1'b0;
  assign r_data_o[1165] = (N3)? \nz.mem [1165] : 
                          (N0)? \nz.mem [2765] : 1'b0;
  assign r_data_o[1164] = (N3)? \nz.mem [1164] : 
                          (N0)? \nz.mem [2764] : 1'b0;
  assign r_data_o[1163] = (N3)? \nz.mem [1163] : 
                          (N0)? \nz.mem [2763] : 1'b0;
  assign r_data_o[1162] = (N3)? \nz.mem [1162] : 
                          (N0)? \nz.mem [2762] : 1'b0;
  assign r_data_o[1161] = (N3)? \nz.mem [1161] : 
                          (N0)? \nz.mem [2761] : 1'b0;
  assign r_data_o[1160] = (N3)? \nz.mem [1160] : 
                          (N0)? \nz.mem [2760] : 1'b0;
  assign r_data_o[1159] = (N3)? \nz.mem [1159] : 
                          (N0)? \nz.mem [2759] : 1'b0;
  assign r_data_o[1158] = (N3)? \nz.mem [1158] : 
                          (N0)? \nz.mem [2758] : 1'b0;
  assign r_data_o[1157] = (N3)? \nz.mem [1157] : 
                          (N0)? \nz.mem [2757] : 1'b0;
  assign r_data_o[1156] = (N3)? \nz.mem [1156] : 
                          (N0)? \nz.mem [2756] : 1'b0;
  assign r_data_o[1155] = (N3)? \nz.mem [1155] : 
                          (N0)? \nz.mem [2755] : 1'b0;
  assign r_data_o[1154] = (N3)? \nz.mem [1154] : 
                          (N0)? \nz.mem [2754] : 1'b0;
  assign r_data_o[1153] = (N3)? \nz.mem [1153] : 
                          (N0)? \nz.mem [2753] : 1'b0;
  assign r_data_o[1152] = (N3)? \nz.mem [1152] : 
                          (N0)? \nz.mem [2752] : 1'b0;
  assign r_data_o[1151] = (N3)? \nz.mem [1151] : 
                          (N0)? \nz.mem [2751] : 1'b0;
  assign r_data_o[1150] = (N3)? \nz.mem [1150] : 
                          (N0)? \nz.mem [2750] : 1'b0;
  assign r_data_o[1149] = (N3)? \nz.mem [1149] : 
                          (N0)? \nz.mem [2749] : 1'b0;
  assign r_data_o[1148] = (N3)? \nz.mem [1148] : 
                          (N0)? \nz.mem [2748] : 1'b0;
  assign r_data_o[1147] = (N3)? \nz.mem [1147] : 
                          (N0)? \nz.mem [2747] : 1'b0;
  assign r_data_o[1146] = (N3)? \nz.mem [1146] : 
                          (N0)? \nz.mem [2746] : 1'b0;
  assign r_data_o[1145] = (N3)? \nz.mem [1145] : 
                          (N0)? \nz.mem [2745] : 1'b0;
  assign r_data_o[1144] = (N3)? \nz.mem [1144] : 
                          (N0)? \nz.mem [2744] : 1'b0;
  assign r_data_o[1143] = (N3)? \nz.mem [1143] : 
                          (N0)? \nz.mem [2743] : 1'b0;
  assign r_data_o[1142] = (N3)? \nz.mem [1142] : 
                          (N0)? \nz.mem [2742] : 1'b0;
  assign r_data_o[1141] = (N3)? \nz.mem [1141] : 
                          (N0)? \nz.mem [2741] : 1'b0;
  assign r_data_o[1140] = (N3)? \nz.mem [1140] : 
                          (N0)? \nz.mem [2740] : 1'b0;
  assign r_data_o[1139] = (N3)? \nz.mem [1139] : 
                          (N0)? \nz.mem [2739] : 1'b0;
  assign r_data_o[1138] = (N3)? \nz.mem [1138] : 
                          (N0)? \nz.mem [2738] : 1'b0;
  assign r_data_o[1137] = (N3)? \nz.mem [1137] : 
                          (N0)? \nz.mem [2737] : 1'b0;
  assign r_data_o[1136] = (N3)? \nz.mem [1136] : 
                          (N0)? \nz.mem [2736] : 1'b0;
  assign r_data_o[1135] = (N3)? \nz.mem [1135] : 
                          (N0)? \nz.mem [2735] : 1'b0;
  assign r_data_o[1134] = (N3)? \nz.mem [1134] : 
                          (N0)? \nz.mem [2734] : 1'b0;
  assign r_data_o[1133] = (N3)? \nz.mem [1133] : 
                          (N0)? \nz.mem [2733] : 1'b0;
  assign r_data_o[1132] = (N3)? \nz.mem [1132] : 
                          (N0)? \nz.mem [2732] : 1'b0;
  assign r_data_o[1131] = (N3)? \nz.mem [1131] : 
                          (N0)? \nz.mem [2731] : 1'b0;
  assign r_data_o[1130] = (N3)? \nz.mem [1130] : 
                          (N0)? \nz.mem [2730] : 1'b0;
  assign r_data_o[1129] = (N3)? \nz.mem [1129] : 
                          (N0)? \nz.mem [2729] : 1'b0;
  assign r_data_o[1128] = (N3)? \nz.mem [1128] : 
                          (N0)? \nz.mem [2728] : 1'b0;
  assign r_data_o[1127] = (N3)? \nz.mem [1127] : 
                          (N0)? \nz.mem [2727] : 1'b0;
  assign r_data_o[1126] = (N3)? \nz.mem [1126] : 
                          (N0)? \nz.mem [2726] : 1'b0;
  assign r_data_o[1125] = (N3)? \nz.mem [1125] : 
                          (N0)? \nz.mem [2725] : 1'b0;
  assign r_data_o[1124] = (N3)? \nz.mem [1124] : 
                          (N0)? \nz.mem [2724] : 1'b0;
  assign r_data_o[1123] = (N3)? \nz.mem [1123] : 
                          (N0)? \nz.mem [2723] : 1'b0;
  assign r_data_o[1122] = (N3)? \nz.mem [1122] : 
                          (N0)? \nz.mem [2722] : 1'b0;
  assign r_data_o[1121] = (N3)? \nz.mem [1121] : 
                          (N0)? \nz.mem [2721] : 1'b0;
  assign r_data_o[1120] = (N3)? \nz.mem [1120] : 
                          (N0)? \nz.mem [2720] : 1'b0;
  assign r_data_o[1119] = (N3)? \nz.mem [1119] : 
                          (N0)? \nz.mem [2719] : 1'b0;
  assign r_data_o[1118] = (N3)? \nz.mem [1118] : 
                          (N0)? \nz.mem [2718] : 1'b0;
  assign r_data_o[1117] = (N3)? \nz.mem [1117] : 
                          (N0)? \nz.mem [2717] : 1'b0;
  assign r_data_o[1116] = (N3)? \nz.mem [1116] : 
                          (N0)? \nz.mem [2716] : 1'b0;
  assign r_data_o[1115] = (N3)? \nz.mem [1115] : 
                          (N0)? \nz.mem [2715] : 1'b0;
  assign r_data_o[1114] = (N3)? \nz.mem [1114] : 
                          (N0)? \nz.mem [2714] : 1'b0;
  assign r_data_o[1113] = (N3)? \nz.mem [1113] : 
                          (N0)? \nz.mem [2713] : 1'b0;
  assign r_data_o[1112] = (N3)? \nz.mem [1112] : 
                          (N0)? \nz.mem [2712] : 1'b0;
  assign r_data_o[1111] = (N3)? \nz.mem [1111] : 
                          (N0)? \nz.mem [2711] : 1'b0;
  assign r_data_o[1110] = (N3)? \nz.mem [1110] : 
                          (N0)? \nz.mem [2710] : 1'b0;
  assign r_data_o[1109] = (N3)? \nz.mem [1109] : 
                          (N0)? \nz.mem [2709] : 1'b0;
  assign r_data_o[1108] = (N3)? \nz.mem [1108] : 
                          (N0)? \nz.mem [2708] : 1'b0;
  assign r_data_o[1107] = (N3)? \nz.mem [1107] : 
                          (N0)? \nz.mem [2707] : 1'b0;
  assign r_data_o[1106] = (N3)? \nz.mem [1106] : 
                          (N0)? \nz.mem [2706] : 1'b0;
  assign r_data_o[1105] = (N3)? \nz.mem [1105] : 
                          (N0)? \nz.mem [2705] : 1'b0;
  assign r_data_o[1104] = (N3)? \nz.mem [1104] : 
                          (N0)? \nz.mem [2704] : 1'b0;
  assign r_data_o[1103] = (N3)? \nz.mem [1103] : 
                          (N0)? \nz.mem [2703] : 1'b0;
  assign r_data_o[1102] = (N3)? \nz.mem [1102] : 
                          (N0)? \nz.mem [2702] : 1'b0;
  assign r_data_o[1101] = (N3)? \nz.mem [1101] : 
                          (N0)? \nz.mem [2701] : 1'b0;
  assign r_data_o[1100] = (N3)? \nz.mem [1100] : 
                          (N0)? \nz.mem [2700] : 1'b0;
  assign r_data_o[1099] = (N3)? \nz.mem [1099] : 
                          (N0)? \nz.mem [2699] : 1'b0;
  assign r_data_o[1098] = (N3)? \nz.mem [1098] : 
                          (N0)? \nz.mem [2698] : 1'b0;
  assign r_data_o[1097] = (N3)? \nz.mem [1097] : 
                          (N0)? \nz.mem [2697] : 1'b0;
  assign r_data_o[1096] = (N3)? \nz.mem [1096] : 
                          (N0)? \nz.mem [2696] : 1'b0;
  assign r_data_o[1095] = (N3)? \nz.mem [1095] : 
                          (N0)? \nz.mem [2695] : 1'b0;
  assign r_data_o[1094] = (N3)? \nz.mem [1094] : 
                          (N0)? \nz.mem [2694] : 1'b0;
  assign r_data_o[1093] = (N3)? \nz.mem [1093] : 
                          (N0)? \nz.mem [2693] : 1'b0;
  assign r_data_o[1092] = (N3)? \nz.mem [1092] : 
                          (N0)? \nz.mem [2692] : 1'b0;
  assign r_data_o[1091] = (N3)? \nz.mem [1091] : 
                          (N0)? \nz.mem [2691] : 1'b0;
  assign r_data_o[1090] = (N3)? \nz.mem [1090] : 
                          (N0)? \nz.mem [2690] : 1'b0;
  assign r_data_o[1089] = (N3)? \nz.mem [1089] : 
                          (N0)? \nz.mem [2689] : 1'b0;
  assign r_data_o[1088] = (N3)? \nz.mem [1088] : 
                          (N0)? \nz.mem [2688] : 1'b0;
  assign r_data_o[1087] = (N3)? \nz.mem [1087] : 
                          (N0)? \nz.mem [2687] : 1'b0;
  assign r_data_o[1086] = (N3)? \nz.mem [1086] : 
                          (N0)? \nz.mem [2686] : 1'b0;
  assign r_data_o[1085] = (N3)? \nz.mem [1085] : 
                          (N0)? \nz.mem [2685] : 1'b0;
  assign r_data_o[1084] = (N3)? \nz.mem [1084] : 
                          (N0)? \nz.mem [2684] : 1'b0;
  assign r_data_o[1083] = (N3)? \nz.mem [1083] : 
                          (N0)? \nz.mem [2683] : 1'b0;
  assign r_data_o[1082] = (N3)? \nz.mem [1082] : 
                          (N0)? \nz.mem [2682] : 1'b0;
  assign r_data_o[1081] = (N3)? \nz.mem [1081] : 
                          (N0)? \nz.mem [2681] : 1'b0;
  assign r_data_o[1080] = (N3)? \nz.mem [1080] : 
                          (N0)? \nz.mem [2680] : 1'b0;
  assign r_data_o[1079] = (N3)? \nz.mem [1079] : 
                          (N0)? \nz.mem [2679] : 1'b0;
  assign r_data_o[1078] = (N3)? \nz.mem [1078] : 
                          (N0)? \nz.mem [2678] : 1'b0;
  assign r_data_o[1077] = (N3)? \nz.mem [1077] : 
                          (N0)? \nz.mem [2677] : 1'b0;
  assign r_data_o[1076] = (N3)? \nz.mem [1076] : 
                          (N0)? \nz.mem [2676] : 1'b0;
  assign r_data_o[1075] = (N3)? \nz.mem [1075] : 
                          (N0)? \nz.mem [2675] : 1'b0;
  assign r_data_o[1074] = (N3)? \nz.mem [1074] : 
                          (N0)? \nz.mem [2674] : 1'b0;
  assign r_data_o[1073] = (N3)? \nz.mem [1073] : 
                          (N0)? \nz.mem [2673] : 1'b0;
  assign r_data_o[1072] = (N3)? \nz.mem [1072] : 
                          (N0)? \nz.mem [2672] : 1'b0;
  assign r_data_o[1071] = (N3)? \nz.mem [1071] : 
                          (N0)? \nz.mem [2671] : 1'b0;
  assign r_data_o[1070] = (N3)? \nz.mem [1070] : 
                          (N0)? \nz.mem [2670] : 1'b0;
  assign r_data_o[1069] = (N3)? \nz.mem [1069] : 
                          (N0)? \nz.mem [2669] : 1'b0;
  assign r_data_o[1068] = (N3)? \nz.mem [1068] : 
                          (N0)? \nz.mem [2668] : 1'b0;
  assign r_data_o[1067] = (N3)? \nz.mem [1067] : 
                          (N0)? \nz.mem [2667] : 1'b0;
  assign r_data_o[1066] = (N3)? \nz.mem [1066] : 
                          (N0)? \nz.mem [2666] : 1'b0;
  assign r_data_o[1065] = (N3)? \nz.mem [1065] : 
                          (N0)? \nz.mem [2665] : 1'b0;
  assign r_data_o[1064] = (N3)? \nz.mem [1064] : 
                          (N0)? \nz.mem [2664] : 1'b0;
  assign r_data_o[1063] = (N3)? \nz.mem [1063] : 
                          (N0)? \nz.mem [2663] : 1'b0;
  assign r_data_o[1062] = (N3)? \nz.mem [1062] : 
                          (N0)? \nz.mem [2662] : 1'b0;
  assign r_data_o[1061] = (N3)? \nz.mem [1061] : 
                          (N0)? \nz.mem [2661] : 1'b0;
  assign r_data_o[1060] = (N3)? \nz.mem [1060] : 
                          (N0)? \nz.mem [2660] : 1'b0;
  assign r_data_o[1059] = (N3)? \nz.mem [1059] : 
                          (N0)? \nz.mem [2659] : 1'b0;
  assign r_data_o[1058] = (N3)? \nz.mem [1058] : 
                          (N0)? \nz.mem [2658] : 1'b0;
  assign r_data_o[1057] = (N3)? \nz.mem [1057] : 
                          (N0)? \nz.mem [2657] : 1'b0;
  assign r_data_o[1056] = (N3)? \nz.mem [1056] : 
                          (N0)? \nz.mem [2656] : 1'b0;
  assign r_data_o[1055] = (N3)? \nz.mem [1055] : 
                          (N0)? \nz.mem [2655] : 1'b0;
  assign r_data_o[1054] = (N3)? \nz.mem [1054] : 
                          (N0)? \nz.mem [2654] : 1'b0;
  assign r_data_o[1053] = (N3)? \nz.mem [1053] : 
                          (N0)? \nz.mem [2653] : 1'b0;
  assign r_data_o[1052] = (N3)? \nz.mem [1052] : 
                          (N0)? \nz.mem [2652] : 1'b0;
  assign r_data_o[1051] = (N3)? \nz.mem [1051] : 
                          (N0)? \nz.mem [2651] : 1'b0;
  assign r_data_o[1050] = (N3)? \nz.mem [1050] : 
                          (N0)? \nz.mem [2650] : 1'b0;
  assign r_data_o[1049] = (N3)? \nz.mem [1049] : 
                          (N0)? \nz.mem [2649] : 1'b0;
  assign r_data_o[1048] = (N3)? \nz.mem [1048] : 
                          (N0)? \nz.mem [2648] : 1'b0;
  assign r_data_o[1047] = (N3)? \nz.mem [1047] : 
                          (N0)? \nz.mem [2647] : 1'b0;
  assign r_data_o[1046] = (N3)? \nz.mem [1046] : 
                          (N0)? \nz.mem [2646] : 1'b0;
  assign r_data_o[1045] = (N3)? \nz.mem [1045] : 
                          (N0)? \nz.mem [2645] : 1'b0;
  assign r_data_o[1044] = (N3)? \nz.mem [1044] : 
                          (N0)? \nz.mem [2644] : 1'b0;
  assign r_data_o[1043] = (N3)? \nz.mem [1043] : 
                          (N0)? \nz.mem [2643] : 1'b0;
  assign r_data_o[1042] = (N3)? \nz.mem [1042] : 
                          (N0)? \nz.mem [2642] : 1'b0;
  assign r_data_o[1041] = (N3)? \nz.mem [1041] : 
                          (N0)? \nz.mem [2641] : 1'b0;
  assign r_data_o[1040] = (N3)? \nz.mem [1040] : 
                          (N0)? \nz.mem [2640] : 1'b0;
  assign r_data_o[1039] = (N3)? \nz.mem [1039] : 
                          (N0)? \nz.mem [2639] : 1'b0;
  assign r_data_o[1038] = (N3)? \nz.mem [1038] : 
                          (N0)? \nz.mem [2638] : 1'b0;
  assign r_data_o[1037] = (N3)? \nz.mem [1037] : 
                          (N0)? \nz.mem [2637] : 1'b0;
  assign r_data_o[1036] = (N3)? \nz.mem [1036] : 
                          (N0)? \nz.mem [2636] : 1'b0;
  assign r_data_o[1035] = (N3)? \nz.mem [1035] : 
                          (N0)? \nz.mem [2635] : 1'b0;
  assign r_data_o[1034] = (N3)? \nz.mem [1034] : 
                          (N0)? \nz.mem [2634] : 1'b0;
  assign r_data_o[1033] = (N3)? \nz.mem [1033] : 
                          (N0)? \nz.mem [2633] : 1'b0;
  assign r_data_o[1032] = (N3)? \nz.mem [1032] : 
                          (N0)? \nz.mem [2632] : 1'b0;
  assign r_data_o[1031] = (N3)? \nz.mem [1031] : 
                          (N0)? \nz.mem [2631] : 1'b0;
  assign r_data_o[1030] = (N3)? \nz.mem [1030] : 
                          (N0)? \nz.mem [2630] : 1'b0;
  assign r_data_o[1029] = (N3)? \nz.mem [1029] : 
                          (N0)? \nz.mem [2629] : 1'b0;
  assign r_data_o[1028] = (N3)? \nz.mem [1028] : 
                          (N0)? \nz.mem [2628] : 1'b0;
  assign r_data_o[1027] = (N3)? \nz.mem [1027] : 
                          (N0)? \nz.mem [2627] : 1'b0;
  assign r_data_o[1026] = (N3)? \nz.mem [1026] : 
                          (N0)? \nz.mem [2626] : 1'b0;
  assign r_data_o[1025] = (N3)? \nz.mem [1025] : 
                          (N0)? \nz.mem [2625] : 1'b0;
  assign r_data_o[1024] = (N3)? \nz.mem [1024] : 
                          (N0)? \nz.mem [2624] : 1'b0;
  assign r_data_o[1023] = (N3)? \nz.mem [1023] : 
                          (N0)? \nz.mem [2623] : 1'b0;
  assign r_data_o[1022] = (N3)? \nz.mem [1022] : 
                          (N0)? \nz.mem [2622] : 1'b0;
  assign r_data_o[1021] = (N3)? \nz.mem [1021] : 
                          (N0)? \nz.mem [2621] : 1'b0;
  assign r_data_o[1020] = (N3)? \nz.mem [1020] : 
                          (N0)? \nz.mem [2620] : 1'b0;
  assign r_data_o[1019] = (N3)? \nz.mem [1019] : 
                          (N0)? \nz.mem [2619] : 1'b0;
  assign r_data_o[1018] = (N3)? \nz.mem [1018] : 
                          (N0)? \nz.mem [2618] : 1'b0;
  assign r_data_o[1017] = (N3)? \nz.mem [1017] : 
                          (N0)? \nz.mem [2617] : 1'b0;
  assign r_data_o[1016] = (N3)? \nz.mem [1016] : 
                          (N0)? \nz.mem [2616] : 1'b0;
  assign r_data_o[1015] = (N3)? \nz.mem [1015] : 
                          (N0)? \nz.mem [2615] : 1'b0;
  assign r_data_o[1014] = (N3)? \nz.mem [1014] : 
                          (N0)? \nz.mem [2614] : 1'b0;
  assign r_data_o[1013] = (N3)? \nz.mem [1013] : 
                          (N0)? \nz.mem [2613] : 1'b0;
  assign r_data_o[1012] = (N3)? \nz.mem [1012] : 
                          (N0)? \nz.mem [2612] : 1'b0;
  assign r_data_o[1011] = (N3)? \nz.mem [1011] : 
                          (N0)? \nz.mem [2611] : 1'b0;
  assign r_data_o[1010] = (N3)? \nz.mem [1010] : 
                          (N0)? \nz.mem [2610] : 1'b0;
  assign r_data_o[1009] = (N3)? \nz.mem [1009] : 
                          (N0)? \nz.mem [2609] : 1'b0;
  assign r_data_o[1008] = (N3)? \nz.mem [1008] : 
                          (N0)? \nz.mem [2608] : 1'b0;
  assign r_data_o[1007] = (N3)? \nz.mem [1007] : 
                          (N0)? \nz.mem [2607] : 1'b0;
  assign r_data_o[1006] = (N3)? \nz.mem [1006] : 
                          (N0)? \nz.mem [2606] : 1'b0;
  assign r_data_o[1005] = (N3)? \nz.mem [1005] : 
                          (N0)? \nz.mem [2605] : 1'b0;
  assign r_data_o[1004] = (N3)? \nz.mem [1004] : 
                          (N0)? \nz.mem [2604] : 1'b0;
  assign r_data_o[1003] = (N3)? \nz.mem [1003] : 
                          (N0)? \nz.mem [2603] : 1'b0;
  assign r_data_o[1002] = (N3)? \nz.mem [1002] : 
                          (N0)? \nz.mem [2602] : 1'b0;
  assign r_data_o[1001] = (N3)? \nz.mem [1001] : 
                          (N0)? \nz.mem [2601] : 1'b0;
  assign r_data_o[1000] = (N3)? \nz.mem [1000] : 
                          (N0)? \nz.mem [2600] : 1'b0;
  assign r_data_o[999] = (N3)? \nz.mem [999] : 
                         (N0)? \nz.mem [2599] : 1'b0;
  assign r_data_o[998] = (N3)? \nz.mem [998] : 
                         (N0)? \nz.mem [2598] : 1'b0;
  assign r_data_o[997] = (N3)? \nz.mem [997] : 
                         (N0)? \nz.mem [2597] : 1'b0;
  assign r_data_o[996] = (N3)? \nz.mem [996] : 
                         (N0)? \nz.mem [2596] : 1'b0;
  assign r_data_o[995] = (N3)? \nz.mem [995] : 
                         (N0)? \nz.mem [2595] : 1'b0;
  assign r_data_o[994] = (N3)? \nz.mem [994] : 
                         (N0)? \nz.mem [2594] : 1'b0;
  assign r_data_o[993] = (N3)? \nz.mem [993] : 
                         (N0)? \nz.mem [2593] : 1'b0;
  assign r_data_o[992] = (N3)? \nz.mem [992] : 
                         (N0)? \nz.mem [2592] : 1'b0;
  assign r_data_o[991] = (N3)? \nz.mem [991] : 
                         (N0)? \nz.mem [2591] : 1'b0;
  assign r_data_o[990] = (N3)? \nz.mem [990] : 
                         (N0)? \nz.mem [2590] : 1'b0;
  assign r_data_o[989] = (N3)? \nz.mem [989] : 
                         (N0)? \nz.mem [2589] : 1'b0;
  assign r_data_o[988] = (N3)? \nz.mem [988] : 
                         (N0)? \nz.mem [2588] : 1'b0;
  assign r_data_o[987] = (N3)? \nz.mem [987] : 
                         (N0)? \nz.mem [2587] : 1'b0;
  assign r_data_o[986] = (N3)? \nz.mem [986] : 
                         (N0)? \nz.mem [2586] : 1'b0;
  assign r_data_o[985] = (N3)? \nz.mem [985] : 
                         (N0)? \nz.mem [2585] : 1'b0;
  assign r_data_o[984] = (N3)? \nz.mem [984] : 
                         (N0)? \nz.mem [2584] : 1'b0;
  assign r_data_o[983] = (N3)? \nz.mem [983] : 
                         (N0)? \nz.mem [2583] : 1'b0;
  assign r_data_o[982] = (N3)? \nz.mem [982] : 
                         (N0)? \nz.mem [2582] : 1'b0;
  assign r_data_o[981] = (N3)? \nz.mem [981] : 
                         (N0)? \nz.mem [2581] : 1'b0;
  assign r_data_o[980] = (N3)? \nz.mem [980] : 
                         (N0)? \nz.mem [2580] : 1'b0;
  assign r_data_o[979] = (N3)? \nz.mem [979] : 
                         (N0)? \nz.mem [2579] : 1'b0;
  assign r_data_o[978] = (N3)? \nz.mem [978] : 
                         (N0)? \nz.mem [2578] : 1'b0;
  assign r_data_o[977] = (N3)? \nz.mem [977] : 
                         (N0)? \nz.mem [2577] : 1'b0;
  assign r_data_o[976] = (N3)? \nz.mem [976] : 
                         (N0)? \nz.mem [2576] : 1'b0;
  assign r_data_o[975] = (N3)? \nz.mem [975] : 
                         (N0)? \nz.mem [2575] : 1'b0;
  assign r_data_o[974] = (N3)? \nz.mem [974] : 
                         (N0)? \nz.mem [2574] : 1'b0;
  assign r_data_o[973] = (N3)? \nz.mem [973] : 
                         (N0)? \nz.mem [2573] : 1'b0;
  assign r_data_o[972] = (N3)? \nz.mem [972] : 
                         (N0)? \nz.mem [2572] : 1'b0;
  assign r_data_o[971] = (N3)? \nz.mem [971] : 
                         (N0)? \nz.mem [2571] : 1'b0;
  assign r_data_o[970] = (N3)? \nz.mem [970] : 
                         (N0)? \nz.mem [2570] : 1'b0;
  assign r_data_o[969] = (N3)? \nz.mem [969] : 
                         (N0)? \nz.mem [2569] : 1'b0;
  assign r_data_o[968] = (N3)? \nz.mem [968] : 
                         (N0)? \nz.mem [2568] : 1'b0;
  assign r_data_o[967] = (N3)? \nz.mem [967] : 
                         (N0)? \nz.mem [2567] : 1'b0;
  assign r_data_o[966] = (N3)? \nz.mem [966] : 
                         (N0)? \nz.mem [2566] : 1'b0;
  assign r_data_o[965] = (N3)? \nz.mem [965] : 
                         (N0)? \nz.mem [2565] : 1'b0;
  assign r_data_o[964] = (N3)? \nz.mem [964] : 
                         (N0)? \nz.mem [2564] : 1'b0;
  assign r_data_o[963] = (N3)? \nz.mem [963] : 
                         (N0)? \nz.mem [2563] : 1'b0;
  assign r_data_o[962] = (N3)? \nz.mem [962] : 
                         (N0)? \nz.mem [2562] : 1'b0;
  assign r_data_o[961] = (N3)? \nz.mem [961] : 
                         (N0)? \nz.mem [2561] : 1'b0;
  assign r_data_o[960] = (N3)? \nz.mem [960] : 
                         (N0)? \nz.mem [2560] : 1'b0;
  assign r_data_o[959] = (N3)? \nz.mem [959] : 
                         (N0)? \nz.mem [2559] : 1'b0;
  assign r_data_o[958] = (N3)? \nz.mem [958] : 
                         (N0)? \nz.mem [2558] : 1'b0;
  assign r_data_o[957] = (N3)? \nz.mem [957] : 
                         (N0)? \nz.mem [2557] : 1'b0;
  assign r_data_o[956] = (N3)? \nz.mem [956] : 
                         (N0)? \nz.mem [2556] : 1'b0;
  assign r_data_o[955] = (N3)? \nz.mem [955] : 
                         (N0)? \nz.mem [2555] : 1'b0;
  assign r_data_o[954] = (N3)? \nz.mem [954] : 
                         (N0)? \nz.mem [2554] : 1'b0;
  assign r_data_o[953] = (N3)? \nz.mem [953] : 
                         (N0)? \nz.mem [2553] : 1'b0;
  assign r_data_o[952] = (N3)? \nz.mem [952] : 
                         (N0)? \nz.mem [2552] : 1'b0;
  assign r_data_o[951] = (N3)? \nz.mem [951] : 
                         (N0)? \nz.mem [2551] : 1'b0;
  assign r_data_o[950] = (N3)? \nz.mem [950] : 
                         (N0)? \nz.mem [2550] : 1'b0;
  assign r_data_o[949] = (N3)? \nz.mem [949] : 
                         (N0)? \nz.mem [2549] : 1'b0;
  assign r_data_o[948] = (N3)? \nz.mem [948] : 
                         (N0)? \nz.mem [2548] : 1'b0;
  assign r_data_o[947] = (N3)? \nz.mem [947] : 
                         (N0)? \nz.mem [2547] : 1'b0;
  assign r_data_o[946] = (N3)? \nz.mem [946] : 
                         (N0)? \nz.mem [2546] : 1'b0;
  assign r_data_o[945] = (N3)? \nz.mem [945] : 
                         (N0)? \nz.mem [2545] : 1'b0;
  assign r_data_o[944] = (N3)? \nz.mem [944] : 
                         (N0)? \nz.mem [2544] : 1'b0;
  assign r_data_o[943] = (N3)? \nz.mem [943] : 
                         (N0)? \nz.mem [2543] : 1'b0;
  assign r_data_o[942] = (N3)? \nz.mem [942] : 
                         (N0)? \nz.mem [2542] : 1'b0;
  assign r_data_o[941] = (N3)? \nz.mem [941] : 
                         (N0)? \nz.mem [2541] : 1'b0;
  assign r_data_o[940] = (N3)? \nz.mem [940] : 
                         (N0)? \nz.mem [2540] : 1'b0;
  assign r_data_o[939] = (N3)? \nz.mem [939] : 
                         (N0)? \nz.mem [2539] : 1'b0;
  assign r_data_o[938] = (N3)? \nz.mem [938] : 
                         (N0)? \nz.mem [2538] : 1'b0;
  assign r_data_o[937] = (N3)? \nz.mem [937] : 
                         (N0)? \nz.mem [2537] : 1'b0;
  assign r_data_o[936] = (N3)? \nz.mem [936] : 
                         (N0)? \nz.mem [2536] : 1'b0;
  assign r_data_o[935] = (N3)? \nz.mem [935] : 
                         (N0)? \nz.mem [2535] : 1'b0;
  assign r_data_o[934] = (N3)? \nz.mem [934] : 
                         (N0)? \nz.mem [2534] : 1'b0;
  assign r_data_o[933] = (N3)? \nz.mem [933] : 
                         (N0)? \nz.mem [2533] : 1'b0;
  assign r_data_o[932] = (N3)? \nz.mem [932] : 
                         (N0)? \nz.mem [2532] : 1'b0;
  assign r_data_o[931] = (N3)? \nz.mem [931] : 
                         (N0)? \nz.mem [2531] : 1'b0;
  assign r_data_o[930] = (N3)? \nz.mem [930] : 
                         (N0)? \nz.mem [2530] : 1'b0;
  assign r_data_o[929] = (N3)? \nz.mem [929] : 
                         (N0)? \nz.mem [2529] : 1'b0;
  assign r_data_o[928] = (N3)? \nz.mem [928] : 
                         (N0)? \nz.mem [2528] : 1'b0;
  assign r_data_o[927] = (N3)? \nz.mem [927] : 
                         (N0)? \nz.mem [2527] : 1'b0;
  assign r_data_o[926] = (N3)? \nz.mem [926] : 
                         (N0)? \nz.mem [2526] : 1'b0;
  assign r_data_o[925] = (N3)? \nz.mem [925] : 
                         (N0)? \nz.mem [2525] : 1'b0;
  assign r_data_o[924] = (N3)? \nz.mem [924] : 
                         (N0)? \nz.mem [2524] : 1'b0;
  assign r_data_o[923] = (N3)? \nz.mem [923] : 
                         (N0)? \nz.mem [2523] : 1'b0;
  assign r_data_o[922] = (N3)? \nz.mem [922] : 
                         (N0)? \nz.mem [2522] : 1'b0;
  assign r_data_o[921] = (N3)? \nz.mem [921] : 
                         (N0)? \nz.mem [2521] : 1'b0;
  assign r_data_o[920] = (N3)? \nz.mem [920] : 
                         (N0)? \nz.mem [2520] : 1'b0;
  assign r_data_o[919] = (N3)? \nz.mem [919] : 
                         (N0)? \nz.mem [2519] : 1'b0;
  assign r_data_o[918] = (N3)? \nz.mem [918] : 
                         (N0)? \nz.mem [2518] : 1'b0;
  assign r_data_o[917] = (N3)? \nz.mem [917] : 
                         (N0)? \nz.mem [2517] : 1'b0;
  assign r_data_o[916] = (N3)? \nz.mem [916] : 
                         (N0)? \nz.mem [2516] : 1'b0;
  assign r_data_o[915] = (N3)? \nz.mem [915] : 
                         (N0)? \nz.mem [2515] : 1'b0;
  assign r_data_o[914] = (N3)? \nz.mem [914] : 
                         (N0)? \nz.mem [2514] : 1'b0;
  assign r_data_o[913] = (N3)? \nz.mem [913] : 
                         (N0)? \nz.mem [2513] : 1'b0;
  assign r_data_o[912] = (N3)? \nz.mem [912] : 
                         (N0)? \nz.mem [2512] : 1'b0;
  assign r_data_o[911] = (N3)? \nz.mem [911] : 
                         (N0)? \nz.mem [2511] : 1'b0;
  assign r_data_o[910] = (N3)? \nz.mem [910] : 
                         (N0)? \nz.mem [2510] : 1'b0;
  assign r_data_o[909] = (N3)? \nz.mem [909] : 
                         (N0)? \nz.mem [2509] : 1'b0;
  assign r_data_o[908] = (N3)? \nz.mem [908] : 
                         (N0)? \nz.mem [2508] : 1'b0;
  assign r_data_o[907] = (N3)? \nz.mem [907] : 
                         (N0)? \nz.mem [2507] : 1'b0;
  assign r_data_o[906] = (N3)? \nz.mem [906] : 
                         (N0)? \nz.mem [2506] : 1'b0;
  assign r_data_o[905] = (N3)? \nz.mem [905] : 
                         (N0)? \nz.mem [2505] : 1'b0;
  assign r_data_o[904] = (N3)? \nz.mem [904] : 
                         (N0)? \nz.mem [2504] : 1'b0;
  assign r_data_o[903] = (N3)? \nz.mem [903] : 
                         (N0)? \nz.mem [2503] : 1'b0;
  assign r_data_o[902] = (N3)? \nz.mem [902] : 
                         (N0)? \nz.mem [2502] : 1'b0;
  assign r_data_o[901] = (N3)? \nz.mem [901] : 
                         (N0)? \nz.mem [2501] : 1'b0;
  assign r_data_o[900] = (N3)? \nz.mem [900] : 
                         (N0)? \nz.mem [2500] : 1'b0;
  assign r_data_o[899] = (N3)? \nz.mem [899] : 
                         (N0)? \nz.mem [2499] : 1'b0;
  assign r_data_o[898] = (N3)? \nz.mem [898] : 
                         (N0)? \nz.mem [2498] : 1'b0;
  assign r_data_o[897] = (N3)? \nz.mem [897] : 
                         (N0)? \nz.mem [2497] : 1'b0;
  assign r_data_o[896] = (N3)? \nz.mem [896] : 
                         (N0)? \nz.mem [2496] : 1'b0;
  assign r_data_o[895] = (N3)? \nz.mem [895] : 
                         (N0)? \nz.mem [2495] : 1'b0;
  assign r_data_o[894] = (N3)? \nz.mem [894] : 
                         (N0)? \nz.mem [2494] : 1'b0;
  assign r_data_o[893] = (N3)? \nz.mem [893] : 
                         (N0)? \nz.mem [2493] : 1'b0;
  assign r_data_o[892] = (N3)? \nz.mem [892] : 
                         (N0)? \nz.mem [2492] : 1'b0;
  assign r_data_o[891] = (N3)? \nz.mem [891] : 
                         (N0)? \nz.mem [2491] : 1'b0;
  assign r_data_o[890] = (N3)? \nz.mem [890] : 
                         (N0)? \nz.mem [2490] : 1'b0;
  assign r_data_o[889] = (N3)? \nz.mem [889] : 
                         (N0)? \nz.mem [2489] : 1'b0;
  assign r_data_o[888] = (N3)? \nz.mem [888] : 
                         (N0)? \nz.mem [2488] : 1'b0;
  assign r_data_o[887] = (N3)? \nz.mem [887] : 
                         (N0)? \nz.mem [2487] : 1'b0;
  assign r_data_o[886] = (N3)? \nz.mem [886] : 
                         (N0)? \nz.mem [2486] : 1'b0;
  assign r_data_o[885] = (N3)? \nz.mem [885] : 
                         (N0)? \nz.mem [2485] : 1'b0;
  assign r_data_o[884] = (N3)? \nz.mem [884] : 
                         (N0)? \nz.mem [2484] : 1'b0;
  assign r_data_o[883] = (N3)? \nz.mem [883] : 
                         (N0)? \nz.mem [2483] : 1'b0;
  assign r_data_o[882] = (N3)? \nz.mem [882] : 
                         (N0)? \nz.mem [2482] : 1'b0;
  assign r_data_o[881] = (N3)? \nz.mem [881] : 
                         (N0)? \nz.mem [2481] : 1'b0;
  assign r_data_o[880] = (N3)? \nz.mem [880] : 
                         (N0)? \nz.mem [2480] : 1'b0;
  assign r_data_o[879] = (N3)? \nz.mem [879] : 
                         (N0)? \nz.mem [2479] : 1'b0;
  assign r_data_o[878] = (N3)? \nz.mem [878] : 
                         (N0)? \nz.mem [2478] : 1'b0;
  assign r_data_o[877] = (N3)? \nz.mem [877] : 
                         (N0)? \nz.mem [2477] : 1'b0;
  assign r_data_o[876] = (N3)? \nz.mem [876] : 
                         (N0)? \nz.mem [2476] : 1'b0;
  assign r_data_o[875] = (N3)? \nz.mem [875] : 
                         (N0)? \nz.mem [2475] : 1'b0;
  assign r_data_o[874] = (N3)? \nz.mem [874] : 
                         (N0)? \nz.mem [2474] : 1'b0;
  assign r_data_o[873] = (N3)? \nz.mem [873] : 
                         (N0)? \nz.mem [2473] : 1'b0;
  assign r_data_o[872] = (N3)? \nz.mem [872] : 
                         (N0)? \nz.mem [2472] : 1'b0;
  assign r_data_o[871] = (N3)? \nz.mem [871] : 
                         (N0)? \nz.mem [2471] : 1'b0;
  assign r_data_o[870] = (N3)? \nz.mem [870] : 
                         (N0)? \nz.mem [2470] : 1'b0;
  assign r_data_o[869] = (N3)? \nz.mem [869] : 
                         (N0)? \nz.mem [2469] : 1'b0;
  assign r_data_o[868] = (N3)? \nz.mem [868] : 
                         (N0)? \nz.mem [2468] : 1'b0;
  assign r_data_o[867] = (N3)? \nz.mem [867] : 
                         (N0)? \nz.mem [2467] : 1'b0;
  assign r_data_o[866] = (N3)? \nz.mem [866] : 
                         (N0)? \nz.mem [2466] : 1'b0;
  assign r_data_o[865] = (N3)? \nz.mem [865] : 
                         (N0)? \nz.mem [2465] : 1'b0;
  assign r_data_o[864] = (N3)? \nz.mem [864] : 
                         (N0)? \nz.mem [2464] : 1'b0;
  assign r_data_o[863] = (N3)? \nz.mem [863] : 
                         (N0)? \nz.mem [2463] : 1'b0;
  assign r_data_o[862] = (N3)? \nz.mem [862] : 
                         (N0)? \nz.mem [2462] : 1'b0;
  assign r_data_o[861] = (N3)? \nz.mem [861] : 
                         (N0)? \nz.mem [2461] : 1'b0;
  assign r_data_o[860] = (N3)? \nz.mem [860] : 
                         (N0)? \nz.mem [2460] : 1'b0;
  assign r_data_o[859] = (N3)? \nz.mem [859] : 
                         (N0)? \nz.mem [2459] : 1'b0;
  assign r_data_o[858] = (N3)? \nz.mem [858] : 
                         (N0)? \nz.mem [2458] : 1'b0;
  assign r_data_o[857] = (N3)? \nz.mem [857] : 
                         (N0)? \nz.mem [2457] : 1'b0;
  assign r_data_o[856] = (N3)? \nz.mem [856] : 
                         (N0)? \nz.mem [2456] : 1'b0;
  assign r_data_o[855] = (N3)? \nz.mem [855] : 
                         (N0)? \nz.mem [2455] : 1'b0;
  assign r_data_o[854] = (N3)? \nz.mem [854] : 
                         (N0)? \nz.mem [2454] : 1'b0;
  assign r_data_o[853] = (N3)? \nz.mem [853] : 
                         (N0)? \nz.mem [2453] : 1'b0;
  assign r_data_o[852] = (N3)? \nz.mem [852] : 
                         (N0)? \nz.mem [2452] : 1'b0;
  assign r_data_o[851] = (N3)? \nz.mem [851] : 
                         (N0)? \nz.mem [2451] : 1'b0;
  assign r_data_o[850] = (N3)? \nz.mem [850] : 
                         (N0)? \nz.mem [2450] : 1'b0;
  assign r_data_o[849] = (N3)? \nz.mem [849] : 
                         (N0)? \nz.mem [2449] : 1'b0;
  assign r_data_o[848] = (N3)? \nz.mem [848] : 
                         (N0)? \nz.mem [2448] : 1'b0;
  assign r_data_o[847] = (N3)? \nz.mem [847] : 
                         (N0)? \nz.mem [2447] : 1'b0;
  assign r_data_o[846] = (N3)? \nz.mem [846] : 
                         (N0)? \nz.mem [2446] : 1'b0;
  assign r_data_o[845] = (N3)? \nz.mem [845] : 
                         (N0)? \nz.mem [2445] : 1'b0;
  assign r_data_o[844] = (N3)? \nz.mem [844] : 
                         (N0)? \nz.mem [2444] : 1'b0;
  assign r_data_o[843] = (N3)? \nz.mem [843] : 
                         (N0)? \nz.mem [2443] : 1'b0;
  assign r_data_o[842] = (N3)? \nz.mem [842] : 
                         (N0)? \nz.mem [2442] : 1'b0;
  assign r_data_o[841] = (N3)? \nz.mem [841] : 
                         (N0)? \nz.mem [2441] : 1'b0;
  assign r_data_o[840] = (N3)? \nz.mem [840] : 
                         (N0)? \nz.mem [2440] : 1'b0;
  assign r_data_o[839] = (N3)? \nz.mem [839] : 
                         (N0)? \nz.mem [2439] : 1'b0;
  assign r_data_o[838] = (N3)? \nz.mem [838] : 
                         (N0)? \nz.mem [2438] : 1'b0;
  assign r_data_o[837] = (N3)? \nz.mem [837] : 
                         (N0)? \nz.mem [2437] : 1'b0;
  assign r_data_o[836] = (N3)? \nz.mem [836] : 
                         (N0)? \nz.mem [2436] : 1'b0;
  assign r_data_o[835] = (N3)? \nz.mem [835] : 
                         (N0)? \nz.mem [2435] : 1'b0;
  assign r_data_o[834] = (N3)? \nz.mem [834] : 
                         (N0)? \nz.mem [2434] : 1'b0;
  assign r_data_o[833] = (N3)? \nz.mem [833] : 
                         (N0)? \nz.mem [2433] : 1'b0;
  assign r_data_o[832] = (N3)? \nz.mem [832] : 
                         (N0)? \nz.mem [2432] : 1'b0;
  assign r_data_o[831] = (N3)? \nz.mem [831] : 
                         (N0)? \nz.mem [2431] : 1'b0;
  assign r_data_o[830] = (N3)? \nz.mem [830] : 
                         (N0)? \nz.mem [2430] : 1'b0;
  assign r_data_o[829] = (N3)? \nz.mem [829] : 
                         (N0)? \nz.mem [2429] : 1'b0;
  assign r_data_o[828] = (N3)? \nz.mem [828] : 
                         (N0)? \nz.mem [2428] : 1'b0;
  assign r_data_o[827] = (N3)? \nz.mem [827] : 
                         (N0)? \nz.mem [2427] : 1'b0;
  assign r_data_o[826] = (N3)? \nz.mem [826] : 
                         (N0)? \nz.mem [2426] : 1'b0;
  assign r_data_o[825] = (N3)? \nz.mem [825] : 
                         (N0)? \nz.mem [2425] : 1'b0;
  assign r_data_o[824] = (N3)? \nz.mem [824] : 
                         (N0)? \nz.mem [2424] : 1'b0;
  assign r_data_o[823] = (N3)? \nz.mem [823] : 
                         (N0)? \nz.mem [2423] : 1'b0;
  assign r_data_o[822] = (N3)? \nz.mem [822] : 
                         (N0)? \nz.mem [2422] : 1'b0;
  assign r_data_o[821] = (N3)? \nz.mem [821] : 
                         (N0)? \nz.mem [2421] : 1'b0;
  assign r_data_o[820] = (N3)? \nz.mem [820] : 
                         (N0)? \nz.mem [2420] : 1'b0;
  assign r_data_o[819] = (N3)? \nz.mem [819] : 
                         (N0)? \nz.mem [2419] : 1'b0;
  assign r_data_o[818] = (N3)? \nz.mem [818] : 
                         (N0)? \nz.mem [2418] : 1'b0;
  assign r_data_o[817] = (N3)? \nz.mem [817] : 
                         (N0)? \nz.mem [2417] : 1'b0;
  assign r_data_o[816] = (N3)? \nz.mem [816] : 
                         (N0)? \nz.mem [2416] : 1'b0;
  assign r_data_o[815] = (N3)? \nz.mem [815] : 
                         (N0)? \nz.mem [2415] : 1'b0;
  assign r_data_o[814] = (N3)? \nz.mem [814] : 
                         (N0)? \nz.mem [2414] : 1'b0;
  assign r_data_o[813] = (N3)? \nz.mem [813] : 
                         (N0)? \nz.mem [2413] : 1'b0;
  assign r_data_o[812] = (N3)? \nz.mem [812] : 
                         (N0)? \nz.mem [2412] : 1'b0;
  assign r_data_o[811] = (N3)? \nz.mem [811] : 
                         (N0)? \nz.mem [2411] : 1'b0;
  assign r_data_o[810] = (N3)? \nz.mem [810] : 
                         (N0)? \nz.mem [2410] : 1'b0;
  assign r_data_o[809] = (N3)? \nz.mem [809] : 
                         (N0)? \nz.mem [2409] : 1'b0;
  assign r_data_o[808] = (N3)? \nz.mem [808] : 
                         (N0)? \nz.mem [2408] : 1'b0;
  assign r_data_o[807] = (N3)? \nz.mem [807] : 
                         (N0)? \nz.mem [2407] : 1'b0;
  assign r_data_o[806] = (N3)? \nz.mem [806] : 
                         (N0)? \nz.mem [2406] : 1'b0;
  assign r_data_o[805] = (N3)? \nz.mem [805] : 
                         (N0)? \nz.mem [2405] : 1'b0;
  assign r_data_o[804] = (N3)? \nz.mem [804] : 
                         (N0)? \nz.mem [2404] : 1'b0;
  assign r_data_o[803] = (N3)? \nz.mem [803] : 
                         (N0)? \nz.mem [2403] : 1'b0;
  assign r_data_o[802] = (N3)? \nz.mem [802] : 
                         (N0)? \nz.mem [2402] : 1'b0;
  assign r_data_o[801] = (N3)? \nz.mem [801] : 
                         (N0)? \nz.mem [2401] : 1'b0;
  assign r_data_o[800] = (N3)? \nz.mem [800] : 
                         (N0)? \nz.mem [2400] : 1'b0;
  assign r_data_o[799] = (N3)? \nz.mem [799] : 
                         (N0)? \nz.mem [2399] : 1'b0;
  assign r_data_o[798] = (N3)? \nz.mem [798] : 
                         (N0)? \nz.mem [2398] : 1'b0;
  assign r_data_o[797] = (N3)? \nz.mem [797] : 
                         (N0)? \nz.mem [2397] : 1'b0;
  assign r_data_o[796] = (N3)? \nz.mem [796] : 
                         (N0)? \nz.mem [2396] : 1'b0;
  assign r_data_o[795] = (N3)? \nz.mem [795] : 
                         (N0)? \nz.mem [2395] : 1'b0;
  assign r_data_o[794] = (N3)? \nz.mem [794] : 
                         (N0)? \nz.mem [2394] : 1'b0;
  assign r_data_o[793] = (N3)? \nz.mem [793] : 
                         (N0)? \nz.mem [2393] : 1'b0;
  assign r_data_o[792] = (N3)? \nz.mem [792] : 
                         (N0)? \nz.mem [2392] : 1'b0;
  assign r_data_o[791] = (N3)? \nz.mem [791] : 
                         (N0)? \nz.mem [2391] : 1'b0;
  assign r_data_o[790] = (N3)? \nz.mem [790] : 
                         (N0)? \nz.mem [2390] : 1'b0;
  assign r_data_o[789] = (N3)? \nz.mem [789] : 
                         (N0)? \nz.mem [2389] : 1'b0;
  assign r_data_o[788] = (N3)? \nz.mem [788] : 
                         (N0)? \nz.mem [2388] : 1'b0;
  assign r_data_o[787] = (N3)? \nz.mem [787] : 
                         (N0)? \nz.mem [2387] : 1'b0;
  assign r_data_o[786] = (N3)? \nz.mem [786] : 
                         (N0)? \nz.mem [2386] : 1'b0;
  assign r_data_o[785] = (N3)? \nz.mem [785] : 
                         (N0)? \nz.mem [2385] : 1'b0;
  assign r_data_o[784] = (N3)? \nz.mem [784] : 
                         (N0)? \nz.mem [2384] : 1'b0;
  assign r_data_o[783] = (N3)? \nz.mem [783] : 
                         (N0)? \nz.mem [2383] : 1'b0;
  assign r_data_o[782] = (N3)? \nz.mem [782] : 
                         (N0)? \nz.mem [2382] : 1'b0;
  assign r_data_o[781] = (N3)? \nz.mem [781] : 
                         (N0)? \nz.mem [2381] : 1'b0;
  assign r_data_o[780] = (N3)? \nz.mem [780] : 
                         (N0)? \nz.mem [2380] : 1'b0;
  assign r_data_o[779] = (N3)? \nz.mem [779] : 
                         (N0)? \nz.mem [2379] : 1'b0;
  assign r_data_o[778] = (N3)? \nz.mem [778] : 
                         (N0)? \nz.mem [2378] : 1'b0;
  assign r_data_o[777] = (N3)? \nz.mem [777] : 
                         (N0)? \nz.mem [2377] : 1'b0;
  assign r_data_o[776] = (N3)? \nz.mem [776] : 
                         (N0)? \nz.mem [2376] : 1'b0;
  assign r_data_o[775] = (N3)? \nz.mem [775] : 
                         (N0)? \nz.mem [2375] : 1'b0;
  assign r_data_o[774] = (N3)? \nz.mem [774] : 
                         (N0)? \nz.mem [2374] : 1'b0;
  assign r_data_o[773] = (N3)? \nz.mem [773] : 
                         (N0)? \nz.mem [2373] : 1'b0;
  assign r_data_o[772] = (N3)? \nz.mem [772] : 
                         (N0)? \nz.mem [2372] : 1'b0;
  assign r_data_o[771] = (N3)? \nz.mem [771] : 
                         (N0)? \nz.mem [2371] : 1'b0;
  assign r_data_o[770] = (N3)? \nz.mem [770] : 
                         (N0)? \nz.mem [2370] : 1'b0;
  assign r_data_o[769] = (N3)? \nz.mem [769] : 
                         (N0)? \nz.mem [2369] : 1'b0;
  assign r_data_o[768] = (N3)? \nz.mem [768] : 
                         (N0)? \nz.mem [2368] : 1'b0;
  assign r_data_o[767] = (N3)? \nz.mem [767] : 
                         (N0)? \nz.mem [2367] : 1'b0;
  assign r_data_o[766] = (N3)? \nz.mem [766] : 
                         (N0)? \nz.mem [2366] : 1'b0;
  assign r_data_o[765] = (N3)? \nz.mem [765] : 
                         (N0)? \nz.mem [2365] : 1'b0;
  assign r_data_o[764] = (N3)? \nz.mem [764] : 
                         (N0)? \nz.mem [2364] : 1'b0;
  assign r_data_o[763] = (N3)? \nz.mem [763] : 
                         (N0)? \nz.mem [2363] : 1'b0;
  assign r_data_o[762] = (N3)? \nz.mem [762] : 
                         (N0)? \nz.mem [2362] : 1'b0;
  assign r_data_o[761] = (N3)? \nz.mem [761] : 
                         (N0)? \nz.mem [2361] : 1'b0;
  assign r_data_o[760] = (N3)? \nz.mem [760] : 
                         (N0)? \nz.mem [2360] : 1'b0;
  assign r_data_o[759] = (N3)? \nz.mem [759] : 
                         (N0)? \nz.mem [2359] : 1'b0;
  assign r_data_o[758] = (N3)? \nz.mem [758] : 
                         (N0)? \nz.mem [2358] : 1'b0;
  assign r_data_o[757] = (N3)? \nz.mem [757] : 
                         (N0)? \nz.mem [2357] : 1'b0;
  assign r_data_o[756] = (N3)? \nz.mem [756] : 
                         (N0)? \nz.mem [2356] : 1'b0;
  assign r_data_o[755] = (N3)? \nz.mem [755] : 
                         (N0)? \nz.mem [2355] : 1'b0;
  assign r_data_o[754] = (N3)? \nz.mem [754] : 
                         (N0)? \nz.mem [2354] : 1'b0;
  assign r_data_o[753] = (N3)? \nz.mem [753] : 
                         (N0)? \nz.mem [2353] : 1'b0;
  assign r_data_o[752] = (N3)? \nz.mem [752] : 
                         (N0)? \nz.mem [2352] : 1'b0;
  assign r_data_o[751] = (N3)? \nz.mem [751] : 
                         (N0)? \nz.mem [2351] : 1'b0;
  assign r_data_o[750] = (N3)? \nz.mem [750] : 
                         (N0)? \nz.mem [2350] : 1'b0;
  assign r_data_o[749] = (N3)? \nz.mem [749] : 
                         (N0)? \nz.mem [2349] : 1'b0;
  assign r_data_o[748] = (N3)? \nz.mem [748] : 
                         (N0)? \nz.mem [2348] : 1'b0;
  assign r_data_o[747] = (N3)? \nz.mem [747] : 
                         (N0)? \nz.mem [2347] : 1'b0;
  assign r_data_o[746] = (N3)? \nz.mem [746] : 
                         (N0)? \nz.mem [2346] : 1'b0;
  assign r_data_o[745] = (N3)? \nz.mem [745] : 
                         (N0)? \nz.mem [2345] : 1'b0;
  assign r_data_o[744] = (N3)? \nz.mem [744] : 
                         (N0)? \nz.mem [2344] : 1'b0;
  assign r_data_o[743] = (N3)? \nz.mem [743] : 
                         (N0)? \nz.mem [2343] : 1'b0;
  assign r_data_o[742] = (N3)? \nz.mem [742] : 
                         (N0)? \nz.mem [2342] : 1'b0;
  assign r_data_o[741] = (N3)? \nz.mem [741] : 
                         (N0)? \nz.mem [2341] : 1'b0;
  assign r_data_o[740] = (N3)? \nz.mem [740] : 
                         (N0)? \nz.mem [2340] : 1'b0;
  assign r_data_o[739] = (N3)? \nz.mem [739] : 
                         (N0)? \nz.mem [2339] : 1'b0;
  assign r_data_o[738] = (N3)? \nz.mem [738] : 
                         (N0)? \nz.mem [2338] : 1'b0;
  assign r_data_o[737] = (N3)? \nz.mem [737] : 
                         (N0)? \nz.mem [2337] : 1'b0;
  assign r_data_o[736] = (N3)? \nz.mem [736] : 
                         (N0)? \nz.mem [2336] : 1'b0;
  assign r_data_o[735] = (N3)? \nz.mem [735] : 
                         (N0)? \nz.mem [2335] : 1'b0;
  assign r_data_o[734] = (N3)? \nz.mem [734] : 
                         (N0)? \nz.mem [2334] : 1'b0;
  assign r_data_o[733] = (N3)? \nz.mem [733] : 
                         (N0)? \nz.mem [2333] : 1'b0;
  assign r_data_o[732] = (N3)? \nz.mem [732] : 
                         (N0)? \nz.mem [2332] : 1'b0;
  assign r_data_o[731] = (N3)? \nz.mem [731] : 
                         (N0)? \nz.mem [2331] : 1'b0;
  assign r_data_o[730] = (N3)? \nz.mem [730] : 
                         (N0)? \nz.mem [2330] : 1'b0;
  assign r_data_o[729] = (N3)? \nz.mem [729] : 
                         (N0)? \nz.mem [2329] : 1'b0;
  assign r_data_o[728] = (N3)? \nz.mem [728] : 
                         (N0)? \nz.mem [2328] : 1'b0;
  assign r_data_o[727] = (N3)? \nz.mem [727] : 
                         (N0)? \nz.mem [2327] : 1'b0;
  assign r_data_o[726] = (N3)? \nz.mem [726] : 
                         (N0)? \nz.mem [2326] : 1'b0;
  assign r_data_o[725] = (N3)? \nz.mem [725] : 
                         (N0)? \nz.mem [2325] : 1'b0;
  assign r_data_o[724] = (N3)? \nz.mem [724] : 
                         (N0)? \nz.mem [2324] : 1'b0;
  assign r_data_o[723] = (N3)? \nz.mem [723] : 
                         (N0)? \nz.mem [2323] : 1'b0;
  assign r_data_o[722] = (N3)? \nz.mem [722] : 
                         (N0)? \nz.mem [2322] : 1'b0;
  assign r_data_o[721] = (N3)? \nz.mem [721] : 
                         (N0)? \nz.mem [2321] : 1'b0;
  assign r_data_o[720] = (N3)? \nz.mem [720] : 
                         (N0)? \nz.mem [2320] : 1'b0;
  assign r_data_o[719] = (N3)? \nz.mem [719] : 
                         (N0)? \nz.mem [2319] : 1'b0;
  assign r_data_o[718] = (N3)? \nz.mem [718] : 
                         (N0)? \nz.mem [2318] : 1'b0;
  assign r_data_o[717] = (N3)? \nz.mem [717] : 
                         (N0)? \nz.mem [2317] : 1'b0;
  assign r_data_o[716] = (N3)? \nz.mem [716] : 
                         (N0)? \nz.mem [2316] : 1'b0;
  assign r_data_o[715] = (N3)? \nz.mem [715] : 
                         (N0)? \nz.mem [2315] : 1'b0;
  assign r_data_o[714] = (N3)? \nz.mem [714] : 
                         (N0)? \nz.mem [2314] : 1'b0;
  assign r_data_o[713] = (N3)? \nz.mem [713] : 
                         (N0)? \nz.mem [2313] : 1'b0;
  assign r_data_o[712] = (N3)? \nz.mem [712] : 
                         (N0)? \nz.mem [2312] : 1'b0;
  assign r_data_o[711] = (N3)? \nz.mem [711] : 
                         (N0)? \nz.mem [2311] : 1'b0;
  assign r_data_o[710] = (N3)? \nz.mem [710] : 
                         (N0)? \nz.mem [2310] : 1'b0;
  assign r_data_o[709] = (N3)? \nz.mem [709] : 
                         (N0)? \nz.mem [2309] : 1'b0;
  assign r_data_o[708] = (N3)? \nz.mem [708] : 
                         (N0)? \nz.mem [2308] : 1'b0;
  assign r_data_o[707] = (N3)? \nz.mem [707] : 
                         (N0)? \nz.mem [2307] : 1'b0;
  assign r_data_o[706] = (N3)? \nz.mem [706] : 
                         (N0)? \nz.mem [2306] : 1'b0;
  assign r_data_o[705] = (N3)? \nz.mem [705] : 
                         (N0)? \nz.mem [2305] : 1'b0;
  assign r_data_o[704] = (N3)? \nz.mem [704] : 
                         (N0)? \nz.mem [2304] : 1'b0;
  assign r_data_o[703] = (N3)? \nz.mem [703] : 
                         (N0)? \nz.mem [2303] : 1'b0;
  assign r_data_o[702] = (N3)? \nz.mem [702] : 
                         (N0)? \nz.mem [2302] : 1'b0;
  assign r_data_o[701] = (N3)? \nz.mem [701] : 
                         (N0)? \nz.mem [2301] : 1'b0;
  assign r_data_o[700] = (N3)? \nz.mem [700] : 
                         (N0)? \nz.mem [2300] : 1'b0;
  assign r_data_o[699] = (N3)? \nz.mem [699] : 
                         (N0)? \nz.mem [2299] : 1'b0;
  assign r_data_o[698] = (N3)? \nz.mem [698] : 
                         (N0)? \nz.mem [2298] : 1'b0;
  assign r_data_o[697] = (N3)? \nz.mem [697] : 
                         (N0)? \nz.mem [2297] : 1'b0;
  assign r_data_o[696] = (N3)? \nz.mem [696] : 
                         (N0)? \nz.mem [2296] : 1'b0;
  assign r_data_o[695] = (N3)? \nz.mem [695] : 
                         (N0)? \nz.mem [2295] : 1'b0;
  assign r_data_o[694] = (N3)? \nz.mem [694] : 
                         (N0)? \nz.mem [2294] : 1'b0;
  assign r_data_o[693] = (N3)? \nz.mem [693] : 
                         (N0)? \nz.mem [2293] : 1'b0;
  assign r_data_o[692] = (N3)? \nz.mem [692] : 
                         (N0)? \nz.mem [2292] : 1'b0;
  assign r_data_o[691] = (N3)? \nz.mem [691] : 
                         (N0)? \nz.mem [2291] : 1'b0;
  assign r_data_o[690] = (N3)? \nz.mem [690] : 
                         (N0)? \nz.mem [2290] : 1'b0;
  assign r_data_o[689] = (N3)? \nz.mem [689] : 
                         (N0)? \nz.mem [2289] : 1'b0;
  assign r_data_o[688] = (N3)? \nz.mem [688] : 
                         (N0)? \nz.mem [2288] : 1'b0;
  assign r_data_o[687] = (N3)? \nz.mem [687] : 
                         (N0)? \nz.mem [2287] : 1'b0;
  assign r_data_o[686] = (N3)? \nz.mem [686] : 
                         (N0)? \nz.mem [2286] : 1'b0;
  assign r_data_o[685] = (N3)? \nz.mem [685] : 
                         (N0)? \nz.mem [2285] : 1'b0;
  assign r_data_o[684] = (N3)? \nz.mem [684] : 
                         (N0)? \nz.mem [2284] : 1'b0;
  assign r_data_o[683] = (N3)? \nz.mem [683] : 
                         (N0)? \nz.mem [2283] : 1'b0;
  assign r_data_o[682] = (N3)? \nz.mem [682] : 
                         (N0)? \nz.mem [2282] : 1'b0;
  assign r_data_o[681] = (N3)? \nz.mem [681] : 
                         (N0)? \nz.mem [2281] : 1'b0;
  assign r_data_o[680] = (N3)? \nz.mem [680] : 
                         (N0)? \nz.mem [2280] : 1'b0;
  assign r_data_o[679] = (N3)? \nz.mem [679] : 
                         (N0)? \nz.mem [2279] : 1'b0;
  assign r_data_o[678] = (N3)? \nz.mem [678] : 
                         (N0)? \nz.mem [2278] : 1'b0;
  assign r_data_o[677] = (N3)? \nz.mem [677] : 
                         (N0)? \nz.mem [2277] : 1'b0;
  assign r_data_o[676] = (N3)? \nz.mem [676] : 
                         (N0)? \nz.mem [2276] : 1'b0;
  assign r_data_o[675] = (N3)? \nz.mem [675] : 
                         (N0)? \nz.mem [2275] : 1'b0;
  assign r_data_o[674] = (N3)? \nz.mem [674] : 
                         (N0)? \nz.mem [2274] : 1'b0;
  assign r_data_o[673] = (N3)? \nz.mem [673] : 
                         (N0)? \nz.mem [2273] : 1'b0;
  assign r_data_o[672] = (N3)? \nz.mem [672] : 
                         (N0)? \nz.mem [2272] : 1'b0;
  assign r_data_o[671] = (N3)? \nz.mem [671] : 
                         (N0)? \nz.mem [2271] : 1'b0;
  assign r_data_o[670] = (N3)? \nz.mem [670] : 
                         (N0)? \nz.mem [2270] : 1'b0;
  assign r_data_o[669] = (N3)? \nz.mem [669] : 
                         (N0)? \nz.mem [2269] : 1'b0;
  assign r_data_o[668] = (N3)? \nz.mem [668] : 
                         (N0)? \nz.mem [2268] : 1'b0;
  assign r_data_o[667] = (N3)? \nz.mem [667] : 
                         (N0)? \nz.mem [2267] : 1'b0;
  assign r_data_o[666] = (N3)? \nz.mem [666] : 
                         (N0)? \nz.mem [2266] : 1'b0;
  assign r_data_o[665] = (N3)? \nz.mem [665] : 
                         (N0)? \nz.mem [2265] : 1'b0;
  assign r_data_o[664] = (N3)? \nz.mem [664] : 
                         (N0)? \nz.mem [2264] : 1'b0;
  assign r_data_o[663] = (N3)? \nz.mem [663] : 
                         (N0)? \nz.mem [2263] : 1'b0;
  assign r_data_o[662] = (N3)? \nz.mem [662] : 
                         (N0)? \nz.mem [2262] : 1'b0;
  assign r_data_o[661] = (N3)? \nz.mem [661] : 
                         (N0)? \nz.mem [2261] : 1'b0;
  assign r_data_o[660] = (N3)? \nz.mem [660] : 
                         (N0)? \nz.mem [2260] : 1'b0;
  assign r_data_o[659] = (N3)? \nz.mem [659] : 
                         (N0)? \nz.mem [2259] : 1'b0;
  assign r_data_o[658] = (N3)? \nz.mem [658] : 
                         (N0)? \nz.mem [2258] : 1'b0;
  assign r_data_o[657] = (N3)? \nz.mem [657] : 
                         (N0)? \nz.mem [2257] : 1'b0;
  assign r_data_o[656] = (N3)? \nz.mem [656] : 
                         (N0)? \nz.mem [2256] : 1'b0;
  assign r_data_o[655] = (N3)? \nz.mem [655] : 
                         (N0)? \nz.mem [2255] : 1'b0;
  assign r_data_o[654] = (N3)? \nz.mem [654] : 
                         (N0)? \nz.mem [2254] : 1'b0;
  assign r_data_o[653] = (N3)? \nz.mem [653] : 
                         (N0)? \nz.mem [2253] : 1'b0;
  assign r_data_o[652] = (N3)? \nz.mem [652] : 
                         (N0)? \nz.mem [2252] : 1'b0;
  assign r_data_o[651] = (N3)? \nz.mem [651] : 
                         (N0)? \nz.mem [2251] : 1'b0;
  assign r_data_o[650] = (N3)? \nz.mem [650] : 
                         (N0)? \nz.mem [2250] : 1'b0;
  assign r_data_o[649] = (N3)? \nz.mem [649] : 
                         (N0)? \nz.mem [2249] : 1'b0;
  assign r_data_o[648] = (N3)? \nz.mem [648] : 
                         (N0)? \nz.mem [2248] : 1'b0;
  assign r_data_o[647] = (N3)? \nz.mem [647] : 
                         (N0)? \nz.mem [2247] : 1'b0;
  assign r_data_o[646] = (N3)? \nz.mem [646] : 
                         (N0)? \nz.mem [2246] : 1'b0;
  assign r_data_o[645] = (N3)? \nz.mem [645] : 
                         (N0)? \nz.mem [2245] : 1'b0;
  assign r_data_o[644] = (N3)? \nz.mem [644] : 
                         (N0)? \nz.mem [2244] : 1'b0;
  assign r_data_o[643] = (N3)? \nz.mem [643] : 
                         (N0)? \nz.mem [2243] : 1'b0;
  assign r_data_o[642] = (N3)? \nz.mem [642] : 
                         (N0)? \nz.mem [2242] : 1'b0;
  assign r_data_o[641] = (N3)? \nz.mem [641] : 
                         (N0)? \nz.mem [2241] : 1'b0;
  assign r_data_o[640] = (N3)? \nz.mem [640] : 
                         (N0)? \nz.mem [2240] : 1'b0;
  assign r_data_o[639] = (N3)? \nz.mem [639] : 
                         (N0)? \nz.mem [2239] : 1'b0;
  assign r_data_o[638] = (N3)? \nz.mem [638] : 
                         (N0)? \nz.mem [2238] : 1'b0;
  assign r_data_o[637] = (N3)? \nz.mem [637] : 
                         (N0)? \nz.mem [2237] : 1'b0;
  assign r_data_o[636] = (N3)? \nz.mem [636] : 
                         (N0)? \nz.mem [2236] : 1'b0;
  assign r_data_o[635] = (N3)? \nz.mem [635] : 
                         (N0)? \nz.mem [2235] : 1'b0;
  assign r_data_o[634] = (N3)? \nz.mem [634] : 
                         (N0)? \nz.mem [2234] : 1'b0;
  assign r_data_o[633] = (N3)? \nz.mem [633] : 
                         (N0)? \nz.mem [2233] : 1'b0;
  assign r_data_o[632] = (N3)? \nz.mem [632] : 
                         (N0)? \nz.mem [2232] : 1'b0;
  assign r_data_o[631] = (N3)? \nz.mem [631] : 
                         (N0)? \nz.mem [2231] : 1'b0;
  assign r_data_o[630] = (N3)? \nz.mem [630] : 
                         (N0)? \nz.mem [2230] : 1'b0;
  assign r_data_o[629] = (N3)? \nz.mem [629] : 
                         (N0)? \nz.mem [2229] : 1'b0;
  assign r_data_o[628] = (N3)? \nz.mem [628] : 
                         (N0)? \nz.mem [2228] : 1'b0;
  assign r_data_o[627] = (N3)? \nz.mem [627] : 
                         (N0)? \nz.mem [2227] : 1'b0;
  assign r_data_o[626] = (N3)? \nz.mem [626] : 
                         (N0)? \nz.mem [2226] : 1'b0;
  assign r_data_o[625] = (N3)? \nz.mem [625] : 
                         (N0)? \nz.mem [2225] : 1'b0;
  assign r_data_o[624] = (N3)? \nz.mem [624] : 
                         (N0)? \nz.mem [2224] : 1'b0;
  assign r_data_o[623] = (N3)? \nz.mem [623] : 
                         (N0)? \nz.mem [2223] : 1'b0;
  assign r_data_o[622] = (N3)? \nz.mem [622] : 
                         (N0)? \nz.mem [2222] : 1'b0;
  assign r_data_o[621] = (N3)? \nz.mem [621] : 
                         (N0)? \nz.mem [2221] : 1'b0;
  assign r_data_o[620] = (N3)? \nz.mem [620] : 
                         (N0)? \nz.mem [2220] : 1'b0;
  assign r_data_o[619] = (N3)? \nz.mem [619] : 
                         (N0)? \nz.mem [2219] : 1'b0;
  assign r_data_o[618] = (N3)? \nz.mem [618] : 
                         (N0)? \nz.mem [2218] : 1'b0;
  assign r_data_o[617] = (N3)? \nz.mem [617] : 
                         (N0)? \nz.mem [2217] : 1'b0;
  assign r_data_o[616] = (N3)? \nz.mem [616] : 
                         (N0)? \nz.mem [2216] : 1'b0;
  assign r_data_o[615] = (N3)? \nz.mem [615] : 
                         (N0)? \nz.mem [2215] : 1'b0;
  assign r_data_o[614] = (N3)? \nz.mem [614] : 
                         (N0)? \nz.mem [2214] : 1'b0;
  assign r_data_o[613] = (N3)? \nz.mem [613] : 
                         (N0)? \nz.mem [2213] : 1'b0;
  assign r_data_o[612] = (N3)? \nz.mem [612] : 
                         (N0)? \nz.mem [2212] : 1'b0;
  assign r_data_o[611] = (N3)? \nz.mem [611] : 
                         (N0)? \nz.mem [2211] : 1'b0;
  assign r_data_o[610] = (N3)? \nz.mem [610] : 
                         (N0)? \nz.mem [2210] : 1'b0;
  assign r_data_o[609] = (N3)? \nz.mem [609] : 
                         (N0)? \nz.mem [2209] : 1'b0;
  assign r_data_o[608] = (N3)? \nz.mem [608] : 
                         (N0)? \nz.mem [2208] : 1'b0;
  assign r_data_o[607] = (N3)? \nz.mem [607] : 
                         (N0)? \nz.mem [2207] : 1'b0;
  assign r_data_o[606] = (N3)? \nz.mem [606] : 
                         (N0)? \nz.mem [2206] : 1'b0;
  assign r_data_o[605] = (N3)? \nz.mem [605] : 
                         (N0)? \nz.mem [2205] : 1'b0;
  assign r_data_o[604] = (N3)? \nz.mem [604] : 
                         (N0)? \nz.mem [2204] : 1'b0;
  assign r_data_o[603] = (N3)? \nz.mem [603] : 
                         (N0)? \nz.mem [2203] : 1'b0;
  assign r_data_o[602] = (N3)? \nz.mem [602] : 
                         (N0)? \nz.mem [2202] : 1'b0;
  assign r_data_o[601] = (N3)? \nz.mem [601] : 
                         (N0)? \nz.mem [2201] : 1'b0;
  assign r_data_o[600] = (N3)? \nz.mem [600] : 
                         (N0)? \nz.mem [2200] : 1'b0;
  assign r_data_o[599] = (N3)? \nz.mem [599] : 
                         (N0)? \nz.mem [2199] : 1'b0;
  assign r_data_o[598] = (N3)? \nz.mem [598] : 
                         (N0)? \nz.mem [2198] : 1'b0;
  assign r_data_o[597] = (N3)? \nz.mem [597] : 
                         (N0)? \nz.mem [2197] : 1'b0;
  assign r_data_o[596] = (N3)? \nz.mem [596] : 
                         (N0)? \nz.mem [2196] : 1'b0;
  assign r_data_o[595] = (N3)? \nz.mem [595] : 
                         (N0)? \nz.mem [2195] : 1'b0;
  assign r_data_o[594] = (N3)? \nz.mem [594] : 
                         (N0)? \nz.mem [2194] : 1'b0;
  assign r_data_o[593] = (N3)? \nz.mem [593] : 
                         (N0)? \nz.mem [2193] : 1'b0;
  assign r_data_o[592] = (N3)? \nz.mem [592] : 
                         (N0)? \nz.mem [2192] : 1'b0;
  assign r_data_o[591] = (N3)? \nz.mem [591] : 
                         (N0)? \nz.mem [2191] : 1'b0;
  assign r_data_o[590] = (N3)? \nz.mem [590] : 
                         (N0)? \nz.mem [2190] : 1'b0;
  assign r_data_o[589] = (N3)? \nz.mem [589] : 
                         (N0)? \nz.mem [2189] : 1'b0;
  assign r_data_o[588] = (N3)? \nz.mem [588] : 
                         (N0)? \nz.mem [2188] : 1'b0;
  assign r_data_o[587] = (N3)? \nz.mem [587] : 
                         (N0)? \nz.mem [2187] : 1'b0;
  assign r_data_o[586] = (N3)? \nz.mem [586] : 
                         (N0)? \nz.mem [2186] : 1'b0;
  assign r_data_o[585] = (N3)? \nz.mem [585] : 
                         (N0)? \nz.mem [2185] : 1'b0;
  assign r_data_o[584] = (N3)? \nz.mem [584] : 
                         (N0)? \nz.mem [2184] : 1'b0;
  assign r_data_o[583] = (N3)? \nz.mem [583] : 
                         (N0)? \nz.mem [2183] : 1'b0;
  assign r_data_o[582] = (N3)? \nz.mem [582] : 
                         (N0)? \nz.mem [2182] : 1'b0;
  assign r_data_o[581] = (N3)? \nz.mem [581] : 
                         (N0)? \nz.mem [2181] : 1'b0;
  assign r_data_o[580] = (N3)? \nz.mem [580] : 
                         (N0)? \nz.mem [2180] : 1'b0;
  assign r_data_o[579] = (N3)? \nz.mem [579] : 
                         (N0)? \nz.mem [2179] : 1'b0;
  assign r_data_o[578] = (N3)? \nz.mem [578] : 
                         (N0)? \nz.mem [2178] : 1'b0;
  assign r_data_o[577] = (N3)? \nz.mem [577] : 
                         (N0)? \nz.mem [2177] : 1'b0;
  assign r_data_o[576] = (N3)? \nz.mem [576] : 
                         (N0)? \nz.mem [2176] : 1'b0;
  assign r_data_o[575] = (N3)? \nz.mem [575] : 
                         (N0)? \nz.mem [2175] : 1'b0;
  assign r_data_o[574] = (N3)? \nz.mem [574] : 
                         (N0)? \nz.mem [2174] : 1'b0;
  assign r_data_o[573] = (N3)? \nz.mem [573] : 
                         (N0)? \nz.mem [2173] : 1'b0;
  assign r_data_o[572] = (N3)? \nz.mem [572] : 
                         (N0)? \nz.mem [2172] : 1'b0;
  assign r_data_o[571] = (N3)? \nz.mem [571] : 
                         (N0)? \nz.mem [2171] : 1'b0;
  assign r_data_o[570] = (N3)? \nz.mem [570] : 
                         (N0)? \nz.mem [2170] : 1'b0;
  assign r_data_o[569] = (N3)? \nz.mem [569] : 
                         (N0)? \nz.mem [2169] : 1'b0;
  assign r_data_o[568] = (N3)? \nz.mem [568] : 
                         (N0)? \nz.mem [2168] : 1'b0;
  assign r_data_o[567] = (N3)? \nz.mem [567] : 
                         (N0)? \nz.mem [2167] : 1'b0;
  assign r_data_o[566] = (N3)? \nz.mem [566] : 
                         (N0)? \nz.mem [2166] : 1'b0;
  assign r_data_o[565] = (N3)? \nz.mem [565] : 
                         (N0)? \nz.mem [2165] : 1'b0;
  assign r_data_o[564] = (N3)? \nz.mem [564] : 
                         (N0)? \nz.mem [2164] : 1'b0;
  assign r_data_o[563] = (N3)? \nz.mem [563] : 
                         (N0)? \nz.mem [2163] : 1'b0;
  assign r_data_o[562] = (N3)? \nz.mem [562] : 
                         (N0)? \nz.mem [2162] : 1'b0;
  assign r_data_o[561] = (N3)? \nz.mem [561] : 
                         (N0)? \nz.mem [2161] : 1'b0;
  assign r_data_o[560] = (N3)? \nz.mem [560] : 
                         (N0)? \nz.mem [2160] : 1'b0;
  assign r_data_o[559] = (N3)? \nz.mem [559] : 
                         (N0)? \nz.mem [2159] : 1'b0;
  assign r_data_o[558] = (N3)? \nz.mem [558] : 
                         (N0)? \nz.mem [2158] : 1'b0;
  assign r_data_o[557] = (N3)? \nz.mem [557] : 
                         (N0)? \nz.mem [2157] : 1'b0;
  assign r_data_o[556] = (N3)? \nz.mem [556] : 
                         (N0)? \nz.mem [2156] : 1'b0;
  assign r_data_o[555] = (N3)? \nz.mem [555] : 
                         (N0)? \nz.mem [2155] : 1'b0;
  assign r_data_o[554] = (N3)? \nz.mem [554] : 
                         (N0)? \nz.mem [2154] : 1'b0;
  assign r_data_o[553] = (N3)? \nz.mem [553] : 
                         (N0)? \nz.mem [2153] : 1'b0;
  assign r_data_o[552] = (N3)? \nz.mem [552] : 
                         (N0)? \nz.mem [2152] : 1'b0;
  assign r_data_o[551] = (N3)? \nz.mem [551] : 
                         (N0)? \nz.mem [2151] : 1'b0;
  assign r_data_o[550] = (N3)? \nz.mem [550] : 
                         (N0)? \nz.mem [2150] : 1'b0;
  assign r_data_o[549] = (N3)? \nz.mem [549] : 
                         (N0)? \nz.mem [2149] : 1'b0;
  assign r_data_o[548] = (N3)? \nz.mem [548] : 
                         (N0)? \nz.mem [2148] : 1'b0;
  assign r_data_o[547] = (N3)? \nz.mem [547] : 
                         (N0)? \nz.mem [2147] : 1'b0;
  assign r_data_o[546] = (N3)? \nz.mem [546] : 
                         (N0)? \nz.mem [2146] : 1'b0;
  assign r_data_o[545] = (N3)? \nz.mem [545] : 
                         (N0)? \nz.mem [2145] : 1'b0;
  assign r_data_o[544] = (N3)? \nz.mem [544] : 
                         (N0)? \nz.mem [2144] : 1'b0;
  assign r_data_o[543] = (N3)? \nz.mem [543] : 
                         (N0)? \nz.mem [2143] : 1'b0;
  assign r_data_o[542] = (N3)? \nz.mem [542] : 
                         (N0)? \nz.mem [2142] : 1'b0;
  assign r_data_o[541] = (N3)? \nz.mem [541] : 
                         (N0)? \nz.mem [2141] : 1'b0;
  assign r_data_o[540] = (N3)? \nz.mem [540] : 
                         (N0)? \nz.mem [2140] : 1'b0;
  assign r_data_o[539] = (N3)? \nz.mem [539] : 
                         (N0)? \nz.mem [2139] : 1'b0;
  assign r_data_o[538] = (N3)? \nz.mem [538] : 
                         (N0)? \nz.mem [2138] : 1'b0;
  assign r_data_o[537] = (N3)? \nz.mem [537] : 
                         (N0)? \nz.mem [2137] : 1'b0;
  assign r_data_o[536] = (N3)? \nz.mem [536] : 
                         (N0)? \nz.mem [2136] : 1'b0;
  assign r_data_o[535] = (N3)? \nz.mem [535] : 
                         (N0)? \nz.mem [2135] : 1'b0;
  assign r_data_o[534] = (N3)? \nz.mem [534] : 
                         (N0)? \nz.mem [2134] : 1'b0;
  assign r_data_o[533] = (N3)? \nz.mem [533] : 
                         (N0)? \nz.mem [2133] : 1'b0;
  assign r_data_o[532] = (N3)? \nz.mem [532] : 
                         (N0)? \nz.mem [2132] : 1'b0;
  assign r_data_o[531] = (N3)? \nz.mem [531] : 
                         (N0)? \nz.mem [2131] : 1'b0;
  assign r_data_o[530] = (N3)? \nz.mem [530] : 
                         (N0)? \nz.mem [2130] : 1'b0;
  assign r_data_o[529] = (N3)? \nz.mem [529] : 
                         (N0)? \nz.mem [2129] : 1'b0;
  assign r_data_o[528] = (N3)? \nz.mem [528] : 
                         (N0)? \nz.mem [2128] : 1'b0;
  assign r_data_o[527] = (N3)? \nz.mem [527] : 
                         (N0)? \nz.mem [2127] : 1'b0;
  assign r_data_o[526] = (N3)? \nz.mem [526] : 
                         (N0)? \nz.mem [2126] : 1'b0;
  assign r_data_o[525] = (N3)? \nz.mem [525] : 
                         (N0)? \nz.mem [2125] : 1'b0;
  assign r_data_o[524] = (N3)? \nz.mem [524] : 
                         (N0)? \nz.mem [2124] : 1'b0;
  assign r_data_o[523] = (N3)? \nz.mem [523] : 
                         (N0)? \nz.mem [2123] : 1'b0;
  assign r_data_o[522] = (N3)? \nz.mem [522] : 
                         (N0)? \nz.mem [2122] : 1'b0;
  assign r_data_o[521] = (N3)? \nz.mem [521] : 
                         (N0)? \nz.mem [2121] : 1'b0;
  assign r_data_o[520] = (N3)? \nz.mem [520] : 
                         (N0)? \nz.mem [2120] : 1'b0;
  assign r_data_o[519] = (N3)? \nz.mem [519] : 
                         (N0)? \nz.mem [2119] : 1'b0;
  assign r_data_o[518] = (N3)? \nz.mem [518] : 
                         (N0)? \nz.mem [2118] : 1'b0;
  assign r_data_o[517] = (N3)? \nz.mem [517] : 
                         (N0)? \nz.mem [2117] : 1'b0;
  assign r_data_o[516] = (N3)? \nz.mem [516] : 
                         (N0)? \nz.mem [2116] : 1'b0;
  assign r_data_o[515] = (N3)? \nz.mem [515] : 
                         (N0)? \nz.mem [2115] : 1'b0;
  assign r_data_o[514] = (N3)? \nz.mem [514] : 
                         (N0)? \nz.mem [2114] : 1'b0;
  assign r_data_o[513] = (N3)? \nz.mem [513] : 
                         (N0)? \nz.mem [2113] : 1'b0;
  assign r_data_o[512] = (N3)? \nz.mem [512] : 
                         (N0)? \nz.mem [2112] : 1'b0;
  assign r_data_o[511] = (N3)? \nz.mem [511] : 
                         (N0)? \nz.mem [2111] : 1'b0;
  assign r_data_o[510] = (N3)? \nz.mem [510] : 
                         (N0)? \nz.mem [2110] : 1'b0;
  assign r_data_o[509] = (N3)? \nz.mem [509] : 
                         (N0)? \nz.mem [2109] : 1'b0;
  assign r_data_o[508] = (N3)? \nz.mem [508] : 
                         (N0)? \nz.mem [2108] : 1'b0;
  assign r_data_o[507] = (N3)? \nz.mem [507] : 
                         (N0)? \nz.mem [2107] : 1'b0;
  assign r_data_o[506] = (N3)? \nz.mem [506] : 
                         (N0)? \nz.mem [2106] : 1'b0;
  assign r_data_o[505] = (N3)? \nz.mem [505] : 
                         (N0)? \nz.mem [2105] : 1'b0;
  assign r_data_o[504] = (N3)? \nz.mem [504] : 
                         (N0)? \nz.mem [2104] : 1'b0;
  assign r_data_o[503] = (N3)? \nz.mem [503] : 
                         (N0)? \nz.mem [2103] : 1'b0;
  assign r_data_o[502] = (N3)? \nz.mem [502] : 
                         (N0)? \nz.mem [2102] : 1'b0;
  assign r_data_o[501] = (N3)? \nz.mem [501] : 
                         (N0)? \nz.mem [2101] : 1'b0;
  assign r_data_o[500] = (N3)? \nz.mem [500] : 
                         (N0)? \nz.mem [2100] : 1'b0;
  assign r_data_o[499] = (N3)? \nz.mem [499] : 
                         (N0)? \nz.mem [2099] : 1'b0;
  assign r_data_o[498] = (N3)? \nz.mem [498] : 
                         (N0)? \nz.mem [2098] : 1'b0;
  assign r_data_o[497] = (N3)? \nz.mem [497] : 
                         (N0)? \nz.mem [2097] : 1'b0;
  assign r_data_o[496] = (N3)? \nz.mem [496] : 
                         (N0)? \nz.mem [2096] : 1'b0;
  assign r_data_o[495] = (N3)? \nz.mem [495] : 
                         (N0)? \nz.mem [2095] : 1'b0;
  assign r_data_o[494] = (N3)? \nz.mem [494] : 
                         (N0)? \nz.mem [2094] : 1'b0;
  assign r_data_o[493] = (N3)? \nz.mem [493] : 
                         (N0)? \nz.mem [2093] : 1'b0;
  assign r_data_o[492] = (N3)? \nz.mem [492] : 
                         (N0)? \nz.mem [2092] : 1'b0;
  assign r_data_o[491] = (N3)? \nz.mem [491] : 
                         (N0)? \nz.mem [2091] : 1'b0;
  assign r_data_o[490] = (N3)? \nz.mem [490] : 
                         (N0)? \nz.mem [2090] : 1'b0;
  assign r_data_o[489] = (N3)? \nz.mem [489] : 
                         (N0)? \nz.mem [2089] : 1'b0;
  assign r_data_o[488] = (N3)? \nz.mem [488] : 
                         (N0)? \nz.mem [2088] : 1'b0;
  assign r_data_o[487] = (N3)? \nz.mem [487] : 
                         (N0)? \nz.mem [2087] : 1'b0;
  assign r_data_o[486] = (N3)? \nz.mem [486] : 
                         (N0)? \nz.mem [2086] : 1'b0;
  assign r_data_o[485] = (N3)? \nz.mem [485] : 
                         (N0)? \nz.mem [2085] : 1'b0;
  assign r_data_o[484] = (N3)? \nz.mem [484] : 
                         (N0)? \nz.mem [2084] : 1'b0;
  assign r_data_o[483] = (N3)? \nz.mem [483] : 
                         (N0)? \nz.mem [2083] : 1'b0;
  assign r_data_o[482] = (N3)? \nz.mem [482] : 
                         (N0)? \nz.mem [2082] : 1'b0;
  assign r_data_o[481] = (N3)? \nz.mem [481] : 
                         (N0)? \nz.mem [2081] : 1'b0;
  assign r_data_o[480] = (N3)? \nz.mem [480] : 
                         (N0)? \nz.mem [2080] : 1'b0;
  assign r_data_o[479] = (N3)? \nz.mem [479] : 
                         (N0)? \nz.mem [2079] : 1'b0;
  assign r_data_o[478] = (N3)? \nz.mem [478] : 
                         (N0)? \nz.mem [2078] : 1'b0;
  assign r_data_o[477] = (N3)? \nz.mem [477] : 
                         (N0)? \nz.mem [2077] : 1'b0;
  assign r_data_o[476] = (N3)? \nz.mem [476] : 
                         (N0)? \nz.mem [2076] : 1'b0;
  assign r_data_o[475] = (N3)? \nz.mem [475] : 
                         (N0)? \nz.mem [2075] : 1'b0;
  assign r_data_o[474] = (N3)? \nz.mem [474] : 
                         (N0)? \nz.mem [2074] : 1'b0;
  assign r_data_o[473] = (N3)? \nz.mem [473] : 
                         (N0)? \nz.mem [2073] : 1'b0;
  assign r_data_o[472] = (N3)? \nz.mem [472] : 
                         (N0)? \nz.mem [2072] : 1'b0;
  assign r_data_o[471] = (N3)? \nz.mem [471] : 
                         (N0)? \nz.mem [2071] : 1'b0;
  assign r_data_o[470] = (N3)? \nz.mem [470] : 
                         (N0)? \nz.mem [2070] : 1'b0;
  assign r_data_o[469] = (N3)? \nz.mem [469] : 
                         (N0)? \nz.mem [2069] : 1'b0;
  assign r_data_o[468] = (N3)? \nz.mem [468] : 
                         (N0)? \nz.mem [2068] : 1'b0;
  assign r_data_o[467] = (N3)? \nz.mem [467] : 
                         (N0)? \nz.mem [2067] : 1'b0;
  assign r_data_o[466] = (N3)? \nz.mem [466] : 
                         (N0)? \nz.mem [2066] : 1'b0;
  assign r_data_o[465] = (N3)? \nz.mem [465] : 
                         (N0)? \nz.mem [2065] : 1'b0;
  assign r_data_o[464] = (N3)? \nz.mem [464] : 
                         (N0)? \nz.mem [2064] : 1'b0;
  assign r_data_o[463] = (N3)? \nz.mem [463] : 
                         (N0)? \nz.mem [2063] : 1'b0;
  assign r_data_o[462] = (N3)? \nz.mem [462] : 
                         (N0)? \nz.mem [2062] : 1'b0;
  assign r_data_o[461] = (N3)? \nz.mem [461] : 
                         (N0)? \nz.mem [2061] : 1'b0;
  assign r_data_o[460] = (N3)? \nz.mem [460] : 
                         (N0)? \nz.mem [2060] : 1'b0;
  assign r_data_o[459] = (N3)? \nz.mem [459] : 
                         (N0)? \nz.mem [2059] : 1'b0;
  assign r_data_o[458] = (N3)? \nz.mem [458] : 
                         (N0)? \nz.mem [2058] : 1'b0;
  assign r_data_o[457] = (N3)? \nz.mem [457] : 
                         (N0)? \nz.mem [2057] : 1'b0;
  assign r_data_o[456] = (N3)? \nz.mem [456] : 
                         (N0)? \nz.mem [2056] : 1'b0;
  assign r_data_o[455] = (N3)? \nz.mem [455] : 
                         (N0)? \nz.mem [2055] : 1'b0;
  assign r_data_o[454] = (N3)? \nz.mem [454] : 
                         (N0)? \nz.mem [2054] : 1'b0;
  assign r_data_o[453] = (N3)? \nz.mem [453] : 
                         (N0)? \nz.mem [2053] : 1'b0;
  assign r_data_o[452] = (N3)? \nz.mem [452] : 
                         (N0)? \nz.mem [2052] : 1'b0;
  assign r_data_o[451] = (N3)? \nz.mem [451] : 
                         (N0)? \nz.mem [2051] : 1'b0;
  assign r_data_o[450] = (N3)? \nz.mem [450] : 
                         (N0)? \nz.mem [2050] : 1'b0;
  assign r_data_o[449] = (N3)? \nz.mem [449] : 
                         (N0)? \nz.mem [2049] : 1'b0;
  assign r_data_o[448] = (N3)? \nz.mem [448] : 
                         (N0)? \nz.mem [2048] : 1'b0;
  assign r_data_o[447] = (N3)? \nz.mem [447] : 
                         (N0)? \nz.mem [2047] : 1'b0;
  assign r_data_o[446] = (N3)? \nz.mem [446] : 
                         (N0)? \nz.mem [2046] : 1'b0;
  assign r_data_o[445] = (N3)? \nz.mem [445] : 
                         (N0)? \nz.mem [2045] : 1'b0;
  assign r_data_o[444] = (N3)? \nz.mem [444] : 
                         (N0)? \nz.mem [2044] : 1'b0;
  assign r_data_o[443] = (N3)? \nz.mem [443] : 
                         (N0)? \nz.mem [2043] : 1'b0;
  assign r_data_o[442] = (N3)? \nz.mem [442] : 
                         (N0)? \nz.mem [2042] : 1'b0;
  assign r_data_o[441] = (N3)? \nz.mem [441] : 
                         (N0)? \nz.mem [2041] : 1'b0;
  assign r_data_o[440] = (N3)? \nz.mem [440] : 
                         (N0)? \nz.mem [2040] : 1'b0;
  assign r_data_o[439] = (N3)? \nz.mem [439] : 
                         (N0)? \nz.mem [2039] : 1'b0;
  assign r_data_o[438] = (N3)? \nz.mem [438] : 
                         (N0)? \nz.mem [2038] : 1'b0;
  assign r_data_o[437] = (N3)? \nz.mem [437] : 
                         (N0)? \nz.mem [2037] : 1'b0;
  assign r_data_o[436] = (N3)? \nz.mem [436] : 
                         (N0)? \nz.mem [2036] : 1'b0;
  assign r_data_o[435] = (N3)? \nz.mem [435] : 
                         (N0)? \nz.mem [2035] : 1'b0;
  assign r_data_o[434] = (N3)? \nz.mem [434] : 
                         (N0)? \nz.mem [2034] : 1'b0;
  assign r_data_o[433] = (N3)? \nz.mem [433] : 
                         (N0)? \nz.mem [2033] : 1'b0;
  assign r_data_o[432] = (N3)? \nz.mem [432] : 
                         (N0)? \nz.mem [2032] : 1'b0;
  assign r_data_o[431] = (N3)? \nz.mem [431] : 
                         (N0)? \nz.mem [2031] : 1'b0;
  assign r_data_o[430] = (N3)? \nz.mem [430] : 
                         (N0)? \nz.mem [2030] : 1'b0;
  assign r_data_o[429] = (N3)? \nz.mem [429] : 
                         (N0)? \nz.mem [2029] : 1'b0;
  assign r_data_o[428] = (N3)? \nz.mem [428] : 
                         (N0)? \nz.mem [2028] : 1'b0;
  assign r_data_o[427] = (N3)? \nz.mem [427] : 
                         (N0)? \nz.mem [2027] : 1'b0;
  assign r_data_o[426] = (N3)? \nz.mem [426] : 
                         (N0)? \nz.mem [2026] : 1'b0;
  assign r_data_o[425] = (N3)? \nz.mem [425] : 
                         (N0)? \nz.mem [2025] : 1'b0;
  assign r_data_o[424] = (N3)? \nz.mem [424] : 
                         (N0)? \nz.mem [2024] : 1'b0;
  assign r_data_o[423] = (N3)? \nz.mem [423] : 
                         (N0)? \nz.mem [2023] : 1'b0;
  assign r_data_o[422] = (N3)? \nz.mem [422] : 
                         (N0)? \nz.mem [2022] : 1'b0;
  assign r_data_o[421] = (N3)? \nz.mem [421] : 
                         (N0)? \nz.mem [2021] : 1'b0;
  assign r_data_o[420] = (N3)? \nz.mem [420] : 
                         (N0)? \nz.mem [2020] : 1'b0;
  assign r_data_o[419] = (N3)? \nz.mem [419] : 
                         (N0)? \nz.mem [2019] : 1'b0;
  assign r_data_o[418] = (N3)? \nz.mem [418] : 
                         (N0)? \nz.mem [2018] : 1'b0;
  assign r_data_o[417] = (N3)? \nz.mem [417] : 
                         (N0)? \nz.mem [2017] : 1'b0;
  assign r_data_o[416] = (N3)? \nz.mem [416] : 
                         (N0)? \nz.mem [2016] : 1'b0;
  assign r_data_o[415] = (N3)? \nz.mem [415] : 
                         (N0)? \nz.mem [2015] : 1'b0;
  assign r_data_o[414] = (N3)? \nz.mem [414] : 
                         (N0)? \nz.mem [2014] : 1'b0;
  assign r_data_o[413] = (N3)? \nz.mem [413] : 
                         (N0)? \nz.mem [2013] : 1'b0;
  assign r_data_o[412] = (N3)? \nz.mem [412] : 
                         (N0)? \nz.mem [2012] : 1'b0;
  assign r_data_o[411] = (N3)? \nz.mem [411] : 
                         (N0)? \nz.mem [2011] : 1'b0;
  assign r_data_o[410] = (N3)? \nz.mem [410] : 
                         (N0)? \nz.mem [2010] : 1'b0;
  assign r_data_o[409] = (N3)? \nz.mem [409] : 
                         (N0)? \nz.mem [2009] : 1'b0;
  assign r_data_o[408] = (N3)? \nz.mem [408] : 
                         (N0)? \nz.mem [2008] : 1'b0;
  assign r_data_o[407] = (N3)? \nz.mem [407] : 
                         (N0)? \nz.mem [2007] : 1'b0;
  assign r_data_o[406] = (N3)? \nz.mem [406] : 
                         (N0)? \nz.mem [2006] : 1'b0;
  assign r_data_o[405] = (N3)? \nz.mem [405] : 
                         (N0)? \nz.mem [2005] : 1'b0;
  assign r_data_o[404] = (N3)? \nz.mem [404] : 
                         (N0)? \nz.mem [2004] : 1'b0;
  assign r_data_o[403] = (N3)? \nz.mem [403] : 
                         (N0)? \nz.mem [2003] : 1'b0;
  assign r_data_o[402] = (N3)? \nz.mem [402] : 
                         (N0)? \nz.mem [2002] : 1'b0;
  assign r_data_o[401] = (N3)? \nz.mem [401] : 
                         (N0)? \nz.mem [2001] : 1'b0;
  assign r_data_o[400] = (N3)? \nz.mem [400] : 
                         (N0)? \nz.mem [2000] : 1'b0;
  assign r_data_o[399] = (N3)? \nz.mem [399] : 
                         (N0)? \nz.mem [1999] : 1'b0;
  assign r_data_o[398] = (N3)? \nz.mem [398] : 
                         (N0)? \nz.mem [1998] : 1'b0;
  assign r_data_o[397] = (N3)? \nz.mem [397] : 
                         (N0)? \nz.mem [1997] : 1'b0;
  assign r_data_o[396] = (N3)? \nz.mem [396] : 
                         (N0)? \nz.mem [1996] : 1'b0;
  assign r_data_o[395] = (N3)? \nz.mem [395] : 
                         (N0)? \nz.mem [1995] : 1'b0;
  assign r_data_o[394] = (N3)? \nz.mem [394] : 
                         (N0)? \nz.mem [1994] : 1'b0;
  assign r_data_o[393] = (N3)? \nz.mem [393] : 
                         (N0)? \nz.mem [1993] : 1'b0;
  assign r_data_o[392] = (N3)? \nz.mem [392] : 
                         (N0)? \nz.mem [1992] : 1'b0;
  assign r_data_o[391] = (N3)? \nz.mem [391] : 
                         (N0)? \nz.mem [1991] : 1'b0;
  assign r_data_o[390] = (N3)? \nz.mem [390] : 
                         (N0)? \nz.mem [1990] : 1'b0;
  assign r_data_o[389] = (N3)? \nz.mem [389] : 
                         (N0)? \nz.mem [1989] : 1'b0;
  assign r_data_o[388] = (N3)? \nz.mem [388] : 
                         (N0)? \nz.mem [1988] : 1'b0;
  assign r_data_o[387] = (N3)? \nz.mem [387] : 
                         (N0)? \nz.mem [1987] : 1'b0;
  assign r_data_o[386] = (N3)? \nz.mem [386] : 
                         (N0)? \nz.mem [1986] : 1'b0;
  assign r_data_o[385] = (N3)? \nz.mem [385] : 
                         (N0)? \nz.mem [1985] : 1'b0;
  assign r_data_o[384] = (N3)? \nz.mem [384] : 
                         (N0)? \nz.mem [1984] : 1'b0;
  assign r_data_o[383] = (N3)? \nz.mem [383] : 
                         (N0)? \nz.mem [1983] : 1'b0;
  assign r_data_o[382] = (N3)? \nz.mem [382] : 
                         (N0)? \nz.mem [1982] : 1'b0;
  assign r_data_o[381] = (N3)? \nz.mem [381] : 
                         (N0)? \nz.mem [1981] : 1'b0;
  assign r_data_o[380] = (N3)? \nz.mem [380] : 
                         (N0)? \nz.mem [1980] : 1'b0;
  assign r_data_o[379] = (N3)? \nz.mem [379] : 
                         (N0)? \nz.mem [1979] : 1'b0;
  assign r_data_o[378] = (N3)? \nz.mem [378] : 
                         (N0)? \nz.mem [1978] : 1'b0;
  assign r_data_o[377] = (N3)? \nz.mem [377] : 
                         (N0)? \nz.mem [1977] : 1'b0;
  assign r_data_o[376] = (N3)? \nz.mem [376] : 
                         (N0)? \nz.mem [1976] : 1'b0;
  assign r_data_o[375] = (N3)? \nz.mem [375] : 
                         (N0)? \nz.mem [1975] : 1'b0;
  assign r_data_o[374] = (N3)? \nz.mem [374] : 
                         (N0)? \nz.mem [1974] : 1'b0;
  assign r_data_o[373] = (N3)? \nz.mem [373] : 
                         (N0)? \nz.mem [1973] : 1'b0;
  assign r_data_o[372] = (N3)? \nz.mem [372] : 
                         (N0)? \nz.mem [1972] : 1'b0;
  assign r_data_o[371] = (N3)? \nz.mem [371] : 
                         (N0)? \nz.mem [1971] : 1'b0;
  assign r_data_o[370] = (N3)? \nz.mem [370] : 
                         (N0)? \nz.mem [1970] : 1'b0;
  assign r_data_o[369] = (N3)? \nz.mem [369] : 
                         (N0)? \nz.mem [1969] : 1'b0;
  assign r_data_o[368] = (N3)? \nz.mem [368] : 
                         (N0)? \nz.mem [1968] : 1'b0;
  assign r_data_o[367] = (N3)? \nz.mem [367] : 
                         (N0)? \nz.mem [1967] : 1'b0;
  assign r_data_o[366] = (N3)? \nz.mem [366] : 
                         (N0)? \nz.mem [1966] : 1'b0;
  assign r_data_o[365] = (N3)? \nz.mem [365] : 
                         (N0)? \nz.mem [1965] : 1'b0;
  assign r_data_o[364] = (N3)? \nz.mem [364] : 
                         (N0)? \nz.mem [1964] : 1'b0;
  assign r_data_o[363] = (N3)? \nz.mem [363] : 
                         (N0)? \nz.mem [1963] : 1'b0;
  assign r_data_o[362] = (N3)? \nz.mem [362] : 
                         (N0)? \nz.mem [1962] : 1'b0;
  assign r_data_o[361] = (N3)? \nz.mem [361] : 
                         (N0)? \nz.mem [1961] : 1'b0;
  assign r_data_o[360] = (N3)? \nz.mem [360] : 
                         (N0)? \nz.mem [1960] : 1'b0;
  assign r_data_o[359] = (N3)? \nz.mem [359] : 
                         (N0)? \nz.mem [1959] : 1'b0;
  assign r_data_o[358] = (N3)? \nz.mem [358] : 
                         (N0)? \nz.mem [1958] : 1'b0;
  assign r_data_o[357] = (N3)? \nz.mem [357] : 
                         (N0)? \nz.mem [1957] : 1'b0;
  assign r_data_o[356] = (N3)? \nz.mem [356] : 
                         (N0)? \nz.mem [1956] : 1'b0;
  assign r_data_o[355] = (N3)? \nz.mem [355] : 
                         (N0)? \nz.mem [1955] : 1'b0;
  assign r_data_o[354] = (N3)? \nz.mem [354] : 
                         (N0)? \nz.mem [1954] : 1'b0;
  assign r_data_o[353] = (N3)? \nz.mem [353] : 
                         (N0)? \nz.mem [1953] : 1'b0;
  assign r_data_o[352] = (N3)? \nz.mem [352] : 
                         (N0)? \nz.mem [1952] : 1'b0;
  assign r_data_o[351] = (N3)? \nz.mem [351] : 
                         (N0)? \nz.mem [1951] : 1'b0;
  assign r_data_o[350] = (N3)? \nz.mem [350] : 
                         (N0)? \nz.mem [1950] : 1'b0;
  assign r_data_o[349] = (N3)? \nz.mem [349] : 
                         (N0)? \nz.mem [1949] : 1'b0;
  assign r_data_o[348] = (N3)? \nz.mem [348] : 
                         (N0)? \nz.mem [1948] : 1'b0;
  assign r_data_o[347] = (N3)? \nz.mem [347] : 
                         (N0)? \nz.mem [1947] : 1'b0;
  assign r_data_o[346] = (N3)? \nz.mem [346] : 
                         (N0)? \nz.mem [1946] : 1'b0;
  assign r_data_o[345] = (N3)? \nz.mem [345] : 
                         (N0)? \nz.mem [1945] : 1'b0;
  assign r_data_o[344] = (N3)? \nz.mem [344] : 
                         (N0)? \nz.mem [1944] : 1'b0;
  assign r_data_o[343] = (N3)? \nz.mem [343] : 
                         (N0)? \nz.mem [1943] : 1'b0;
  assign r_data_o[342] = (N3)? \nz.mem [342] : 
                         (N0)? \nz.mem [1942] : 1'b0;
  assign r_data_o[341] = (N3)? \nz.mem [341] : 
                         (N0)? \nz.mem [1941] : 1'b0;
  assign r_data_o[340] = (N3)? \nz.mem [340] : 
                         (N0)? \nz.mem [1940] : 1'b0;
  assign r_data_o[339] = (N3)? \nz.mem [339] : 
                         (N0)? \nz.mem [1939] : 1'b0;
  assign r_data_o[338] = (N3)? \nz.mem [338] : 
                         (N0)? \nz.mem [1938] : 1'b0;
  assign r_data_o[337] = (N3)? \nz.mem [337] : 
                         (N0)? \nz.mem [1937] : 1'b0;
  assign r_data_o[336] = (N3)? \nz.mem [336] : 
                         (N0)? \nz.mem [1936] : 1'b0;
  assign r_data_o[335] = (N3)? \nz.mem [335] : 
                         (N0)? \nz.mem [1935] : 1'b0;
  assign r_data_o[334] = (N3)? \nz.mem [334] : 
                         (N0)? \nz.mem [1934] : 1'b0;
  assign r_data_o[333] = (N3)? \nz.mem [333] : 
                         (N0)? \nz.mem [1933] : 1'b0;
  assign r_data_o[332] = (N3)? \nz.mem [332] : 
                         (N0)? \nz.mem [1932] : 1'b0;
  assign r_data_o[331] = (N3)? \nz.mem [331] : 
                         (N0)? \nz.mem [1931] : 1'b0;
  assign r_data_o[330] = (N3)? \nz.mem [330] : 
                         (N0)? \nz.mem [1930] : 1'b0;
  assign r_data_o[329] = (N3)? \nz.mem [329] : 
                         (N0)? \nz.mem [1929] : 1'b0;
  assign r_data_o[328] = (N3)? \nz.mem [328] : 
                         (N0)? \nz.mem [1928] : 1'b0;
  assign r_data_o[327] = (N3)? \nz.mem [327] : 
                         (N0)? \nz.mem [1927] : 1'b0;
  assign r_data_o[326] = (N3)? \nz.mem [326] : 
                         (N0)? \nz.mem [1926] : 1'b0;
  assign r_data_o[325] = (N3)? \nz.mem [325] : 
                         (N0)? \nz.mem [1925] : 1'b0;
  assign r_data_o[324] = (N3)? \nz.mem [324] : 
                         (N0)? \nz.mem [1924] : 1'b0;
  assign r_data_o[323] = (N3)? \nz.mem [323] : 
                         (N0)? \nz.mem [1923] : 1'b0;
  assign r_data_o[322] = (N3)? \nz.mem [322] : 
                         (N0)? \nz.mem [1922] : 1'b0;
  assign r_data_o[321] = (N3)? \nz.mem [321] : 
                         (N0)? \nz.mem [1921] : 1'b0;
  assign r_data_o[320] = (N3)? \nz.mem [320] : 
                         (N0)? \nz.mem [1920] : 1'b0;
  assign r_data_o[319] = (N3)? \nz.mem [319] : 
                         (N0)? \nz.mem [1919] : 1'b0;
  assign r_data_o[318] = (N3)? \nz.mem [318] : 
                         (N0)? \nz.mem [1918] : 1'b0;
  assign r_data_o[317] = (N3)? \nz.mem [317] : 
                         (N0)? \nz.mem [1917] : 1'b0;
  assign r_data_o[316] = (N3)? \nz.mem [316] : 
                         (N0)? \nz.mem [1916] : 1'b0;
  assign r_data_o[315] = (N3)? \nz.mem [315] : 
                         (N0)? \nz.mem [1915] : 1'b0;
  assign r_data_o[314] = (N3)? \nz.mem [314] : 
                         (N0)? \nz.mem [1914] : 1'b0;
  assign r_data_o[313] = (N3)? \nz.mem [313] : 
                         (N0)? \nz.mem [1913] : 1'b0;
  assign r_data_o[312] = (N3)? \nz.mem [312] : 
                         (N0)? \nz.mem [1912] : 1'b0;
  assign r_data_o[311] = (N3)? \nz.mem [311] : 
                         (N0)? \nz.mem [1911] : 1'b0;
  assign r_data_o[310] = (N3)? \nz.mem [310] : 
                         (N0)? \nz.mem [1910] : 1'b0;
  assign r_data_o[309] = (N3)? \nz.mem [309] : 
                         (N0)? \nz.mem [1909] : 1'b0;
  assign r_data_o[308] = (N3)? \nz.mem [308] : 
                         (N0)? \nz.mem [1908] : 1'b0;
  assign r_data_o[307] = (N3)? \nz.mem [307] : 
                         (N0)? \nz.mem [1907] : 1'b0;
  assign r_data_o[306] = (N3)? \nz.mem [306] : 
                         (N0)? \nz.mem [1906] : 1'b0;
  assign r_data_o[305] = (N3)? \nz.mem [305] : 
                         (N0)? \nz.mem [1905] : 1'b0;
  assign r_data_o[304] = (N3)? \nz.mem [304] : 
                         (N0)? \nz.mem [1904] : 1'b0;
  assign r_data_o[303] = (N3)? \nz.mem [303] : 
                         (N0)? \nz.mem [1903] : 1'b0;
  assign r_data_o[302] = (N3)? \nz.mem [302] : 
                         (N0)? \nz.mem [1902] : 1'b0;
  assign r_data_o[301] = (N3)? \nz.mem [301] : 
                         (N0)? \nz.mem [1901] : 1'b0;
  assign r_data_o[300] = (N3)? \nz.mem [300] : 
                         (N0)? \nz.mem [1900] : 1'b0;
  assign r_data_o[299] = (N3)? \nz.mem [299] : 
                         (N0)? \nz.mem [1899] : 1'b0;
  assign r_data_o[298] = (N3)? \nz.mem [298] : 
                         (N0)? \nz.mem [1898] : 1'b0;
  assign r_data_o[297] = (N3)? \nz.mem [297] : 
                         (N0)? \nz.mem [1897] : 1'b0;
  assign r_data_o[296] = (N3)? \nz.mem [296] : 
                         (N0)? \nz.mem [1896] : 1'b0;
  assign r_data_o[295] = (N3)? \nz.mem [295] : 
                         (N0)? \nz.mem [1895] : 1'b0;
  assign r_data_o[294] = (N3)? \nz.mem [294] : 
                         (N0)? \nz.mem [1894] : 1'b0;
  assign r_data_o[293] = (N3)? \nz.mem [293] : 
                         (N0)? \nz.mem [1893] : 1'b0;
  assign r_data_o[292] = (N3)? \nz.mem [292] : 
                         (N0)? \nz.mem [1892] : 1'b0;
  assign r_data_o[291] = (N3)? \nz.mem [291] : 
                         (N0)? \nz.mem [1891] : 1'b0;
  assign r_data_o[290] = (N3)? \nz.mem [290] : 
                         (N0)? \nz.mem [1890] : 1'b0;
  assign r_data_o[289] = (N3)? \nz.mem [289] : 
                         (N0)? \nz.mem [1889] : 1'b0;
  assign r_data_o[288] = (N3)? \nz.mem [288] : 
                         (N0)? \nz.mem [1888] : 1'b0;
  assign r_data_o[287] = (N3)? \nz.mem [287] : 
                         (N0)? \nz.mem [1887] : 1'b0;
  assign r_data_o[286] = (N3)? \nz.mem [286] : 
                         (N0)? \nz.mem [1886] : 1'b0;
  assign r_data_o[285] = (N3)? \nz.mem [285] : 
                         (N0)? \nz.mem [1885] : 1'b0;
  assign r_data_o[284] = (N3)? \nz.mem [284] : 
                         (N0)? \nz.mem [1884] : 1'b0;
  assign r_data_o[283] = (N3)? \nz.mem [283] : 
                         (N0)? \nz.mem [1883] : 1'b0;
  assign r_data_o[282] = (N3)? \nz.mem [282] : 
                         (N0)? \nz.mem [1882] : 1'b0;
  assign r_data_o[281] = (N3)? \nz.mem [281] : 
                         (N0)? \nz.mem [1881] : 1'b0;
  assign r_data_o[280] = (N3)? \nz.mem [280] : 
                         (N0)? \nz.mem [1880] : 1'b0;
  assign r_data_o[279] = (N3)? \nz.mem [279] : 
                         (N0)? \nz.mem [1879] : 1'b0;
  assign r_data_o[278] = (N3)? \nz.mem [278] : 
                         (N0)? \nz.mem [1878] : 1'b0;
  assign r_data_o[277] = (N3)? \nz.mem [277] : 
                         (N0)? \nz.mem [1877] : 1'b0;
  assign r_data_o[276] = (N3)? \nz.mem [276] : 
                         (N0)? \nz.mem [1876] : 1'b0;
  assign r_data_o[275] = (N3)? \nz.mem [275] : 
                         (N0)? \nz.mem [1875] : 1'b0;
  assign r_data_o[274] = (N3)? \nz.mem [274] : 
                         (N0)? \nz.mem [1874] : 1'b0;
  assign r_data_o[273] = (N3)? \nz.mem [273] : 
                         (N0)? \nz.mem [1873] : 1'b0;
  assign r_data_o[272] = (N3)? \nz.mem [272] : 
                         (N0)? \nz.mem [1872] : 1'b0;
  assign r_data_o[271] = (N3)? \nz.mem [271] : 
                         (N0)? \nz.mem [1871] : 1'b0;
  assign r_data_o[270] = (N3)? \nz.mem [270] : 
                         (N0)? \nz.mem [1870] : 1'b0;
  assign r_data_o[269] = (N3)? \nz.mem [269] : 
                         (N0)? \nz.mem [1869] : 1'b0;
  assign r_data_o[268] = (N3)? \nz.mem [268] : 
                         (N0)? \nz.mem [1868] : 1'b0;
  assign r_data_o[267] = (N3)? \nz.mem [267] : 
                         (N0)? \nz.mem [1867] : 1'b0;
  assign r_data_o[266] = (N3)? \nz.mem [266] : 
                         (N0)? \nz.mem [1866] : 1'b0;
  assign r_data_o[265] = (N3)? \nz.mem [265] : 
                         (N0)? \nz.mem [1865] : 1'b0;
  assign r_data_o[264] = (N3)? \nz.mem [264] : 
                         (N0)? \nz.mem [1864] : 1'b0;
  assign r_data_o[263] = (N3)? \nz.mem [263] : 
                         (N0)? \nz.mem [1863] : 1'b0;
  assign r_data_o[262] = (N3)? \nz.mem [262] : 
                         (N0)? \nz.mem [1862] : 1'b0;
  assign r_data_o[261] = (N3)? \nz.mem [261] : 
                         (N0)? \nz.mem [1861] : 1'b0;
  assign r_data_o[260] = (N3)? \nz.mem [260] : 
                         (N0)? \nz.mem [1860] : 1'b0;
  assign r_data_o[259] = (N3)? \nz.mem [259] : 
                         (N0)? \nz.mem [1859] : 1'b0;
  assign r_data_o[258] = (N3)? \nz.mem [258] : 
                         (N0)? \nz.mem [1858] : 1'b0;
  assign r_data_o[257] = (N3)? \nz.mem [257] : 
                         (N0)? \nz.mem [1857] : 1'b0;
  assign r_data_o[256] = (N3)? \nz.mem [256] : 
                         (N0)? \nz.mem [1856] : 1'b0;
  assign r_data_o[255] = (N3)? \nz.mem [255] : 
                         (N0)? \nz.mem [1855] : 1'b0;
  assign r_data_o[254] = (N3)? \nz.mem [254] : 
                         (N0)? \nz.mem [1854] : 1'b0;
  assign r_data_o[253] = (N3)? \nz.mem [253] : 
                         (N0)? \nz.mem [1853] : 1'b0;
  assign r_data_o[252] = (N3)? \nz.mem [252] : 
                         (N0)? \nz.mem [1852] : 1'b0;
  assign r_data_o[251] = (N3)? \nz.mem [251] : 
                         (N0)? \nz.mem [1851] : 1'b0;
  assign r_data_o[250] = (N3)? \nz.mem [250] : 
                         (N0)? \nz.mem [1850] : 1'b0;
  assign r_data_o[249] = (N3)? \nz.mem [249] : 
                         (N0)? \nz.mem [1849] : 1'b0;
  assign r_data_o[248] = (N3)? \nz.mem [248] : 
                         (N0)? \nz.mem [1848] : 1'b0;
  assign r_data_o[247] = (N3)? \nz.mem [247] : 
                         (N0)? \nz.mem [1847] : 1'b0;
  assign r_data_o[246] = (N3)? \nz.mem [246] : 
                         (N0)? \nz.mem [1846] : 1'b0;
  assign r_data_o[245] = (N3)? \nz.mem [245] : 
                         (N0)? \nz.mem [1845] : 1'b0;
  assign r_data_o[244] = (N3)? \nz.mem [244] : 
                         (N0)? \nz.mem [1844] : 1'b0;
  assign r_data_o[243] = (N3)? \nz.mem [243] : 
                         (N0)? \nz.mem [1843] : 1'b0;
  assign r_data_o[242] = (N3)? \nz.mem [242] : 
                         (N0)? \nz.mem [1842] : 1'b0;
  assign r_data_o[241] = (N3)? \nz.mem [241] : 
                         (N0)? \nz.mem [1841] : 1'b0;
  assign r_data_o[240] = (N3)? \nz.mem [240] : 
                         (N0)? \nz.mem [1840] : 1'b0;
  assign r_data_o[239] = (N3)? \nz.mem [239] : 
                         (N0)? \nz.mem [1839] : 1'b0;
  assign r_data_o[238] = (N3)? \nz.mem [238] : 
                         (N0)? \nz.mem [1838] : 1'b0;
  assign r_data_o[237] = (N3)? \nz.mem [237] : 
                         (N0)? \nz.mem [1837] : 1'b0;
  assign r_data_o[236] = (N3)? \nz.mem [236] : 
                         (N0)? \nz.mem [1836] : 1'b0;
  assign r_data_o[235] = (N3)? \nz.mem [235] : 
                         (N0)? \nz.mem [1835] : 1'b0;
  assign r_data_o[234] = (N3)? \nz.mem [234] : 
                         (N0)? \nz.mem [1834] : 1'b0;
  assign r_data_o[233] = (N3)? \nz.mem [233] : 
                         (N0)? \nz.mem [1833] : 1'b0;
  assign r_data_o[232] = (N3)? \nz.mem [232] : 
                         (N0)? \nz.mem [1832] : 1'b0;
  assign r_data_o[231] = (N3)? \nz.mem [231] : 
                         (N0)? \nz.mem [1831] : 1'b0;
  assign r_data_o[230] = (N3)? \nz.mem [230] : 
                         (N0)? \nz.mem [1830] : 1'b0;
  assign r_data_o[229] = (N3)? \nz.mem [229] : 
                         (N0)? \nz.mem [1829] : 1'b0;
  assign r_data_o[228] = (N3)? \nz.mem [228] : 
                         (N0)? \nz.mem [1828] : 1'b0;
  assign r_data_o[227] = (N3)? \nz.mem [227] : 
                         (N0)? \nz.mem [1827] : 1'b0;
  assign r_data_o[226] = (N3)? \nz.mem [226] : 
                         (N0)? \nz.mem [1826] : 1'b0;
  assign r_data_o[225] = (N3)? \nz.mem [225] : 
                         (N0)? \nz.mem [1825] : 1'b0;
  assign r_data_o[224] = (N3)? \nz.mem [224] : 
                         (N0)? \nz.mem [1824] : 1'b0;
  assign r_data_o[223] = (N3)? \nz.mem [223] : 
                         (N0)? \nz.mem [1823] : 1'b0;
  assign r_data_o[222] = (N3)? \nz.mem [222] : 
                         (N0)? \nz.mem [1822] : 1'b0;
  assign r_data_o[221] = (N3)? \nz.mem [221] : 
                         (N0)? \nz.mem [1821] : 1'b0;
  assign r_data_o[220] = (N3)? \nz.mem [220] : 
                         (N0)? \nz.mem [1820] : 1'b0;
  assign r_data_o[219] = (N3)? \nz.mem [219] : 
                         (N0)? \nz.mem [1819] : 1'b0;
  assign r_data_o[218] = (N3)? \nz.mem [218] : 
                         (N0)? \nz.mem [1818] : 1'b0;
  assign r_data_o[217] = (N3)? \nz.mem [217] : 
                         (N0)? \nz.mem [1817] : 1'b0;
  assign r_data_o[216] = (N3)? \nz.mem [216] : 
                         (N0)? \nz.mem [1816] : 1'b0;
  assign r_data_o[215] = (N3)? \nz.mem [215] : 
                         (N0)? \nz.mem [1815] : 1'b0;
  assign r_data_o[214] = (N3)? \nz.mem [214] : 
                         (N0)? \nz.mem [1814] : 1'b0;
  assign r_data_o[213] = (N3)? \nz.mem [213] : 
                         (N0)? \nz.mem [1813] : 1'b0;
  assign r_data_o[212] = (N3)? \nz.mem [212] : 
                         (N0)? \nz.mem [1812] : 1'b0;
  assign r_data_o[211] = (N3)? \nz.mem [211] : 
                         (N0)? \nz.mem [1811] : 1'b0;
  assign r_data_o[210] = (N3)? \nz.mem [210] : 
                         (N0)? \nz.mem [1810] : 1'b0;
  assign r_data_o[209] = (N3)? \nz.mem [209] : 
                         (N0)? \nz.mem [1809] : 1'b0;
  assign r_data_o[208] = (N3)? \nz.mem [208] : 
                         (N0)? \nz.mem [1808] : 1'b0;
  assign r_data_o[207] = (N3)? \nz.mem [207] : 
                         (N0)? \nz.mem [1807] : 1'b0;
  assign r_data_o[206] = (N3)? \nz.mem [206] : 
                         (N0)? \nz.mem [1806] : 1'b0;
  assign r_data_o[205] = (N3)? \nz.mem [205] : 
                         (N0)? \nz.mem [1805] : 1'b0;
  assign r_data_o[204] = (N3)? \nz.mem [204] : 
                         (N0)? \nz.mem [1804] : 1'b0;
  assign r_data_o[203] = (N3)? \nz.mem [203] : 
                         (N0)? \nz.mem [1803] : 1'b0;
  assign r_data_o[202] = (N3)? \nz.mem [202] : 
                         (N0)? \nz.mem [1802] : 1'b0;
  assign r_data_o[201] = (N3)? \nz.mem [201] : 
                         (N0)? \nz.mem [1801] : 1'b0;
  assign r_data_o[200] = (N3)? \nz.mem [200] : 
                         (N0)? \nz.mem [1800] : 1'b0;
  assign r_data_o[199] = (N3)? \nz.mem [199] : 
                         (N0)? \nz.mem [1799] : 1'b0;
  assign r_data_o[198] = (N3)? \nz.mem [198] : 
                         (N0)? \nz.mem [1798] : 1'b0;
  assign r_data_o[197] = (N3)? \nz.mem [197] : 
                         (N0)? \nz.mem [1797] : 1'b0;
  assign r_data_o[196] = (N3)? \nz.mem [196] : 
                         (N0)? \nz.mem [1796] : 1'b0;
  assign r_data_o[195] = (N3)? \nz.mem [195] : 
                         (N0)? \nz.mem [1795] : 1'b0;
  assign r_data_o[194] = (N3)? \nz.mem [194] : 
                         (N0)? \nz.mem [1794] : 1'b0;
  assign r_data_o[193] = (N3)? \nz.mem [193] : 
                         (N0)? \nz.mem [1793] : 1'b0;
  assign r_data_o[192] = (N3)? \nz.mem [192] : 
                         (N0)? \nz.mem [1792] : 1'b0;
  assign r_data_o[191] = (N3)? \nz.mem [191] : 
                         (N0)? \nz.mem [1791] : 1'b0;
  assign r_data_o[190] = (N3)? \nz.mem [190] : 
                         (N0)? \nz.mem [1790] : 1'b0;
  assign r_data_o[189] = (N3)? \nz.mem [189] : 
                         (N0)? \nz.mem [1789] : 1'b0;
  assign r_data_o[188] = (N3)? \nz.mem [188] : 
                         (N0)? \nz.mem [1788] : 1'b0;
  assign r_data_o[187] = (N3)? \nz.mem [187] : 
                         (N0)? \nz.mem [1787] : 1'b0;
  assign r_data_o[186] = (N3)? \nz.mem [186] : 
                         (N0)? \nz.mem [1786] : 1'b0;
  assign r_data_o[185] = (N3)? \nz.mem [185] : 
                         (N0)? \nz.mem [1785] : 1'b0;
  assign r_data_o[184] = (N3)? \nz.mem [184] : 
                         (N0)? \nz.mem [1784] : 1'b0;
  assign r_data_o[183] = (N3)? \nz.mem [183] : 
                         (N0)? \nz.mem [1783] : 1'b0;
  assign r_data_o[182] = (N3)? \nz.mem [182] : 
                         (N0)? \nz.mem [1782] : 1'b0;
  assign r_data_o[181] = (N3)? \nz.mem [181] : 
                         (N0)? \nz.mem [1781] : 1'b0;
  assign r_data_o[180] = (N3)? \nz.mem [180] : 
                         (N0)? \nz.mem [1780] : 1'b0;
  assign r_data_o[179] = (N3)? \nz.mem [179] : 
                         (N0)? \nz.mem [1779] : 1'b0;
  assign r_data_o[178] = (N3)? \nz.mem [178] : 
                         (N0)? \nz.mem [1778] : 1'b0;
  assign r_data_o[177] = (N3)? \nz.mem [177] : 
                         (N0)? \nz.mem [1777] : 1'b0;
  assign r_data_o[176] = (N3)? \nz.mem [176] : 
                         (N0)? \nz.mem [1776] : 1'b0;
  assign r_data_o[175] = (N3)? \nz.mem [175] : 
                         (N0)? \nz.mem [1775] : 1'b0;
  assign r_data_o[174] = (N3)? \nz.mem [174] : 
                         (N0)? \nz.mem [1774] : 1'b0;
  assign r_data_o[173] = (N3)? \nz.mem [173] : 
                         (N0)? \nz.mem [1773] : 1'b0;
  assign r_data_o[172] = (N3)? \nz.mem [172] : 
                         (N0)? \nz.mem [1772] : 1'b0;
  assign r_data_o[171] = (N3)? \nz.mem [171] : 
                         (N0)? \nz.mem [1771] : 1'b0;
  assign r_data_o[170] = (N3)? \nz.mem [170] : 
                         (N0)? \nz.mem [1770] : 1'b0;
  assign r_data_o[169] = (N3)? \nz.mem [169] : 
                         (N0)? \nz.mem [1769] : 1'b0;
  assign r_data_o[168] = (N3)? \nz.mem [168] : 
                         (N0)? \nz.mem [1768] : 1'b0;
  assign r_data_o[167] = (N3)? \nz.mem [167] : 
                         (N0)? \nz.mem [1767] : 1'b0;
  assign r_data_o[166] = (N3)? \nz.mem [166] : 
                         (N0)? \nz.mem [1766] : 1'b0;
  assign r_data_o[165] = (N3)? \nz.mem [165] : 
                         (N0)? \nz.mem [1765] : 1'b0;
  assign r_data_o[164] = (N3)? \nz.mem [164] : 
                         (N0)? \nz.mem [1764] : 1'b0;
  assign r_data_o[163] = (N3)? \nz.mem [163] : 
                         (N0)? \nz.mem [1763] : 1'b0;
  assign r_data_o[162] = (N3)? \nz.mem [162] : 
                         (N0)? \nz.mem [1762] : 1'b0;
  assign r_data_o[161] = (N3)? \nz.mem [161] : 
                         (N0)? \nz.mem [1761] : 1'b0;
  assign r_data_o[160] = (N3)? \nz.mem [160] : 
                         (N0)? \nz.mem [1760] : 1'b0;
  assign r_data_o[159] = (N3)? \nz.mem [159] : 
                         (N0)? \nz.mem [1759] : 1'b0;
  assign r_data_o[158] = (N3)? \nz.mem [158] : 
                         (N0)? \nz.mem [1758] : 1'b0;
  assign r_data_o[157] = (N3)? \nz.mem [157] : 
                         (N0)? \nz.mem [1757] : 1'b0;
  assign r_data_o[156] = (N3)? \nz.mem [156] : 
                         (N0)? \nz.mem [1756] : 1'b0;
  assign r_data_o[155] = (N3)? \nz.mem [155] : 
                         (N0)? \nz.mem [1755] : 1'b0;
  assign r_data_o[154] = (N3)? \nz.mem [154] : 
                         (N0)? \nz.mem [1754] : 1'b0;
  assign r_data_o[153] = (N3)? \nz.mem [153] : 
                         (N0)? \nz.mem [1753] : 1'b0;
  assign r_data_o[152] = (N3)? \nz.mem [152] : 
                         (N0)? \nz.mem [1752] : 1'b0;
  assign r_data_o[151] = (N3)? \nz.mem [151] : 
                         (N0)? \nz.mem [1751] : 1'b0;
  assign r_data_o[150] = (N3)? \nz.mem [150] : 
                         (N0)? \nz.mem [1750] : 1'b0;
  assign r_data_o[149] = (N3)? \nz.mem [149] : 
                         (N0)? \nz.mem [1749] : 1'b0;
  assign r_data_o[148] = (N3)? \nz.mem [148] : 
                         (N0)? \nz.mem [1748] : 1'b0;
  assign r_data_o[147] = (N3)? \nz.mem [147] : 
                         (N0)? \nz.mem [1747] : 1'b0;
  assign r_data_o[146] = (N3)? \nz.mem [146] : 
                         (N0)? \nz.mem [1746] : 1'b0;
  assign r_data_o[145] = (N3)? \nz.mem [145] : 
                         (N0)? \nz.mem [1745] : 1'b0;
  assign r_data_o[144] = (N3)? \nz.mem [144] : 
                         (N0)? \nz.mem [1744] : 1'b0;
  assign r_data_o[143] = (N3)? \nz.mem [143] : 
                         (N0)? \nz.mem [1743] : 1'b0;
  assign r_data_o[142] = (N3)? \nz.mem [142] : 
                         (N0)? \nz.mem [1742] : 1'b0;
  assign r_data_o[141] = (N3)? \nz.mem [141] : 
                         (N0)? \nz.mem [1741] : 1'b0;
  assign r_data_o[140] = (N3)? \nz.mem [140] : 
                         (N0)? \nz.mem [1740] : 1'b0;
  assign r_data_o[139] = (N3)? \nz.mem [139] : 
                         (N0)? \nz.mem [1739] : 1'b0;
  assign r_data_o[138] = (N3)? \nz.mem [138] : 
                         (N0)? \nz.mem [1738] : 1'b0;
  assign r_data_o[137] = (N3)? \nz.mem [137] : 
                         (N0)? \nz.mem [1737] : 1'b0;
  assign r_data_o[136] = (N3)? \nz.mem [136] : 
                         (N0)? \nz.mem [1736] : 1'b0;
  assign r_data_o[135] = (N3)? \nz.mem [135] : 
                         (N0)? \nz.mem [1735] : 1'b0;
  assign r_data_o[134] = (N3)? \nz.mem [134] : 
                         (N0)? \nz.mem [1734] : 1'b0;
  assign r_data_o[133] = (N3)? \nz.mem [133] : 
                         (N0)? \nz.mem [1733] : 1'b0;
  assign r_data_o[132] = (N3)? \nz.mem [132] : 
                         (N0)? \nz.mem [1732] : 1'b0;
  assign r_data_o[131] = (N3)? \nz.mem [131] : 
                         (N0)? \nz.mem [1731] : 1'b0;
  assign r_data_o[130] = (N3)? \nz.mem [130] : 
                         (N0)? \nz.mem [1730] : 1'b0;
  assign r_data_o[129] = (N3)? \nz.mem [129] : 
                         (N0)? \nz.mem [1729] : 1'b0;
  assign r_data_o[128] = (N3)? \nz.mem [128] : 
                         (N0)? \nz.mem [1728] : 1'b0;
  assign r_data_o[127] = (N3)? \nz.mem [127] : 
                         (N0)? \nz.mem [1727] : 1'b0;
  assign r_data_o[126] = (N3)? \nz.mem [126] : 
                         (N0)? \nz.mem [1726] : 1'b0;
  assign r_data_o[125] = (N3)? \nz.mem [125] : 
                         (N0)? \nz.mem [1725] : 1'b0;
  assign r_data_o[124] = (N3)? \nz.mem [124] : 
                         (N0)? \nz.mem [1724] : 1'b0;
  assign r_data_o[123] = (N3)? \nz.mem [123] : 
                         (N0)? \nz.mem [1723] : 1'b0;
  assign r_data_o[122] = (N3)? \nz.mem [122] : 
                         (N0)? \nz.mem [1722] : 1'b0;
  assign r_data_o[121] = (N3)? \nz.mem [121] : 
                         (N0)? \nz.mem [1721] : 1'b0;
  assign r_data_o[120] = (N3)? \nz.mem [120] : 
                         (N0)? \nz.mem [1720] : 1'b0;
  assign r_data_o[119] = (N3)? \nz.mem [119] : 
                         (N0)? \nz.mem [1719] : 1'b0;
  assign r_data_o[118] = (N3)? \nz.mem [118] : 
                         (N0)? \nz.mem [1718] : 1'b0;
  assign r_data_o[117] = (N3)? \nz.mem [117] : 
                         (N0)? \nz.mem [1717] : 1'b0;
  assign r_data_o[116] = (N3)? \nz.mem [116] : 
                         (N0)? \nz.mem [1716] : 1'b0;
  assign r_data_o[115] = (N3)? \nz.mem [115] : 
                         (N0)? \nz.mem [1715] : 1'b0;
  assign r_data_o[114] = (N3)? \nz.mem [114] : 
                         (N0)? \nz.mem [1714] : 1'b0;
  assign r_data_o[113] = (N3)? \nz.mem [113] : 
                         (N0)? \nz.mem [1713] : 1'b0;
  assign r_data_o[112] = (N3)? \nz.mem [112] : 
                         (N0)? \nz.mem [1712] : 1'b0;
  assign r_data_o[111] = (N3)? \nz.mem [111] : 
                         (N0)? \nz.mem [1711] : 1'b0;
  assign r_data_o[110] = (N3)? \nz.mem [110] : 
                         (N0)? \nz.mem [1710] : 1'b0;
  assign r_data_o[109] = (N3)? \nz.mem [109] : 
                         (N0)? \nz.mem [1709] : 1'b0;
  assign r_data_o[108] = (N3)? \nz.mem [108] : 
                         (N0)? \nz.mem [1708] : 1'b0;
  assign r_data_o[107] = (N3)? \nz.mem [107] : 
                         (N0)? \nz.mem [1707] : 1'b0;
  assign r_data_o[106] = (N3)? \nz.mem [106] : 
                         (N0)? \nz.mem [1706] : 1'b0;
  assign r_data_o[105] = (N3)? \nz.mem [105] : 
                         (N0)? \nz.mem [1705] : 1'b0;
  assign r_data_o[104] = (N3)? \nz.mem [104] : 
                         (N0)? \nz.mem [1704] : 1'b0;
  assign r_data_o[103] = (N3)? \nz.mem [103] : 
                         (N0)? \nz.mem [1703] : 1'b0;
  assign r_data_o[102] = (N3)? \nz.mem [102] : 
                         (N0)? \nz.mem [1702] : 1'b0;
  assign r_data_o[101] = (N3)? \nz.mem [101] : 
                         (N0)? \nz.mem [1701] : 1'b0;
  assign r_data_o[100] = (N3)? \nz.mem [100] : 
                         (N0)? \nz.mem [1700] : 1'b0;
  assign r_data_o[99] = (N3)? \nz.mem [99] : 
                        (N0)? \nz.mem [1699] : 1'b0;
  assign r_data_o[98] = (N3)? \nz.mem [98] : 
                        (N0)? \nz.mem [1698] : 1'b0;
  assign r_data_o[97] = (N3)? \nz.mem [97] : 
                        (N0)? \nz.mem [1697] : 1'b0;
  assign r_data_o[96] = (N3)? \nz.mem [96] : 
                        (N0)? \nz.mem [1696] : 1'b0;
  assign r_data_o[95] = (N3)? \nz.mem [95] : 
                        (N0)? \nz.mem [1695] : 1'b0;
  assign r_data_o[94] = (N3)? \nz.mem [94] : 
                        (N0)? \nz.mem [1694] : 1'b0;
  assign r_data_o[93] = (N3)? \nz.mem [93] : 
                        (N0)? \nz.mem [1693] : 1'b0;
  assign r_data_o[92] = (N3)? \nz.mem [92] : 
                        (N0)? \nz.mem [1692] : 1'b0;
  assign r_data_o[91] = (N3)? \nz.mem [91] : 
                        (N0)? \nz.mem [1691] : 1'b0;
  assign r_data_o[90] = (N3)? \nz.mem [90] : 
                        (N0)? \nz.mem [1690] : 1'b0;
  assign r_data_o[89] = (N3)? \nz.mem [89] : 
                        (N0)? \nz.mem [1689] : 1'b0;
  assign r_data_o[88] = (N3)? \nz.mem [88] : 
                        (N0)? \nz.mem [1688] : 1'b0;
  assign r_data_o[87] = (N3)? \nz.mem [87] : 
                        (N0)? \nz.mem [1687] : 1'b0;
  assign r_data_o[86] = (N3)? \nz.mem [86] : 
                        (N0)? \nz.mem [1686] : 1'b0;
  assign r_data_o[85] = (N3)? \nz.mem [85] : 
                        (N0)? \nz.mem [1685] : 1'b0;
  assign r_data_o[84] = (N3)? \nz.mem [84] : 
                        (N0)? \nz.mem [1684] : 1'b0;
  assign r_data_o[83] = (N3)? \nz.mem [83] : 
                        (N0)? \nz.mem [1683] : 1'b0;
  assign r_data_o[82] = (N3)? \nz.mem [82] : 
                        (N0)? \nz.mem [1682] : 1'b0;
  assign r_data_o[81] = (N3)? \nz.mem [81] : 
                        (N0)? \nz.mem [1681] : 1'b0;
  assign r_data_o[80] = (N3)? \nz.mem [80] : 
                        (N0)? \nz.mem [1680] : 1'b0;
  assign r_data_o[79] = (N3)? \nz.mem [79] : 
                        (N0)? \nz.mem [1679] : 1'b0;
  assign r_data_o[78] = (N3)? \nz.mem [78] : 
                        (N0)? \nz.mem [1678] : 1'b0;
  assign r_data_o[77] = (N3)? \nz.mem [77] : 
                        (N0)? \nz.mem [1677] : 1'b0;
  assign r_data_o[76] = (N3)? \nz.mem [76] : 
                        (N0)? \nz.mem [1676] : 1'b0;
  assign r_data_o[75] = (N3)? \nz.mem [75] : 
                        (N0)? \nz.mem [1675] : 1'b0;
  assign r_data_o[74] = (N3)? \nz.mem [74] : 
                        (N0)? \nz.mem [1674] : 1'b0;
  assign r_data_o[73] = (N3)? \nz.mem [73] : 
                        (N0)? \nz.mem [1673] : 1'b0;
  assign r_data_o[72] = (N3)? \nz.mem [72] : 
                        (N0)? \nz.mem [1672] : 1'b0;
  assign r_data_o[71] = (N3)? \nz.mem [71] : 
                        (N0)? \nz.mem [1671] : 1'b0;
  assign r_data_o[70] = (N3)? \nz.mem [70] : 
                        (N0)? \nz.mem [1670] : 1'b0;
  assign r_data_o[69] = (N3)? \nz.mem [69] : 
                        (N0)? \nz.mem [1669] : 1'b0;
  assign r_data_o[68] = (N3)? \nz.mem [68] : 
                        (N0)? \nz.mem [1668] : 1'b0;
  assign r_data_o[67] = (N3)? \nz.mem [67] : 
                        (N0)? \nz.mem [1667] : 1'b0;
  assign r_data_o[66] = (N3)? \nz.mem [66] : 
                        (N0)? \nz.mem [1666] : 1'b0;
  assign r_data_o[65] = (N3)? \nz.mem [65] : 
                        (N0)? \nz.mem [1665] : 1'b0;
  assign r_data_o[64] = (N3)? \nz.mem [64] : 
                        (N0)? \nz.mem [1664] : 1'b0;
  assign r_data_o[63] = (N3)? \nz.mem [63] : 
                        (N0)? \nz.mem [1663] : 1'b0;
  assign r_data_o[62] = (N3)? \nz.mem [62] : 
                        (N0)? \nz.mem [1662] : 1'b0;
  assign r_data_o[61] = (N3)? \nz.mem [61] : 
                        (N0)? \nz.mem [1661] : 1'b0;
  assign r_data_o[60] = (N3)? \nz.mem [60] : 
                        (N0)? \nz.mem [1660] : 1'b0;
  assign r_data_o[59] = (N3)? \nz.mem [59] : 
                        (N0)? \nz.mem [1659] : 1'b0;
  assign r_data_o[58] = (N3)? \nz.mem [58] : 
                        (N0)? \nz.mem [1658] : 1'b0;
  assign r_data_o[57] = (N3)? \nz.mem [57] : 
                        (N0)? \nz.mem [1657] : 1'b0;
  assign r_data_o[56] = (N3)? \nz.mem [56] : 
                        (N0)? \nz.mem [1656] : 1'b0;
  assign r_data_o[55] = (N3)? \nz.mem [55] : 
                        (N0)? \nz.mem [1655] : 1'b0;
  assign r_data_o[54] = (N3)? \nz.mem [54] : 
                        (N0)? \nz.mem [1654] : 1'b0;
  assign r_data_o[53] = (N3)? \nz.mem [53] : 
                        (N0)? \nz.mem [1653] : 1'b0;
  assign r_data_o[52] = (N3)? \nz.mem [52] : 
                        (N0)? \nz.mem [1652] : 1'b0;
  assign r_data_o[51] = (N3)? \nz.mem [51] : 
                        (N0)? \nz.mem [1651] : 1'b0;
  assign r_data_o[50] = (N3)? \nz.mem [50] : 
                        (N0)? \nz.mem [1650] : 1'b0;
  assign r_data_o[49] = (N3)? \nz.mem [49] : 
                        (N0)? \nz.mem [1649] : 1'b0;
  assign r_data_o[48] = (N3)? \nz.mem [48] : 
                        (N0)? \nz.mem [1648] : 1'b0;
  assign r_data_o[47] = (N3)? \nz.mem [47] : 
                        (N0)? \nz.mem [1647] : 1'b0;
  assign r_data_o[46] = (N3)? \nz.mem [46] : 
                        (N0)? \nz.mem [1646] : 1'b0;
  assign r_data_o[45] = (N3)? \nz.mem [45] : 
                        (N0)? \nz.mem [1645] : 1'b0;
  assign r_data_o[44] = (N3)? \nz.mem [44] : 
                        (N0)? \nz.mem [1644] : 1'b0;
  assign r_data_o[43] = (N3)? \nz.mem [43] : 
                        (N0)? \nz.mem [1643] : 1'b0;
  assign r_data_o[42] = (N3)? \nz.mem [42] : 
                        (N0)? \nz.mem [1642] : 1'b0;
  assign r_data_o[41] = (N3)? \nz.mem [41] : 
                        (N0)? \nz.mem [1641] : 1'b0;
  assign r_data_o[40] = (N3)? \nz.mem [40] : 
                        (N0)? \nz.mem [1640] : 1'b0;
  assign r_data_o[39] = (N3)? \nz.mem [39] : 
                        (N0)? \nz.mem [1639] : 1'b0;
  assign r_data_o[38] = (N3)? \nz.mem [38] : 
                        (N0)? \nz.mem [1638] : 1'b0;
  assign r_data_o[37] = (N3)? \nz.mem [37] : 
                        (N0)? \nz.mem [1637] : 1'b0;
  assign r_data_o[36] = (N3)? \nz.mem [36] : 
                        (N0)? \nz.mem [1636] : 1'b0;
  assign r_data_o[35] = (N3)? \nz.mem [35] : 
                        (N0)? \nz.mem [1635] : 1'b0;
  assign r_data_o[34] = (N3)? \nz.mem [34] : 
                        (N0)? \nz.mem [1634] : 1'b0;
  assign r_data_o[33] = (N3)? \nz.mem [33] : 
                        (N0)? \nz.mem [1633] : 1'b0;
  assign r_data_o[32] = (N3)? \nz.mem [32] : 
                        (N0)? \nz.mem [1632] : 1'b0;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [1631] : 1'b0;
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [1630] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [1629] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [1628] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [1627] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [1626] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [1625] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [1624] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [1623] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [1622] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [1621] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [1620] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [1619] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [1618] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [1617] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [1616] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [1615] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [1614] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [1613] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [1612] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [1611] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [1610] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [1609] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [1608] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [1607] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [1606] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [1605] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [1604] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [1603] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [1602] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [1601] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [1600] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5 } : 
                                                                                                                                                                           (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N23) begin
      \nz.mem_3199_sv2v_reg  <= w_data_i[1599];
      \nz.mem_3198_sv2v_reg  <= w_data_i[1598];
      \nz.mem_3197_sv2v_reg  <= w_data_i[1597];
      \nz.mem_3196_sv2v_reg  <= w_data_i[1596];
      \nz.mem_3195_sv2v_reg  <= w_data_i[1595];
      \nz.mem_3194_sv2v_reg  <= w_data_i[1594];
      \nz.mem_3193_sv2v_reg  <= w_data_i[1593];
      \nz.mem_3192_sv2v_reg  <= w_data_i[1592];
      \nz.mem_3191_sv2v_reg  <= w_data_i[1591];
      \nz.mem_3190_sv2v_reg  <= w_data_i[1590];
      \nz.mem_3189_sv2v_reg  <= w_data_i[1589];
      \nz.mem_3188_sv2v_reg  <= w_data_i[1588];
      \nz.mem_3187_sv2v_reg  <= w_data_i[1587];
      \nz.mem_3186_sv2v_reg  <= w_data_i[1586];
      \nz.mem_3185_sv2v_reg  <= w_data_i[1585];
      \nz.mem_3184_sv2v_reg  <= w_data_i[1584];
      \nz.mem_3183_sv2v_reg  <= w_data_i[1583];
      \nz.mem_3182_sv2v_reg  <= w_data_i[1582];
      \nz.mem_3181_sv2v_reg  <= w_data_i[1581];
      \nz.mem_3180_sv2v_reg  <= w_data_i[1580];
      \nz.mem_3179_sv2v_reg  <= w_data_i[1579];
      \nz.mem_3178_sv2v_reg  <= w_data_i[1578];
      \nz.mem_3177_sv2v_reg  <= w_data_i[1577];
      \nz.mem_3176_sv2v_reg  <= w_data_i[1576];
      \nz.mem_3175_sv2v_reg  <= w_data_i[1575];
      \nz.mem_3174_sv2v_reg  <= w_data_i[1574];
      \nz.mem_3173_sv2v_reg  <= w_data_i[1573];
      \nz.mem_3172_sv2v_reg  <= w_data_i[1572];
      \nz.mem_3171_sv2v_reg  <= w_data_i[1571];
      \nz.mem_3170_sv2v_reg  <= w_data_i[1570];
      \nz.mem_3169_sv2v_reg  <= w_data_i[1569];
      \nz.mem_3168_sv2v_reg  <= w_data_i[1568];
      \nz.mem_3167_sv2v_reg  <= w_data_i[1567];
      \nz.mem_3166_sv2v_reg  <= w_data_i[1566];
      \nz.mem_3165_sv2v_reg  <= w_data_i[1565];
      \nz.mem_3164_sv2v_reg  <= w_data_i[1564];
      \nz.mem_3163_sv2v_reg  <= w_data_i[1563];
      \nz.mem_3162_sv2v_reg  <= w_data_i[1562];
      \nz.mem_3161_sv2v_reg  <= w_data_i[1561];
      \nz.mem_3160_sv2v_reg  <= w_data_i[1560];
      \nz.mem_3159_sv2v_reg  <= w_data_i[1559];
      \nz.mem_3158_sv2v_reg  <= w_data_i[1558];
      \nz.mem_3157_sv2v_reg  <= w_data_i[1557];
      \nz.mem_3156_sv2v_reg  <= w_data_i[1556];
      \nz.mem_3155_sv2v_reg  <= w_data_i[1555];
      \nz.mem_3154_sv2v_reg  <= w_data_i[1554];
      \nz.mem_3153_sv2v_reg  <= w_data_i[1553];
      \nz.mem_3152_sv2v_reg  <= w_data_i[1552];
      \nz.mem_3151_sv2v_reg  <= w_data_i[1551];
      \nz.mem_3150_sv2v_reg  <= w_data_i[1550];
      \nz.mem_3149_sv2v_reg  <= w_data_i[1549];
      \nz.mem_3148_sv2v_reg  <= w_data_i[1548];
      \nz.mem_3147_sv2v_reg  <= w_data_i[1547];
      \nz.mem_3146_sv2v_reg  <= w_data_i[1546];
      \nz.mem_3145_sv2v_reg  <= w_data_i[1545];
      \nz.mem_3144_sv2v_reg  <= w_data_i[1544];
      \nz.mem_3143_sv2v_reg  <= w_data_i[1543];
      \nz.mem_3142_sv2v_reg  <= w_data_i[1542];
      \nz.mem_3141_sv2v_reg  <= w_data_i[1541];
      \nz.mem_3140_sv2v_reg  <= w_data_i[1540];
      \nz.mem_3139_sv2v_reg  <= w_data_i[1539];
      \nz.mem_3138_sv2v_reg  <= w_data_i[1538];
      \nz.mem_3137_sv2v_reg  <= w_data_i[1537];
      \nz.mem_3136_sv2v_reg  <= w_data_i[1536];
      \nz.mem_3135_sv2v_reg  <= w_data_i[1535];
      \nz.mem_3134_sv2v_reg  <= w_data_i[1534];
      \nz.mem_3133_sv2v_reg  <= w_data_i[1533];
      \nz.mem_3132_sv2v_reg  <= w_data_i[1532];
      \nz.mem_3131_sv2v_reg  <= w_data_i[1531];
      \nz.mem_3130_sv2v_reg  <= w_data_i[1530];
      \nz.mem_3129_sv2v_reg  <= w_data_i[1529];
      \nz.mem_3128_sv2v_reg  <= w_data_i[1528];
      \nz.mem_3127_sv2v_reg  <= w_data_i[1527];
      \nz.mem_3126_sv2v_reg  <= w_data_i[1526];
      \nz.mem_3125_sv2v_reg  <= w_data_i[1525];
      \nz.mem_3124_sv2v_reg  <= w_data_i[1524];
      \nz.mem_3123_sv2v_reg  <= w_data_i[1523];
      \nz.mem_3122_sv2v_reg  <= w_data_i[1522];
      \nz.mem_3121_sv2v_reg  <= w_data_i[1521];
      \nz.mem_3120_sv2v_reg  <= w_data_i[1520];
      \nz.mem_3119_sv2v_reg  <= w_data_i[1519];
      \nz.mem_3118_sv2v_reg  <= w_data_i[1518];
      \nz.mem_3117_sv2v_reg  <= w_data_i[1517];
      \nz.mem_3116_sv2v_reg  <= w_data_i[1516];
      \nz.mem_3115_sv2v_reg  <= w_data_i[1515];
      \nz.mem_3114_sv2v_reg  <= w_data_i[1514];
      \nz.mem_3113_sv2v_reg  <= w_data_i[1513];
      \nz.mem_3112_sv2v_reg  <= w_data_i[1512];
      \nz.mem_3111_sv2v_reg  <= w_data_i[1511];
      \nz.mem_3110_sv2v_reg  <= w_data_i[1510];
      \nz.mem_3109_sv2v_reg  <= w_data_i[1509];
      \nz.mem_3108_sv2v_reg  <= w_data_i[1508];
      \nz.mem_3107_sv2v_reg  <= w_data_i[1507];
      \nz.mem_3106_sv2v_reg  <= w_data_i[1506];
      \nz.mem_3105_sv2v_reg  <= w_data_i[1505];
      \nz.mem_3104_sv2v_reg  <= w_data_i[1504];
      \nz.mem_3103_sv2v_reg  <= w_data_i[1503];
      \nz.mem_3102_sv2v_reg  <= w_data_i[1502];
      \nz.mem_3101_sv2v_reg  <= w_data_i[1501];
      \nz.mem_1600_sv2v_reg  <= w_data_i[0];
    end 
    if(N24) begin
      \nz.mem_3100_sv2v_reg  <= w_data_i[1500];
      \nz.mem_3099_sv2v_reg  <= w_data_i[1499];
      \nz.mem_3098_sv2v_reg  <= w_data_i[1498];
      \nz.mem_3097_sv2v_reg  <= w_data_i[1497];
      \nz.mem_3096_sv2v_reg  <= w_data_i[1496];
      \nz.mem_3095_sv2v_reg  <= w_data_i[1495];
      \nz.mem_3094_sv2v_reg  <= w_data_i[1494];
      \nz.mem_3093_sv2v_reg  <= w_data_i[1493];
      \nz.mem_3092_sv2v_reg  <= w_data_i[1492];
      \nz.mem_3091_sv2v_reg  <= w_data_i[1491];
      \nz.mem_3090_sv2v_reg  <= w_data_i[1490];
      \nz.mem_3089_sv2v_reg  <= w_data_i[1489];
      \nz.mem_3088_sv2v_reg  <= w_data_i[1488];
      \nz.mem_3087_sv2v_reg  <= w_data_i[1487];
      \nz.mem_3086_sv2v_reg  <= w_data_i[1486];
      \nz.mem_3085_sv2v_reg  <= w_data_i[1485];
      \nz.mem_3084_sv2v_reg  <= w_data_i[1484];
      \nz.mem_3083_sv2v_reg  <= w_data_i[1483];
      \nz.mem_3082_sv2v_reg  <= w_data_i[1482];
      \nz.mem_3081_sv2v_reg  <= w_data_i[1481];
      \nz.mem_3080_sv2v_reg  <= w_data_i[1480];
      \nz.mem_3079_sv2v_reg  <= w_data_i[1479];
      \nz.mem_3078_sv2v_reg  <= w_data_i[1478];
      \nz.mem_3077_sv2v_reg  <= w_data_i[1477];
      \nz.mem_3076_sv2v_reg  <= w_data_i[1476];
      \nz.mem_3075_sv2v_reg  <= w_data_i[1475];
      \nz.mem_3074_sv2v_reg  <= w_data_i[1474];
      \nz.mem_3073_sv2v_reg  <= w_data_i[1473];
      \nz.mem_3072_sv2v_reg  <= w_data_i[1472];
      \nz.mem_3071_sv2v_reg  <= w_data_i[1471];
      \nz.mem_3070_sv2v_reg  <= w_data_i[1470];
      \nz.mem_3069_sv2v_reg  <= w_data_i[1469];
      \nz.mem_3068_sv2v_reg  <= w_data_i[1468];
      \nz.mem_3067_sv2v_reg  <= w_data_i[1467];
      \nz.mem_3066_sv2v_reg  <= w_data_i[1466];
      \nz.mem_3065_sv2v_reg  <= w_data_i[1465];
      \nz.mem_3064_sv2v_reg  <= w_data_i[1464];
      \nz.mem_3063_sv2v_reg  <= w_data_i[1463];
      \nz.mem_3062_sv2v_reg  <= w_data_i[1462];
      \nz.mem_3061_sv2v_reg  <= w_data_i[1461];
      \nz.mem_3060_sv2v_reg  <= w_data_i[1460];
      \nz.mem_3059_sv2v_reg  <= w_data_i[1459];
      \nz.mem_3058_sv2v_reg  <= w_data_i[1458];
      \nz.mem_3057_sv2v_reg  <= w_data_i[1457];
      \nz.mem_3056_sv2v_reg  <= w_data_i[1456];
      \nz.mem_3055_sv2v_reg  <= w_data_i[1455];
      \nz.mem_3054_sv2v_reg  <= w_data_i[1454];
      \nz.mem_3053_sv2v_reg  <= w_data_i[1453];
      \nz.mem_3052_sv2v_reg  <= w_data_i[1452];
      \nz.mem_3051_sv2v_reg  <= w_data_i[1451];
      \nz.mem_3050_sv2v_reg  <= w_data_i[1450];
      \nz.mem_3049_sv2v_reg  <= w_data_i[1449];
      \nz.mem_3048_sv2v_reg  <= w_data_i[1448];
      \nz.mem_3047_sv2v_reg  <= w_data_i[1447];
      \nz.mem_3046_sv2v_reg  <= w_data_i[1446];
      \nz.mem_3045_sv2v_reg  <= w_data_i[1445];
      \nz.mem_3044_sv2v_reg  <= w_data_i[1444];
      \nz.mem_3043_sv2v_reg  <= w_data_i[1443];
      \nz.mem_3042_sv2v_reg  <= w_data_i[1442];
      \nz.mem_3041_sv2v_reg  <= w_data_i[1441];
      \nz.mem_3040_sv2v_reg  <= w_data_i[1440];
      \nz.mem_3039_sv2v_reg  <= w_data_i[1439];
      \nz.mem_3038_sv2v_reg  <= w_data_i[1438];
      \nz.mem_3037_sv2v_reg  <= w_data_i[1437];
      \nz.mem_3036_sv2v_reg  <= w_data_i[1436];
      \nz.mem_3035_sv2v_reg  <= w_data_i[1435];
      \nz.mem_3034_sv2v_reg  <= w_data_i[1434];
      \nz.mem_3033_sv2v_reg  <= w_data_i[1433];
      \nz.mem_3032_sv2v_reg  <= w_data_i[1432];
      \nz.mem_3031_sv2v_reg  <= w_data_i[1431];
      \nz.mem_3030_sv2v_reg  <= w_data_i[1430];
      \nz.mem_3029_sv2v_reg  <= w_data_i[1429];
      \nz.mem_3028_sv2v_reg  <= w_data_i[1428];
      \nz.mem_3027_sv2v_reg  <= w_data_i[1427];
      \nz.mem_3026_sv2v_reg  <= w_data_i[1426];
      \nz.mem_3025_sv2v_reg  <= w_data_i[1425];
      \nz.mem_3024_sv2v_reg  <= w_data_i[1424];
      \nz.mem_3023_sv2v_reg  <= w_data_i[1423];
      \nz.mem_3022_sv2v_reg  <= w_data_i[1422];
      \nz.mem_3021_sv2v_reg  <= w_data_i[1421];
      \nz.mem_3020_sv2v_reg  <= w_data_i[1420];
      \nz.mem_3019_sv2v_reg  <= w_data_i[1419];
      \nz.mem_3018_sv2v_reg  <= w_data_i[1418];
      \nz.mem_3017_sv2v_reg  <= w_data_i[1417];
      \nz.mem_3016_sv2v_reg  <= w_data_i[1416];
      \nz.mem_3015_sv2v_reg  <= w_data_i[1415];
      \nz.mem_3014_sv2v_reg  <= w_data_i[1414];
      \nz.mem_3013_sv2v_reg  <= w_data_i[1413];
      \nz.mem_3012_sv2v_reg  <= w_data_i[1412];
      \nz.mem_3011_sv2v_reg  <= w_data_i[1411];
      \nz.mem_3010_sv2v_reg  <= w_data_i[1410];
      \nz.mem_3009_sv2v_reg  <= w_data_i[1409];
      \nz.mem_3008_sv2v_reg  <= w_data_i[1408];
      \nz.mem_3007_sv2v_reg  <= w_data_i[1407];
      \nz.mem_3006_sv2v_reg  <= w_data_i[1406];
      \nz.mem_3005_sv2v_reg  <= w_data_i[1405];
      \nz.mem_3004_sv2v_reg  <= w_data_i[1404];
      \nz.mem_3003_sv2v_reg  <= w_data_i[1403];
      \nz.mem_3002_sv2v_reg  <= w_data_i[1402];
      \nz.mem_1601_sv2v_reg  <= w_data_i[1];
    end 
    if(N25) begin
      \nz.mem_3001_sv2v_reg  <= w_data_i[1401];
      \nz.mem_3000_sv2v_reg  <= w_data_i[1400];
      \nz.mem_2999_sv2v_reg  <= w_data_i[1399];
      \nz.mem_2998_sv2v_reg  <= w_data_i[1398];
      \nz.mem_2997_sv2v_reg  <= w_data_i[1397];
      \nz.mem_2996_sv2v_reg  <= w_data_i[1396];
      \nz.mem_2995_sv2v_reg  <= w_data_i[1395];
      \nz.mem_2994_sv2v_reg  <= w_data_i[1394];
      \nz.mem_2993_sv2v_reg  <= w_data_i[1393];
      \nz.mem_2992_sv2v_reg  <= w_data_i[1392];
      \nz.mem_2991_sv2v_reg  <= w_data_i[1391];
      \nz.mem_2990_sv2v_reg  <= w_data_i[1390];
      \nz.mem_2989_sv2v_reg  <= w_data_i[1389];
      \nz.mem_2988_sv2v_reg  <= w_data_i[1388];
      \nz.mem_2987_sv2v_reg  <= w_data_i[1387];
      \nz.mem_2986_sv2v_reg  <= w_data_i[1386];
      \nz.mem_2985_sv2v_reg  <= w_data_i[1385];
      \nz.mem_2984_sv2v_reg  <= w_data_i[1384];
      \nz.mem_2983_sv2v_reg  <= w_data_i[1383];
      \nz.mem_2982_sv2v_reg  <= w_data_i[1382];
      \nz.mem_2981_sv2v_reg  <= w_data_i[1381];
      \nz.mem_2980_sv2v_reg  <= w_data_i[1380];
      \nz.mem_2979_sv2v_reg  <= w_data_i[1379];
      \nz.mem_2978_sv2v_reg  <= w_data_i[1378];
      \nz.mem_2977_sv2v_reg  <= w_data_i[1377];
      \nz.mem_2976_sv2v_reg  <= w_data_i[1376];
      \nz.mem_2975_sv2v_reg  <= w_data_i[1375];
      \nz.mem_2974_sv2v_reg  <= w_data_i[1374];
      \nz.mem_2973_sv2v_reg  <= w_data_i[1373];
      \nz.mem_2972_sv2v_reg  <= w_data_i[1372];
      \nz.mem_2971_sv2v_reg  <= w_data_i[1371];
      \nz.mem_2970_sv2v_reg  <= w_data_i[1370];
      \nz.mem_2969_sv2v_reg  <= w_data_i[1369];
      \nz.mem_2968_sv2v_reg  <= w_data_i[1368];
      \nz.mem_2967_sv2v_reg  <= w_data_i[1367];
      \nz.mem_2966_sv2v_reg  <= w_data_i[1366];
      \nz.mem_2965_sv2v_reg  <= w_data_i[1365];
      \nz.mem_2964_sv2v_reg  <= w_data_i[1364];
      \nz.mem_2963_sv2v_reg  <= w_data_i[1363];
      \nz.mem_2962_sv2v_reg  <= w_data_i[1362];
      \nz.mem_2961_sv2v_reg  <= w_data_i[1361];
      \nz.mem_2960_sv2v_reg  <= w_data_i[1360];
      \nz.mem_2959_sv2v_reg  <= w_data_i[1359];
      \nz.mem_2958_sv2v_reg  <= w_data_i[1358];
      \nz.mem_2957_sv2v_reg  <= w_data_i[1357];
      \nz.mem_2956_sv2v_reg  <= w_data_i[1356];
      \nz.mem_2955_sv2v_reg  <= w_data_i[1355];
      \nz.mem_2954_sv2v_reg  <= w_data_i[1354];
      \nz.mem_2953_sv2v_reg  <= w_data_i[1353];
      \nz.mem_2952_sv2v_reg  <= w_data_i[1352];
      \nz.mem_2951_sv2v_reg  <= w_data_i[1351];
      \nz.mem_2950_sv2v_reg  <= w_data_i[1350];
      \nz.mem_2949_sv2v_reg  <= w_data_i[1349];
      \nz.mem_2948_sv2v_reg  <= w_data_i[1348];
      \nz.mem_2947_sv2v_reg  <= w_data_i[1347];
      \nz.mem_2946_sv2v_reg  <= w_data_i[1346];
      \nz.mem_2945_sv2v_reg  <= w_data_i[1345];
      \nz.mem_2944_sv2v_reg  <= w_data_i[1344];
      \nz.mem_2943_sv2v_reg  <= w_data_i[1343];
      \nz.mem_2942_sv2v_reg  <= w_data_i[1342];
      \nz.mem_2941_sv2v_reg  <= w_data_i[1341];
      \nz.mem_2940_sv2v_reg  <= w_data_i[1340];
      \nz.mem_2939_sv2v_reg  <= w_data_i[1339];
      \nz.mem_2938_sv2v_reg  <= w_data_i[1338];
      \nz.mem_2937_sv2v_reg  <= w_data_i[1337];
      \nz.mem_2936_sv2v_reg  <= w_data_i[1336];
      \nz.mem_2935_sv2v_reg  <= w_data_i[1335];
      \nz.mem_2934_sv2v_reg  <= w_data_i[1334];
      \nz.mem_2933_sv2v_reg  <= w_data_i[1333];
      \nz.mem_2932_sv2v_reg  <= w_data_i[1332];
      \nz.mem_2931_sv2v_reg  <= w_data_i[1331];
      \nz.mem_2930_sv2v_reg  <= w_data_i[1330];
      \nz.mem_2929_sv2v_reg  <= w_data_i[1329];
      \nz.mem_2928_sv2v_reg  <= w_data_i[1328];
      \nz.mem_2927_sv2v_reg  <= w_data_i[1327];
      \nz.mem_2926_sv2v_reg  <= w_data_i[1326];
      \nz.mem_2925_sv2v_reg  <= w_data_i[1325];
      \nz.mem_2924_sv2v_reg  <= w_data_i[1324];
      \nz.mem_2923_sv2v_reg  <= w_data_i[1323];
      \nz.mem_2922_sv2v_reg  <= w_data_i[1322];
      \nz.mem_2921_sv2v_reg  <= w_data_i[1321];
      \nz.mem_2920_sv2v_reg  <= w_data_i[1320];
      \nz.mem_2919_sv2v_reg  <= w_data_i[1319];
      \nz.mem_2918_sv2v_reg  <= w_data_i[1318];
      \nz.mem_2917_sv2v_reg  <= w_data_i[1317];
      \nz.mem_2916_sv2v_reg  <= w_data_i[1316];
      \nz.mem_2915_sv2v_reg  <= w_data_i[1315];
      \nz.mem_2914_sv2v_reg  <= w_data_i[1314];
      \nz.mem_2913_sv2v_reg  <= w_data_i[1313];
      \nz.mem_2912_sv2v_reg  <= w_data_i[1312];
      \nz.mem_2911_sv2v_reg  <= w_data_i[1311];
      \nz.mem_2910_sv2v_reg  <= w_data_i[1310];
      \nz.mem_2909_sv2v_reg  <= w_data_i[1309];
      \nz.mem_2908_sv2v_reg  <= w_data_i[1308];
      \nz.mem_2907_sv2v_reg  <= w_data_i[1307];
      \nz.mem_2906_sv2v_reg  <= w_data_i[1306];
      \nz.mem_2905_sv2v_reg  <= w_data_i[1305];
      \nz.mem_2904_sv2v_reg  <= w_data_i[1304];
      \nz.mem_2903_sv2v_reg  <= w_data_i[1303];
      \nz.mem_1602_sv2v_reg  <= w_data_i[2];
    end 
    if(N26) begin
      \nz.mem_2902_sv2v_reg  <= w_data_i[1302];
      \nz.mem_2901_sv2v_reg  <= w_data_i[1301];
      \nz.mem_2900_sv2v_reg  <= w_data_i[1300];
      \nz.mem_2899_sv2v_reg  <= w_data_i[1299];
      \nz.mem_2898_sv2v_reg  <= w_data_i[1298];
      \nz.mem_2897_sv2v_reg  <= w_data_i[1297];
      \nz.mem_2896_sv2v_reg  <= w_data_i[1296];
      \nz.mem_2895_sv2v_reg  <= w_data_i[1295];
      \nz.mem_2894_sv2v_reg  <= w_data_i[1294];
      \nz.mem_2893_sv2v_reg  <= w_data_i[1293];
      \nz.mem_2892_sv2v_reg  <= w_data_i[1292];
      \nz.mem_2891_sv2v_reg  <= w_data_i[1291];
      \nz.mem_2890_sv2v_reg  <= w_data_i[1290];
      \nz.mem_2889_sv2v_reg  <= w_data_i[1289];
      \nz.mem_2888_sv2v_reg  <= w_data_i[1288];
      \nz.mem_2887_sv2v_reg  <= w_data_i[1287];
      \nz.mem_2886_sv2v_reg  <= w_data_i[1286];
      \nz.mem_2885_sv2v_reg  <= w_data_i[1285];
      \nz.mem_2884_sv2v_reg  <= w_data_i[1284];
      \nz.mem_2883_sv2v_reg  <= w_data_i[1283];
      \nz.mem_2882_sv2v_reg  <= w_data_i[1282];
      \nz.mem_2881_sv2v_reg  <= w_data_i[1281];
      \nz.mem_2880_sv2v_reg  <= w_data_i[1280];
      \nz.mem_2879_sv2v_reg  <= w_data_i[1279];
      \nz.mem_2878_sv2v_reg  <= w_data_i[1278];
      \nz.mem_2877_sv2v_reg  <= w_data_i[1277];
      \nz.mem_2876_sv2v_reg  <= w_data_i[1276];
      \nz.mem_2875_sv2v_reg  <= w_data_i[1275];
      \nz.mem_2874_sv2v_reg  <= w_data_i[1274];
      \nz.mem_2873_sv2v_reg  <= w_data_i[1273];
      \nz.mem_2872_sv2v_reg  <= w_data_i[1272];
      \nz.mem_2871_sv2v_reg  <= w_data_i[1271];
      \nz.mem_2870_sv2v_reg  <= w_data_i[1270];
      \nz.mem_2869_sv2v_reg  <= w_data_i[1269];
      \nz.mem_2868_sv2v_reg  <= w_data_i[1268];
      \nz.mem_2867_sv2v_reg  <= w_data_i[1267];
      \nz.mem_2866_sv2v_reg  <= w_data_i[1266];
      \nz.mem_2865_sv2v_reg  <= w_data_i[1265];
      \nz.mem_2864_sv2v_reg  <= w_data_i[1264];
      \nz.mem_2863_sv2v_reg  <= w_data_i[1263];
      \nz.mem_2862_sv2v_reg  <= w_data_i[1262];
      \nz.mem_2861_sv2v_reg  <= w_data_i[1261];
      \nz.mem_2860_sv2v_reg  <= w_data_i[1260];
      \nz.mem_2859_sv2v_reg  <= w_data_i[1259];
      \nz.mem_2858_sv2v_reg  <= w_data_i[1258];
      \nz.mem_2857_sv2v_reg  <= w_data_i[1257];
      \nz.mem_2856_sv2v_reg  <= w_data_i[1256];
      \nz.mem_2855_sv2v_reg  <= w_data_i[1255];
      \nz.mem_2854_sv2v_reg  <= w_data_i[1254];
      \nz.mem_2853_sv2v_reg  <= w_data_i[1253];
      \nz.mem_2852_sv2v_reg  <= w_data_i[1252];
      \nz.mem_2851_sv2v_reg  <= w_data_i[1251];
      \nz.mem_2850_sv2v_reg  <= w_data_i[1250];
      \nz.mem_2849_sv2v_reg  <= w_data_i[1249];
      \nz.mem_2848_sv2v_reg  <= w_data_i[1248];
      \nz.mem_2847_sv2v_reg  <= w_data_i[1247];
      \nz.mem_2846_sv2v_reg  <= w_data_i[1246];
      \nz.mem_2845_sv2v_reg  <= w_data_i[1245];
      \nz.mem_2844_sv2v_reg  <= w_data_i[1244];
      \nz.mem_2843_sv2v_reg  <= w_data_i[1243];
      \nz.mem_2842_sv2v_reg  <= w_data_i[1242];
      \nz.mem_2841_sv2v_reg  <= w_data_i[1241];
      \nz.mem_2840_sv2v_reg  <= w_data_i[1240];
      \nz.mem_2839_sv2v_reg  <= w_data_i[1239];
      \nz.mem_2838_sv2v_reg  <= w_data_i[1238];
      \nz.mem_2837_sv2v_reg  <= w_data_i[1237];
      \nz.mem_2836_sv2v_reg  <= w_data_i[1236];
      \nz.mem_2835_sv2v_reg  <= w_data_i[1235];
      \nz.mem_2834_sv2v_reg  <= w_data_i[1234];
      \nz.mem_2833_sv2v_reg  <= w_data_i[1233];
      \nz.mem_2832_sv2v_reg  <= w_data_i[1232];
      \nz.mem_2831_sv2v_reg  <= w_data_i[1231];
      \nz.mem_2830_sv2v_reg  <= w_data_i[1230];
      \nz.mem_2829_sv2v_reg  <= w_data_i[1229];
      \nz.mem_2828_sv2v_reg  <= w_data_i[1228];
      \nz.mem_2827_sv2v_reg  <= w_data_i[1227];
      \nz.mem_2826_sv2v_reg  <= w_data_i[1226];
      \nz.mem_2825_sv2v_reg  <= w_data_i[1225];
      \nz.mem_2824_sv2v_reg  <= w_data_i[1224];
      \nz.mem_2823_sv2v_reg  <= w_data_i[1223];
      \nz.mem_2822_sv2v_reg  <= w_data_i[1222];
      \nz.mem_2821_sv2v_reg  <= w_data_i[1221];
      \nz.mem_2820_sv2v_reg  <= w_data_i[1220];
      \nz.mem_2819_sv2v_reg  <= w_data_i[1219];
      \nz.mem_2818_sv2v_reg  <= w_data_i[1218];
      \nz.mem_2817_sv2v_reg  <= w_data_i[1217];
      \nz.mem_2816_sv2v_reg  <= w_data_i[1216];
      \nz.mem_2815_sv2v_reg  <= w_data_i[1215];
      \nz.mem_2814_sv2v_reg  <= w_data_i[1214];
      \nz.mem_2813_sv2v_reg  <= w_data_i[1213];
      \nz.mem_2812_sv2v_reg  <= w_data_i[1212];
      \nz.mem_2811_sv2v_reg  <= w_data_i[1211];
      \nz.mem_2810_sv2v_reg  <= w_data_i[1210];
      \nz.mem_2809_sv2v_reg  <= w_data_i[1209];
      \nz.mem_2808_sv2v_reg  <= w_data_i[1208];
      \nz.mem_2807_sv2v_reg  <= w_data_i[1207];
      \nz.mem_2806_sv2v_reg  <= w_data_i[1206];
      \nz.mem_2805_sv2v_reg  <= w_data_i[1205];
      \nz.mem_2804_sv2v_reg  <= w_data_i[1204];
      \nz.mem_1603_sv2v_reg  <= w_data_i[3];
    end 
    if(N27) begin
      \nz.mem_2803_sv2v_reg  <= w_data_i[1203];
      \nz.mem_2802_sv2v_reg  <= w_data_i[1202];
      \nz.mem_2801_sv2v_reg  <= w_data_i[1201];
      \nz.mem_2800_sv2v_reg  <= w_data_i[1200];
      \nz.mem_2799_sv2v_reg  <= w_data_i[1199];
      \nz.mem_2798_sv2v_reg  <= w_data_i[1198];
      \nz.mem_2797_sv2v_reg  <= w_data_i[1197];
      \nz.mem_2796_sv2v_reg  <= w_data_i[1196];
      \nz.mem_2795_sv2v_reg  <= w_data_i[1195];
      \nz.mem_2794_sv2v_reg  <= w_data_i[1194];
      \nz.mem_2793_sv2v_reg  <= w_data_i[1193];
      \nz.mem_2792_sv2v_reg  <= w_data_i[1192];
      \nz.mem_2791_sv2v_reg  <= w_data_i[1191];
      \nz.mem_2790_sv2v_reg  <= w_data_i[1190];
      \nz.mem_2789_sv2v_reg  <= w_data_i[1189];
      \nz.mem_2788_sv2v_reg  <= w_data_i[1188];
      \nz.mem_2787_sv2v_reg  <= w_data_i[1187];
      \nz.mem_2786_sv2v_reg  <= w_data_i[1186];
      \nz.mem_2785_sv2v_reg  <= w_data_i[1185];
      \nz.mem_2784_sv2v_reg  <= w_data_i[1184];
      \nz.mem_2783_sv2v_reg  <= w_data_i[1183];
      \nz.mem_2782_sv2v_reg  <= w_data_i[1182];
      \nz.mem_2781_sv2v_reg  <= w_data_i[1181];
      \nz.mem_2780_sv2v_reg  <= w_data_i[1180];
      \nz.mem_2779_sv2v_reg  <= w_data_i[1179];
      \nz.mem_2778_sv2v_reg  <= w_data_i[1178];
      \nz.mem_2777_sv2v_reg  <= w_data_i[1177];
      \nz.mem_2776_sv2v_reg  <= w_data_i[1176];
      \nz.mem_2775_sv2v_reg  <= w_data_i[1175];
      \nz.mem_2774_sv2v_reg  <= w_data_i[1174];
      \nz.mem_2773_sv2v_reg  <= w_data_i[1173];
      \nz.mem_2772_sv2v_reg  <= w_data_i[1172];
      \nz.mem_2771_sv2v_reg  <= w_data_i[1171];
      \nz.mem_2770_sv2v_reg  <= w_data_i[1170];
      \nz.mem_2769_sv2v_reg  <= w_data_i[1169];
      \nz.mem_2768_sv2v_reg  <= w_data_i[1168];
      \nz.mem_2767_sv2v_reg  <= w_data_i[1167];
      \nz.mem_2766_sv2v_reg  <= w_data_i[1166];
      \nz.mem_2765_sv2v_reg  <= w_data_i[1165];
      \nz.mem_2764_sv2v_reg  <= w_data_i[1164];
      \nz.mem_2763_sv2v_reg  <= w_data_i[1163];
      \nz.mem_2762_sv2v_reg  <= w_data_i[1162];
      \nz.mem_2761_sv2v_reg  <= w_data_i[1161];
      \nz.mem_2760_sv2v_reg  <= w_data_i[1160];
      \nz.mem_2759_sv2v_reg  <= w_data_i[1159];
      \nz.mem_2758_sv2v_reg  <= w_data_i[1158];
      \nz.mem_2757_sv2v_reg  <= w_data_i[1157];
      \nz.mem_2756_sv2v_reg  <= w_data_i[1156];
      \nz.mem_2755_sv2v_reg  <= w_data_i[1155];
      \nz.mem_2754_sv2v_reg  <= w_data_i[1154];
      \nz.mem_2753_sv2v_reg  <= w_data_i[1153];
      \nz.mem_2752_sv2v_reg  <= w_data_i[1152];
      \nz.mem_2751_sv2v_reg  <= w_data_i[1151];
      \nz.mem_2750_sv2v_reg  <= w_data_i[1150];
      \nz.mem_2749_sv2v_reg  <= w_data_i[1149];
      \nz.mem_2748_sv2v_reg  <= w_data_i[1148];
      \nz.mem_2747_sv2v_reg  <= w_data_i[1147];
      \nz.mem_2746_sv2v_reg  <= w_data_i[1146];
      \nz.mem_2745_sv2v_reg  <= w_data_i[1145];
      \nz.mem_2744_sv2v_reg  <= w_data_i[1144];
      \nz.mem_2743_sv2v_reg  <= w_data_i[1143];
      \nz.mem_2742_sv2v_reg  <= w_data_i[1142];
      \nz.mem_2741_sv2v_reg  <= w_data_i[1141];
      \nz.mem_2740_sv2v_reg  <= w_data_i[1140];
      \nz.mem_2739_sv2v_reg  <= w_data_i[1139];
      \nz.mem_2738_sv2v_reg  <= w_data_i[1138];
      \nz.mem_2737_sv2v_reg  <= w_data_i[1137];
      \nz.mem_2736_sv2v_reg  <= w_data_i[1136];
      \nz.mem_2735_sv2v_reg  <= w_data_i[1135];
      \nz.mem_2734_sv2v_reg  <= w_data_i[1134];
      \nz.mem_2733_sv2v_reg  <= w_data_i[1133];
      \nz.mem_2732_sv2v_reg  <= w_data_i[1132];
      \nz.mem_2731_sv2v_reg  <= w_data_i[1131];
      \nz.mem_2730_sv2v_reg  <= w_data_i[1130];
      \nz.mem_2729_sv2v_reg  <= w_data_i[1129];
      \nz.mem_2728_sv2v_reg  <= w_data_i[1128];
      \nz.mem_2727_sv2v_reg  <= w_data_i[1127];
      \nz.mem_2726_sv2v_reg  <= w_data_i[1126];
      \nz.mem_2725_sv2v_reg  <= w_data_i[1125];
      \nz.mem_2724_sv2v_reg  <= w_data_i[1124];
      \nz.mem_2723_sv2v_reg  <= w_data_i[1123];
      \nz.mem_2722_sv2v_reg  <= w_data_i[1122];
      \nz.mem_2721_sv2v_reg  <= w_data_i[1121];
      \nz.mem_2720_sv2v_reg  <= w_data_i[1120];
      \nz.mem_2719_sv2v_reg  <= w_data_i[1119];
      \nz.mem_2718_sv2v_reg  <= w_data_i[1118];
      \nz.mem_2717_sv2v_reg  <= w_data_i[1117];
      \nz.mem_2716_sv2v_reg  <= w_data_i[1116];
      \nz.mem_2715_sv2v_reg  <= w_data_i[1115];
      \nz.mem_2714_sv2v_reg  <= w_data_i[1114];
      \nz.mem_2713_sv2v_reg  <= w_data_i[1113];
      \nz.mem_2712_sv2v_reg  <= w_data_i[1112];
      \nz.mem_2711_sv2v_reg  <= w_data_i[1111];
      \nz.mem_2710_sv2v_reg  <= w_data_i[1110];
      \nz.mem_2709_sv2v_reg  <= w_data_i[1109];
      \nz.mem_2708_sv2v_reg  <= w_data_i[1108];
      \nz.mem_2707_sv2v_reg  <= w_data_i[1107];
      \nz.mem_2706_sv2v_reg  <= w_data_i[1106];
      \nz.mem_2705_sv2v_reg  <= w_data_i[1105];
      \nz.mem_1604_sv2v_reg  <= w_data_i[4];
    end 
    if(N28) begin
      \nz.mem_2704_sv2v_reg  <= w_data_i[1104];
      \nz.mem_2703_sv2v_reg  <= w_data_i[1103];
      \nz.mem_2702_sv2v_reg  <= w_data_i[1102];
      \nz.mem_2701_sv2v_reg  <= w_data_i[1101];
      \nz.mem_2700_sv2v_reg  <= w_data_i[1100];
      \nz.mem_2699_sv2v_reg  <= w_data_i[1099];
      \nz.mem_2698_sv2v_reg  <= w_data_i[1098];
      \nz.mem_2697_sv2v_reg  <= w_data_i[1097];
      \nz.mem_2696_sv2v_reg  <= w_data_i[1096];
      \nz.mem_2695_sv2v_reg  <= w_data_i[1095];
      \nz.mem_2694_sv2v_reg  <= w_data_i[1094];
      \nz.mem_2693_sv2v_reg  <= w_data_i[1093];
      \nz.mem_2692_sv2v_reg  <= w_data_i[1092];
      \nz.mem_2691_sv2v_reg  <= w_data_i[1091];
      \nz.mem_2690_sv2v_reg  <= w_data_i[1090];
      \nz.mem_2689_sv2v_reg  <= w_data_i[1089];
      \nz.mem_2688_sv2v_reg  <= w_data_i[1088];
      \nz.mem_2687_sv2v_reg  <= w_data_i[1087];
      \nz.mem_2686_sv2v_reg  <= w_data_i[1086];
      \nz.mem_2685_sv2v_reg  <= w_data_i[1085];
      \nz.mem_2684_sv2v_reg  <= w_data_i[1084];
      \nz.mem_2683_sv2v_reg  <= w_data_i[1083];
      \nz.mem_2682_sv2v_reg  <= w_data_i[1082];
      \nz.mem_2681_sv2v_reg  <= w_data_i[1081];
      \nz.mem_2680_sv2v_reg  <= w_data_i[1080];
      \nz.mem_2679_sv2v_reg  <= w_data_i[1079];
      \nz.mem_2678_sv2v_reg  <= w_data_i[1078];
      \nz.mem_2677_sv2v_reg  <= w_data_i[1077];
      \nz.mem_2676_sv2v_reg  <= w_data_i[1076];
      \nz.mem_2675_sv2v_reg  <= w_data_i[1075];
      \nz.mem_2674_sv2v_reg  <= w_data_i[1074];
      \nz.mem_2673_sv2v_reg  <= w_data_i[1073];
      \nz.mem_2672_sv2v_reg  <= w_data_i[1072];
      \nz.mem_2671_sv2v_reg  <= w_data_i[1071];
      \nz.mem_2670_sv2v_reg  <= w_data_i[1070];
      \nz.mem_2669_sv2v_reg  <= w_data_i[1069];
      \nz.mem_2668_sv2v_reg  <= w_data_i[1068];
      \nz.mem_2667_sv2v_reg  <= w_data_i[1067];
      \nz.mem_2666_sv2v_reg  <= w_data_i[1066];
      \nz.mem_2665_sv2v_reg  <= w_data_i[1065];
      \nz.mem_2664_sv2v_reg  <= w_data_i[1064];
      \nz.mem_2663_sv2v_reg  <= w_data_i[1063];
      \nz.mem_2662_sv2v_reg  <= w_data_i[1062];
      \nz.mem_2661_sv2v_reg  <= w_data_i[1061];
      \nz.mem_2660_sv2v_reg  <= w_data_i[1060];
      \nz.mem_2659_sv2v_reg  <= w_data_i[1059];
      \nz.mem_2658_sv2v_reg  <= w_data_i[1058];
      \nz.mem_2657_sv2v_reg  <= w_data_i[1057];
      \nz.mem_2656_sv2v_reg  <= w_data_i[1056];
      \nz.mem_2655_sv2v_reg  <= w_data_i[1055];
      \nz.mem_2654_sv2v_reg  <= w_data_i[1054];
      \nz.mem_2653_sv2v_reg  <= w_data_i[1053];
      \nz.mem_2652_sv2v_reg  <= w_data_i[1052];
      \nz.mem_2651_sv2v_reg  <= w_data_i[1051];
      \nz.mem_2650_sv2v_reg  <= w_data_i[1050];
      \nz.mem_2649_sv2v_reg  <= w_data_i[1049];
      \nz.mem_2648_sv2v_reg  <= w_data_i[1048];
      \nz.mem_2647_sv2v_reg  <= w_data_i[1047];
      \nz.mem_2646_sv2v_reg  <= w_data_i[1046];
      \nz.mem_2645_sv2v_reg  <= w_data_i[1045];
      \nz.mem_2644_sv2v_reg  <= w_data_i[1044];
      \nz.mem_2643_sv2v_reg  <= w_data_i[1043];
      \nz.mem_2642_sv2v_reg  <= w_data_i[1042];
      \nz.mem_2641_sv2v_reg  <= w_data_i[1041];
      \nz.mem_2640_sv2v_reg  <= w_data_i[1040];
      \nz.mem_2639_sv2v_reg  <= w_data_i[1039];
      \nz.mem_2638_sv2v_reg  <= w_data_i[1038];
      \nz.mem_2637_sv2v_reg  <= w_data_i[1037];
      \nz.mem_2636_sv2v_reg  <= w_data_i[1036];
      \nz.mem_2635_sv2v_reg  <= w_data_i[1035];
      \nz.mem_2634_sv2v_reg  <= w_data_i[1034];
      \nz.mem_2633_sv2v_reg  <= w_data_i[1033];
      \nz.mem_2632_sv2v_reg  <= w_data_i[1032];
      \nz.mem_2631_sv2v_reg  <= w_data_i[1031];
      \nz.mem_2630_sv2v_reg  <= w_data_i[1030];
      \nz.mem_2629_sv2v_reg  <= w_data_i[1029];
      \nz.mem_2628_sv2v_reg  <= w_data_i[1028];
      \nz.mem_2627_sv2v_reg  <= w_data_i[1027];
      \nz.mem_2626_sv2v_reg  <= w_data_i[1026];
      \nz.mem_2625_sv2v_reg  <= w_data_i[1025];
      \nz.mem_2624_sv2v_reg  <= w_data_i[1024];
      \nz.mem_2623_sv2v_reg  <= w_data_i[1023];
      \nz.mem_2622_sv2v_reg  <= w_data_i[1022];
      \nz.mem_2621_sv2v_reg  <= w_data_i[1021];
      \nz.mem_2620_sv2v_reg  <= w_data_i[1020];
      \nz.mem_2619_sv2v_reg  <= w_data_i[1019];
      \nz.mem_2618_sv2v_reg  <= w_data_i[1018];
      \nz.mem_2617_sv2v_reg  <= w_data_i[1017];
      \nz.mem_2616_sv2v_reg  <= w_data_i[1016];
      \nz.mem_2615_sv2v_reg  <= w_data_i[1015];
      \nz.mem_2614_sv2v_reg  <= w_data_i[1014];
      \nz.mem_2613_sv2v_reg  <= w_data_i[1013];
      \nz.mem_2612_sv2v_reg  <= w_data_i[1012];
      \nz.mem_2611_sv2v_reg  <= w_data_i[1011];
      \nz.mem_2610_sv2v_reg  <= w_data_i[1010];
      \nz.mem_2609_sv2v_reg  <= w_data_i[1009];
      \nz.mem_2608_sv2v_reg  <= w_data_i[1008];
      \nz.mem_2607_sv2v_reg  <= w_data_i[1007];
      \nz.mem_2606_sv2v_reg  <= w_data_i[1006];
      \nz.mem_1605_sv2v_reg  <= w_data_i[5];
    end 
    if(N29) begin
      \nz.mem_2605_sv2v_reg  <= w_data_i[1005];
      \nz.mem_2604_sv2v_reg  <= w_data_i[1004];
      \nz.mem_2603_sv2v_reg  <= w_data_i[1003];
      \nz.mem_2602_sv2v_reg  <= w_data_i[1002];
      \nz.mem_2601_sv2v_reg  <= w_data_i[1001];
      \nz.mem_2600_sv2v_reg  <= w_data_i[1000];
      \nz.mem_2599_sv2v_reg  <= w_data_i[999];
      \nz.mem_2598_sv2v_reg  <= w_data_i[998];
      \nz.mem_2597_sv2v_reg  <= w_data_i[997];
      \nz.mem_2596_sv2v_reg  <= w_data_i[996];
      \nz.mem_2595_sv2v_reg  <= w_data_i[995];
      \nz.mem_2594_sv2v_reg  <= w_data_i[994];
      \nz.mem_2593_sv2v_reg  <= w_data_i[993];
      \nz.mem_2592_sv2v_reg  <= w_data_i[992];
      \nz.mem_2591_sv2v_reg  <= w_data_i[991];
      \nz.mem_2590_sv2v_reg  <= w_data_i[990];
      \nz.mem_2589_sv2v_reg  <= w_data_i[989];
      \nz.mem_2588_sv2v_reg  <= w_data_i[988];
      \nz.mem_2587_sv2v_reg  <= w_data_i[987];
      \nz.mem_2586_sv2v_reg  <= w_data_i[986];
      \nz.mem_2585_sv2v_reg  <= w_data_i[985];
      \nz.mem_2584_sv2v_reg  <= w_data_i[984];
      \nz.mem_2583_sv2v_reg  <= w_data_i[983];
      \nz.mem_2582_sv2v_reg  <= w_data_i[982];
      \nz.mem_2581_sv2v_reg  <= w_data_i[981];
      \nz.mem_2580_sv2v_reg  <= w_data_i[980];
      \nz.mem_2579_sv2v_reg  <= w_data_i[979];
      \nz.mem_2578_sv2v_reg  <= w_data_i[978];
      \nz.mem_2577_sv2v_reg  <= w_data_i[977];
      \nz.mem_2576_sv2v_reg  <= w_data_i[976];
      \nz.mem_2575_sv2v_reg  <= w_data_i[975];
      \nz.mem_2574_sv2v_reg  <= w_data_i[974];
      \nz.mem_2573_sv2v_reg  <= w_data_i[973];
      \nz.mem_2572_sv2v_reg  <= w_data_i[972];
      \nz.mem_2571_sv2v_reg  <= w_data_i[971];
      \nz.mem_2570_sv2v_reg  <= w_data_i[970];
      \nz.mem_2569_sv2v_reg  <= w_data_i[969];
      \nz.mem_2568_sv2v_reg  <= w_data_i[968];
      \nz.mem_2567_sv2v_reg  <= w_data_i[967];
      \nz.mem_2566_sv2v_reg  <= w_data_i[966];
      \nz.mem_2565_sv2v_reg  <= w_data_i[965];
      \nz.mem_2564_sv2v_reg  <= w_data_i[964];
      \nz.mem_2563_sv2v_reg  <= w_data_i[963];
      \nz.mem_2562_sv2v_reg  <= w_data_i[962];
      \nz.mem_2561_sv2v_reg  <= w_data_i[961];
      \nz.mem_2560_sv2v_reg  <= w_data_i[960];
      \nz.mem_2559_sv2v_reg  <= w_data_i[959];
      \nz.mem_2558_sv2v_reg  <= w_data_i[958];
      \nz.mem_2557_sv2v_reg  <= w_data_i[957];
      \nz.mem_2556_sv2v_reg  <= w_data_i[956];
      \nz.mem_2555_sv2v_reg  <= w_data_i[955];
      \nz.mem_2554_sv2v_reg  <= w_data_i[954];
      \nz.mem_2553_sv2v_reg  <= w_data_i[953];
      \nz.mem_2552_sv2v_reg  <= w_data_i[952];
      \nz.mem_2551_sv2v_reg  <= w_data_i[951];
      \nz.mem_2550_sv2v_reg  <= w_data_i[950];
      \nz.mem_2549_sv2v_reg  <= w_data_i[949];
      \nz.mem_2548_sv2v_reg  <= w_data_i[948];
      \nz.mem_2547_sv2v_reg  <= w_data_i[947];
      \nz.mem_2546_sv2v_reg  <= w_data_i[946];
      \nz.mem_2545_sv2v_reg  <= w_data_i[945];
      \nz.mem_2544_sv2v_reg  <= w_data_i[944];
      \nz.mem_2543_sv2v_reg  <= w_data_i[943];
      \nz.mem_2542_sv2v_reg  <= w_data_i[942];
      \nz.mem_2541_sv2v_reg  <= w_data_i[941];
      \nz.mem_2540_sv2v_reg  <= w_data_i[940];
      \nz.mem_2539_sv2v_reg  <= w_data_i[939];
      \nz.mem_2538_sv2v_reg  <= w_data_i[938];
      \nz.mem_2537_sv2v_reg  <= w_data_i[937];
      \nz.mem_2536_sv2v_reg  <= w_data_i[936];
      \nz.mem_2535_sv2v_reg  <= w_data_i[935];
      \nz.mem_2534_sv2v_reg  <= w_data_i[934];
      \nz.mem_2533_sv2v_reg  <= w_data_i[933];
      \nz.mem_2532_sv2v_reg  <= w_data_i[932];
      \nz.mem_2531_sv2v_reg  <= w_data_i[931];
      \nz.mem_2530_sv2v_reg  <= w_data_i[930];
      \nz.mem_2529_sv2v_reg  <= w_data_i[929];
      \nz.mem_2528_sv2v_reg  <= w_data_i[928];
      \nz.mem_2527_sv2v_reg  <= w_data_i[927];
      \nz.mem_2526_sv2v_reg  <= w_data_i[926];
      \nz.mem_2525_sv2v_reg  <= w_data_i[925];
      \nz.mem_2524_sv2v_reg  <= w_data_i[924];
      \nz.mem_2523_sv2v_reg  <= w_data_i[923];
      \nz.mem_2522_sv2v_reg  <= w_data_i[922];
      \nz.mem_2521_sv2v_reg  <= w_data_i[921];
      \nz.mem_2520_sv2v_reg  <= w_data_i[920];
      \nz.mem_2519_sv2v_reg  <= w_data_i[919];
      \nz.mem_2518_sv2v_reg  <= w_data_i[918];
      \nz.mem_2517_sv2v_reg  <= w_data_i[917];
      \nz.mem_2516_sv2v_reg  <= w_data_i[916];
      \nz.mem_2515_sv2v_reg  <= w_data_i[915];
      \nz.mem_2514_sv2v_reg  <= w_data_i[914];
      \nz.mem_2513_sv2v_reg  <= w_data_i[913];
      \nz.mem_2512_sv2v_reg  <= w_data_i[912];
      \nz.mem_2511_sv2v_reg  <= w_data_i[911];
      \nz.mem_2510_sv2v_reg  <= w_data_i[910];
      \nz.mem_2509_sv2v_reg  <= w_data_i[909];
      \nz.mem_2508_sv2v_reg  <= w_data_i[908];
      \nz.mem_2507_sv2v_reg  <= w_data_i[907];
      \nz.mem_1606_sv2v_reg  <= w_data_i[6];
    end 
    if(N30) begin
      \nz.mem_2506_sv2v_reg  <= w_data_i[906];
      \nz.mem_2505_sv2v_reg  <= w_data_i[905];
      \nz.mem_2504_sv2v_reg  <= w_data_i[904];
      \nz.mem_2503_sv2v_reg  <= w_data_i[903];
      \nz.mem_2502_sv2v_reg  <= w_data_i[902];
      \nz.mem_2501_sv2v_reg  <= w_data_i[901];
      \nz.mem_2500_sv2v_reg  <= w_data_i[900];
      \nz.mem_2499_sv2v_reg  <= w_data_i[899];
      \nz.mem_2498_sv2v_reg  <= w_data_i[898];
      \nz.mem_2497_sv2v_reg  <= w_data_i[897];
      \nz.mem_2496_sv2v_reg  <= w_data_i[896];
      \nz.mem_2495_sv2v_reg  <= w_data_i[895];
      \nz.mem_2494_sv2v_reg  <= w_data_i[894];
      \nz.mem_2493_sv2v_reg  <= w_data_i[893];
      \nz.mem_2492_sv2v_reg  <= w_data_i[892];
      \nz.mem_2491_sv2v_reg  <= w_data_i[891];
      \nz.mem_2490_sv2v_reg  <= w_data_i[890];
      \nz.mem_2489_sv2v_reg  <= w_data_i[889];
      \nz.mem_2488_sv2v_reg  <= w_data_i[888];
      \nz.mem_2487_sv2v_reg  <= w_data_i[887];
      \nz.mem_2486_sv2v_reg  <= w_data_i[886];
      \nz.mem_2485_sv2v_reg  <= w_data_i[885];
      \nz.mem_2484_sv2v_reg  <= w_data_i[884];
      \nz.mem_2483_sv2v_reg  <= w_data_i[883];
      \nz.mem_2482_sv2v_reg  <= w_data_i[882];
      \nz.mem_2481_sv2v_reg  <= w_data_i[881];
      \nz.mem_2480_sv2v_reg  <= w_data_i[880];
      \nz.mem_2479_sv2v_reg  <= w_data_i[879];
      \nz.mem_2478_sv2v_reg  <= w_data_i[878];
      \nz.mem_2477_sv2v_reg  <= w_data_i[877];
      \nz.mem_2476_sv2v_reg  <= w_data_i[876];
      \nz.mem_2475_sv2v_reg  <= w_data_i[875];
      \nz.mem_2474_sv2v_reg  <= w_data_i[874];
      \nz.mem_2473_sv2v_reg  <= w_data_i[873];
      \nz.mem_2472_sv2v_reg  <= w_data_i[872];
      \nz.mem_2471_sv2v_reg  <= w_data_i[871];
      \nz.mem_2470_sv2v_reg  <= w_data_i[870];
      \nz.mem_2469_sv2v_reg  <= w_data_i[869];
      \nz.mem_2468_sv2v_reg  <= w_data_i[868];
      \nz.mem_2467_sv2v_reg  <= w_data_i[867];
      \nz.mem_2466_sv2v_reg  <= w_data_i[866];
      \nz.mem_2465_sv2v_reg  <= w_data_i[865];
      \nz.mem_2464_sv2v_reg  <= w_data_i[864];
      \nz.mem_2463_sv2v_reg  <= w_data_i[863];
      \nz.mem_2462_sv2v_reg  <= w_data_i[862];
      \nz.mem_2461_sv2v_reg  <= w_data_i[861];
      \nz.mem_2460_sv2v_reg  <= w_data_i[860];
      \nz.mem_2459_sv2v_reg  <= w_data_i[859];
      \nz.mem_2458_sv2v_reg  <= w_data_i[858];
      \nz.mem_2457_sv2v_reg  <= w_data_i[857];
      \nz.mem_2456_sv2v_reg  <= w_data_i[856];
      \nz.mem_2455_sv2v_reg  <= w_data_i[855];
      \nz.mem_2454_sv2v_reg  <= w_data_i[854];
      \nz.mem_2453_sv2v_reg  <= w_data_i[853];
      \nz.mem_2452_sv2v_reg  <= w_data_i[852];
      \nz.mem_2451_sv2v_reg  <= w_data_i[851];
      \nz.mem_2450_sv2v_reg  <= w_data_i[850];
      \nz.mem_2449_sv2v_reg  <= w_data_i[849];
      \nz.mem_2448_sv2v_reg  <= w_data_i[848];
      \nz.mem_2447_sv2v_reg  <= w_data_i[847];
      \nz.mem_2446_sv2v_reg  <= w_data_i[846];
      \nz.mem_2445_sv2v_reg  <= w_data_i[845];
      \nz.mem_2444_sv2v_reg  <= w_data_i[844];
      \nz.mem_2443_sv2v_reg  <= w_data_i[843];
      \nz.mem_2442_sv2v_reg  <= w_data_i[842];
      \nz.mem_2441_sv2v_reg  <= w_data_i[841];
      \nz.mem_2440_sv2v_reg  <= w_data_i[840];
      \nz.mem_2439_sv2v_reg  <= w_data_i[839];
      \nz.mem_2438_sv2v_reg  <= w_data_i[838];
      \nz.mem_2437_sv2v_reg  <= w_data_i[837];
      \nz.mem_2436_sv2v_reg  <= w_data_i[836];
      \nz.mem_2435_sv2v_reg  <= w_data_i[835];
      \nz.mem_2434_sv2v_reg  <= w_data_i[834];
      \nz.mem_2433_sv2v_reg  <= w_data_i[833];
      \nz.mem_2432_sv2v_reg  <= w_data_i[832];
      \nz.mem_2431_sv2v_reg  <= w_data_i[831];
      \nz.mem_2430_sv2v_reg  <= w_data_i[830];
      \nz.mem_2429_sv2v_reg  <= w_data_i[829];
      \nz.mem_2428_sv2v_reg  <= w_data_i[828];
      \nz.mem_2427_sv2v_reg  <= w_data_i[827];
      \nz.mem_2426_sv2v_reg  <= w_data_i[826];
      \nz.mem_2425_sv2v_reg  <= w_data_i[825];
      \nz.mem_2424_sv2v_reg  <= w_data_i[824];
      \nz.mem_2423_sv2v_reg  <= w_data_i[823];
      \nz.mem_2422_sv2v_reg  <= w_data_i[822];
      \nz.mem_2421_sv2v_reg  <= w_data_i[821];
      \nz.mem_2420_sv2v_reg  <= w_data_i[820];
      \nz.mem_2419_sv2v_reg  <= w_data_i[819];
      \nz.mem_2418_sv2v_reg  <= w_data_i[818];
      \nz.mem_2417_sv2v_reg  <= w_data_i[817];
      \nz.mem_2416_sv2v_reg  <= w_data_i[816];
      \nz.mem_2415_sv2v_reg  <= w_data_i[815];
      \nz.mem_2414_sv2v_reg  <= w_data_i[814];
      \nz.mem_2413_sv2v_reg  <= w_data_i[813];
      \nz.mem_2412_sv2v_reg  <= w_data_i[812];
      \nz.mem_2411_sv2v_reg  <= w_data_i[811];
      \nz.mem_2410_sv2v_reg  <= w_data_i[810];
      \nz.mem_2409_sv2v_reg  <= w_data_i[809];
      \nz.mem_2408_sv2v_reg  <= w_data_i[808];
      \nz.mem_1607_sv2v_reg  <= w_data_i[7];
    end 
    if(N31) begin
      \nz.mem_2407_sv2v_reg  <= w_data_i[807];
      \nz.mem_2406_sv2v_reg  <= w_data_i[806];
      \nz.mem_2405_sv2v_reg  <= w_data_i[805];
      \nz.mem_2404_sv2v_reg  <= w_data_i[804];
      \nz.mem_2403_sv2v_reg  <= w_data_i[803];
      \nz.mem_2402_sv2v_reg  <= w_data_i[802];
      \nz.mem_2401_sv2v_reg  <= w_data_i[801];
      \nz.mem_2400_sv2v_reg  <= w_data_i[800];
      \nz.mem_2399_sv2v_reg  <= w_data_i[799];
      \nz.mem_2398_sv2v_reg  <= w_data_i[798];
      \nz.mem_2397_sv2v_reg  <= w_data_i[797];
      \nz.mem_2396_sv2v_reg  <= w_data_i[796];
      \nz.mem_2395_sv2v_reg  <= w_data_i[795];
      \nz.mem_2394_sv2v_reg  <= w_data_i[794];
      \nz.mem_2393_sv2v_reg  <= w_data_i[793];
      \nz.mem_2392_sv2v_reg  <= w_data_i[792];
      \nz.mem_2391_sv2v_reg  <= w_data_i[791];
      \nz.mem_2390_sv2v_reg  <= w_data_i[790];
      \nz.mem_2389_sv2v_reg  <= w_data_i[789];
      \nz.mem_2388_sv2v_reg  <= w_data_i[788];
      \nz.mem_2387_sv2v_reg  <= w_data_i[787];
      \nz.mem_2386_sv2v_reg  <= w_data_i[786];
      \nz.mem_2385_sv2v_reg  <= w_data_i[785];
      \nz.mem_2384_sv2v_reg  <= w_data_i[784];
      \nz.mem_2383_sv2v_reg  <= w_data_i[783];
      \nz.mem_2382_sv2v_reg  <= w_data_i[782];
      \nz.mem_2381_sv2v_reg  <= w_data_i[781];
      \nz.mem_2380_sv2v_reg  <= w_data_i[780];
      \nz.mem_2379_sv2v_reg  <= w_data_i[779];
      \nz.mem_2378_sv2v_reg  <= w_data_i[778];
      \nz.mem_2377_sv2v_reg  <= w_data_i[777];
      \nz.mem_2376_sv2v_reg  <= w_data_i[776];
      \nz.mem_2375_sv2v_reg  <= w_data_i[775];
      \nz.mem_2374_sv2v_reg  <= w_data_i[774];
      \nz.mem_2373_sv2v_reg  <= w_data_i[773];
      \nz.mem_2372_sv2v_reg  <= w_data_i[772];
      \nz.mem_2371_sv2v_reg  <= w_data_i[771];
      \nz.mem_2370_sv2v_reg  <= w_data_i[770];
      \nz.mem_2369_sv2v_reg  <= w_data_i[769];
      \nz.mem_2368_sv2v_reg  <= w_data_i[768];
      \nz.mem_2367_sv2v_reg  <= w_data_i[767];
      \nz.mem_2366_sv2v_reg  <= w_data_i[766];
      \nz.mem_2365_sv2v_reg  <= w_data_i[765];
      \nz.mem_2364_sv2v_reg  <= w_data_i[764];
      \nz.mem_2363_sv2v_reg  <= w_data_i[763];
      \nz.mem_2362_sv2v_reg  <= w_data_i[762];
      \nz.mem_2361_sv2v_reg  <= w_data_i[761];
      \nz.mem_2360_sv2v_reg  <= w_data_i[760];
      \nz.mem_2359_sv2v_reg  <= w_data_i[759];
      \nz.mem_2358_sv2v_reg  <= w_data_i[758];
      \nz.mem_2357_sv2v_reg  <= w_data_i[757];
      \nz.mem_2356_sv2v_reg  <= w_data_i[756];
      \nz.mem_2355_sv2v_reg  <= w_data_i[755];
      \nz.mem_2354_sv2v_reg  <= w_data_i[754];
      \nz.mem_2353_sv2v_reg  <= w_data_i[753];
      \nz.mem_2352_sv2v_reg  <= w_data_i[752];
      \nz.mem_2351_sv2v_reg  <= w_data_i[751];
      \nz.mem_2350_sv2v_reg  <= w_data_i[750];
      \nz.mem_2349_sv2v_reg  <= w_data_i[749];
      \nz.mem_2348_sv2v_reg  <= w_data_i[748];
      \nz.mem_2347_sv2v_reg  <= w_data_i[747];
      \nz.mem_2346_sv2v_reg  <= w_data_i[746];
      \nz.mem_2345_sv2v_reg  <= w_data_i[745];
      \nz.mem_2344_sv2v_reg  <= w_data_i[744];
      \nz.mem_2343_sv2v_reg  <= w_data_i[743];
      \nz.mem_2342_sv2v_reg  <= w_data_i[742];
      \nz.mem_2341_sv2v_reg  <= w_data_i[741];
      \nz.mem_2340_sv2v_reg  <= w_data_i[740];
      \nz.mem_2339_sv2v_reg  <= w_data_i[739];
      \nz.mem_2338_sv2v_reg  <= w_data_i[738];
      \nz.mem_2337_sv2v_reg  <= w_data_i[737];
      \nz.mem_2336_sv2v_reg  <= w_data_i[736];
      \nz.mem_2335_sv2v_reg  <= w_data_i[735];
      \nz.mem_2334_sv2v_reg  <= w_data_i[734];
      \nz.mem_2333_sv2v_reg  <= w_data_i[733];
      \nz.mem_2332_sv2v_reg  <= w_data_i[732];
      \nz.mem_2331_sv2v_reg  <= w_data_i[731];
      \nz.mem_2330_sv2v_reg  <= w_data_i[730];
      \nz.mem_2329_sv2v_reg  <= w_data_i[729];
      \nz.mem_2328_sv2v_reg  <= w_data_i[728];
      \nz.mem_2327_sv2v_reg  <= w_data_i[727];
      \nz.mem_2326_sv2v_reg  <= w_data_i[726];
      \nz.mem_2325_sv2v_reg  <= w_data_i[725];
      \nz.mem_2324_sv2v_reg  <= w_data_i[724];
      \nz.mem_2323_sv2v_reg  <= w_data_i[723];
      \nz.mem_2322_sv2v_reg  <= w_data_i[722];
      \nz.mem_2321_sv2v_reg  <= w_data_i[721];
      \nz.mem_2320_sv2v_reg  <= w_data_i[720];
      \nz.mem_2319_sv2v_reg  <= w_data_i[719];
      \nz.mem_2318_sv2v_reg  <= w_data_i[718];
      \nz.mem_2317_sv2v_reg  <= w_data_i[717];
      \nz.mem_2316_sv2v_reg  <= w_data_i[716];
      \nz.mem_2315_sv2v_reg  <= w_data_i[715];
      \nz.mem_2314_sv2v_reg  <= w_data_i[714];
      \nz.mem_2313_sv2v_reg  <= w_data_i[713];
      \nz.mem_2312_sv2v_reg  <= w_data_i[712];
      \nz.mem_2311_sv2v_reg  <= w_data_i[711];
      \nz.mem_2310_sv2v_reg  <= w_data_i[710];
      \nz.mem_2309_sv2v_reg  <= w_data_i[709];
      \nz.mem_1608_sv2v_reg  <= w_data_i[8];
    end 
    if(N32) begin
      \nz.mem_2308_sv2v_reg  <= w_data_i[708];
      \nz.mem_2307_sv2v_reg  <= w_data_i[707];
      \nz.mem_2306_sv2v_reg  <= w_data_i[706];
      \nz.mem_2305_sv2v_reg  <= w_data_i[705];
      \nz.mem_2304_sv2v_reg  <= w_data_i[704];
      \nz.mem_2303_sv2v_reg  <= w_data_i[703];
      \nz.mem_2302_sv2v_reg  <= w_data_i[702];
      \nz.mem_2301_sv2v_reg  <= w_data_i[701];
      \nz.mem_2300_sv2v_reg  <= w_data_i[700];
      \nz.mem_2299_sv2v_reg  <= w_data_i[699];
      \nz.mem_2298_sv2v_reg  <= w_data_i[698];
      \nz.mem_2297_sv2v_reg  <= w_data_i[697];
      \nz.mem_2296_sv2v_reg  <= w_data_i[696];
      \nz.mem_2295_sv2v_reg  <= w_data_i[695];
      \nz.mem_2294_sv2v_reg  <= w_data_i[694];
      \nz.mem_2293_sv2v_reg  <= w_data_i[693];
      \nz.mem_2292_sv2v_reg  <= w_data_i[692];
      \nz.mem_2291_sv2v_reg  <= w_data_i[691];
      \nz.mem_2290_sv2v_reg  <= w_data_i[690];
      \nz.mem_2289_sv2v_reg  <= w_data_i[689];
      \nz.mem_2288_sv2v_reg  <= w_data_i[688];
      \nz.mem_2287_sv2v_reg  <= w_data_i[687];
      \nz.mem_2286_sv2v_reg  <= w_data_i[686];
      \nz.mem_2285_sv2v_reg  <= w_data_i[685];
      \nz.mem_2284_sv2v_reg  <= w_data_i[684];
      \nz.mem_2283_sv2v_reg  <= w_data_i[683];
      \nz.mem_2282_sv2v_reg  <= w_data_i[682];
      \nz.mem_2281_sv2v_reg  <= w_data_i[681];
      \nz.mem_2280_sv2v_reg  <= w_data_i[680];
      \nz.mem_2279_sv2v_reg  <= w_data_i[679];
      \nz.mem_2278_sv2v_reg  <= w_data_i[678];
      \nz.mem_2277_sv2v_reg  <= w_data_i[677];
      \nz.mem_2276_sv2v_reg  <= w_data_i[676];
      \nz.mem_2275_sv2v_reg  <= w_data_i[675];
      \nz.mem_2274_sv2v_reg  <= w_data_i[674];
      \nz.mem_2273_sv2v_reg  <= w_data_i[673];
      \nz.mem_2272_sv2v_reg  <= w_data_i[672];
      \nz.mem_2271_sv2v_reg  <= w_data_i[671];
      \nz.mem_2270_sv2v_reg  <= w_data_i[670];
      \nz.mem_2269_sv2v_reg  <= w_data_i[669];
      \nz.mem_2268_sv2v_reg  <= w_data_i[668];
      \nz.mem_2267_sv2v_reg  <= w_data_i[667];
      \nz.mem_2266_sv2v_reg  <= w_data_i[666];
      \nz.mem_2265_sv2v_reg  <= w_data_i[665];
      \nz.mem_2264_sv2v_reg  <= w_data_i[664];
      \nz.mem_2263_sv2v_reg  <= w_data_i[663];
      \nz.mem_2262_sv2v_reg  <= w_data_i[662];
      \nz.mem_2261_sv2v_reg  <= w_data_i[661];
      \nz.mem_2260_sv2v_reg  <= w_data_i[660];
      \nz.mem_2259_sv2v_reg  <= w_data_i[659];
      \nz.mem_2258_sv2v_reg  <= w_data_i[658];
      \nz.mem_2257_sv2v_reg  <= w_data_i[657];
      \nz.mem_2256_sv2v_reg  <= w_data_i[656];
      \nz.mem_2255_sv2v_reg  <= w_data_i[655];
      \nz.mem_2254_sv2v_reg  <= w_data_i[654];
      \nz.mem_2253_sv2v_reg  <= w_data_i[653];
      \nz.mem_2252_sv2v_reg  <= w_data_i[652];
      \nz.mem_2251_sv2v_reg  <= w_data_i[651];
      \nz.mem_2250_sv2v_reg  <= w_data_i[650];
      \nz.mem_2249_sv2v_reg  <= w_data_i[649];
      \nz.mem_2248_sv2v_reg  <= w_data_i[648];
      \nz.mem_2247_sv2v_reg  <= w_data_i[647];
      \nz.mem_2246_sv2v_reg  <= w_data_i[646];
      \nz.mem_2245_sv2v_reg  <= w_data_i[645];
      \nz.mem_2244_sv2v_reg  <= w_data_i[644];
      \nz.mem_2243_sv2v_reg  <= w_data_i[643];
      \nz.mem_2242_sv2v_reg  <= w_data_i[642];
      \nz.mem_2241_sv2v_reg  <= w_data_i[641];
      \nz.mem_2240_sv2v_reg  <= w_data_i[640];
      \nz.mem_2239_sv2v_reg  <= w_data_i[639];
      \nz.mem_2238_sv2v_reg  <= w_data_i[638];
      \nz.mem_2237_sv2v_reg  <= w_data_i[637];
      \nz.mem_2236_sv2v_reg  <= w_data_i[636];
      \nz.mem_2235_sv2v_reg  <= w_data_i[635];
      \nz.mem_2234_sv2v_reg  <= w_data_i[634];
      \nz.mem_2233_sv2v_reg  <= w_data_i[633];
      \nz.mem_2232_sv2v_reg  <= w_data_i[632];
      \nz.mem_2231_sv2v_reg  <= w_data_i[631];
      \nz.mem_2230_sv2v_reg  <= w_data_i[630];
      \nz.mem_2229_sv2v_reg  <= w_data_i[629];
      \nz.mem_2228_sv2v_reg  <= w_data_i[628];
      \nz.mem_2227_sv2v_reg  <= w_data_i[627];
      \nz.mem_2226_sv2v_reg  <= w_data_i[626];
      \nz.mem_2225_sv2v_reg  <= w_data_i[625];
      \nz.mem_2224_sv2v_reg  <= w_data_i[624];
      \nz.mem_2223_sv2v_reg  <= w_data_i[623];
      \nz.mem_2222_sv2v_reg  <= w_data_i[622];
      \nz.mem_2221_sv2v_reg  <= w_data_i[621];
      \nz.mem_2220_sv2v_reg  <= w_data_i[620];
      \nz.mem_2219_sv2v_reg  <= w_data_i[619];
      \nz.mem_2218_sv2v_reg  <= w_data_i[618];
      \nz.mem_2217_sv2v_reg  <= w_data_i[617];
      \nz.mem_2216_sv2v_reg  <= w_data_i[616];
      \nz.mem_2215_sv2v_reg  <= w_data_i[615];
      \nz.mem_2214_sv2v_reg  <= w_data_i[614];
      \nz.mem_2213_sv2v_reg  <= w_data_i[613];
      \nz.mem_2212_sv2v_reg  <= w_data_i[612];
      \nz.mem_2211_sv2v_reg  <= w_data_i[611];
      \nz.mem_2210_sv2v_reg  <= w_data_i[610];
      \nz.mem_1609_sv2v_reg  <= w_data_i[9];
    end 
    if(N33) begin
      \nz.mem_2209_sv2v_reg  <= w_data_i[609];
      \nz.mem_2208_sv2v_reg  <= w_data_i[608];
      \nz.mem_2207_sv2v_reg  <= w_data_i[607];
      \nz.mem_2206_sv2v_reg  <= w_data_i[606];
      \nz.mem_2205_sv2v_reg  <= w_data_i[605];
      \nz.mem_2204_sv2v_reg  <= w_data_i[604];
      \nz.mem_2203_sv2v_reg  <= w_data_i[603];
      \nz.mem_2202_sv2v_reg  <= w_data_i[602];
      \nz.mem_2201_sv2v_reg  <= w_data_i[601];
      \nz.mem_2200_sv2v_reg  <= w_data_i[600];
      \nz.mem_2199_sv2v_reg  <= w_data_i[599];
      \nz.mem_2198_sv2v_reg  <= w_data_i[598];
      \nz.mem_2197_sv2v_reg  <= w_data_i[597];
      \nz.mem_2196_sv2v_reg  <= w_data_i[596];
      \nz.mem_2195_sv2v_reg  <= w_data_i[595];
      \nz.mem_2194_sv2v_reg  <= w_data_i[594];
      \nz.mem_2193_sv2v_reg  <= w_data_i[593];
      \nz.mem_2192_sv2v_reg  <= w_data_i[592];
      \nz.mem_2191_sv2v_reg  <= w_data_i[591];
      \nz.mem_2190_sv2v_reg  <= w_data_i[590];
      \nz.mem_2189_sv2v_reg  <= w_data_i[589];
      \nz.mem_2188_sv2v_reg  <= w_data_i[588];
      \nz.mem_2187_sv2v_reg  <= w_data_i[587];
      \nz.mem_2186_sv2v_reg  <= w_data_i[586];
      \nz.mem_2185_sv2v_reg  <= w_data_i[585];
      \nz.mem_2184_sv2v_reg  <= w_data_i[584];
      \nz.mem_2183_sv2v_reg  <= w_data_i[583];
      \nz.mem_2182_sv2v_reg  <= w_data_i[582];
      \nz.mem_2181_sv2v_reg  <= w_data_i[581];
      \nz.mem_2180_sv2v_reg  <= w_data_i[580];
      \nz.mem_2179_sv2v_reg  <= w_data_i[579];
      \nz.mem_2178_sv2v_reg  <= w_data_i[578];
      \nz.mem_2177_sv2v_reg  <= w_data_i[577];
      \nz.mem_2176_sv2v_reg  <= w_data_i[576];
      \nz.mem_2175_sv2v_reg  <= w_data_i[575];
      \nz.mem_2174_sv2v_reg  <= w_data_i[574];
      \nz.mem_2173_sv2v_reg  <= w_data_i[573];
      \nz.mem_2172_sv2v_reg  <= w_data_i[572];
      \nz.mem_2171_sv2v_reg  <= w_data_i[571];
      \nz.mem_2170_sv2v_reg  <= w_data_i[570];
      \nz.mem_2169_sv2v_reg  <= w_data_i[569];
      \nz.mem_2168_sv2v_reg  <= w_data_i[568];
      \nz.mem_2167_sv2v_reg  <= w_data_i[567];
      \nz.mem_2166_sv2v_reg  <= w_data_i[566];
      \nz.mem_2165_sv2v_reg  <= w_data_i[565];
      \nz.mem_2164_sv2v_reg  <= w_data_i[564];
      \nz.mem_2163_sv2v_reg  <= w_data_i[563];
      \nz.mem_2162_sv2v_reg  <= w_data_i[562];
      \nz.mem_2161_sv2v_reg  <= w_data_i[561];
      \nz.mem_2160_sv2v_reg  <= w_data_i[560];
      \nz.mem_2159_sv2v_reg  <= w_data_i[559];
      \nz.mem_2158_sv2v_reg  <= w_data_i[558];
      \nz.mem_2157_sv2v_reg  <= w_data_i[557];
      \nz.mem_2156_sv2v_reg  <= w_data_i[556];
      \nz.mem_2155_sv2v_reg  <= w_data_i[555];
      \nz.mem_2154_sv2v_reg  <= w_data_i[554];
      \nz.mem_2153_sv2v_reg  <= w_data_i[553];
      \nz.mem_2152_sv2v_reg  <= w_data_i[552];
      \nz.mem_2151_sv2v_reg  <= w_data_i[551];
      \nz.mem_2150_sv2v_reg  <= w_data_i[550];
      \nz.mem_2149_sv2v_reg  <= w_data_i[549];
      \nz.mem_2148_sv2v_reg  <= w_data_i[548];
      \nz.mem_2147_sv2v_reg  <= w_data_i[547];
      \nz.mem_2146_sv2v_reg  <= w_data_i[546];
      \nz.mem_2145_sv2v_reg  <= w_data_i[545];
      \nz.mem_2144_sv2v_reg  <= w_data_i[544];
      \nz.mem_2143_sv2v_reg  <= w_data_i[543];
      \nz.mem_2142_sv2v_reg  <= w_data_i[542];
      \nz.mem_2141_sv2v_reg  <= w_data_i[541];
      \nz.mem_2140_sv2v_reg  <= w_data_i[540];
      \nz.mem_2139_sv2v_reg  <= w_data_i[539];
      \nz.mem_2138_sv2v_reg  <= w_data_i[538];
      \nz.mem_2137_sv2v_reg  <= w_data_i[537];
      \nz.mem_2136_sv2v_reg  <= w_data_i[536];
      \nz.mem_2135_sv2v_reg  <= w_data_i[535];
      \nz.mem_2134_sv2v_reg  <= w_data_i[534];
      \nz.mem_2133_sv2v_reg  <= w_data_i[533];
      \nz.mem_2132_sv2v_reg  <= w_data_i[532];
      \nz.mem_2131_sv2v_reg  <= w_data_i[531];
      \nz.mem_2130_sv2v_reg  <= w_data_i[530];
      \nz.mem_2129_sv2v_reg  <= w_data_i[529];
      \nz.mem_2128_sv2v_reg  <= w_data_i[528];
      \nz.mem_2127_sv2v_reg  <= w_data_i[527];
      \nz.mem_2126_sv2v_reg  <= w_data_i[526];
      \nz.mem_2125_sv2v_reg  <= w_data_i[525];
      \nz.mem_2124_sv2v_reg  <= w_data_i[524];
      \nz.mem_2123_sv2v_reg  <= w_data_i[523];
      \nz.mem_2122_sv2v_reg  <= w_data_i[522];
      \nz.mem_2121_sv2v_reg  <= w_data_i[521];
      \nz.mem_2120_sv2v_reg  <= w_data_i[520];
      \nz.mem_2119_sv2v_reg  <= w_data_i[519];
      \nz.mem_2118_sv2v_reg  <= w_data_i[518];
      \nz.mem_2117_sv2v_reg  <= w_data_i[517];
      \nz.mem_2116_sv2v_reg  <= w_data_i[516];
      \nz.mem_2115_sv2v_reg  <= w_data_i[515];
      \nz.mem_2114_sv2v_reg  <= w_data_i[514];
      \nz.mem_2113_sv2v_reg  <= w_data_i[513];
      \nz.mem_2112_sv2v_reg  <= w_data_i[512];
      \nz.mem_2111_sv2v_reg  <= w_data_i[511];
      \nz.mem_1610_sv2v_reg  <= w_data_i[10];
    end 
    if(N34) begin
      \nz.mem_2110_sv2v_reg  <= w_data_i[510];
      \nz.mem_2109_sv2v_reg  <= w_data_i[509];
      \nz.mem_2108_sv2v_reg  <= w_data_i[508];
      \nz.mem_2107_sv2v_reg  <= w_data_i[507];
      \nz.mem_2106_sv2v_reg  <= w_data_i[506];
      \nz.mem_2105_sv2v_reg  <= w_data_i[505];
      \nz.mem_2104_sv2v_reg  <= w_data_i[504];
      \nz.mem_2103_sv2v_reg  <= w_data_i[503];
      \nz.mem_2102_sv2v_reg  <= w_data_i[502];
      \nz.mem_2101_sv2v_reg  <= w_data_i[501];
      \nz.mem_2100_sv2v_reg  <= w_data_i[500];
      \nz.mem_2099_sv2v_reg  <= w_data_i[499];
      \nz.mem_2098_sv2v_reg  <= w_data_i[498];
      \nz.mem_2097_sv2v_reg  <= w_data_i[497];
      \nz.mem_2096_sv2v_reg  <= w_data_i[496];
      \nz.mem_2095_sv2v_reg  <= w_data_i[495];
      \nz.mem_2094_sv2v_reg  <= w_data_i[494];
      \nz.mem_2093_sv2v_reg  <= w_data_i[493];
      \nz.mem_2092_sv2v_reg  <= w_data_i[492];
      \nz.mem_2091_sv2v_reg  <= w_data_i[491];
      \nz.mem_2090_sv2v_reg  <= w_data_i[490];
      \nz.mem_2089_sv2v_reg  <= w_data_i[489];
      \nz.mem_2088_sv2v_reg  <= w_data_i[488];
      \nz.mem_2087_sv2v_reg  <= w_data_i[487];
      \nz.mem_2086_sv2v_reg  <= w_data_i[486];
      \nz.mem_2085_sv2v_reg  <= w_data_i[485];
      \nz.mem_2084_sv2v_reg  <= w_data_i[484];
      \nz.mem_2083_sv2v_reg  <= w_data_i[483];
      \nz.mem_2082_sv2v_reg  <= w_data_i[482];
      \nz.mem_2081_sv2v_reg  <= w_data_i[481];
      \nz.mem_2080_sv2v_reg  <= w_data_i[480];
      \nz.mem_2079_sv2v_reg  <= w_data_i[479];
      \nz.mem_2078_sv2v_reg  <= w_data_i[478];
      \nz.mem_2077_sv2v_reg  <= w_data_i[477];
      \nz.mem_2076_sv2v_reg  <= w_data_i[476];
      \nz.mem_2075_sv2v_reg  <= w_data_i[475];
      \nz.mem_2074_sv2v_reg  <= w_data_i[474];
      \nz.mem_2073_sv2v_reg  <= w_data_i[473];
      \nz.mem_2072_sv2v_reg  <= w_data_i[472];
      \nz.mem_2071_sv2v_reg  <= w_data_i[471];
      \nz.mem_2070_sv2v_reg  <= w_data_i[470];
      \nz.mem_2069_sv2v_reg  <= w_data_i[469];
      \nz.mem_2068_sv2v_reg  <= w_data_i[468];
      \nz.mem_2067_sv2v_reg  <= w_data_i[467];
      \nz.mem_2066_sv2v_reg  <= w_data_i[466];
      \nz.mem_2065_sv2v_reg  <= w_data_i[465];
      \nz.mem_2064_sv2v_reg  <= w_data_i[464];
      \nz.mem_2063_sv2v_reg  <= w_data_i[463];
      \nz.mem_2062_sv2v_reg  <= w_data_i[462];
      \nz.mem_2061_sv2v_reg  <= w_data_i[461];
      \nz.mem_2060_sv2v_reg  <= w_data_i[460];
      \nz.mem_2059_sv2v_reg  <= w_data_i[459];
      \nz.mem_2058_sv2v_reg  <= w_data_i[458];
      \nz.mem_2057_sv2v_reg  <= w_data_i[457];
      \nz.mem_2056_sv2v_reg  <= w_data_i[456];
      \nz.mem_2055_sv2v_reg  <= w_data_i[455];
      \nz.mem_2054_sv2v_reg  <= w_data_i[454];
      \nz.mem_2053_sv2v_reg  <= w_data_i[453];
      \nz.mem_2052_sv2v_reg  <= w_data_i[452];
      \nz.mem_2051_sv2v_reg  <= w_data_i[451];
      \nz.mem_2050_sv2v_reg  <= w_data_i[450];
      \nz.mem_2049_sv2v_reg  <= w_data_i[449];
      \nz.mem_2048_sv2v_reg  <= w_data_i[448];
      \nz.mem_2047_sv2v_reg  <= w_data_i[447];
      \nz.mem_2046_sv2v_reg  <= w_data_i[446];
      \nz.mem_2045_sv2v_reg  <= w_data_i[445];
      \nz.mem_2044_sv2v_reg  <= w_data_i[444];
      \nz.mem_2043_sv2v_reg  <= w_data_i[443];
      \nz.mem_2042_sv2v_reg  <= w_data_i[442];
      \nz.mem_2041_sv2v_reg  <= w_data_i[441];
      \nz.mem_2040_sv2v_reg  <= w_data_i[440];
      \nz.mem_2039_sv2v_reg  <= w_data_i[439];
      \nz.mem_2038_sv2v_reg  <= w_data_i[438];
      \nz.mem_2037_sv2v_reg  <= w_data_i[437];
      \nz.mem_2036_sv2v_reg  <= w_data_i[436];
      \nz.mem_2035_sv2v_reg  <= w_data_i[435];
      \nz.mem_2034_sv2v_reg  <= w_data_i[434];
      \nz.mem_2033_sv2v_reg  <= w_data_i[433];
      \nz.mem_2032_sv2v_reg  <= w_data_i[432];
      \nz.mem_2031_sv2v_reg  <= w_data_i[431];
      \nz.mem_2030_sv2v_reg  <= w_data_i[430];
      \nz.mem_2029_sv2v_reg  <= w_data_i[429];
      \nz.mem_2028_sv2v_reg  <= w_data_i[428];
      \nz.mem_2027_sv2v_reg  <= w_data_i[427];
      \nz.mem_2026_sv2v_reg  <= w_data_i[426];
      \nz.mem_2025_sv2v_reg  <= w_data_i[425];
      \nz.mem_2024_sv2v_reg  <= w_data_i[424];
      \nz.mem_2023_sv2v_reg  <= w_data_i[423];
      \nz.mem_2022_sv2v_reg  <= w_data_i[422];
      \nz.mem_2021_sv2v_reg  <= w_data_i[421];
      \nz.mem_2020_sv2v_reg  <= w_data_i[420];
      \nz.mem_2019_sv2v_reg  <= w_data_i[419];
      \nz.mem_2018_sv2v_reg  <= w_data_i[418];
      \nz.mem_2017_sv2v_reg  <= w_data_i[417];
      \nz.mem_2016_sv2v_reg  <= w_data_i[416];
      \nz.mem_2015_sv2v_reg  <= w_data_i[415];
      \nz.mem_2014_sv2v_reg  <= w_data_i[414];
      \nz.mem_2013_sv2v_reg  <= w_data_i[413];
      \nz.mem_2012_sv2v_reg  <= w_data_i[412];
      \nz.mem_1611_sv2v_reg  <= w_data_i[11];
    end 
    if(N35) begin
      \nz.mem_2011_sv2v_reg  <= w_data_i[411];
      \nz.mem_2010_sv2v_reg  <= w_data_i[410];
      \nz.mem_2009_sv2v_reg  <= w_data_i[409];
      \nz.mem_2008_sv2v_reg  <= w_data_i[408];
      \nz.mem_2007_sv2v_reg  <= w_data_i[407];
      \nz.mem_2006_sv2v_reg  <= w_data_i[406];
      \nz.mem_2005_sv2v_reg  <= w_data_i[405];
      \nz.mem_2004_sv2v_reg  <= w_data_i[404];
      \nz.mem_2003_sv2v_reg  <= w_data_i[403];
      \nz.mem_2002_sv2v_reg  <= w_data_i[402];
      \nz.mem_2001_sv2v_reg  <= w_data_i[401];
      \nz.mem_2000_sv2v_reg  <= w_data_i[400];
      \nz.mem_1999_sv2v_reg  <= w_data_i[399];
      \nz.mem_1998_sv2v_reg  <= w_data_i[398];
      \nz.mem_1997_sv2v_reg  <= w_data_i[397];
      \nz.mem_1996_sv2v_reg  <= w_data_i[396];
      \nz.mem_1995_sv2v_reg  <= w_data_i[395];
      \nz.mem_1994_sv2v_reg  <= w_data_i[394];
      \nz.mem_1993_sv2v_reg  <= w_data_i[393];
      \nz.mem_1992_sv2v_reg  <= w_data_i[392];
      \nz.mem_1991_sv2v_reg  <= w_data_i[391];
      \nz.mem_1990_sv2v_reg  <= w_data_i[390];
      \nz.mem_1989_sv2v_reg  <= w_data_i[389];
      \nz.mem_1988_sv2v_reg  <= w_data_i[388];
      \nz.mem_1987_sv2v_reg  <= w_data_i[387];
      \nz.mem_1986_sv2v_reg  <= w_data_i[386];
      \nz.mem_1985_sv2v_reg  <= w_data_i[385];
      \nz.mem_1984_sv2v_reg  <= w_data_i[384];
      \nz.mem_1983_sv2v_reg  <= w_data_i[383];
      \nz.mem_1982_sv2v_reg  <= w_data_i[382];
      \nz.mem_1981_sv2v_reg  <= w_data_i[381];
      \nz.mem_1980_sv2v_reg  <= w_data_i[380];
      \nz.mem_1979_sv2v_reg  <= w_data_i[379];
      \nz.mem_1978_sv2v_reg  <= w_data_i[378];
      \nz.mem_1977_sv2v_reg  <= w_data_i[377];
      \nz.mem_1976_sv2v_reg  <= w_data_i[376];
      \nz.mem_1975_sv2v_reg  <= w_data_i[375];
      \nz.mem_1974_sv2v_reg  <= w_data_i[374];
      \nz.mem_1973_sv2v_reg  <= w_data_i[373];
      \nz.mem_1972_sv2v_reg  <= w_data_i[372];
      \nz.mem_1971_sv2v_reg  <= w_data_i[371];
      \nz.mem_1970_sv2v_reg  <= w_data_i[370];
      \nz.mem_1969_sv2v_reg  <= w_data_i[369];
      \nz.mem_1968_sv2v_reg  <= w_data_i[368];
      \nz.mem_1967_sv2v_reg  <= w_data_i[367];
      \nz.mem_1966_sv2v_reg  <= w_data_i[366];
      \nz.mem_1965_sv2v_reg  <= w_data_i[365];
      \nz.mem_1964_sv2v_reg  <= w_data_i[364];
      \nz.mem_1963_sv2v_reg  <= w_data_i[363];
      \nz.mem_1962_sv2v_reg  <= w_data_i[362];
      \nz.mem_1961_sv2v_reg  <= w_data_i[361];
      \nz.mem_1960_sv2v_reg  <= w_data_i[360];
      \nz.mem_1959_sv2v_reg  <= w_data_i[359];
      \nz.mem_1958_sv2v_reg  <= w_data_i[358];
      \nz.mem_1957_sv2v_reg  <= w_data_i[357];
      \nz.mem_1956_sv2v_reg  <= w_data_i[356];
      \nz.mem_1955_sv2v_reg  <= w_data_i[355];
      \nz.mem_1954_sv2v_reg  <= w_data_i[354];
      \nz.mem_1953_sv2v_reg  <= w_data_i[353];
      \nz.mem_1952_sv2v_reg  <= w_data_i[352];
      \nz.mem_1951_sv2v_reg  <= w_data_i[351];
      \nz.mem_1950_sv2v_reg  <= w_data_i[350];
      \nz.mem_1949_sv2v_reg  <= w_data_i[349];
      \nz.mem_1948_sv2v_reg  <= w_data_i[348];
      \nz.mem_1947_sv2v_reg  <= w_data_i[347];
      \nz.mem_1946_sv2v_reg  <= w_data_i[346];
      \nz.mem_1945_sv2v_reg  <= w_data_i[345];
      \nz.mem_1944_sv2v_reg  <= w_data_i[344];
      \nz.mem_1943_sv2v_reg  <= w_data_i[343];
      \nz.mem_1942_sv2v_reg  <= w_data_i[342];
      \nz.mem_1941_sv2v_reg  <= w_data_i[341];
      \nz.mem_1940_sv2v_reg  <= w_data_i[340];
      \nz.mem_1939_sv2v_reg  <= w_data_i[339];
      \nz.mem_1938_sv2v_reg  <= w_data_i[338];
      \nz.mem_1937_sv2v_reg  <= w_data_i[337];
      \nz.mem_1936_sv2v_reg  <= w_data_i[336];
      \nz.mem_1935_sv2v_reg  <= w_data_i[335];
      \nz.mem_1934_sv2v_reg  <= w_data_i[334];
      \nz.mem_1933_sv2v_reg  <= w_data_i[333];
      \nz.mem_1932_sv2v_reg  <= w_data_i[332];
      \nz.mem_1931_sv2v_reg  <= w_data_i[331];
      \nz.mem_1930_sv2v_reg  <= w_data_i[330];
      \nz.mem_1929_sv2v_reg  <= w_data_i[329];
      \nz.mem_1928_sv2v_reg  <= w_data_i[328];
      \nz.mem_1927_sv2v_reg  <= w_data_i[327];
      \nz.mem_1926_sv2v_reg  <= w_data_i[326];
      \nz.mem_1925_sv2v_reg  <= w_data_i[325];
      \nz.mem_1924_sv2v_reg  <= w_data_i[324];
      \nz.mem_1923_sv2v_reg  <= w_data_i[323];
      \nz.mem_1922_sv2v_reg  <= w_data_i[322];
      \nz.mem_1921_sv2v_reg  <= w_data_i[321];
      \nz.mem_1920_sv2v_reg  <= w_data_i[320];
      \nz.mem_1919_sv2v_reg  <= w_data_i[319];
      \nz.mem_1918_sv2v_reg  <= w_data_i[318];
      \nz.mem_1917_sv2v_reg  <= w_data_i[317];
      \nz.mem_1916_sv2v_reg  <= w_data_i[316];
      \nz.mem_1915_sv2v_reg  <= w_data_i[315];
      \nz.mem_1914_sv2v_reg  <= w_data_i[314];
      \nz.mem_1913_sv2v_reg  <= w_data_i[313];
      \nz.mem_1612_sv2v_reg  <= w_data_i[12];
    end 
    if(N36) begin
      \nz.mem_1912_sv2v_reg  <= w_data_i[312];
      \nz.mem_1911_sv2v_reg  <= w_data_i[311];
      \nz.mem_1910_sv2v_reg  <= w_data_i[310];
      \nz.mem_1909_sv2v_reg  <= w_data_i[309];
      \nz.mem_1908_sv2v_reg  <= w_data_i[308];
      \nz.mem_1907_sv2v_reg  <= w_data_i[307];
      \nz.mem_1906_sv2v_reg  <= w_data_i[306];
      \nz.mem_1905_sv2v_reg  <= w_data_i[305];
      \nz.mem_1904_sv2v_reg  <= w_data_i[304];
      \nz.mem_1903_sv2v_reg  <= w_data_i[303];
      \nz.mem_1902_sv2v_reg  <= w_data_i[302];
      \nz.mem_1901_sv2v_reg  <= w_data_i[301];
      \nz.mem_1900_sv2v_reg  <= w_data_i[300];
      \nz.mem_1899_sv2v_reg  <= w_data_i[299];
      \nz.mem_1898_sv2v_reg  <= w_data_i[298];
      \nz.mem_1897_sv2v_reg  <= w_data_i[297];
      \nz.mem_1896_sv2v_reg  <= w_data_i[296];
      \nz.mem_1895_sv2v_reg  <= w_data_i[295];
      \nz.mem_1894_sv2v_reg  <= w_data_i[294];
      \nz.mem_1893_sv2v_reg  <= w_data_i[293];
      \nz.mem_1892_sv2v_reg  <= w_data_i[292];
      \nz.mem_1891_sv2v_reg  <= w_data_i[291];
      \nz.mem_1890_sv2v_reg  <= w_data_i[290];
      \nz.mem_1889_sv2v_reg  <= w_data_i[289];
      \nz.mem_1888_sv2v_reg  <= w_data_i[288];
      \nz.mem_1887_sv2v_reg  <= w_data_i[287];
      \nz.mem_1886_sv2v_reg  <= w_data_i[286];
      \nz.mem_1885_sv2v_reg  <= w_data_i[285];
      \nz.mem_1884_sv2v_reg  <= w_data_i[284];
      \nz.mem_1883_sv2v_reg  <= w_data_i[283];
      \nz.mem_1882_sv2v_reg  <= w_data_i[282];
      \nz.mem_1881_sv2v_reg  <= w_data_i[281];
      \nz.mem_1880_sv2v_reg  <= w_data_i[280];
      \nz.mem_1879_sv2v_reg  <= w_data_i[279];
      \nz.mem_1878_sv2v_reg  <= w_data_i[278];
      \nz.mem_1877_sv2v_reg  <= w_data_i[277];
      \nz.mem_1876_sv2v_reg  <= w_data_i[276];
      \nz.mem_1875_sv2v_reg  <= w_data_i[275];
      \nz.mem_1874_sv2v_reg  <= w_data_i[274];
      \nz.mem_1873_sv2v_reg  <= w_data_i[273];
      \nz.mem_1872_sv2v_reg  <= w_data_i[272];
      \nz.mem_1871_sv2v_reg  <= w_data_i[271];
      \nz.mem_1870_sv2v_reg  <= w_data_i[270];
      \nz.mem_1869_sv2v_reg  <= w_data_i[269];
      \nz.mem_1868_sv2v_reg  <= w_data_i[268];
      \nz.mem_1867_sv2v_reg  <= w_data_i[267];
      \nz.mem_1866_sv2v_reg  <= w_data_i[266];
      \nz.mem_1865_sv2v_reg  <= w_data_i[265];
      \nz.mem_1864_sv2v_reg  <= w_data_i[264];
      \nz.mem_1863_sv2v_reg  <= w_data_i[263];
      \nz.mem_1862_sv2v_reg  <= w_data_i[262];
      \nz.mem_1861_sv2v_reg  <= w_data_i[261];
      \nz.mem_1860_sv2v_reg  <= w_data_i[260];
      \nz.mem_1859_sv2v_reg  <= w_data_i[259];
      \nz.mem_1858_sv2v_reg  <= w_data_i[258];
      \nz.mem_1857_sv2v_reg  <= w_data_i[257];
      \nz.mem_1856_sv2v_reg  <= w_data_i[256];
      \nz.mem_1855_sv2v_reg  <= w_data_i[255];
      \nz.mem_1854_sv2v_reg  <= w_data_i[254];
      \nz.mem_1853_sv2v_reg  <= w_data_i[253];
      \nz.mem_1852_sv2v_reg  <= w_data_i[252];
      \nz.mem_1851_sv2v_reg  <= w_data_i[251];
      \nz.mem_1850_sv2v_reg  <= w_data_i[250];
      \nz.mem_1849_sv2v_reg  <= w_data_i[249];
      \nz.mem_1848_sv2v_reg  <= w_data_i[248];
      \nz.mem_1847_sv2v_reg  <= w_data_i[247];
      \nz.mem_1846_sv2v_reg  <= w_data_i[246];
      \nz.mem_1845_sv2v_reg  <= w_data_i[245];
      \nz.mem_1844_sv2v_reg  <= w_data_i[244];
      \nz.mem_1843_sv2v_reg  <= w_data_i[243];
      \nz.mem_1842_sv2v_reg  <= w_data_i[242];
      \nz.mem_1841_sv2v_reg  <= w_data_i[241];
      \nz.mem_1840_sv2v_reg  <= w_data_i[240];
      \nz.mem_1839_sv2v_reg  <= w_data_i[239];
      \nz.mem_1838_sv2v_reg  <= w_data_i[238];
      \nz.mem_1837_sv2v_reg  <= w_data_i[237];
      \nz.mem_1836_sv2v_reg  <= w_data_i[236];
      \nz.mem_1835_sv2v_reg  <= w_data_i[235];
      \nz.mem_1834_sv2v_reg  <= w_data_i[234];
      \nz.mem_1833_sv2v_reg  <= w_data_i[233];
      \nz.mem_1832_sv2v_reg  <= w_data_i[232];
      \nz.mem_1831_sv2v_reg  <= w_data_i[231];
      \nz.mem_1830_sv2v_reg  <= w_data_i[230];
      \nz.mem_1829_sv2v_reg  <= w_data_i[229];
      \nz.mem_1828_sv2v_reg  <= w_data_i[228];
      \nz.mem_1827_sv2v_reg  <= w_data_i[227];
      \nz.mem_1826_sv2v_reg  <= w_data_i[226];
      \nz.mem_1825_sv2v_reg  <= w_data_i[225];
      \nz.mem_1824_sv2v_reg  <= w_data_i[224];
      \nz.mem_1823_sv2v_reg  <= w_data_i[223];
      \nz.mem_1822_sv2v_reg  <= w_data_i[222];
      \nz.mem_1821_sv2v_reg  <= w_data_i[221];
      \nz.mem_1820_sv2v_reg  <= w_data_i[220];
      \nz.mem_1819_sv2v_reg  <= w_data_i[219];
      \nz.mem_1818_sv2v_reg  <= w_data_i[218];
      \nz.mem_1817_sv2v_reg  <= w_data_i[217];
      \nz.mem_1816_sv2v_reg  <= w_data_i[216];
      \nz.mem_1815_sv2v_reg  <= w_data_i[215];
      \nz.mem_1814_sv2v_reg  <= w_data_i[214];
      \nz.mem_1613_sv2v_reg  <= w_data_i[13];
    end 
    if(N37) begin
      \nz.mem_1813_sv2v_reg  <= w_data_i[213];
      \nz.mem_1812_sv2v_reg  <= w_data_i[212];
      \nz.mem_1811_sv2v_reg  <= w_data_i[211];
      \nz.mem_1810_sv2v_reg  <= w_data_i[210];
      \nz.mem_1809_sv2v_reg  <= w_data_i[209];
      \nz.mem_1808_sv2v_reg  <= w_data_i[208];
      \nz.mem_1807_sv2v_reg  <= w_data_i[207];
      \nz.mem_1806_sv2v_reg  <= w_data_i[206];
      \nz.mem_1805_sv2v_reg  <= w_data_i[205];
      \nz.mem_1804_sv2v_reg  <= w_data_i[204];
      \nz.mem_1803_sv2v_reg  <= w_data_i[203];
      \nz.mem_1802_sv2v_reg  <= w_data_i[202];
      \nz.mem_1801_sv2v_reg  <= w_data_i[201];
      \nz.mem_1800_sv2v_reg  <= w_data_i[200];
      \nz.mem_1799_sv2v_reg  <= w_data_i[199];
      \nz.mem_1798_sv2v_reg  <= w_data_i[198];
      \nz.mem_1797_sv2v_reg  <= w_data_i[197];
      \nz.mem_1796_sv2v_reg  <= w_data_i[196];
      \nz.mem_1795_sv2v_reg  <= w_data_i[195];
      \nz.mem_1794_sv2v_reg  <= w_data_i[194];
      \nz.mem_1793_sv2v_reg  <= w_data_i[193];
      \nz.mem_1792_sv2v_reg  <= w_data_i[192];
      \nz.mem_1791_sv2v_reg  <= w_data_i[191];
      \nz.mem_1790_sv2v_reg  <= w_data_i[190];
      \nz.mem_1789_sv2v_reg  <= w_data_i[189];
      \nz.mem_1788_sv2v_reg  <= w_data_i[188];
      \nz.mem_1787_sv2v_reg  <= w_data_i[187];
      \nz.mem_1786_sv2v_reg  <= w_data_i[186];
      \nz.mem_1785_sv2v_reg  <= w_data_i[185];
      \nz.mem_1784_sv2v_reg  <= w_data_i[184];
      \nz.mem_1783_sv2v_reg  <= w_data_i[183];
      \nz.mem_1782_sv2v_reg  <= w_data_i[182];
      \nz.mem_1781_sv2v_reg  <= w_data_i[181];
      \nz.mem_1780_sv2v_reg  <= w_data_i[180];
      \nz.mem_1779_sv2v_reg  <= w_data_i[179];
      \nz.mem_1778_sv2v_reg  <= w_data_i[178];
      \nz.mem_1777_sv2v_reg  <= w_data_i[177];
      \nz.mem_1776_sv2v_reg  <= w_data_i[176];
      \nz.mem_1775_sv2v_reg  <= w_data_i[175];
      \nz.mem_1774_sv2v_reg  <= w_data_i[174];
      \nz.mem_1773_sv2v_reg  <= w_data_i[173];
      \nz.mem_1772_sv2v_reg  <= w_data_i[172];
      \nz.mem_1771_sv2v_reg  <= w_data_i[171];
      \nz.mem_1770_sv2v_reg  <= w_data_i[170];
      \nz.mem_1769_sv2v_reg  <= w_data_i[169];
      \nz.mem_1768_sv2v_reg  <= w_data_i[168];
      \nz.mem_1767_sv2v_reg  <= w_data_i[167];
      \nz.mem_1766_sv2v_reg  <= w_data_i[166];
      \nz.mem_1765_sv2v_reg  <= w_data_i[165];
      \nz.mem_1764_sv2v_reg  <= w_data_i[164];
      \nz.mem_1763_sv2v_reg  <= w_data_i[163];
      \nz.mem_1762_sv2v_reg  <= w_data_i[162];
      \nz.mem_1761_sv2v_reg  <= w_data_i[161];
      \nz.mem_1760_sv2v_reg  <= w_data_i[160];
      \nz.mem_1759_sv2v_reg  <= w_data_i[159];
      \nz.mem_1758_sv2v_reg  <= w_data_i[158];
      \nz.mem_1757_sv2v_reg  <= w_data_i[157];
      \nz.mem_1756_sv2v_reg  <= w_data_i[156];
      \nz.mem_1755_sv2v_reg  <= w_data_i[155];
      \nz.mem_1754_sv2v_reg  <= w_data_i[154];
      \nz.mem_1753_sv2v_reg  <= w_data_i[153];
      \nz.mem_1752_sv2v_reg  <= w_data_i[152];
      \nz.mem_1751_sv2v_reg  <= w_data_i[151];
      \nz.mem_1750_sv2v_reg  <= w_data_i[150];
      \nz.mem_1749_sv2v_reg  <= w_data_i[149];
      \nz.mem_1748_sv2v_reg  <= w_data_i[148];
      \nz.mem_1747_sv2v_reg  <= w_data_i[147];
      \nz.mem_1746_sv2v_reg  <= w_data_i[146];
      \nz.mem_1745_sv2v_reg  <= w_data_i[145];
      \nz.mem_1744_sv2v_reg  <= w_data_i[144];
      \nz.mem_1743_sv2v_reg  <= w_data_i[143];
      \nz.mem_1742_sv2v_reg  <= w_data_i[142];
      \nz.mem_1741_sv2v_reg  <= w_data_i[141];
      \nz.mem_1740_sv2v_reg  <= w_data_i[140];
      \nz.mem_1739_sv2v_reg  <= w_data_i[139];
      \nz.mem_1738_sv2v_reg  <= w_data_i[138];
      \nz.mem_1737_sv2v_reg  <= w_data_i[137];
      \nz.mem_1736_sv2v_reg  <= w_data_i[136];
      \nz.mem_1735_sv2v_reg  <= w_data_i[135];
      \nz.mem_1734_sv2v_reg  <= w_data_i[134];
      \nz.mem_1733_sv2v_reg  <= w_data_i[133];
      \nz.mem_1732_sv2v_reg  <= w_data_i[132];
      \nz.mem_1731_sv2v_reg  <= w_data_i[131];
      \nz.mem_1730_sv2v_reg  <= w_data_i[130];
      \nz.mem_1729_sv2v_reg  <= w_data_i[129];
      \nz.mem_1728_sv2v_reg  <= w_data_i[128];
      \nz.mem_1727_sv2v_reg  <= w_data_i[127];
      \nz.mem_1726_sv2v_reg  <= w_data_i[126];
      \nz.mem_1725_sv2v_reg  <= w_data_i[125];
      \nz.mem_1724_sv2v_reg  <= w_data_i[124];
      \nz.mem_1723_sv2v_reg  <= w_data_i[123];
      \nz.mem_1722_sv2v_reg  <= w_data_i[122];
      \nz.mem_1721_sv2v_reg  <= w_data_i[121];
      \nz.mem_1720_sv2v_reg  <= w_data_i[120];
      \nz.mem_1719_sv2v_reg  <= w_data_i[119];
      \nz.mem_1718_sv2v_reg  <= w_data_i[118];
      \nz.mem_1717_sv2v_reg  <= w_data_i[117];
      \nz.mem_1716_sv2v_reg  <= w_data_i[116];
      \nz.mem_1715_sv2v_reg  <= w_data_i[115];
      \nz.mem_1614_sv2v_reg  <= w_data_i[14];
    end 
    if(N38) begin
      \nz.mem_1714_sv2v_reg  <= w_data_i[114];
      \nz.mem_1713_sv2v_reg  <= w_data_i[113];
      \nz.mem_1712_sv2v_reg  <= w_data_i[112];
      \nz.mem_1711_sv2v_reg  <= w_data_i[111];
      \nz.mem_1710_sv2v_reg  <= w_data_i[110];
      \nz.mem_1709_sv2v_reg  <= w_data_i[109];
      \nz.mem_1708_sv2v_reg  <= w_data_i[108];
      \nz.mem_1707_sv2v_reg  <= w_data_i[107];
      \nz.mem_1706_sv2v_reg  <= w_data_i[106];
      \nz.mem_1705_sv2v_reg  <= w_data_i[105];
      \nz.mem_1704_sv2v_reg  <= w_data_i[104];
      \nz.mem_1703_sv2v_reg  <= w_data_i[103];
      \nz.mem_1702_sv2v_reg  <= w_data_i[102];
      \nz.mem_1701_sv2v_reg  <= w_data_i[101];
      \nz.mem_1700_sv2v_reg  <= w_data_i[100];
      \nz.mem_1699_sv2v_reg  <= w_data_i[99];
      \nz.mem_1698_sv2v_reg  <= w_data_i[98];
      \nz.mem_1697_sv2v_reg  <= w_data_i[97];
      \nz.mem_1696_sv2v_reg  <= w_data_i[96];
      \nz.mem_1695_sv2v_reg  <= w_data_i[95];
      \nz.mem_1694_sv2v_reg  <= w_data_i[94];
      \nz.mem_1693_sv2v_reg  <= w_data_i[93];
      \nz.mem_1692_sv2v_reg  <= w_data_i[92];
      \nz.mem_1691_sv2v_reg  <= w_data_i[91];
      \nz.mem_1690_sv2v_reg  <= w_data_i[90];
      \nz.mem_1689_sv2v_reg  <= w_data_i[89];
      \nz.mem_1688_sv2v_reg  <= w_data_i[88];
      \nz.mem_1687_sv2v_reg  <= w_data_i[87];
      \nz.mem_1686_sv2v_reg  <= w_data_i[86];
      \nz.mem_1685_sv2v_reg  <= w_data_i[85];
      \nz.mem_1684_sv2v_reg  <= w_data_i[84];
      \nz.mem_1683_sv2v_reg  <= w_data_i[83];
      \nz.mem_1682_sv2v_reg  <= w_data_i[82];
      \nz.mem_1681_sv2v_reg  <= w_data_i[81];
      \nz.mem_1680_sv2v_reg  <= w_data_i[80];
      \nz.mem_1679_sv2v_reg  <= w_data_i[79];
      \nz.mem_1678_sv2v_reg  <= w_data_i[78];
      \nz.mem_1677_sv2v_reg  <= w_data_i[77];
      \nz.mem_1676_sv2v_reg  <= w_data_i[76];
      \nz.mem_1675_sv2v_reg  <= w_data_i[75];
      \nz.mem_1674_sv2v_reg  <= w_data_i[74];
      \nz.mem_1673_sv2v_reg  <= w_data_i[73];
      \nz.mem_1672_sv2v_reg  <= w_data_i[72];
      \nz.mem_1671_sv2v_reg  <= w_data_i[71];
      \nz.mem_1670_sv2v_reg  <= w_data_i[70];
      \nz.mem_1669_sv2v_reg  <= w_data_i[69];
      \nz.mem_1668_sv2v_reg  <= w_data_i[68];
      \nz.mem_1667_sv2v_reg  <= w_data_i[67];
      \nz.mem_1666_sv2v_reg  <= w_data_i[66];
      \nz.mem_1665_sv2v_reg  <= w_data_i[65];
      \nz.mem_1664_sv2v_reg  <= w_data_i[64];
      \nz.mem_1663_sv2v_reg  <= w_data_i[63];
      \nz.mem_1662_sv2v_reg  <= w_data_i[62];
      \nz.mem_1661_sv2v_reg  <= w_data_i[61];
      \nz.mem_1660_sv2v_reg  <= w_data_i[60];
      \nz.mem_1659_sv2v_reg  <= w_data_i[59];
      \nz.mem_1658_sv2v_reg  <= w_data_i[58];
      \nz.mem_1657_sv2v_reg  <= w_data_i[57];
      \nz.mem_1656_sv2v_reg  <= w_data_i[56];
      \nz.mem_1655_sv2v_reg  <= w_data_i[55];
      \nz.mem_1654_sv2v_reg  <= w_data_i[54];
      \nz.mem_1653_sv2v_reg  <= w_data_i[53];
      \nz.mem_1652_sv2v_reg  <= w_data_i[52];
      \nz.mem_1651_sv2v_reg  <= w_data_i[51];
      \nz.mem_1650_sv2v_reg  <= w_data_i[50];
      \nz.mem_1649_sv2v_reg  <= w_data_i[49];
      \nz.mem_1648_sv2v_reg  <= w_data_i[48];
      \nz.mem_1647_sv2v_reg  <= w_data_i[47];
      \nz.mem_1646_sv2v_reg  <= w_data_i[46];
      \nz.mem_1645_sv2v_reg  <= w_data_i[45];
      \nz.mem_1644_sv2v_reg  <= w_data_i[44];
      \nz.mem_1643_sv2v_reg  <= w_data_i[43];
      \nz.mem_1642_sv2v_reg  <= w_data_i[42];
      \nz.mem_1641_sv2v_reg  <= w_data_i[41];
      \nz.mem_1640_sv2v_reg  <= w_data_i[40];
      \nz.mem_1639_sv2v_reg  <= w_data_i[39];
      \nz.mem_1638_sv2v_reg  <= w_data_i[38];
      \nz.mem_1637_sv2v_reg  <= w_data_i[37];
      \nz.mem_1636_sv2v_reg  <= w_data_i[36];
      \nz.mem_1635_sv2v_reg  <= w_data_i[35];
      \nz.mem_1634_sv2v_reg  <= w_data_i[34];
      \nz.mem_1633_sv2v_reg  <= w_data_i[33];
      \nz.mem_1632_sv2v_reg  <= w_data_i[32];
      \nz.mem_1631_sv2v_reg  <= w_data_i[31];
      \nz.mem_1630_sv2v_reg  <= w_data_i[30];
      \nz.mem_1629_sv2v_reg  <= w_data_i[29];
      \nz.mem_1628_sv2v_reg  <= w_data_i[28];
      \nz.mem_1627_sv2v_reg  <= w_data_i[27];
      \nz.mem_1626_sv2v_reg  <= w_data_i[26];
      \nz.mem_1625_sv2v_reg  <= w_data_i[25];
      \nz.mem_1624_sv2v_reg  <= w_data_i[24];
      \nz.mem_1623_sv2v_reg  <= w_data_i[23];
      \nz.mem_1622_sv2v_reg  <= w_data_i[22];
      \nz.mem_1621_sv2v_reg  <= w_data_i[21];
      \nz.mem_1620_sv2v_reg  <= w_data_i[20];
      \nz.mem_1619_sv2v_reg  <= w_data_i[19];
      \nz.mem_1618_sv2v_reg  <= w_data_i[18];
      \nz.mem_1617_sv2v_reg  <= w_data_i[17];
      \nz.mem_1616_sv2v_reg  <= w_data_i[16];
      \nz.mem_1615_sv2v_reg  <= w_data_i[15];
    end 
    if(N7) begin
      \nz.mem_1599_sv2v_reg  <= w_data_i[1599];
      \nz.mem_1598_sv2v_reg  <= w_data_i[1598];
      \nz.mem_1597_sv2v_reg  <= w_data_i[1597];
      \nz.mem_1596_sv2v_reg  <= w_data_i[1596];
      \nz.mem_1595_sv2v_reg  <= w_data_i[1595];
      \nz.mem_1594_sv2v_reg  <= w_data_i[1594];
      \nz.mem_1593_sv2v_reg  <= w_data_i[1593];
      \nz.mem_1592_sv2v_reg  <= w_data_i[1592];
      \nz.mem_1591_sv2v_reg  <= w_data_i[1591];
      \nz.mem_1590_sv2v_reg  <= w_data_i[1590];
      \nz.mem_1589_sv2v_reg  <= w_data_i[1589];
      \nz.mem_1588_sv2v_reg  <= w_data_i[1588];
      \nz.mem_1587_sv2v_reg  <= w_data_i[1587];
      \nz.mem_1586_sv2v_reg  <= w_data_i[1586];
      \nz.mem_1585_sv2v_reg  <= w_data_i[1585];
      \nz.mem_1584_sv2v_reg  <= w_data_i[1584];
      \nz.mem_1583_sv2v_reg  <= w_data_i[1583];
      \nz.mem_1582_sv2v_reg  <= w_data_i[1582];
      \nz.mem_1581_sv2v_reg  <= w_data_i[1581];
      \nz.mem_1580_sv2v_reg  <= w_data_i[1580];
      \nz.mem_1579_sv2v_reg  <= w_data_i[1579];
      \nz.mem_1578_sv2v_reg  <= w_data_i[1578];
      \nz.mem_1577_sv2v_reg  <= w_data_i[1577];
      \nz.mem_1576_sv2v_reg  <= w_data_i[1576];
      \nz.mem_1575_sv2v_reg  <= w_data_i[1575];
      \nz.mem_1574_sv2v_reg  <= w_data_i[1574];
      \nz.mem_1573_sv2v_reg  <= w_data_i[1573];
      \nz.mem_1572_sv2v_reg  <= w_data_i[1572];
      \nz.mem_1571_sv2v_reg  <= w_data_i[1571];
      \nz.mem_1570_sv2v_reg  <= w_data_i[1570];
      \nz.mem_1569_sv2v_reg  <= w_data_i[1569];
      \nz.mem_1568_sv2v_reg  <= w_data_i[1568];
      \nz.mem_1567_sv2v_reg  <= w_data_i[1567];
      \nz.mem_1566_sv2v_reg  <= w_data_i[1566];
      \nz.mem_1565_sv2v_reg  <= w_data_i[1565];
      \nz.mem_1564_sv2v_reg  <= w_data_i[1564];
      \nz.mem_1563_sv2v_reg  <= w_data_i[1563];
      \nz.mem_1562_sv2v_reg  <= w_data_i[1562];
      \nz.mem_1561_sv2v_reg  <= w_data_i[1561];
      \nz.mem_1560_sv2v_reg  <= w_data_i[1560];
      \nz.mem_1559_sv2v_reg  <= w_data_i[1559];
      \nz.mem_1558_sv2v_reg  <= w_data_i[1558];
      \nz.mem_1557_sv2v_reg  <= w_data_i[1557];
      \nz.mem_1556_sv2v_reg  <= w_data_i[1556];
      \nz.mem_1555_sv2v_reg  <= w_data_i[1555];
      \nz.mem_1554_sv2v_reg  <= w_data_i[1554];
      \nz.mem_1553_sv2v_reg  <= w_data_i[1553];
      \nz.mem_1552_sv2v_reg  <= w_data_i[1552];
      \nz.mem_1551_sv2v_reg  <= w_data_i[1551];
      \nz.mem_1550_sv2v_reg  <= w_data_i[1550];
      \nz.mem_1549_sv2v_reg  <= w_data_i[1549];
      \nz.mem_1548_sv2v_reg  <= w_data_i[1548];
      \nz.mem_1547_sv2v_reg  <= w_data_i[1547];
      \nz.mem_1546_sv2v_reg  <= w_data_i[1546];
      \nz.mem_1545_sv2v_reg  <= w_data_i[1545];
      \nz.mem_1544_sv2v_reg  <= w_data_i[1544];
      \nz.mem_1543_sv2v_reg  <= w_data_i[1543];
      \nz.mem_1542_sv2v_reg  <= w_data_i[1542];
      \nz.mem_1541_sv2v_reg  <= w_data_i[1541];
      \nz.mem_1540_sv2v_reg  <= w_data_i[1540];
      \nz.mem_1539_sv2v_reg  <= w_data_i[1539];
      \nz.mem_1538_sv2v_reg  <= w_data_i[1538];
      \nz.mem_1537_sv2v_reg  <= w_data_i[1537];
      \nz.mem_1536_sv2v_reg  <= w_data_i[1536];
      \nz.mem_1535_sv2v_reg  <= w_data_i[1535];
      \nz.mem_1534_sv2v_reg  <= w_data_i[1534];
      \nz.mem_1533_sv2v_reg  <= w_data_i[1533];
      \nz.mem_1532_sv2v_reg  <= w_data_i[1532];
      \nz.mem_1531_sv2v_reg  <= w_data_i[1531];
      \nz.mem_1530_sv2v_reg  <= w_data_i[1530];
      \nz.mem_1529_sv2v_reg  <= w_data_i[1529];
      \nz.mem_1528_sv2v_reg  <= w_data_i[1528];
      \nz.mem_1527_sv2v_reg  <= w_data_i[1527];
      \nz.mem_1526_sv2v_reg  <= w_data_i[1526];
      \nz.mem_1525_sv2v_reg  <= w_data_i[1525];
      \nz.mem_1524_sv2v_reg  <= w_data_i[1524];
      \nz.mem_1523_sv2v_reg  <= w_data_i[1523];
      \nz.mem_1522_sv2v_reg  <= w_data_i[1522];
      \nz.mem_1521_sv2v_reg  <= w_data_i[1521];
      \nz.mem_1520_sv2v_reg  <= w_data_i[1520];
      \nz.mem_1519_sv2v_reg  <= w_data_i[1519];
      \nz.mem_1518_sv2v_reg  <= w_data_i[1518];
      \nz.mem_1517_sv2v_reg  <= w_data_i[1517];
      \nz.mem_1516_sv2v_reg  <= w_data_i[1516];
      \nz.mem_1515_sv2v_reg  <= w_data_i[1515];
      \nz.mem_1514_sv2v_reg  <= w_data_i[1514];
      \nz.mem_1513_sv2v_reg  <= w_data_i[1513];
      \nz.mem_1512_sv2v_reg  <= w_data_i[1512];
      \nz.mem_1511_sv2v_reg  <= w_data_i[1511];
      \nz.mem_1510_sv2v_reg  <= w_data_i[1510];
      \nz.mem_1509_sv2v_reg  <= w_data_i[1509];
      \nz.mem_1508_sv2v_reg  <= w_data_i[1508];
      \nz.mem_1507_sv2v_reg  <= w_data_i[1507];
      \nz.mem_1506_sv2v_reg  <= w_data_i[1506];
      \nz.mem_1505_sv2v_reg  <= w_data_i[1505];
      \nz.mem_1504_sv2v_reg  <= w_data_i[1504];
      \nz.mem_1503_sv2v_reg  <= w_data_i[1503];
      \nz.mem_1502_sv2v_reg  <= w_data_i[1502];
      \nz.mem_1501_sv2v_reg  <= w_data_i[1501];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
    if(N8) begin
      \nz.mem_1500_sv2v_reg  <= w_data_i[1500];
      \nz.mem_1499_sv2v_reg  <= w_data_i[1499];
      \nz.mem_1498_sv2v_reg  <= w_data_i[1498];
      \nz.mem_1497_sv2v_reg  <= w_data_i[1497];
      \nz.mem_1496_sv2v_reg  <= w_data_i[1496];
      \nz.mem_1495_sv2v_reg  <= w_data_i[1495];
      \nz.mem_1494_sv2v_reg  <= w_data_i[1494];
      \nz.mem_1493_sv2v_reg  <= w_data_i[1493];
      \nz.mem_1492_sv2v_reg  <= w_data_i[1492];
      \nz.mem_1491_sv2v_reg  <= w_data_i[1491];
      \nz.mem_1490_sv2v_reg  <= w_data_i[1490];
      \nz.mem_1489_sv2v_reg  <= w_data_i[1489];
      \nz.mem_1488_sv2v_reg  <= w_data_i[1488];
      \nz.mem_1487_sv2v_reg  <= w_data_i[1487];
      \nz.mem_1486_sv2v_reg  <= w_data_i[1486];
      \nz.mem_1485_sv2v_reg  <= w_data_i[1485];
      \nz.mem_1484_sv2v_reg  <= w_data_i[1484];
      \nz.mem_1483_sv2v_reg  <= w_data_i[1483];
      \nz.mem_1482_sv2v_reg  <= w_data_i[1482];
      \nz.mem_1481_sv2v_reg  <= w_data_i[1481];
      \nz.mem_1480_sv2v_reg  <= w_data_i[1480];
      \nz.mem_1479_sv2v_reg  <= w_data_i[1479];
      \nz.mem_1478_sv2v_reg  <= w_data_i[1478];
      \nz.mem_1477_sv2v_reg  <= w_data_i[1477];
      \nz.mem_1476_sv2v_reg  <= w_data_i[1476];
      \nz.mem_1475_sv2v_reg  <= w_data_i[1475];
      \nz.mem_1474_sv2v_reg  <= w_data_i[1474];
      \nz.mem_1473_sv2v_reg  <= w_data_i[1473];
      \nz.mem_1472_sv2v_reg  <= w_data_i[1472];
      \nz.mem_1471_sv2v_reg  <= w_data_i[1471];
      \nz.mem_1470_sv2v_reg  <= w_data_i[1470];
      \nz.mem_1469_sv2v_reg  <= w_data_i[1469];
      \nz.mem_1468_sv2v_reg  <= w_data_i[1468];
      \nz.mem_1467_sv2v_reg  <= w_data_i[1467];
      \nz.mem_1466_sv2v_reg  <= w_data_i[1466];
      \nz.mem_1465_sv2v_reg  <= w_data_i[1465];
      \nz.mem_1464_sv2v_reg  <= w_data_i[1464];
      \nz.mem_1463_sv2v_reg  <= w_data_i[1463];
      \nz.mem_1462_sv2v_reg  <= w_data_i[1462];
      \nz.mem_1461_sv2v_reg  <= w_data_i[1461];
      \nz.mem_1460_sv2v_reg  <= w_data_i[1460];
      \nz.mem_1459_sv2v_reg  <= w_data_i[1459];
      \nz.mem_1458_sv2v_reg  <= w_data_i[1458];
      \nz.mem_1457_sv2v_reg  <= w_data_i[1457];
      \nz.mem_1456_sv2v_reg  <= w_data_i[1456];
      \nz.mem_1455_sv2v_reg  <= w_data_i[1455];
      \nz.mem_1454_sv2v_reg  <= w_data_i[1454];
      \nz.mem_1453_sv2v_reg  <= w_data_i[1453];
      \nz.mem_1452_sv2v_reg  <= w_data_i[1452];
      \nz.mem_1451_sv2v_reg  <= w_data_i[1451];
      \nz.mem_1450_sv2v_reg  <= w_data_i[1450];
      \nz.mem_1449_sv2v_reg  <= w_data_i[1449];
      \nz.mem_1448_sv2v_reg  <= w_data_i[1448];
      \nz.mem_1447_sv2v_reg  <= w_data_i[1447];
      \nz.mem_1446_sv2v_reg  <= w_data_i[1446];
      \nz.mem_1445_sv2v_reg  <= w_data_i[1445];
      \nz.mem_1444_sv2v_reg  <= w_data_i[1444];
      \nz.mem_1443_sv2v_reg  <= w_data_i[1443];
      \nz.mem_1442_sv2v_reg  <= w_data_i[1442];
      \nz.mem_1441_sv2v_reg  <= w_data_i[1441];
      \nz.mem_1440_sv2v_reg  <= w_data_i[1440];
      \nz.mem_1439_sv2v_reg  <= w_data_i[1439];
      \nz.mem_1438_sv2v_reg  <= w_data_i[1438];
      \nz.mem_1437_sv2v_reg  <= w_data_i[1437];
      \nz.mem_1436_sv2v_reg  <= w_data_i[1436];
      \nz.mem_1435_sv2v_reg  <= w_data_i[1435];
      \nz.mem_1434_sv2v_reg  <= w_data_i[1434];
      \nz.mem_1433_sv2v_reg  <= w_data_i[1433];
      \nz.mem_1432_sv2v_reg  <= w_data_i[1432];
      \nz.mem_1431_sv2v_reg  <= w_data_i[1431];
      \nz.mem_1430_sv2v_reg  <= w_data_i[1430];
      \nz.mem_1429_sv2v_reg  <= w_data_i[1429];
      \nz.mem_1428_sv2v_reg  <= w_data_i[1428];
      \nz.mem_1427_sv2v_reg  <= w_data_i[1427];
      \nz.mem_1426_sv2v_reg  <= w_data_i[1426];
      \nz.mem_1425_sv2v_reg  <= w_data_i[1425];
      \nz.mem_1424_sv2v_reg  <= w_data_i[1424];
      \nz.mem_1423_sv2v_reg  <= w_data_i[1423];
      \nz.mem_1422_sv2v_reg  <= w_data_i[1422];
      \nz.mem_1421_sv2v_reg  <= w_data_i[1421];
      \nz.mem_1420_sv2v_reg  <= w_data_i[1420];
      \nz.mem_1419_sv2v_reg  <= w_data_i[1419];
      \nz.mem_1418_sv2v_reg  <= w_data_i[1418];
      \nz.mem_1417_sv2v_reg  <= w_data_i[1417];
      \nz.mem_1416_sv2v_reg  <= w_data_i[1416];
      \nz.mem_1415_sv2v_reg  <= w_data_i[1415];
      \nz.mem_1414_sv2v_reg  <= w_data_i[1414];
      \nz.mem_1413_sv2v_reg  <= w_data_i[1413];
      \nz.mem_1412_sv2v_reg  <= w_data_i[1412];
      \nz.mem_1411_sv2v_reg  <= w_data_i[1411];
      \nz.mem_1410_sv2v_reg  <= w_data_i[1410];
      \nz.mem_1409_sv2v_reg  <= w_data_i[1409];
      \nz.mem_1408_sv2v_reg  <= w_data_i[1408];
      \nz.mem_1407_sv2v_reg  <= w_data_i[1407];
      \nz.mem_1406_sv2v_reg  <= w_data_i[1406];
      \nz.mem_1405_sv2v_reg  <= w_data_i[1405];
      \nz.mem_1404_sv2v_reg  <= w_data_i[1404];
      \nz.mem_1403_sv2v_reg  <= w_data_i[1403];
      \nz.mem_1402_sv2v_reg  <= w_data_i[1402];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
    end 
    if(N9) begin
      \nz.mem_1401_sv2v_reg  <= w_data_i[1401];
      \nz.mem_1400_sv2v_reg  <= w_data_i[1400];
      \nz.mem_1399_sv2v_reg  <= w_data_i[1399];
      \nz.mem_1398_sv2v_reg  <= w_data_i[1398];
      \nz.mem_1397_sv2v_reg  <= w_data_i[1397];
      \nz.mem_1396_sv2v_reg  <= w_data_i[1396];
      \nz.mem_1395_sv2v_reg  <= w_data_i[1395];
      \nz.mem_1394_sv2v_reg  <= w_data_i[1394];
      \nz.mem_1393_sv2v_reg  <= w_data_i[1393];
      \nz.mem_1392_sv2v_reg  <= w_data_i[1392];
      \nz.mem_1391_sv2v_reg  <= w_data_i[1391];
      \nz.mem_1390_sv2v_reg  <= w_data_i[1390];
      \nz.mem_1389_sv2v_reg  <= w_data_i[1389];
      \nz.mem_1388_sv2v_reg  <= w_data_i[1388];
      \nz.mem_1387_sv2v_reg  <= w_data_i[1387];
      \nz.mem_1386_sv2v_reg  <= w_data_i[1386];
      \nz.mem_1385_sv2v_reg  <= w_data_i[1385];
      \nz.mem_1384_sv2v_reg  <= w_data_i[1384];
      \nz.mem_1383_sv2v_reg  <= w_data_i[1383];
      \nz.mem_1382_sv2v_reg  <= w_data_i[1382];
      \nz.mem_1381_sv2v_reg  <= w_data_i[1381];
      \nz.mem_1380_sv2v_reg  <= w_data_i[1380];
      \nz.mem_1379_sv2v_reg  <= w_data_i[1379];
      \nz.mem_1378_sv2v_reg  <= w_data_i[1378];
      \nz.mem_1377_sv2v_reg  <= w_data_i[1377];
      \nz.mem_1376_sv2v_reg  <= w_data_i[1376];
      \nz.mem_1375_sv2v_reg  <= w_data_i[1375];
      \nz.mem_1374_sv2v_reg  <= w_data_i[1374];
      \nz.mem_1373_sv2v_reg  <= w_data_i[1373];
      \nz.mem_1372_sv2v_reg  <= w_data_i[1372];
      \nz.mem_1371_sv2v_reg  <= w_data_i[1371];
      \nz.mem_1370_sv2v_reg  <= w_data_i[1370];
      \nz.mem_1369_sv2v_reg  <= w_data_i[1369];
      \nz.mem_1368_sv2v_reg  <= w_data_i[1368];
      \nz.mem_1367_sv2v_reg  <= w_data_i[1367];
      \nz.mem_1366_sv2v_reg  <= w_data_i[1366];
      \nz.mem_1365_sv2v_reg  <= w_data_i[1365];
      \nz.mem_1364_sv2v_reg  <= w_data_i[1364];
      \nz.mem_1363_sv2v_reg  <= w_data_i[1363];
      \nz.mem_1362_sv2v_reg  <= w_data_i[1362];
      \nz.mem_1361_sv2v_reg  <= w_data_i[1361];
      \nz.mem_1360_sv2v_reg  <= w_data_i[1360];
      \nz.mem_1359_sv2v_reg  <= w_data_i[1359];
      \nz.mem_1358_sv2v_reg  <= w_data_i[1358];
      \nz.mem_1357_sv2v_reg  <= w_data_i[1357];
      \nz.mem_1356_sv2v_reg  <= w_data_i[1356];
      \nz.mem_1355_sv2v_reg  <= w_data_i[1355];
      \nz.mem_1354_sv2v_reg  <= w_data_i[1354];
      \nz.mem_1353_sv2v_reg  <= w_data_i[1353];
      \nz.mem_1352_sv2v_reg  <= w_data_i[1352];
      \nz.mem_1351_sv2v_reg  <= w_data_i[1351];
      \nz.mem_1350_sv2v_reg  <= w_data_i[1350];
      \nz.mem_1349_sv2v_reg  <= w_data_i[1349];
      \nz.mem_1348_sv2v_reg  <= w_data_i[1348];
      \nz.mem_1347_sv2v_reg  <= w_data_i[1347];
      \nz.mem_1346_sv2v_reg  <= w_data_i[1346];
      \nz.mem_1345_sv2v_reg  <= w_data_i[1345];
      \nz.mem_1344_sv2v_reg  <= w_data_i[1344];
      \nz.mem_1343_sv2v_reg  <= w_data_i[1343];
      \nz.mem_1342_sv2v_reg  <= w_data_i[1342];
      \nz.mem_1341_sv2v_reg  <= w_data_i[1341];
      \nz.mem_1340_sv2v_reg  <= w_data_i[1340];
      \nz.mem_1339_sv2v_reg  <= w_data_i[1339];
      \nz.mem_1338_sv2v_reg  <= w_data_i[1338];
      \nz.mem_1337_sv2v_reg  <= w_data_i[1337];
      \nz.mem_1336_sv2v_reg  <= w_data_i[1336];
      \nz.mem_1335_sv2v_reg  <= w_data_i[1335];
      \nz.mem_1334_sv2v_reg  <= w_data_i[1334];
      \nz.mem_1333_sv2v_reg  <= w_data_i[1333];
      \nz.mem_1332_sv2v_reg  <= w_data_i[1332];
      \nz.mem_1331_sv2v_reg  <= w_data_i[1331];
      \nz.mem_1330_sv2v_reg  <= w_data_i[1330];
      \nz.mem_1329_sv2v_reg  <= w_data_i[1329];
      \nz.mem_1328_sv2v_reg  <= w_data_i[1328];
      \nz.mem_1327_sv2v_reg  <= w_data_i[1327];
      \nz.mem_1326_sv2v_reg  <= w_data_i[1326];
      \nz.mem_1325_sv2v_reg  <= w_data_i[1325];
      \nz.mem_1324_sv2v_reg  <= w_data_i[1324];
      \nz.mem_1323_sv2v_reg  <= w_data_i[1323];
      \nz.mem_1322_sv2v_reg  <= w_data_i[1322];
      \nz.mem_1321_sv2v_reg  <= w_data_i[1321];
      \nz.mem_1320_sv2v_reg  <= w_data_i[1320];
      \nz.mem_1319_sv2v_reg  <= w_data_i[1319];
      \nz.mem_1318_sv2v_reg  <= w_data_i[1318];
      \nz.mem_1317_sv2v_reg  <= w_data_i[1317];
      \nz.mem_1316_sv2v_reg  <= w_data_i[1316];
      \nz.mem_1315_sv2v_reg  <= w_data_i[1315];
      \nz.mem_1314_sv2v_reg  <= w_data_i[1314];
      \nz.mem_1313_sv2v_reg  <= w_data_i[1313];
      \nz.mem_1312_sv2v_reg  <= w_data_i[1312];
      \nz.mem_1311_sv2v_reg  <= w_data_i[1311];
      \nz.mem_1310_sv2v_reg  <= w_data_i[1310];
      \nz.mem_1309_sv2v_reg  <= w_data_i[1309];
      \nz.mem_1308_sv2v_reg  <= w_data_i[1308];
      \nz.mem_1307_sv2v_reg  <= w_data_i[1307];
      \nz.mem_1306_sv2v_reg  <= w_data_i[1306];
      \nz.mem_1305_sv2v_reg  <= w_data_i[1305];
      \nz.mem_1304_sv2v_reg  <= w_data_i[1304];
      \nz.mem_1303_sv2v_reg  <= w_data_i[1303];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
    end 
    if(N10) begin
      \nz.mem_1302_sv2v_reg  <= w_data_i[1302];
      \nz.mem_1301_sv2v_reg  <= w_data_i[1301];
      \nz.mem_1300_sv2v_reg  <= w_data_i[1300];
      \nz.mem_1299_sv2v_reg  <= w_data_i[1299];
      \nz.mem_1298_sv2v_reg  <= w_data_i[1298];
      \nz.mem_1297_sv2v_reg  <= w_data_i[1297];
      \nz.mem_1296_sv2v_reg  <= w_data_i[1296];
      \nz.mem_1295_sv2v_reg  <= w_data_i[1295];
      \nz.mem_1294_sv2v_reg  <= w_data_i[1294];
      \nz.mem_1293_sv2v_reg  <= w_data_i[1293];
      \nz.mem_1292_sv2v_reg  <= w_data_i[1292];
      \nz.mem_1291_sv2v_reg  <= w_data_i[1291];
      \nz.mem_1290_sv2v_reg  <= w_data_i[1290];
      \nz.mem_1289_sv2v_reg  <= w_data_i[1289];
      \nz.mem_1288_sv2v_reg  <= w_data_i[1288];
      \nz.mem_1287_sv2v_reg  <= w_data_i[1287];
      \nz.mem_1286_sv2v_reg  <= w_data_i[1286];
      \nz.mem_1285_sv2v_reg  <= w_data_i[1285];
      \nz.mem_1284_sv2v_reg  <= w_data_i[1284];
      \nz.mem_1283_sv2v_reg  <= w_data_i[1283];
      \nz.mem_1282_sv2v_reg  <= w_data_i[1282];
      \nz.mem_1281_sv2v_reg  <= w_data_i[1281];
      \nz.mem_1280_sv2v_reg  <= w_data_i[1280];
      \nz.mem_1279_sv2v_reg  <= w_data_i[1279];
      \nz.mem_1278_sv2v_reg  <= w_data_i[1278];
      \nz.mem_1277_sv2v_reg  <= w_data_i[1277];
      \nz.mem_1276_sv2v_reg  <= w_data_i[1276];
      \nz.mem_1275_sv2v_reg  <= w_data_i[1275];
      \nz.mem_1274_sv2v_reg  <= w_data_i[1274];
      \nz.mem_1273_sv2v_reg  <= w_data_i[1273];
      \nz.mem_1272_sv2v_reg  <= w_data_i[1272];
      \nz.mem_1271_sv2v_reg  <= w_data_i[1271];
      \nz.mem_1270_sv2v_reg  <= w_data_i[1270];
      \nz.mem_1269_sv2v_reg  <= w_data_i[1269];
      \nz.mem_1268_sv2v_reg  <= w_data_i[1268];
      \nz.mem_1267_sv2v_reg  <= w_data_i[1267];
      \nz.mem_1266_sv2v_reg  <= w_data_i[1266];
      \nz.mem_1265_sv2v_reg  <= w_data_i[1265];
      \nz.mem_1264_sv2v_reg  <= w_data_i[1264];
      \nz.mem_1263_sv2v_reg  <= w_data_i[1263];
      \nz.mem_1262_sv2v_reg  <= w_data_i[1262];
      \nz.mem_1261_sv2v_reg  <= w_data_i[1261];
      \nz.mem_1260_sv2v_reg  <= w_data_i[1260];
      \nz.mem_1259_sv2v_reg  <= w_data_i[1259];
      \nz.mem_1258_sv2v_reg  <= w_data_i[1258];
      \nz.mem_1257_sv2v_reg  <= w_data_i[1257];
      \nz.mem_1256_sv2v_reg  <= w_data_i[1256];
      \nz.mem_1255_sv2v_reg  <= w_data_i[1255];
      \nz.mem_1254_sv2v_reg  <= w_data_i[1254];
      \nz.mem_1253_sv2v_reg  <= w_data_i[1253];
      \nz.mem_1252_sv2v_reg  <= w_data_i[1252];
      \nz.mem_1251_sv2v_reg  <= w_data_i[1251];
      \nz.mem_1250_sv2v_reg  <= w_data_i[1250];
      \nz.mem_1249_sv2v_reg  <= w_data_i[1249];
      \nz.mem_1248_sv2v_reg  <= w_data_i[1248];
      \nz.mem_1247_sv2v_reg  <= w_data_i[1247];
      \nz.mem_1246_sv2v_reg  <= w_data_i[1246];
      \nz.mem_1245_sv2v_reg  <= w_data_i[1245];
      \nz.mem_1244_sv2v_reg  <= w_data_i[1244];
      \nz.mem_1243_sv2v_reg  <= w_data_i[1243];
      \nz.mem_1242_sv2v_reg  <= w_data_i[1242];
      \nz.mem_1241_sv2v_reg  <= w_data_i[1241];
      \nz.mem_1240_sv2v_reg  <= w_data_i[1240];
      \nz.mem_1239_sv2v_reg  <= w_data_i[1239];
      \nz.mem_1238_sv2v_reg  <= w_data_i[1238];
      \nz.mem_1237_sv2v_reg  <= w_data_i[1237];
      \nz.mem_1236_sv2v_reg  <= w_data_i[1236];
      \nz.mem_1235_sv2v_reg  <= w_data_i[1235];
      \nz.mem_1234_sv2v_reg  <= w_data_i[1234];
      \nz.mem_1233_sv2v_reg  <= w_data_i[1233];
      \nz.mem_1232_sv2v_reg  <= w_data_i[1232];
      \nz.mem_1231_sv2v_reg  <= w_data_i[1231];
      \nz.mem_1230_sv2v_reg  <= w_data_i[1230];
      \nz.mem_1229_sv2v_reg  <= w_data_i[1229];
      \nz.mem_1228_sv2v_reg  <= w_data_i[1228];
      \nz.mem_1227_sv2v_reg  <= w_data_i[1227];
      \nz.mem_1226_sv2v_reg  <= w_data_i[1226];
      \nz.mem_1225_sv2v_reg  <= w_data_i[1225];
      \nz.mem_1224_sv2v_reg  <= w_data_i[1224];
      \nz.mem_1223_sv2v_reg  <= w_data_i[1223];
      \nz.mem_1222_sv2v_reg  <= w_data_i[1222];
      \nz.mem_1221_sv2v_reg  <= w_data_i[1221];
      \nz.mem_1220_sv2v_reg  <= w_data_i[1220];
      \nz.mem_1219_sv2v_reg  <= w_data_i[1219];
      \nz.mem_1218_sv2v_reg  <= w_data_i[1218];
      \nz.mem_1217_sv2v_reg  <= w_data_i[1217];
      \nz.mem_1216_sv2v_reg  <= w_data_i[1216];
      \nz.mem_1215_sv2v_reg  <= w_data_i[1215];
      \nz.mem_1214_sv2v_reg  <= w_data_i[1214];
      \nz.mem_1213_sv2v_reg  <= w_data_i[1213];
      \nz.mem_1212_sv2v_reg  <= w_data_i[1212];
      \nz.mem_1211_sv2v_reg  <= w_data_i[1211];
      \nz.mem_1210_sv2v_reg  <= w_data_i[1210];
      \nz.mem_1209_sv2v_reg  <= w_data_i[1209];
      \nz.mem_1208_sv2v_reg  <= w_data_i[1208];
      \nz.mem_1207_sv2v_reg  <= w_data_i[1207];
      \nz.mem_1206_sv2v_reg  <= w_data_i[1206];
      \nz.mem_1205_sv2v_reg  <= w_data_i[1205];
      \nz.mem_1204_sv2v_reg  <= w_data_i[1204];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
    end 
    if(N11) begin
      \nz.mem_1203_sv2v_reg  <= w_data_i[1203];
      \nz.mem_1202_sv2v_reg  <= w_data_i[1202];
      \nz.mem_1201_sv2v_reg  <= w_data_i[1201];
      \nz.mem_1200_sv2v_reg  <= w_data_i[1200];
      \nz.mem_1199_sv2v_reg  <= w_data_i[1199];
      \nz.mem_1198_sv2v_reg  <= w_data_i[1198];
      \nz.mem_1197_sv2v_reg  <= w_data_i[1197];
      \nz.mem_1196_sv2v_reg  <= w_data_i[1196];
      \nz.mem_1195_sv2v_reg  <= w_data_i[1195];
      \nz.mem_1194_sv2v_reg  <= w_data_i[1194];
      \nz.mem_1193_sv2v_reg  <= w_data_i[1193];
      \nz.mem_1192_sv2v_reg  <= w_data_i[1192];
      \nz.mem_1191_sv2v_reg  <= w_data_i[1191];
      \nz.mem_1190_sv2v_reg  <= w_data_i[1190];
      \nz.mem_1189_sv2v_reg  <= w_data_i[1189];
      \nz.mem_1188_sv2v_reg  <= w_data_i[1188];
      \nz.mem_1187_sv2v_reg  <= w_data_i[1187];
      \nz.mem_1186_sv2v_reg  <= w_data_i[1186];
      \nz.mem_1185_sv2v_reg  <= w_data_i[1185];
      \nz.mem_1184_sv2v_reg  <= w_data_i[1184];
      \nz.mem_1183_sv2v_reg  <= w_data_i[1183];
      \nz.mem_1182_sv2v_reg  <= w_data_i[1182];
      \nz.mem_1181_sv2v_reg  <= w_data_i[1181];
      \nz.mem_1180_sv2v_reg  <= w_data_i[1180];
      \nz.mem_1179_sv2v_reg  <= w_data_i[1179];
      \nz.mem_1178_sv2v_reg  <= w_data_i[1178];
      \nz.mem_1177_sv2v_reg  <= w_data_i[1177];
      \nz.mem_1176_sv2v_reg  <= w_data_i[1176];
      \nz.mem_1175_sv2v_reg  <= w_data_i[1175];
      \nz.mem_1174_sv2v_reg  <= w_data_i[1174];
      \nz.mem_1173_sv2v_reg  <= w_data_i[1173];
      \nz.mem_1172_sv2v_reg  <= w_data_i[1172];
      \nz.mem_1171_sv2v_reg  <= w_data_i[1171];
      \nz.mem_1170_sv2v_reg  <= w_data_i[1170];
      \nz.mem_1169_sv2v_reg  <= w_data_i[1169];
      \nz.mem_1168_sv2v_reg  <= w_data_i[1168];
      \nz.mem_1167_sv2v_reg  <= w_data_i[1167];
      \nz.mem_1166_sv2v_reg  <= w_data_i[1166];
      \nz.mem_1165_sv2v_reg  <= w_data_i[1165];
      \nz.mem_1164_sv2v_reg  <= w_data_i[1164];
      \nz.mem_1163_sv2v_reg  <= w_data_i[1163];
      \nz.mem_1162_sv2v_reg  <= w_data_i[1162];
      \nz.mem_1161_sv2v_reg  <= w_data_i[1161];
      \nz.mem_1160_sv2v_reg  <= w_data_i[1160];
      \nz.mem_1159_sv2v_reg  <= w_data_i[1159];
      \nz.mem_1158_sv2v_reg  <= w_data_i[1158];
      \nz.mem_1157_sv2v_reg  <= w_data_i[1157];
      \nz.mem_1156_sv2v_reg  <= w_data_i[1156];
      \nz.mem_1155_sv2v_reg  <= w_data_i[1155];
      \nz.mem_1154_sv2v_reg  <= w_data_i[1154];
      \nz.mem_1153_sv2v_reg  <= w_data_i[1153];
      \nz.mem_1152_sv2v_reg  <= w_data_i[1152];
      \nz.mem_1151_sv2v_reg  <= w_data_i[1151];
      \nz.mem_1150_sv2v_reg  <= w_data_i[1150];
      \nz.mem_1149_sv2v_reg  <= w_data_i[1149];
      \nz.mem_1148_sv2v_reg  <= w_data_i[1148];
      \nz.mem_1147_sv2v_reg  <= w_data_i[1147];
      \nz.mem_1146_sv2v_reg  <= w_data_i[1146];
      \nz.mem_1145_sv2v_reg  <= w_data_i[1145];
      \nz.mem_1144_sv2v_reg  <= w_data_i[1144];
      \nz.mem_1143_sv2v_reg  <= w_data_i[1143];
      \nz.mem_1142_sv2v_reg  <= w_data_i[1142];
      \nz.mem_1141_sv2v_reg  <= w_data_i[1141];
      \nz.mem_1140_sv2v_reg  <= w_data_i[1140];
      \nz.mem_1139_sv2v_reg  <= w_data_i[1139];
      \nz.mem_1138_sv2v_reg  <= w_data_i[1138];
      \nz.mem_1137_sv2v_reg  <= w_data_i[1137];
      \nz.mem_1136_sv2v_reg  <= w_data_i[1136];
      \nz.mem_1135_sv2v_reg  <= w_data_i[1135];
      \nz.mem_1134_sv2v_reg  <= w_data_i[1134];
      \nz.mem_1133_sv2v_reg  <= w_data_i[1133];
      \nz.mem_1132_sv2v_reg  <= w_data_i[1132];
      \nz.mem_1131_sv2v_reg  <= w_data_i[1131];
      \nz.mem_1130_sv2v_reg  <= w_data_i[1130];
      \nz.mem_1129_sv2v_reg  <= w_data_i[1129];
      \nz.mem_1128_sv2v_reg  <= w_data_i[1128];
      \nz.mem_1127_sv2v_reg  <= w_data_i[1127];
      \nz.mem_1126_sv2v_reg  <= w_data_i[1126];
      \nz.mem_1125_sv2v_reg  <= w_data_i[1125];
      \nz.mem_1124_sv2v_reg  <= w_data_i[1124];
      \nz.mem_1123_sv2v_reg  <= w_data_i[1123];
      \nz.mem_1122_sv2v_reg  <= w_data_i[1122];
      \nz.mem_1121_sv2v_reg  <= w_data_i[1121];
      \nz.mem_1120_sv2v_reg  <= w_data_i[1120];
      \nz.mem_1119_sv2v_reg  <= w_data_i[1119];
      \nz.mem_1118_sv2v_reg  <= w_data_i[1118];
      \nz.mem_1117_sv2v_reg  <= w_data_i[1117];
      \nz.mem_1116_sv2v_reg  <= w_data_i[1116];
      \nz.mem_1115_sv2v_reg  <= w_data_i[1115];
      \nz.mem_1114_sv2v_reg  <= w_data_i[1114];
      \nz.mem_1113_sv2v_reg  <= w_data_i[1113];
      \nz.mem_1112_sv2v_reg  <= w_data_i[1112];
      \nz.mem_1111_sv2v_reg  <= w_data_i[1111];
      \nz.mem_1110_sv2v_reg  <= w_data_i[1110];
      \nz.mem_1109_sv2v_reg  <= w_data_i[1109];
      \nz.mem_1108_sv2v_reg  <= w_data_i[1108];
      \nz.mem_1107_sv2v_reg  <= w_data_i[1107];
      \nz.mem_1106_sv2v_reg  <= w_data_i[1106];
      \nz.mem_1105_sv2v_reg  <= w_data_i[1105];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
    end 
    if(N12) begin
      \nz.mem_1104_sv2v_reg  <= w_data_i[1104];
      \nz.mem_1103_sv2v_reg  <= w_data_i[1103];
      \nz.mem_1102_sv2v_reg  <= w_data_i[1102];
      \nz.mem_1101_sv2v_reg  <= w_data_i[1101];
      \nz.mem_1100_sv2v_reg  <= w_data_i[1100];
      \nz.mem_1099_sv2v_reg  <= w_data_i[1099];
      \nz.mem_1098_sv2v_reg  <= w_data_i[1098];
      \nz.mem_1097_sv2v_reg  <= w_data_i[1097];
      \nz.mem_1096_sv2v_reg  <= w_data_i[1096];
      \nz.mem_1095_sv2v_reg  <= w_data_i[1095];
      \nz.mem_1094_sv2v_reg  <= w_data_i[1094];
      \nz.mem_1093_sv2v_reg  <= w_data_i[1093];
      \nz.mem_1092_sv2v_reg  <= w_data_i[1092];
      \nz.mem_1091_sv2v_reg  <= w_data_i[1091];
      \nz.mem_1090_sv2v_reg  <= w_data_i[1090];
      \nz.mem_1089_sv2v_reg  <= w_data_i[1089];
      \nz.mem_1088_sv2v_reg  <= w_data_i[1088];
      \nz.mem_1087_sv2v_reg  <= w_data_i[1087];
      \nz.mem_1086_sv2v_reg  <= w_data_i[1086];
      \nz.mem_1085_sv2v_reg  <= w_data_i[1085];
      \nz.mem_1084_sv2v_reg  <= w_data_i[1084];
      \nz.mem_1083_sv2v_reg  <= w_data_i[1083];
      \nz.mem_1082_sv2v_reg  <= w_data_i[1082];
      \nz.mem_1081_sv2v_reg  <= w_data_i[1081];
      \nz.mem_1080_sv2v_reg  <= w_data_i[1080];
      \nz.mem_1079_sv2v_reg  <= w_data_i[1079];
      \nz.mem_1078_sv2v_reg  <= w_data_i[1078];
      \nz.mem_1077_sv2v_reg  <= w_data_i[1077];
      \nz.mem_1076_sv2v_reg  <= w_data_i[1076];
      \nz.mem_1075_sv2v_reg  <= w_data_i[1075];
      \nz.mem_1074_sv2v_reg  <= w_data_i[1074];
      \nz.mem_1073_sv2v_reg  <= w_data_i[1073];
      \nz.mem_1072_sv2v_reg  <= w_data_i[1072];
      \nz.mem_1071_sv2v_reg  <= w_data_i[1071];
      \nz.mem_1070_sv2v_reg  <= w_data_i[1070];
      \nz.mem_1069_sv2v_reg  <= w_data_i[1069];
      \nz.mem_1068_sv2v_reg  <= w_data_i[1068];
      \nz.mem_1067_sv2v_reg  <= w_data_i[1067];
      \nz.mem_1066_sv2v_reg  <= w_data_i[1066];
      \nz.mem_1065_sv2v_reg  <= w_data_i[1065];
      \nz.mem_1064_sv2v_reg  <= w_data_i[1064];
      \nz.mem_1063_sv2v_reg  <= w_data_i[1063];
      \nz.mem_1062_sv2v_reg  <= w_data_i[1062];
      \nz.mem_1061_sv2v_reg  <= w_data_i[1061];
      \nz.mem_1060_sv2v_reg  <= w_data_i[1060];
      \nz.mem_1059_sv2v_reg  <= w_data_i[1059];
      \nz.mem_1058_sv2v_reg  <= w_data_i[1058];
      \nz.mem_1057_sv2v_reg  <= w_data_i[1057];
      \nz.mem_1056_sv2v_reg  <= w_data_i[1056];
      \nz.mem_1055_sv2v_reg  <= w_data_i[1055];
      \nz.mem_1054_sv2v_reg  <= w_data_i[1054];
      \nz.mem_1053_sv2v_reg  <= w_data_i[1053];
      \nz.mem_1052_sv2v_reg  <= w_data_i[1052];
      \nz.mem_1051_sv2v_reg  <= w_data_i[1051];
      \nz.mem_1050_sv2v_reg  <= w_data_i[1050];
      \nz.mem_1049_sv2v_reg  <= w_data_i[1049];
      \nz.mem_1048_sv2v_reg  <= w_data_i[1048];
      \nz.mem_1047_sv2v_reg  <= w_data_i[1047];
      \nz.mem_1046_sv2v_reg  <= w_data_i[1046];
      \nz.mem_1045_sv2v_reg  <= w_data_i[1045];
      \nz.mem_1044_sv2v_reg  <= w_data_i[1044];
      \nz.mem_1043_sv2v_reg  <= w_data_i[1043];
      \nz.mem_1042_sv2v_reg  <= w_data_i[1042];
      \nz.mem_1041_sv2v_reg  <= w_data_i[1041];
      \nz.mem_1040_sv2v_reg  <= w_data_i[1040];
      \nz.mem_1039_sv2v_reg  <= w_data_i[1039];
      \nz.mem_1038_sv2v_reg  <= w_data_i[1038];
      \nz.mem_1037_sv2v_reg  <= w_data_i[1037];
      \nz.mem_1036_sv2v_reg  <= w_data_i[1036];
      \nz.mem_1035_sv2v_reg  <= w_data_i[1035];
      \nz.mem_1034_sv2v_reg  <= w_data_i[1034];
      \nz.mem_1033_sv2v_reg  <= w_data_i[1033];
      \nz.mem_1032_sv2v_reg  <= w_data_i[1032];
      \nz.mem_1031_sv2v_reg  <= w_data_i[1031];
      \nz.mem_1030_sv2v_reg  <= w_data_i[1030];
      \nz.mem_1029_sv2v_reg  <= w_data_i[1029];
      \nz.mem_1028_sv2v_reg  <= w_data_i[1028];
      \nz.mem_1027_sv2v_reg  <= w_data_i[1027];
      \nz.mem_1026_sv2v_reg  <= w_data_i[1026];
      \nz.mem_1025_sv2v_reg  <= w_data_i[1025];
      \nz.mem_1024_sv2v_reg  <= w_data_i[1024];
      \nz.mem_1023_sv2v_reg  <= w_data_i[1023];
      \nz.mem_1022_sv2v_reg  <= w_data_i[1022];
      \nz.mem_1021_sv2v_reg  <= w_data_i[1021];
      \nz.mem_1020_sv2v_reg  <= w_data_i[1020];
      \nz.mem_1019_sv2v_reg  <= w_data_i[1019];
      \nz.mem_1018_sv2v_reg  <= w_data_i[1018];
      \nz.mem_1017_sv2v_reg  <= w_data_i[1017];
      \nz.mem_1016_sv2v_reg  <= w_data_i[1016];
      \nz.mem_1015_sv2v_reg  <= w_data_i[1015];
      \nz.mem_1014_sv2v_reg  <= w_data_i[1014];
      \nz.mem_1013_sv2v_reg  <= w_data_i[1013];
      \nz.mem_1012_sv2v_reg  <= w_data_i[1012];
      \nz.mem_1011_sv2v_reg  <= w_data_i[1011];
      \nz.mem_1010_sv2v_reg  <= w_data_i[1010];
      \nz.mem_1009_sv2v_reg  <= w_data_i[1009];
      \nz.mem_1008_sv2v_reg  <= w_data_i[1008];
      \nz.mem_1007_sv2v_reg  <= w_data_i[1007];
      \nz.mem_1006_sv2v_reg  <= w_data_i[1006];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
    end 
    if(N13) begin
      \nz.mem_1005_sv2v_reg  <= w_data_i[1005];
      \nz.mem_1004_sv2v_reg  <= w_data_i[1004];
      \nz.mem_1003_sv2v_reg  <= w_data_i[1003];
      \nz.mem_1002_sv2v_reg  <= w_data_i[1002];
      \nz.mem_1001_sv2v_reg  <= w_data_i[1001];
      \nz.mem_1000_sv2v_reg  <= w_data_i[1000];
      \nz.mem_999_sv2v_reg  <= w_data_i[999];
      \nz.mem_998_sv2v_reg  <= w_data_i[998];
      \nz.mem_997_sv2v_reg  <= w_data_i[997];
      \nz.mem_996_sv2v_reg  <= w_data_i[996];
      \nz.mem_995_sv2v_reg  <= w_data_i[995];
      \nz.mem_994_sv2v_reg  <= w_data_i[994];
      \nz.mem_993_sv2v_reg  <= w_data_i[993];
      \nz.mem_992_sv2v_reg  <= w_data_i[992];
      \nz.mem_991_sv2v_reg  <= w_data_i[991];
      \nz.mem_990_sv2v_reg  <= w_data_i[990];
      \nz.mem_989_sv2v_reg  <= w_data_i[989];
      \nz.mem_988_sv2v_reg  <= w_data_i[988];
      \nz.mem_987_sv2v_reg  <= w_data_i[987];
      \nz.mem_986_sv2v_reg  <= w_data_i[986];
      \nz.mem_985_sv2v_reg  <= w_data_i[985];
      \nz.mem_984_sv2v_reg  <= w_data_i[984];
      \nz.mem_983_sv2v_reg  <= w_data_i[983];
      \nz.mem_982_sv2v_reg  <= w_data_i[982];
      \nz.mem_981_sv2v_reg  <= w_data_i[981];
      \nz.mem_980_sv2v_reg  <= w_data_i[980];
      \nz.mem_979_sv2v_reg  <= w_data_i[979];
      \nz.mem_978_sv2v_reg  <= w_data_i[978];
      \nz.mem_977_sv2v_reg  <= w_data_i[977];
      \nz.mem_976_sv2v_reg  <= w_data_i[976];
      \nz.mem_975_sv2v_reg  <= w_data_i[975];
      \nz.mem_974_sv2v_reg  <= w_data_i[974];
      \nz.mem_973_sv2v_reg  <= w_data_i[973];
      \nz.mem_972_sv2v_reg  <= w_data_i[972];
      \nz.mem_971_sv2v_reg  <= w_data_i[971];
      \nz.mem_970_sv2v_reg  <= w_data_i[970];
      \nz.mem_969_sv2v_reg  <= w_data_i[969];
      \nz.mem_968_sv2v_reg  <= w_data_i[968];
      \nz.mem_967_sv2v_reg  <= w_data_i[967];
      \nz.mem_966_sv2v_reg  <= w_data_i[966];
      \nz.mem_965_sv2v_reg  <= w_data_i[965];
      \nz.mem_964_sv2v_reg  <= w_data_i[964];
      \nz.mem_963_sv2v_reg  <= w_data_i[963];
      \nz.mem_962_sv2v_reg  <= w_data_i[962];
      \nz.mem_961_sv2v_reg  <= w_data_i[961];
      \nz.mem_960_sv2v_reg  <= w_data_i[960];
      \nz.mem_959_sv2v_reg  <= w_data_i[959];
      \nz.mem_958_sv2v_reg  <= w_data_i[958];
      \nz.mem_957_sv2v_reg  <= w_data_i[957];
      \nz.mem_956_sv2v_reg  <= w_data_i[956];
      \nz.mem_955_sv2v_reg  <= w_data_i[955];
      \nz.mem_954_sv2v_reg  <= w_data_i[954];
      \nz.mem_953_sv2v_reg  <= w_data_i[953];
      \nz.mem_952_sv2v_reg  <= w_data_i[952];
      \nz.mem_951_sv2v_reg  <= w_data_i[951];
      \nz.mem_950_sv2v_reg  <= w_data_i[950];
      \nz.mem_949_sv2v_reg  <= w_data_i[949];
      \nz.mem_948_sv2v_reg  <= w_data_i[948];
      \nz.mem_947_sv2v_reg  <= w_data_i[947];
      \nz.mem_946_sv2v_reg  <= w_data_i[946];
      \nz.mem_945_sv2v_reg  <= w_data_i[945];
      \nz.mem_944_sv2v_reg  <= w_data_i[944];
      \nz.mem_943_sv2v_reg  <= w_data_i[943];
      \nz.mem_942_sv2v_reg  <= w_data_i[942];
      \nz.mem_941_sv2v_reg  <= w_data_i[941];
      \nz.mem_940_sv2v_reg  <= w_data_i[940];
      \nz.mem_939_sv2v_reg  <= w_data_i[939];
      \nz.mem_938_sv2v_reg  <= w_data_i[938];
      \nz.mem_937_sv2v_reg  <= w_data_i[937];
      \nz.mem_936_sv2v_reg  <= w_data_i[936];
      \nz.mem_935_sv2v_reg  <= w_data_i[935];
      \nz.mem_934_sv2v_reg  <= w_data_i[934];
      \nz.mem_933_sv2v_reg  <= w_data_i[933];
      \nz.mem_932_sv2v_reg  <= w_data_i[932];
      \nz.mem_931_sv2v_reg  <= w_data_i[931];
      \nz.mem_930_sv2v_reg  <= w_data_i[930];
      \nz.mem_929_sv2v_reg  <= w_data_i[929];
      \nz.mem_928_sv2v_reg  <= w_data_i[928];
      \nz.mem_927_sv2v_reg  <= w_data_i[927];
      \nz.mem_926_sv2v_reg  <= w_data_i[926];
      \nz.mem_925_sv2v_reg  <= w_data_i[925];
      \nz.mem_924_sv2v_reg  <= w_data_i[924];
      \nz.mem_923_sv2v_reg  <= w_data_i[923];
      \nz.mem_922_sv2v_reg  <= w_data_i[922];
      \nz.mem_921_sv2v_reg  <= w_data_i[921];
      \nz.mem_920_sv2v_reg  <= w_data_i[920];
      \nz.mem_919_sv2v_reg  <= w_data_i[919];
      \nz.mem_918_sv2v_reg  <= w_data_i[918];
      \nz.mem_917_sv2v_reg  <= w_data_i[917];
      \nz.mem_916_sv2v_reg  <= w_data_i[916];
      \nz.mem_915_sv2v_reg  <= w_data_i[915];
      \nz.mem_914_sv2v_reg  <= w_data_i[914];
      \nz.mem_913_sv2v_reg  <= w_data_i[913];
      \nz.mem_912_sv2v_reg  <= w_data_i[912];
      \nz.mem_911_sv2v_reg  <= w_data_i[911];
      \nz.mem_910_sv2v_reg  <= w_data_i[910];
      \nz.mem_909_sv2v_reg  <= w_data_i[909];
      \nz.mem_908_sv2v_reg  <= w_data_i[908];
      \nz.mem_907_sv2v_reg  <= w_data_i[907];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
    end 
    if(N14) begin
      \nz.mem_906_sv2v_reg  <= w_data_i[906];
      \nz.mem_905_sv2v_reg  <= w_data_i[905];
      \nz.mem_904_sv2v_reg  <= w_data_i[904];
      \nz.mem_903_sv2v_reg  <= w_data_i[903];
      \nz.mem_902_sv2v_reg  <= w_data_i[902];
      \nz.mem_901_sv2v_reg  <= w_data_i[901];
      \nz.mem_900_sv2v_reg  <= w_data_i[900];
      \nz.mem_899_sv2v_reg  <= w_data_i[899];
      \nz.mem_898_sv2v_reg  <= w_data_i[898];
      \nz.mem_897_sv2v_reg  <= w_data_i[897];
      \nz.mem_896_sv2v_reg  <= w_data_i[896];
      \nz.mem_895_sv2v_reg  <= w_data_i[895];
      \nz.mem_894_sv2v_reg  <= w_data_i[894];
      \nz.mem_893_sv2v_reg  <= w_data_i[893];
      \nz.mem_892_sv2v_reg  <= w_data_i[892];
      \nz.mem_891_sv2v_reg  <= w_data_i[891];
      \nz.mem_890_sv2v_reg  <= w_data_i[890];
      \nz.mem_889_sv2v_reg  <= w_data_i[889];
      \nz.mem_888_sv2v_reg  <= w_data_i[888];
      \nz.mem_887_sv2v_reg  <= w_data_i[887];
      \nz.mem_886_sv2v_reg  <= w_data_i[886];
      \nz.mem_885_sv2v_reg  <= w_data_i[885];
      \nz.mem_884_sv2v_reg  <= w_data_i[884];
      \nz.mem_883_sv2v_reg  <= w_data_i[883];
      \nz.mem_882_sv2v_reg  <= w_data_i[882];
      \nz.mem_881_sv2v_reg  <= w_data_i[881];
      \nz.mem_880_sv2v_reg  <= w_data_i[880];
      \nz.mem_879_sv2v_reg  <= w_data_i[879];
      \nz.mem_878_sv2v_reg  <= w_data_i[878];
      \nz.mem_877_sv2v_reg  <= w_data_i[877];
      \nz.mem_876_sv2v_reg  <= w_data_i[876];
      \nz.mem_875_sv2v_reg  <= w_data_i[875];
      \nz.mem_874_sv2v_reg  <= w_data_i[874];
      \nz.mem_873_sv2v_reg  <= w_data_i[873];
      \nz.mem_872_sv2v_reg  <= w_data_i[872];
      \nz.mem_871_sv2v_reg  <= w_data_i[871];
      \nz.mem_870_sv2v_reg  <= w_data_i[870];
      \nz.mem_869_sv2v_reg  <= w_data_i[869];
      \nz.mem_868_sv2v_reg  <= w_data_i[868];
      \nz.mem_867_sv2v_reg  <= w_data_i[867];
      \nz.mem_866_sv2v_reg  <= w_data_i[866];
      \nz.mem_865_sv2v_reg  <= w_data_i[865];
      \nz.mem_864_sv2v_reg  <= w_data_i[864];
      \nz.mem_863_sv2v_reg  <= w_data_i[863];
      \nz.mem_862_sv2v_reg  <= w_data_i[862];
      \nz.mem_861_sv2v_reg  <= w_data_i[861];
      \nz.mem_860_sv2v_reg  <= w_data_i[860];
      \nz.mem_859_sv2v_reg  <= w_data_i[859];
      \nz.mem_858_sv2v_reg  <= w_data_i[858];
      \nz.mem_857_sv2v_reg  <= w_data_i[857];
      \nz.mem_856_sv2v_reg  <= w_data_i[856];
      \nz.mem_855_sv2v_reg  <= w_data_i[855];
      \nz.mem_854_sv2v_reg  <= w_data_i[854];
      \nz.mem_853_sv2v_reg  <= w_data_i[853];
      \nz.mem_852_sv2v_reg  <= w_data_i[852];
      \nz.mem_851_sv2v_reg  <= w_data_i[851];
      \nz.mem_850_sv2v_reg  <= w_data_i[850];
      \nz.mem_849_sv2v_reg  <= w_data_i[849];
      \nz.mem_848_sv2v_reg  <= w_data_i[848];
      \nz.mem_847_sv2v_reg  <= w_data_i[847];
      \nz.mem_846_sv2v_reg  <= w_data_i[846];
      \nz.mem_845_sv2v_reg  <= w_data_i[845];
      \nz.mem_844_sv2v_reg  <= w_data_i[844];
      \nz.mem_843_sv2v_reg  <= w_data_i[843];
      \nz.mem_842_sv2v_reg  <= w_data_i[842];
      \nz.mem_841_sv2v_reg  <= w_data_i[841];
      \nz.mem_840_sv2v_reg  <= w_data_i[840];
      \nz.mem_839_sv2v_reg  <= w_data_i[839];
      \nz.mem_838_sv2v_reg  <= w_data_i[838];
      \nz.mem_837_sv2v_reg  <= w_data_i[837];
      \nz.mem_836_sv2v_reg  <= w_data_i[836];
      \nz.mem_835_sv2v_reg  <= w_data_i[835];
      \nz.mem_834_sv2v_reg  <= w_data_i[834];
      \nz.mem_833_sv2v_reg  <= w_data_i[833];
      \nz.mem_832_sv2v_reg  <= w_data_i[832];
      \nz.mem_831_sv2v_reg  <= w_data_i[831];
      \nz.mem_830_sv2v_reg  <= w_data_i[830];
      \nz.mem_829_sv2v_reg  <= w_data_i[829];
      \nz.mem_828_sv2v_reg  <= w_data_i[828];
      \nz.mem_827_sv2v_reg  <= w_data_i[827];
      \nz.mem_826_sv2v_reg  <= w_data_i[826];
      \nz.mem_825_sv2v_reg  <= w_data_i[825];
      \nz.mem_824_sv2v_reg  <= w_data_i[824];
      \nz.mem_823_sv2v_reg  <= w_data_i[823];
      \nz.mem_822_sv2v_reg  <= w_data_i[822];
      \nz.mem_821_sv2v_reg  <= w_data_i[821];
      \nz.mem_820_sv2v_reg  <= w_data_i[820];
      \nz.mem_819_sv2v_reg  <= w_data_i[819];
      \nz.mem_818_sv2v_reg  <= w_data_i[818];
      \nz.mem_817_sv2v_reg  <= w_data_i[817];
      \nz.mem_816_sv2v_reg  <= w_data_i[816];
      \nz.mem_815_sv2v_reg  <= w_data_i[815];
      \nz.mem_814_sv2v_reg  <= w_data_i[814];
      \nz.mem_813_sv2v_reg  <= w_data_i[813];
      \nz.mem_812_sv2v_reg  <= w_data_i[812];
      \nz.mem_811_sv2v_reg  <= w_data_i[811];
      \nz.mem_810_sv2v_reg  <= w_data_i[810];
      \nz.mem_809_sv2v_reg  <= w_data_i[809];
      \nz.mem_808_sv2v_reg  <= w_data_i[808];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
    end 
    if(N15) begin
      \nz.mem_807_sv2v_reg  <= w_data_i[807];
      \nz.mem_806_sv2v_reg  <= w_data_i[806];
      \nz.mem_805_sv2v_reg  <= w_data_i[805];
      \nz.mem_804_sv2v_reg  <= w_data_i[804];
      \nz.mem_803_sv2v_reg  <= w_data_i[803];
      \nz.mem_802_sv2v_reg  <= w_data_i[802];
      \nz.mem_801_sv2v_reg  <= w_data_i[801];
      \nz.mem_800_sv2v_reg  <= w_data_i[800];
      \nz.mem_799_sv2v_reg  <= w_data_i[799];
      \nz.mem_798_sv2v_reg  <= w_data_i[798];
      \nz.mem_797_sv2v_reg  <= w_data_i[797];
      \nz.mem_796_sv2v_reg  <= w_data_i[796];
      \nz.mem_795_sv2v_reg  <= w_data_i[795];
      \nz.mem_794_sv2v_reg  <= w_data_i[794];
      \nz.mem_793_sv2v_reg  <= w_data_i[793];
      \nz.mem_792_sv2v_reg  <= w_data_i[792];
      \nz.mem_791_sv2v_reg  <= w_data_i[791];
      \nz.mem_790_sv2v_reg  <= w_data_i[790];
      \nz.mem_789_sv2v_reg  <= w_data_i[789];
      \nz.mem_788_sv2v_reg  <= w_data_i[788];
      \nz.mem_787_sv2v_reg  <= w_data_i[787];
      \nz.mem_786_sv2v_reg  <= w_data_i[786];
      \nz.mem_785_sv2v_reg  <= w_data_i[785];
      \nz.mem_784_sv2v_reg  <= w_data_i[784];
      \nz.mem_783_sv2v_reg  <= w_data_i[783];
      \nz.mem_782_sv2v_reg  <= w_data_i[782];
      \nz.mem_781_sv2v_reg  <= w_data_i[781];
      \nz.mem_780_sv2v_reg  <= w_data_i[780];
      \nz.mem_779_sv2v_reg  <= w_data_i[779];
      \nz.mem_778_sv2v_reg  <= w_data_i[778];
      \nz.mem_777_sv2v_reg  <= w_data_i[777];
      \nz.mem_776_sv2v_reg  <= w_data_i[776];
      \nz.mem_775_sv2v_reg  <= w_data_i[775];
      \nz.mem_774_sv2v_reg  <= w_data_i[774];
      \nz.mem_773_sv2v_reg  <= w_data_i[773];
      \nz.mem_772_sv2v_reg  <= w_data_i[772];
      \nz.mem_771_sv2v_reg  <= w_data_i[771];
      \nz.mem_770_sv2v_reg  <= w_data_i[770];
      \nz.mem_769_sv2v_reg  <= w_data_i[769];
      \nz.mem_768_sv2v_reg  <= w_data_i[768];
      \nz.mem_767_sv2v_reg  <= w_data_i[767];
      \nz.mem_766_sv2v_reg  <= w_data_i[766];
      \nz.mem_765_sv2v_reg  <= w_data_i[765];
      \nz.mem_764_sv2v_reg  <= w_data_i[764];
      \nz.mem_763_sv2v_reg  <= w_data_i[763];
      \nz.mem_762_sv2v_reg  <= w_data_i[762];
      \nz.mem_761_sv2v_reg  <= w_data_i[761];
      \nz.mem_760_sv2v_reg  <= w_data_i[760];
      \nz.mem_759_sv2v_reg  <= w_data_i[759];
      \nz.mem_758_sv2v_reg  <= w_data_i[758];
      \nz.mem_757_sv2v_reg  <= w_data_i[757];
      \nz.mem_756_sv2v_reg  <= w_data_i[756];
      \nz.mem_755_sv2v_reg  <= w_data_i[755];
      \nz.mem_754_sv2v_reg  <= w_data_i[754];
      \nz.mem_753_sv2v_reg  <= w_data_i[753];
      \nz.mem_752_sv2v_reg  <= w_data_i[752];
      \nz.mem_751_sv2v_reg  <= w_data_i[751];
      \nz.mem_750_sv2v_reg  <= w_data_i[750];
      \nz.mem_749_sv2v_reg  <= w_data_i[749];
      \nz.mem_748_sv2v_reg  <= w_data_i[748];
      \nz.mem_747_sv2v_reg  <= w_data_i[747];
      \nz.mem_746_sv2v_reg  <= w_data_i[746];
      \nz.mem_745_sv2v_reg  <= w_data_i[745];
      \nz.mem_744_sv2v_reg  <= w_data_i[744];
      \nz.mem_743_sv2v_reg  <= w_data_i[743];
      \nz.mem_742_sv2v_reg  <= w_data_i[742];
      \nz.mem_741_sv2v_reg  <= w_data_i[741];
      \nz.mem_740_sv2v_reg  <= w_data_i[740];
      \nz.mem_739_sv2v_reg  <= w_data_i[739];
      \nz.mem_738_sv2v_reg  <= w_data_i[738];
      \nz.mem_737_sv2v_reg  <= w_data_i[737];
      \nz.mem_736_sv2v_reg  <= w_data_i[736];
      \nz.mem_735_sv2v_reg  <= w_data_i[735];
      \nz.mem_734_sv2v_reg  <= w_data_i[734];
      \nz.mem_733_sv2v_reg  <= w_data_i[733];
      \nz.mem_732_sv2v_reg  <= w_data_i[732];
      \nz.mem_731_sv2v_reg  <= w_data_i[731];
      \nz.mem_730_sv2v_reg  <= w_data_i[730];
      \nz.mem_729_sv2v_reg  <= w_data_i[729];
      \nz.mem_728_sv2v_reg  <= w_data_i[728];
      \nz.mem_727_sv2v_reg  <= w_data_i[727];
      \nz.mem_726_sv2v_reg  <= w_data_i[726];
      \nz.mem_725_sv2v_reg  <= w_data_i[725];
      \nz.mem_724_sv2v_reg  <= w_data_i[724];
      \nz.mem_723_sv2v_reg  <= w_data_i[723];
      \nz.mem_722_sv2v_reg  <= w_data_i[722];
      \nz.mem_721_sv2v_reg  <= w_data_i[721];
      \nz.mem_720_sv2v_reg  <= w_data_i[720];
      \nz.mem_719_sv2v_reg  <= w_data_i[719];
      \nz.mem_718_sv2v_reg  <= w_data_i[718];
      \nz.mem_717_sv2v_reg  <= w_data_i[717];
      \nz.mem_716_sv2v_reg  <= w_data_i[716];
      \nz.mem_715_sv2v_reg  <= w_data_i[715];
      \nz.mem_714_sv2v_reg  <= w_data_i[714];
      \nz.mem_713_sv2v_reg  <= w_data_i[713];
      \nz.mem_712_sv2v_reg  <= w_data_i[712];
      \nz.mem_711_sv2v_reg  <= w_data_i[711];
      \nz.mem_710_sv2v_reg  <= w_data_i[710];
      \nz.mem_709_sv2v_reg  <= w_data_i[709];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
    end 
    if(N16) begin
      \nz.mem_708_sv2v_reg  <= w_data_i[708];
      \nz.mem_707_sv2v_reg  <= w_data_i[707];
      \nz.mem_706_sv2v_reg  <= w_data_i[706];
      \nz.mem_705_sv2v_reg  <= w_data_i[705];
      \nz.mem_704_sv2v_reg  <= w_data_i[704];
      \nz.mem_703_sv2v_reg  <= w_data_i[703];
      \nz.mem_702_sv2v_reg  <= w_data_i[702];
      \nz.mem_701_sv2v_reg  <= w_data_i[701];
      \nz.mem_700_sv2v_reg  <= w_data_i[700];
      \nz.mem_699_sv2v_reg  <= w_data_i[699];
      \nz.mem_698_sv2v_reg  <= w_data_i[698];
      \nz.mem_697_sv2v_reg  <= w_data_i[697];
      \nz.mem_696_sv2v_reg  <= w_data_i[696];
      \nz.mem_695_sv2v_reg  <= w_data_i[695];
      \nz.mem_694_sv2v_reg  <= w_data_i[694];
      \nz.mem_693_sv2v_reg  <= w_data_i[693];
      \nz.mem_692_sv2v_reg  <= w_data_i[692];
      \nz.mem_691_sv2v_reg  <= w_data_i[691];
      \nz.mem_690_sv2v_reg  <= w_data_i[690];
      \nz.mem_689_sv2v_reg  <= w_data_i[689];
      \nz.mem_688_sv2v_reg  <= w_data_i[688];
      \nz.mem_687_sv2v_reg  <= w_data_i[687];
      \nz.mem_686_sv2v_reg  <= w_data_i[686];
      \nz.mem_685_sv2v_reg  <= w_data_i[685];
      \nz.mem_684_sv2v_reg  <= w_data_i[684];
      \nz.mem_683_sv2v_reg  <= w_data_i[683];
      \nz.mem_682_sv2v_reg  <= w_data_i[682];
      \nz.mem_681_sv2v_reg  <= w_data_i[681];
      \nz.mem_680_sv2v_reg  <= w_data_i[680];
      \nz.mem_679_sv2v_reg  <= w_data_i[679];
      \nz.mem_678_sv2v_reg  <= w_data_i[678];
      \nz.mem_677_sv2v_reg  <= w_data_i[677];
      \nz.mem_676_sv2v_reg  <= w_data_i[676];
      \nz.mem_675_sv2v_reg  <= w_data_i[675];
      \nz.mem_674_sv2v_reg  <= w_data_i[674];
      \nz.mem_673_sv2v_reg  <= w_data_i[673];
      \nz.mem_672_sv2v_reg  <= w_data_i[672];
      \nz.mem_671_sv2v_reg  <= w_data_i[671];
      \nz.mem_670_sv2v_reg  <= w_data_i[670];
      \nz.mem_669_sv2v_reg  <= w_data_i[669];
      \nz.mem_668_sv2v_reg  <= w_data_i[668];
      \nz.mem_667_sv2v_reg  <= w_data_i[667];
      \nz.mem_666_sv2v_reg  <= w_data_i[666];
      \nz.mem_665_sv2v_reg  <= w_data_i[665];
      \nz.mem_664_sv2v_reg  <= w_data_i[664];
      \nz.mem_663_sv2v_reg  <= w_data_i[663];
      \nz.mem_662_sv2v_reg  <= w_data_i[662];
      \nz.mem_661_sv2v_reg  <= w_data_i[661];
      \nz.mem_660_sv2v_reg  <= w_data_i[660];
      \nz.mem_659_sv2v_reg  <= w_data_i[659];
      \nz.mem_658_sv2v_reg  <= w_data_i[658];
      \nz.mem_657_sv2v_reg  <= w_data_i[657];
      \nz.mem_656_sv2v_reg  <= w_data_i[656];
      \nz.mem_655_sv2v_reg  <= w_data_i[655];
      \nz.mem_654_sv2v_reg  <= w_data_i[654];
      \nz.mem_653_sv2v_reg  <= w_data_i[653];
      \nz.mem_652_sv2v_reg  <= w_data_i[652];
      \nz.mem_651_sv2v_reg  <= w_data_i[651];
      \nz.mem_650_sv2v_reg  <= w_data_i[650];
      \nz.mem_649_sv2v_reg  <= w_data_i[649];
      \nz.mem_648_sv2v_reg  <= w_data_i[648];
      \nz.mem_647_sv2v_reg  <= w_data_i[647];
      \nz.mem_646_sv2v_reg  <= w_data_i[646];
      \nz.mem_645_sv2v_reg  <= w_data_i[645];
      \nz.mem_644_sv2v_reg  <= w_data_i[644];
      \nz.mem_643_sv2v_reg  <= w_data_i[643];
      \nz.mem_642_sv2v_reg  <= w_data_i[642];
      \nz.mem_641_sv2v_reg  <= w_data_i[641];
      \nz.mem_640_sv2v_reg  <= w_data_i[640];
      \nz.mem_639_sv2v_reg  <= w_data_i[639];
      \nz.mem_638_sv2v_reg  <= w_data_i[638];
      \nz.mem_637_sv2v_reg  <= w_data_i[637];
      \nz.mem_636_sv2v_reg  <= w_data_i[636];
      \nz.mem_635_sv2v_reg  <= w_data_i[635];
      \nz.mem_634_sv2v_reg  <= w_data_i[634];
      \nz.mem_633_sv2v_reg  <= w_data_i[633];
      \nz.mem_632_sv2v_reg  <= w_data_i[632];
      \nz.mem_631_sv2v_reg  <= w_data_i[631];
      \nz.mem_630_sv2v_reg  <= w_data_i[630];
      \nz.mem_629_sv2v_reg  <= w_data_i[629];
      \nz.mem_628_sv2v_reg  <= w_data_i[628];
      \nz.mem_627_sv2v_reg  <= w_data_i[627];
      \nz.mem_626_sv2v_reg  <= w_data_i[626];
      \nz.mem_625_sv2v_reg  <= w_data_i[625];
      \nz.mem_624_sv2v_reg  <= w_data_i[624];
      \nz.mem_623_sv2v_reg  <= w_data_i[623];
      \nz.mem_622_sv2v_reg  <= w_data_i[622];
      \nz.mem_621_sv2v_reg  <= w_data_i[621];
      \nz.mem_620_sv2v_reg  <= w_data_i[620];
      \nz.mem_619_sv2v_reg  <= w_data_i[619];
      \nz.mem_618_sv2v_reg  <= w_data_i[618];
      \nz.mem_617_sv2v_reg  <= w_data_i[617];
      \nz.mem_616_sv2v_reg  <= w_data_i[616];
      \nz.mem_615_sv2v_reg  <= w_data_i[615];
      \nz.mem_614_sv2v_reg  <= w_data_i[614];
      \nz.mem_613_sv2v_reg  <= w_data_i[613];
      \nz.mem_612_sv2v_reg  <= w_data_i[612];
      \nz.mem_611_sv2v_reg  <= w_data_i[611];
      \nz.mem_610_sv2v_reg  <= w_data_i[610];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
    end 
    if(N17) begin
      \nz.mem_609_sv2v_reg  <= w_data_i[609];
      \nz.mem_608_sv2v_reg  <= w_data_i[608];
      \nz.mem_607_sv2v_reg  <= w_data_i[607];
      \nz.mem_606_sv2v_reg  <= w_data_i[606];
      \nz.mem_605_sv2v_reg  <= w_data_i[605];
      \nz.mem_604_sv2v_reg  <= w_data_i[604];
      \nz.mem_603_sv2v_reg  <= w_data_i[603];
      \nz.mem_602_sv2v_reg  <= w_data_i[602];
      \nz.mem_601_sv2v_reg  <= w_data_i[601];
      \nz.mem_600_sv2v_reg  <= w_data_i[600];
      \nz.mem_599_sv2v_reg  <= w_data_i[599];
      \nz.mem_598_sv2v_reg  <= w_data_i[598];
      \nz.mem_597_sv2v_reg  <= w_data_i[597];
      \nz.mem_596_sv2v_reg  <= w_data_i[596];
      \nz.mem_595_sv2v_reg  <= w_data_i[595];
      \nz.mem_594_sv2v_reg  <= w_data_i[594];
      \nz.mem_593_sv2v_reg  <= w_data_i[593];
      \nz.mem_592_sv2v_reg  <= w_data_i[592];
      \nz.mem_591_sv2v_reg  <= w_data_i[591];
      \nz.mem_590_sv2v_reg  <= w_data_i[590];
      \nz.mem_589_sv2v_reg  <= w_data_i[589];
      \nz.mem_588_sv2v_reg  <= w_data_i[588];
      \nz.mem_587_sv2v_reg  <= w_data_i[587];
      \nz.mem_586_sv2v_reg  <= w_data_i[586];
      \nz.mem_585_sv2v_reg  <= w_data_i[585];
      \nz.mem_584_sv2v_reg  <= w_data_i[584];
      \nz.mem_583_sv2v_reg  <= w_data_i[583];
      \nz.mem_582_sv2v_reg  <= w_data_i[582];
      \nz.mem_581_sv2v_reg  <= w_data_i[581];
      \nz.mem_580_sv2v_reg  <= w_data_i[580];
      \nz.mem_579_sv2v_reg  <= w_data_i[579];
      \nz.mem_578_sv2v_reg  <= w_data_i[578];
      \nz.mem_577_sv2v_reg  <= w_data_i[577];
      \nz.mem_576_sv2v_reg  <= w_data_i[576];
      \nz.mem_575_sv2v_reg  <= w_data_i[575];
      \nz.mem_574_sv2v_reg  <= w_data_i[574];
      \nz.mem_573_sv2v_reg  <= w_data_i[573];
      \nz.mem_572_sv2v_reg  <= w_data_i[572];
      \nz.mem_571_sv2v_reg  <= w_data_i[571];
      \nz.mem_570_sv2v_reg  <= w_data_i[570];
      \nz.mem_569_sv2v_reg  <= w_data_i[569];
      \nz.mem_568_sv2v_reg  <= w_data_i[568];
      \nz.mem_567_sv2v_reg  <= w_data_i[567];
      \nz.mem_566_sv2v_reg  <= w_data_i[566];
      \nz.mem_565_sv2v_reg  <= w_data_i[565];
      \nz.mem_564_sv2v_reg  <= w_data_i[564];
      \nz.mem_563_sv2v_reg  <= w_data_i[563];
      \nz.mem_562_sv2v_reg  <= w_data_i[562];
      \nz.mem_561_sv2v_reg  <= w_data_i[561];
      \nz.mem_560_sv2v_reg  <= w_data_i[560];
      \nz.mem_559_sv2v_reg  <= w_data_i[559];
      \nz.mem_558_sv2v_reg  <= w_data_i[558];
      \nz.mem_557_sv2v_reg  <= w_data_i[557];
      \nz.mem_556_sv2v_reg  <= w_data_i[556];
      \nz.mem_555_sv2v_reg  <= w_data_i[555];
      \nz.mem_554_sv2v_reg  <= w_data_i[554];
      \nz.mem_553_sv2v_reg  <= w_data_i[553];
      \nz.mem_552_sv2v_reg  <= w_data_i[552];
      \nz.mem_551_sv2v_reg  <= w_data_i[551];
      \nz.mem_550_sv2v_reg  <= w_data_i[550];
      \nz.mem_549_sv2v_reg  <= w_data_i[549];
      \nz.mem_548_sv2v_reg  <= w_data_i[548];
      \nz.mem_547_sv2v_reg  <= w_data_i[547];
      \nz.mem_546_sv2v_reg  <= w_data_i[546];
      \nz.mem_545_sv2v_reg  <= w_data_i[545];
      \nz.mem_544_sv2v_reg  <= w_data_i[544];
      \nz.mem_543_sv2v_reg  <= w_data_i[543];
      \nz.mem_542_sv2v_reg  <= w_data_i[542];
      \nz.mem_541_sv2v_reg  <= w_data_i[541];
      \nz.mem_540_sv2v_reg  <= w_data_i[540];
      \nz.mem_539_sv2v_reg  <= w_data_i[539];
      \nz.mem_538_sv2v_reg  <= w_data_i[538];
      \nz.mem_537_sv2v_reg  <= w_data_i[537];
      \nz.mem_536_sv2v_reg  <= w_data_i[536];
      \nz.mem_535_sv2v_reg  <= w_data_i[535];
      \nz.mem_534_sv2v_reg  <= w_data_i[534];
      \nz.mem_533_sv2v_reg  <= w_data_i[533];
      \nz.mem_532_sv2v_reg  <= w_data_i[532];
      \nz.mem_531_sv2v_reg  <= w_data_i[531];
      \nz.mem_530_sv2v_reg  <= w_data_i[530];
      \nz.mem_529_sv2v_reg  <= w_data_i[529];
      \nz.mem_528_sv2v_reg  <= w_data_i[528];
      \nz.mem_527_sv2v_reg  <= w_data_i[527];
      \nz.mem_526_sv2v_reg  <= w_data_i[526];
      \nz.mem_525_sv2v_reg  <= w_data_i[525];
      \nz.mem_524_sv2v_reg  <= w_data_i[524];
      \nz.mem_523_sv2v_reg  <= w_data_i[523];
      \nz.mem_522_sv2v_reg  <= w_data_i[522];
      \nz.mem_521_sv2v_reg  <= w_data_i[521];
      \nz.mem_520_sv2v_reg  <= w_data_i[520];
      \nz.mem_519_sv2v_reg  <= w_data_i[519];
      \nz.mem_518_sv2v_reg  <= w_data_i[518];
      \nz.mem_517_sv2v_reg  <= w_data_i[517];
      \nz.mem_516_sv2v_reg  <= w_data_i[516];
      \nz.mem_515_sv2v_reg  <= w_data_i[515];
      \nz.mem_514_sv2v_reg  <= w_data_i[514];
      \nz.mem_513_sv2v_reg  <= w_data_i[513];
      \nz.mem_512_sv2v_reg  <= w_data_i[512];
      \nz.mem_511_sv2v_reg  <= w_data_i[511];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
    end 
    if(N18) begin
      \nz.mem_510_sv2v_reg  <= w_data_i[510];
      \nz.mem_509_sv2v_reg  <= w_data_i[509];
      \nz.mem_508_sv2v_reg  <= w_data_i[508];
      \nz.mem_507_sv2v_reg  <= w_data_i[507];
      \nz.mem_506_sv2v_reg  <= w_data_i[506];
      \nz.mem_505_sv2v_reg  <= w_data_i[505];
      \nz.mem_504_sv2v_reg  <= w_data_i[504];
      \nz.mem_503_sv2v_reg  <= w_data_i[503];
      \nz.mem_502_sv2v_reg  <= w_data_i[502];
      \nz.mem_501_sv2v_reg  <= w_data_i[501];
      \nz.mem_500_sv2v_reg  <= w_data_i[500];
      \nz.mem_499_sv2v_reg  <= w_data_i[499];
      \nz.mem_498_sv2v_reg  <= w_data_i[498];
      \nz.mem_497_sv2v_reg  <= w_data_i[497];
      \nz.mem_496_sv2v_reg  <= w_data_i[496];
      \nz.mem_495_sv2v_reg  <= w_data_i[495];
      \nz.mem_494_sv2v_reg  <= w_data_i[494];
      \nz.mem_493_sv2v_reg  <= w_data_i[493];
      \nz.mem_492_sv2v_reg  <= w_data_i[492];
      \nz.mem_491_sv2v_reg  <= w_data_i[491];
      \nz.mem_490_sv2v_reg  <= w_data_i[490];
      \nz.mem_489_sv2v_reg  <= w_data_i[489];
      \nz.mem_488_sv2v_reg  <= w_data_i[488];
      \nz.mem_487_sv2v_reg  <= w_data_i[487];
      \nz.mem_486_sv2v_reg  <= w_data_i[486];
      \nz.mem_485_sv2v_reg  <= w_data_i[485];
      \nz.mem_484_sv2v_reg  <= w_data_i[484];
      \nz.mem_483_sv2v_reg  <= w_data_i[483];
      \nz.mem_482_sv2v_reg  <= w_data_i[482];
      \nz.mem_481_sv2v_reg  <= w_data_i[481];
      \nz.mem_480_sv2v_reg  <= w_data_i[480];
      \nz.mem_479_sv2v_reg  <= w_data_i[479];
      \nz.mem_478_sv2v_reg  <= w_data_i[478];
      \nz.mem_477_sv2v_reg  <= w_data_i[477];
      \nz.mem_476_sv2v_reg  <= w_data_i[476];
      \nz.mem_475_sv2v_reg  <= w_data_i[475];
      \nz.mem_474_sv2v_reg  <= w_data_i[474];
      \nz.mem_473_sv2v_reg  <= w_data_i[473];
      \nz.mem_472_sv2v_reg  <= w_data_i[472];
      \nz.mem_471_sv2v_reg  <= w_data_i[471];
      \nz.mem_470_sv2v_reg  <= w_data_i[470];
      \nz.mem_469_sv2v_reg  <= w_data_i[469];
      \nz.mem_468_sv2v_reg  <= w_data_i[468];
      \nz.mem_467_sv2v_reg  <= w_data_i[467];
      \nz.mem_466_sv2v_reg  <= w_data_i[466];
      \nz.mem_465_sv2v_reg  <= w_data_i[465];
      \nz.mem_464_sv2v_reg  <= w_data_i[464];
      \nz.mem_463_sv2v_reg  <= w_data_i[463];
      \nz.mem_462_sv2v_reg  <= w_data_i[462];
      \nz.mem_461_sv2v_reg  <= w_data_i[461];
      \nz.mem_460_sv2v_reg  <= w_data_i[460];
      \nz.mem_459_sv2v_reg  <= w_data_i[459];
      \nz.mem_458_sv2v_reg  <= w_data_i[458];
      \nz.mem_457_sv2v_reg  <= w_data_i[457];
      \nz.mem_456_sv2v_reg  <= w_data_i[456];
      \nz.mem_455_sv2v_reg  <= w_data_i[455];
      \nz.mem_454_sv2v_reg  <= w_data_i[454];
      \nz.mem_453_sv2v_reg  <= w_data_i[453];
      \nz.mem_452_sv2v_reg  <= w_data_i[452];
      \nz.mem_451_sv2v_reg  <= w_data_i[451];
      \nz.mem_450_sv2v_reg  <= w_data_i[450];
      \nz.mem_449_sv2v_reg  <= w_data_i[449];
      \nz.mem_448_sv2v_reg  <= w_data_i[448];
      \nz.mem_447_sv2v_reg  <= w_data_i[447];
      \nz.mem_446_sv2v_reg  <= w_data_i[446];
      \nz.mem_445_sv2v_reg  <= w_data_i[445];
      \nz.mem_444_sv2v_reg  <= w_data_i[444];
      \nz.mem_443_sv2v_reg  <= w_data_i[443];
      \nz.mem_442_sv2v_reg  <= w_data_i[442];
      \nz.mem_441_sv2v_reg  <= w_data_i[441];
      \nz.mem_440_sv2v_reg  <= w_data_i[440];
      \nz.mem_439_sv2v_reg  <= w_data_i[439];
      \nz.mem_438_sv2v_reg  <= w_data_i[438];
      \nz.mem_437_sv2v_reg  <= w_data_i[437];
      \nz.mem_436_sv2v_reg  <= w_data_i[436];
      \nz.mem_435_sv2v_reg  <= w_data_i[435];
      \nz.mem_434_sv2v_reg  <= w_data_i[434];
      \nz.mem_433_sv2v_reg  <= w_data_i[433];
      \nz.mem_432_sv2v_reg  <= w_data_i[432];
      \nz.mem_431_sv2v_reg  <= w_data_i[431];
      \nz.mem_430_sv2v_reg  <= w_data_i[430];
      \nz.mem_429_sv2v_reg  <= w_data_i[429];
      \nz.mem_428_sv2v_reg  <= w_data_i[428];
      \nz.mem_427_sv2v_reg  <= w_data_i[427];
      \nz.mem_426_sv2v_reg  <= w_data_i[426];
      \nz.mem_425_sv2v_reg  <= w_data_i[425];
      \nz.mem_424_sv2v_reg  <= w_data_i[424];
      \nz.mem_423_sv2v_reg  <= w_data_i[423];
      \nz.mem_422_sv2v_reg  <= w_data_i[422];
      \nz.mem_421_sv2v_reg  <= w_data_i[421];
      \nz.mem_420_sv2v_reg  <= w_data_i[420];
      \nz.mem_419_sv2v_reg  <= w_data_i[419];
      \nz.mem_418_sv2v_reg  <= w_data_i[418];
      \nz.mem_417_sv2v_reg  <= w_data_i[417];
      \nz.mem_416_sv2v_reg  <= w_data_i[416];
      \nz.mem_415_sv2v_reg  <= w_data_i[415];
      \nz.mem_414_sv2v_reg  <= w_data_i[414];
      \nz.mem_413_sv2v_reg  <= w_data_i[413];
      \nz.mem_412_sv2v_reg  <= w_data_i[412];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
    end 
    if(N19) begin
      \nz.mem_411_sv2v_reg  <= w_data_i[411];
      \nz.mem_410_sv2v_reg  <= w_data_i[410];
      \nz.mem_409_sv2v_reg  <= w_data_i[409];
      \nz.mem_408_sv2v_reg  <= w_data_i[408];
      \nz.mem_407_sv2v_reg  <= w_data_i[407];
      \nz.mem_406_sv2v_reg  <= w_data_i[406];
      \nz.mem_405_sv2v_reg  <= w_data_i[405];
      \nz.mem_404_sv2v_reg  <= w_data_i[404];
      \nz.mem_403_sv2v_reg  <= w_data_i[403];
      \nz.mem_402_sv2v_reg  <= w_data_i[402];
      \nz.mem_401_sv2v_reg  <= w_data_i[401];
      \nz.mem_400_sv2v_reg  <= w_data_i[400];
      \nz.mem_399_sv2v_reg  <= w_data_i[399];
      \nz.mem_398_sv2v_reg  <= w_data_i[398];
      \nz.mem_397_sv2v_reg  <= w_data_i[397];
      \nz.mem_396_sv2v_reg  <= w_data_i[396];
      \nz.mem_395_sv2v_reg  <= w_data_i[395];
      \nz.mem_394_sv2v_reg  <= w_data_i[394];
      \nz.mem_393_sv2v_reg  <= w_data_i[393];
      \nz.mem_392_sv2v_reg  <= w_data_i[392];
      \nz.mem_391_sv2v_reg  <= w_data_i[391];
      \nz.mem_390_sv2v_reg  <= w_data_i[390];
      \nz.mem_389_sv2v_reg  <= w_data_i[389];
      \nz.mem_388_sv2v_reg  <= w_data_i[388];
      \nz.mem_387_sv2v_reg  <= w_data_i[387];
      \nz.mem_386_sv2v_reg  <= w_data_i[386];
      \nz.mem_385_sv2v_reg  <= w_data_i[385];
      \nz.mem_384_sv2v_reg  <= w_data_i[384];
      \nz.mem_383_sv2v_reg  <= w_data_i[383];
      \nz.mem_382_sv2v_reg  <= w_data_i[382];
      \nz.mem_381_sv2v_reg  <= w_data_i[381];
      \nz.mem_380_sv2v_reg  <= w_data_i[380];
      \nz.mem_379_sv2v_reg  <= w_data_i[379];
      \nz.mem_378_sv2v_reg  <= w_data_i[378];
      \nz.mem_377_sv2v_reg  <= w_data_i[377];
      \nz.mem_376_sv2v_reg  <= w_data_i[376];
      \nz.mem_375_sv2v_reg  <= w_data_i[375];
      \nz.mem_374_sv2v_reg  <= w_data_i[374];
      \nz.mem_373_sv2v_reg  <= w_data_i[373];
      \nz.mem_372_sv2v_reg  <= w_data_i[372];
      \nz.mem_371_sv2v_reg  <= w_data_i[371];
      \nz.mem_370_sv2v_reg  <= w_data_i[370];
      \nz.mem_369_sv2v_reg  <= w_data_i[369];
      \nz.mem_368_sv2v_reg  <= w_data_i[368];
      \nz.mem_367_sv2v_reg  <= w_data_i[367];
      \nz.mem_366_sv2v_reg  <= w_data_i[366];
      \nz.mem_365_sv2v_reg  <= w_data_i[365];
      \nz.mem_364_sv2v_reg  <= w_data_i[364];
      \nz.mem_363_sv2v_reg  <= w_data_i[363];
      \nz.mem_362_sv2v_reg  <= w_data_i[362];
      \nz.mem_361_sv2v_reg  <= w_data_i[361];
      \nz.mem_360_sv2v_reg  <= w_data_i[360];
      \nz.mem_359_sv2v_reg  <= w_data_i[359];
      \nz.mem_358_sv2v_reg  <= w_data_i[358];
      \nz.mem_357_sv2v_reg  <= w_data_i[357];
      \nz.mem_356_sv2v_reg  <= w_data_i[356];
      \nz.mem_355_sv2v_reg  <= w_data_i[355];
      \nz.mem_354_sv2v_reg  <= w_data_i[354];
      \nz.mem_353_sv2v_reg  <= w_data_i[353];
      \nz.mem_352_sv2v_reg  <= w_data_i[352];
      \nz.mem_351_sv2v_reg  <= w_data_i[351];
      \nz.mem_350_sv2v_reg  <= w_data_i[350];
      \nz.mem_349_sv2v_reg  <= w_data_i[349];
      \nz.mem_348_sv2v_reg  <= w_data_i[348];
      \nz.mem_347_sv2v_reg  <= w_data_i[347];
      \nz.mem_346_sv2v_reg  <= w_data_i[346];
      \nz.mem_345_sv2v_reg  <= w_data_i[345];
      \nz.mem_344_sv2v_reg  <= w_data_i[344];
      \nz.mem_343_sv2v_reg  <= w_data_i[343];
      \nz.mem_342_sv2v_reg  <= w_data_i[342];
      \nz.mem_341_sv2v_reg  <= w_data_i[341];
      \nz.mem_340_sv2v_reg  <= w_data_i[340];
      \nz.mem_339_sv2v_reg  <= w_data_i[339];
      \nz.mem_338_sv2v_reg  <= w_data_i[338];
      \nz.mem_337_sv2v_reg  <= w_data_i[337];
      \nz.mem_336_sv2v_reg  <= w_data_i[336];
      \nz.mem_335_sv2v_reg  <= w_data_i[335];
      \nz.mem_334_sv2v_reg  <= w_data_i[334];
      \nz.mem_333_sv2v_reg  <= w_data_i[333];
      \nz.mem_332_sv2v_reg  <= w_data_i[332];
      \nz.mem_331_sv2v_reg  <= w_data_i[331];
      \nz.mem_330_sv2v_reg  <= w_data_i[330];
      \nz.mem_329_sv2v_reg  <= w_data_i[329];
      \nz.mem_328_sv2v_reg  <= w_data_i[328];
      \nz.mem_327_sv2v_reg  <= w_data_i[327];
      \nz.mem_326_sv2v_reg  <= w_data_i[326];
      \nz.mem_325_sv2v_reg  <= w_data_i[325];
      \nz.mem_324_sv2v_reg  <= w_data_i[324];
      \nz.mem_323_sv2v_reg  <= w_data_i[323];
      \nz.mem_322_sv2v_reg  <= w_data_i[322];
      \nz.mem_321_sv2v_reg  <= w_data_i[321];
      \nz.mem_320_sv2v_reg  <= w_data_i[320];
      \nz.mem_319_sv2v_reg  <= w_data_i[319];
      \nz.mem_318_sv2v_reg  <= w_data_i[318];
      \nz.mem_317_sv2v_reg  <= w_data_i[317];
      \nz.mem_316_sv2v_reg  <= w_data_i[316];
      \nz.mem_315_sv2v_reg  <= w_data_i[315];
      \nz.mem_314_sv2v_reg  <= w_data_i[314];
      \nz.mem_313_sv2v_reg  <= w_data_i[313];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
    end 
    if(N20) begin
      \nz.mem_312_sv2v_reg  <= w_data_i[312];
      \nz.mem_311_sv2v_reg  <= w_data_i[311];
      \nz.mem_310_sv2v_reg  <= w_data_i[310];
      \nz.mem_309_sv2v_reg  <= w_data_i[309];
      \nz.mem_308_sv2v_reg  <= w_data_i[308];
      \nz.mem_307_sv2v_reg  <= w_data_i[307];
      \nz.mem_306_sv2v_reg  <= w_data_i[306];
      \nz.mem_305_sv2v_reg  <= w_data_i[305];
      \nz.mem_304_sv2v_reg  <= w_data_i[304];
      \nz.mem_303_sv2v_reg  <= w_data_i[303];
      \nz.mem_302_sv2v_reg  <= w_data_i[302];
      \nz.mem_301_sv2v_reg  <= w_data_i[301];
      \nz.mem_300_sv2v_reg  <= w_data_i[300];
      \nz.mem_299_sv2v_reg  <= w_data_i[299];
      \nz.mem_298_sv2v_reg  <= w_data_i[298];
      \nz.mem_297_sv2v_reg  <= w_data_i[297];
      \nz.mem_296_sv2v_reg  <= w_data_i[296];
      \nz.mem_295_sv2v_reg  <= w_data_i[295];
      \nz.mem_294_sv2v_reg  <= w_data_i[294];
      \nz.mem_293_sv2v_reg  <= w_data_i[293];
      \nz.mem_292_sv2v_reg  <= w_data_i[292];
      \nz.mem_291_sv2v_reg  <= w_data_i[291];
      \nz.mem_290_sv2v_reg  <= w_data_i[290];
      \nz.mem_289_sv2v_reg  <= w_data_i[289];
      \nz.mem_288_sv2v_reg  <= w_data_i[288];
      \nz.mem_287_sv2v_reg  <= w_data_i[287];
      \nz.mem_286_sv2v_reg  <= w_data_i[286];
      \nz.mem_285_sv2v_reg  <= w_data_i[285];
      \nz.mem_284_sv2v_reg  <= w_data_i[284];
      \nz.mem_283_sv2v_reg  <= w_data_i[283];
      \nz.mem_282_sv2v_reg  <= w_data_i[282];
      \nz.mem_281_sv2v_reg  <= w_data_i[281];
      \nz.mem_280_sv2v_reg  <= w_data_i[280];
      \nz.mem_279_sv2v_reg  <= w_data_i[279];
      \nz.mem_278_sv2v_reg  <= w_data_i[278];
      \nz.mem_277_sv2v_reg  <= w_data_i[277];
      \nz.mem_276_sv2v_reg  <= w_data_i[276];
      \nz.mem_275_sv2v_reg  <= w_data_i[275];
      \nz.mem_274_sv2v_reg  <= w_data_i[274];
      \nz.mem_273_sv2v_reg  <= w_data_i[273];
      \nz.mem_272_sv2v_reg  <= w_data_i[272];
      \nz.mem_271_sv2v_reg  <= w_data_i[271];
      \nz.mem_270_sv2v_reg  <= w_data_i[270];
      \nz.mem_269_sv2v_reg  <= w_data_i[269];
      \nz.mem_268_sv2v_reg  <= w_data_i[268];
      \nz.mem_267_sv2v_reg  <= w_data_i[267];
      \nz.mem_266_sv2v_reg  <= w_data_i[266];
      \nz.mem_265_sv2v_reg  <= w_data_i[265];
      \nz.mem_264_sv2v_reg  <= w_data_i[264];
      \nz.mem_263_sv2v_reg  <= w_data_i[263];
      \nz.mem_262_sv2v_reg  <= w_data_i[262];
      \nz.mem_261_sv2v_reg  <= w_data_i[261];
      \nz.mem_260_sv2v_reg  <= w_data_i[260];
      \nz.mem_259_sv2v_reg  <= w_data_i[259];
      \nz.mem_258_sv2v_reg  <= w_data_i[258];
      \nz.mem_257_sv2v_reg  <= w_data_i[257];
      \nz.mem_256_sv2v_reg  <= w_data_i[256];
      \nz.mem_255_sv2v_reg  <= w_data_i[255];
      \nz.mem_254_sv2v_reg  <= w_data_i[254];
      \nz.mem_253_sv2v_reg  <= w_data_i[253];
      \nz.mem_252_sv2v_reg  <= w_data_i[252];
      \nz.mem_251_sv2v_reg  <= w_data_i[251];
      \nz.mem_250_sv2v_reg  <= w_data_i[250];
      \nz.mem_249_sv2v_reg  <= w_data_i[249];
      \nz.mem_248_sv2v_reg  <= w_data_i[248];
      \nz.mem_247_sv2v_reg  <= w_data_i[247];
      \nz.mem_246_sv2v_reg  <= w_data_i[246];
      \nz.mem_245_sv2v_reg  <= w_data_i[245];
      \nz.mem_244_sv2v_reg  <= w_data_i[244];
      \nz.mem_243_sv2v_reg  <= w_data_i[243];
      \nz.mem_242_sv2v_reg  <= w_data_i[242];
      \nz.mem_241_sv2v_reg  <= w_data_i[241];
      \nz.mem_240_sv2v_reg  <= w_data_i[240];
      \nz.mem_239_sv2v_reg  <= w_data_i[239];
      \nz.mem_238_sv2v_reg  <= w_data_i[238];
      \nz.mem_237_sv2v_reg  <= w_data_i[237];
      \nz.mem_236_sv2v_reg  <= w_data_i[236];
      \nz.mem_235_sv2v_reg  <= w_data_i[235];
      \nz.mem_234_sv2v_reg  <= w_data_i[234];
      \nz.mem_233_sv2v_reg  <= w_data_i[233];
      \nz.mem_232_sv2v_reg  <= w_data_i[232];
      \nz.mem_231_sv2v_reg  <= w_data_i[231];
      \nz.mem_230_sv2v_reg  <= w_data_i[230];
      \nz.mem_229_sv2v_reg  <= w_data_i[229];
      \nz.mem_228_sv2v_reg  <= w_data_i[228];
      \nz.mem_227_sv2v_reg  <= w_data_i[227];
      \nz.mem_226_sv2v_reg  <= w_data_i[226];
      \nz.mem_225_sv2v_reg  <= w_data_i[225];
      \nz.mem_224_sv2v_reg  <= w_data_i[224];
      \nz.mem_223_sv2v_reg  <= w_data_i[223];
      \nz.mem_222_sv2v_reg  <= w_data_i[222];
      \nz.mem_221_sv2v_reg  <= w_data_i[221];
      \nz.mem_220_sv2v_reg  <= w_data_i[220];
      \nz.mem_219_sv2v_reg  <= w_data_i[219];
      \nz.mem_218_sv2v_reg  <= w_data_i[218];
      \nz.mem_217_sv2v_reg  <= w_data_i[217];
      \nz.mem_216_sv2v_reg  <= w_data_i[216];
      \nz.mem_215_sv2v_reg  <= w_data_i[215];
      \nz.mem_214_sv2v_reg  <= w_data_i[214];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
    end 
    if(N21) begin
      \nz.mem_213_sv2v_reg  <= w_data_i[213];
      \nz.mem_212_sv2v_reg  <= w_data_i[212];
      \nz.mem_211_sv2v_reg  <= w_data_i[211];
      \nz.mem_210_sv2v_reg  <= w_data_i[210];
      \nz.mem_209_sv2v_reg  <= w_data_i[209];
      \nz.mem_208_sv2v_reg  <= w_data_i[208];
      \nz.mem_207_sv2v_reg  <= w_data_i[207];
      \nz.mem_206_sv2v_reg  <= w_data_i[206];
      \nz.mem_205_sv2v_reg  <= w_data_i[205];
      \nz.mem_204_sv2v_reg  <= w_data_i[204];
      \nz.mem_203_sv2v_reg  <= w_data_i[203];
      \nz.mem_202_sv2v_reg  <= w_data_i[202];
      \nz.mem_201_sv2v_reg  <= w_data_i[201];
      \nz.mem_200_sv2v_reg  <= w_data_i[200];
      \nz.mem_199_sv2v_reg  <= w_data_i[199];
      \nz.mem_198_sv2v_reg  <= w_data_i[198];
      \nz.mem_197_sv2v_reg  <= w_data_i[197];
      \nz.mem_196_sv2v_reg  <= w_data_i[196];
      \nz.mem_195_sv2v_reg  <= w_data_i[195];
      \nz.mem_194_sv2v_reg  <= w_data_i[194];
      \nz.mem_193_sv2v_reg  <= w_data_i[193];
      \nz.mem_192_sv2v_reg  <= w_data_i[192];
      \nz.mem_191_sv2v_reg  <= w_data_i[191];
      \nz.mem_190_sv2v_reg  <= w_data_i[190];
      \nz.mem_189_sv2v_reg  <= w_data_i[189];
      \nz.mem_188_sv2v_reg  <= w_data_i[188];
      \nz.mem_187_sv2v_reg  <= w_data_i[187];
      \nz.mem_186_sv2v_reg  <= w_data_i[186];
      \nz.mem_185_sv2v_reg  <= w_data_i[185];
      \nz.mem_184_sv2v_reg  <= w_data_i[184];
      \nz.mem_183_sv2v_reg  <= w_data_i[183];
      \nz.mem_182_sv2v_reg  <= w_data_i[182];
      \nz.mem_181_sv2v_reg  <= w_data_i[181];
      \nz.mem_180_sv2v_reg  <= w_data_i[180];
      \nz.mem_179_sv2v_reg  <= w_data_i[179];
      \nz.mem_178_sv2v_reg  <= w_data_i[178];
      \nz.mem_177_sv2v_reg  <= w_data_i[177];
      \nz.mem_176_sv2v_reg  <= w_data_i[176];
      \nz.mem_175_sv2v_reg  <= w_data_i[175];
      \nz.mem_174_sv2v_reg  <= w_data_i[174];
      \nz.mem_173_sv2v_reg  <= w_data_i[173];
      \nz.mem_172_sv2v_reg  <= w_data_i[172];
      \nz.mem_171_sv2v_reg  <= w_data_i[171];
      \nz.mem_170_sv2v_reg  <= w_data_i[170];
      \nz.mem_169_sv2v_reg  <= w_data_i[169];
      \nz.mem_168_sv2v_reg  <= w_data_i[168];
      \nz.mem_167_sv2v_reg  <= w_data_i[167];
      \nz.mem_166_sv2v_reg  <= w_data_i[166];
      \nz.mem_165_sv2v_reg  <= w_data_i[165];
      \nz.mem_164_sv2v_reg  <= w_data_i[164];
      \nz.mem_163_sv2v_reg  <= w_data_i[163];
      \nz.mem_162_sv2v_reg  <= w_data_i[162];
      \nz.mem_161_sv2v_reg  <= w_data_i[161];
      \nz.mem_160_sv2v_reg  <= w_data_i[160];
      \nz.mem_159_sv2v_reg  <= w_data_i[159];
      \nz.mem_158_sv2v_reg  <= w_data_i[158];
      \nz.mem_157_sv2v_reg  <= w_data_i[157];
      \nz.mem_156_sv2v_reg  <= w_data_i[156];
      \nz.mem_155_sv2v_reg  <= w_data_i[155];
      \nz.mem_154_sv2v_reg  <= w_data_i[154];
      \nz.mem_153_sv2v_reg  <= w_data_i[153];
      \nz.mem_152_sv2v_reg  <= w_data_i[152];
      \nz.mem_151_sv2v_reg  <= w_data_i[151];
      \nz.mem_150_sv2v_reg  <= w_data_i[150];
      \nz.mem_149_sv2v_reg  <= w_data_i[149];
      \nz.mem_148_sv2v_reg  <= w_data_i[148];
      \nz.mem_147_sv2v_reg  <= w_data_i[147];
      \nz.mem_146_sv2v_reg  <= w_data_i[146];
      \nz.mem_145_sv2v_reg  <= w_data_i[145];
      \nz.mem_144_sv2v_reg  <= w_data_i[144];
      \nz.mem_143_sv2v_reg  <= w_data_i[143];
      \nz.mem_142_sv2v_reg  <= w_data_i[142];
      \nz.mem_141_sv2v_reg  <= w_data_i[141];
      \nz.mem_140_sv2v_reg  <= w_data_i[140];
      \nz.mem_139_sv2v_reg  <= w_data_i[139];
      \nz.mem_138_sv2v_reg  <= w_data_i[138];
      \nz.mem_137_sv2v_reg  <= w_data_i[137];
      \nz.mem_136_sv2v_reg  <= w_data_i[136];
      \nz.mem_135_sv2v_reg  <= w_data_i[135];
      \nz.mem_134_sv2v_reg  <= w_data_i[134];
      \nz.mem_133_sv2v_reg  <= w_data_i[133];
      \nz.mem_132_sv2v_reg  <= w_data_i[132];
      \nz.mem_131_sv2v_reg  <= w_data_i[131];
      \nz.mem_130_sv2v_reg  <= w_data_i[130];
      \nz.mem_129_sv2v_reg  <= w_data_i[129];
      \nz.mem_128_sv2v_reg  <= w_data_i[128];
      \nz.mem_127_sv2v_reg  <= w_data_i[127];
      \nz.mem_126_sv2v_reg  <= w_data_i[126];
      \nz.mem_125_sv2v_reg  <= w_data_i[125];
      \nz.mem_124_sv2v_reg  <= w_data_i[124];
      \nz.mem_123_sv2v_reg  <= w_data_i[123];
      \nz.mem_122_sv2v_reg  <= w_data_i[122];
      \nz.mem_121_sv2v_reg  <= w_data_i[121];
      \nz.mem_120_sv2v_reg  <= w_data_i[120];
      \nz.mem_119_sv2v_reg  <= w_data_i[119];
      \nz.mem_118_sv2v_reg  <= w_data_i[118];
      \nz.mem_117_sv2v_reg  <= w_data_i[117];
      \nz.mem_116_sv2v_reg  <= w_data_i[116];
      \nz.mem_115_sv2v_reg  <= w_data_i[115];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
    end 
    if(N22) begin
      \nz.mem_114_sv2v_reg  <= w_data_i[114];
      \nz.mem_113_sv2v_reg  <= w_data_i[113];
      \nz.mem_112_sv2v_reg  <= w_data_i[112];
      \nz.mem_111_sv2v_reg  <= w_data_i[111];
      \nz.mem_110_sv2v_reg  <= w_data_i[110];
      \nz.mem_109_sv2v_reg  <= w_data_i[109];
      \nz.mem_108_sv2v_reg  <= w_data_i[108];
      \nz.mem_107_sv2v_reg  <= w_data_i[107];
      \nz.mem_106_sv2v_reg  <= w_data_i[106];
      \nz.mem_105_sv2v_reg  <= w_data_i[105];
      \nz.mem_104_sv2v_reg  <= w_data_i[104];
      \nz.mem_103_sv2v_reg  <= w_data_i[103];
      \nz.mem_102_sv2v_reg  <= w_data_i[102];
      \nz.mem_101_sv2v_reg  <= w_data_i[101];
      \nz.mem_100_sv2v_reg  <= w_data_i[100];
      \nz.mem_99_sv2v_reg  <= w_data_i[99];
      \nz.mem_98_sv2v_reg  <= w_data_i[98];
      \nz.mem_97_sv2v_reg  <= w_data_i[97];
      \nz.mem_96_sv2v_reg  <= w_data_i[96];
      \nz.mem_95_sv2v_reg  <= w_data_i[95];
      \nz.mem_94_sv2v_reg  <= w_data_i[94];
      \nz.mem_93_sv2v_reg  <= w_data_i[93];
      \nz.mem_92_sv2v_reg  <= w_data_i[92];
      \nz.mem_91_sv2v_reg  <= w_data_i[91];
      \nz.mem_90_sv2v_reg  <= w_data_i[90];
      \nz.mem_89_sv2v_reg  <= w_data_i[89];
      \nz.mem_88_sv2v_reg  <= w_data_i[88];
      \nz.mem_87_sv2v_reg  <= w_data_i[87];
      \nz.mem_86_sv2v_reg  <= w_data_i[86];
      \nz.mem_85_sv2v_reg  <= w_data_i[85];
      \nz.mem_84_sv2v_reg  <= w_data_i[84];
      \nz.mem_83_sv2v_reg  <= w_data_i[83];
      \nz.mem_82_sv2v_reg  <= w_data_i[82];
      \nz.mem_81_sv2v_reg  <= w_data_i[81];
      \nz.mem_80_sv2v_reg  <= w_data_i[80];
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p1600_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [1599:0] w_data_i;
  input [0:0] r_addr_i;
  output [1599:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [1599:0] r_data_o;

  bsg_mem_1r1w_synth_width_p1600_els_p2_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p1600
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [1599:0] data_i;
  output [1599:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [1599:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p1600_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p49_init_val_p0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [5:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [5:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N2,N3,N7,N30,N19;
  reg count_o_5_sv2v_reg,count_o_4_sv2v_reg,count_o_3_sv2v_reg,count_o_2_sv2v_reg,
  count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[5] = count_o_5_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N19 = reset_i | clear_i;
  assign { N11, N10, N9, N8, N6, N5 } = count_o + 1'b1;
  assign N12 = (N0)? 1'b1 : 
               (N7)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N14 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N13 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N18;
  assign N15 = ~reset_i;
  assign N16 = ~clear_i;
  assign N17 = N15 & N16;
  assign N18 = up_i & N17;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N16;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N19) begin
      count_o_5_sv2v_reg <= 1'b0;
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N14) begin
      count_o_5_sv2v_reg <= N11;
      count_o_4_sv2v_reg <= N10;
      count_o_3_sv2v_reg <= N9;
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N12) begin
      count_o_0_sv2v_reg <= N13;
    end 
  end


endmodule



module bsg_mux_width_p32_els_p50
(
  data_i,
  sel_i,
  data_o
);

  input [1599:0] data_i;
  input [5:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312;
  assign N0 = N4 & N5;
  assign N1 = N0 & N6;
  assign N2 = N1 & N7;
  assign N3 = N2 & N8;
  assign N263 = N3 & N9;
  assign N4 = ~sel_i[5];
  assign N5 = ~sel_i[4];
  assign N6 = ~sel_i[3];
  assign N7 = ~sel_i[2];
  assign N8 = ~sel_i[0];
  assign N9 = ~sel_i[1];
  assign N10 = sel_i[5] & N14;
  assign N11 = N10 & N15;
  assign N12 = N11 & N16;
  assign N13 = N12 & N17;
  assign N264 = N13 & N18;
  assign N14 = ~sel_i[4];
  assign N15 = ~sel_i[3];
  assign N16 = ~sel_i[2];
  assign N17 = ~sel_i[0];
  assign N18 = ~sel_i[1];
  assign N19 = N23 & N24;
  assign N20 = N19 & N25;
  assign N21 = N20 & N26;
  assign N22 = N21 & sel_i[0];
  assign N265 = N22 & N27;
  assign N23 = ~sel_i[5];
  assign N24 = ~sel_i[4];
  assign N25 = ~sel_i[3];
  assign N26 = ~sel_i[2];
  assign N27 = ~sel_i[1];
  assign N28 = N32 & N33;
  assign N29 = N28 & N34;
  assign N30 = N29 & N35;
  assign N31 = N30 & N36;
  assign N267 = N31 & sel_i[1];
  assign N32 = ~sel_i[5];
  assign N33 = ~sel_i[4];
  assign N34 = ~sel_i[3];
  assign N35 = ~sel_i[2];
  assign N36 = ~sel_i[0];
  assign N37 = N41 & N42;
  assign N38 = N37 & N43;
  assign N39 = N38 & N44;
  assign N40 = N39 & sel_i[0];
  assign N269 = N40 & sel_i[1];
  assign N41 = ~sel_i[5];
  assign N42 = ~sel_i[4];
  assign N43 = ~sel_i[3];
  assign N44 = ~sel_i[2];
  assign N45 = N49 & N50;
  assign N46 = N45 & N51;
  assign N47 = N46 & sel_i[2];
  assign N48 = N47 & N52;
  assign N271 = N48 & N53;
  assign N49 = ~sel_i[5];
  assign N50 = ~sel_i[4];
  assign N51 = ~sel_i[3];
  assign N52 = ~sel_i[0];
  assign N53 = ~sel_i[1];
  assign N54 = N58 & N59;
  assign N55 = N54 & N60;
  assign N56 = N55 & sel_i[2];
  assign N57 = N56 & sel_i[0];
  assign N273 = N57 & N61;
  assign N58 = ~sel_i[5];
  assign N59 = ~sel_i[4];
  assign N60 = ~sel_i[3];
  assign N61 = ~sel_i[1];
  assign N62 = N66 & N67;
  assign N63 = N62 & N68;
  assign N64 = N63 & sel_i[2];
  assign N65 = N64 & N69;
  assign N275 = N65 & sel_i[1];
  assign N66 = ~sel_i[5];
  assign N67 = ~sel_i[4];
  assign N68 = ~sel_i[3];
  assign N69 = ~sel_i[0];
  assign N70 = N74 & N75;
  assign N71 = N70 & N76;
  assign N72 = N71 & sel_i[2];
  assign N73 = N72 & sel_i[0];
  assign N277 = N73 & sel_i[1];
  assign N74 = ~sel_i[5];
  assign N75 = ~sel_i[4];
  assign N76 = ~sel_i[3];
  assign N77 = N81 & N82;
  assign N78 = N77 & sel_i[3];
  assign N79 = N78 & N83;
  assign N80 = N79 & N84;
  assign N279 = N80 & N85;
  assign N81 = ~sel_i[5];
  assign N82 = ~sel_i[4];
  assign N83 = ~sel_i[2];
  assign N84 = ~sel_i[0];
  assign N85 = ~sel_i[1];
  assign N86 = N90 & N91;
  assign N87 = N86 & sel_i[3];
  assign N88 = N87 & N92;
  assign N89 = N88 & sel_i[0];
  assign N281 = N89 & N93;
  assign N90 = ~sel_i[5];
  assign N91 = ~sel_i[4];
  assign N92 = ~sel_i[2];
  assign N93 = ~sel_i[1];
  assign N94 = N98 & N99;
  assign N95 = N94 & sel_i[3];
  assign N96 = N95 & N100;
  assign N97 = N96 & N101;
  assign N283 = N97 & sel_i[1];
  assign N98 = ~sel_i[5];
  assign N99 = ~sel_i[4];
  assign N100 = ~sel_i[2];
  assign N101 = ~sel_i[0];
  assign N102 = N106 & N107;
  assign N103 = N102 & sel_i[3];
  assign N104 = N103 & N108;
  assign N105 = N104 & sel_i[0];
  assign N285 = N105 & sel_i[1];
  assign N106 = ~sel_i[5];
  assign N107 = ~sel_i[4];
  assign N108 = ~sel_i[2];
  assign N109 = N113 & N114;
  assign N110 = N109 & sel_i[3];
  assign N111 = N110 & sel_i[2];
  assign N112 = N111 & N115;
  assign N287 = N112 & N116;
  assign N113 = ~sel_i[5];
  assign N114 = ~sel_i[4];
  assign N115 = ~sel_i[0];
  assign N116 = ~sel_i[1];
  assign N117 = N121 & N122;
  assign N118 = N117 & sel_i[3];
  assign N119 = N118 & sel_i[2];
  assign N120 = N119 & sel_i[0];
  assign N289 = N120 & N123;
  assign N121 = ~sel_i[5];
  assign N122 = ~sel_i[4];
  assign N123 = ~sel_i[1];
  assign N124 = N128 & N129;
  assign N125 = N124 & sel_i[3];
  assign N126 = N125 & sel_i[2];
  assign N127 = N126 & N130;
  assign N291 = N127 & sel_i[1];
  assign N128 = ~sel_i[5];
  assign N129 = ~sel_i[4];
  assign N130 = ~sel_i[0];
  assign N131 = N135 & N136;
  assign N132 = N131 & sel_i[3];
  assign N133 = N132 & sel_i[2];
  assign N134 = N133 & sel_i[0];
  assign N293 = N134 & sel_i[1];
  assign N135 = ~sel_i[5];
  assign N136 = ~sel_i[4];
  assign N137 = N141 & sel_i[4];
  assign N138 = N137 & N142;
  assign N139 = N138 & N143;
  assign N140 = N139 & N144;
  assign N295 = N140 & N145;
  assign N141 = ~sel_i[5];
  assign N142 = ~sel_i[3];
  assign N143 = ~sel_i[2];
  assign N144 = ~sel_i[0];
  assign N145 = ~sel_i[1];
  assign N146 = N150 & sel_i[4];
  assign N147 = N146 & N151;
  assign N148 = N147 & N152;
  assign N149 = N148 & sel_i[0];
  assign N297 = N149 & N153;
  assign N150 = ~sel_i[5];
  assign N151 = ~sel_i[3];
  assign N152 = ~sel_i[2];
  assign N153 = ~sel_i[1];
  assign N299 = sel_i[4] & N154 & (N155 & N156) & sel_i[1];
  assign N154 = ~sel_i[3];
  assign N155 = ~sel_i[2];
  assign N156 = ~sel_i[0];
  assign N300 = sel_i[4] & N157 & (N158 & sel_i[0]) & sel_i[1];
  assign N157 = ~sel_i[3];
  assign N158 = ~sel_i[2];
  assign N301 = sel_i[4] & N159 & (sel_i[2] & N160) & N161;
  assign N159 = ~sel_i[3];
  assign N160 = ~sel_i[0];
  assign N161 = ~sel_i[1];
  assign N302 = sel_i[4] & N162 & (sel_i[2] & sel_i[0]) & N163;
  assign N162 = ~sel_i[3];
  assign N163 = ~sel_i[1];
  assign N303 = sel_i[4] & N164 & (sel_i[2] & N165) & sel_i[1];
  assign N164 = ~sel_i[3];
  assign N165 = ~sel_i[0];
  assign N304 = sel_i[4] & N166 & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N166 = ~sel_i[3];
  assign N305 = sel_i[4] & sel_i[3] & (N167 & N168) & N169;
  assign N167 = ~sel_i[2];
  assign N168 = ~sel_i[0];
  assign N169 = ~sel_i[1];
  assign N306 = sel_i[4] & sel_i[3] & (N170 & sel_i[0]) & N171;
  assign N170 = ~sel_i[2];
  assign N171 = ~sel_i[1];
  assign N307 = sel_i[4] & sel_i[3] & (N172 & N173) & sel_i[1];
  assign N172 = ~sel_i[2];
  assign N173 = ~sel_i[0];
  assign N308 = sel_i[4] & sel_i[3] & (N174 & sel_i[0]) & sel_i[1];
  assign N174 = ~sel_i[2];
  assign N309 = sel_i[4] & sel_i[3] & (sel_i[2] & N175) & N176;
  assign N175 = ~sel_i[0];
  assign N176 = ~sel_i[1];
  assign N310 = sel_i[4] & sel_i[3] & (sel_i[2] & sel_i[0]) & N177;
  assign N177 = ~sel_i[1];
  assign N311 = sel_i[4] & sel_i[3] & (sel_i[2] & N178) & sel_i[1];
  assign N178 = ~sel_i[0];
  assign N312 = sel_i[4] & sel_i[3] & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N179 = sel_i[5] & N183;
  assign N180 = N179 & N184;
  assign N181 = N180 & N185;
  assign N182 = N181 & sel_i[0];
  assign N266 = N182 & N186;
  assign N183 = ~sel_i[4];
  assign N184 = ~sel_i[3];
  assign N185 = ~sel_i[2];
  assign N186 = ~sel_i[1];
  assign N268 = sel_i[5] & N187 & (N188 & N189) & sel_i[1];
  assign N187 = ~sel_i[3];
  assign N188 = ~sel_i[2];
  assign N189 = ~sel_i[0];
  assign N270 = sel_i[5] & N190 & (N191 & sel_i[0]) & sel_i[1];
  assign N190 = ~sel_i[3];
  assign N191 = ~sel_i[2];
  assign N272 = sel_i[5] & N192 & (sel_i[2] & N193) & N194;
  assign N192 = ~sel_i[3];
  assign N193 = ~sel_i[0];
  assign N194 = ~sel_i[1];
  assign N274 = sel_i[5] & N195 & (sel_i[2] & sel_i[0]) & N196;
  assign N195 = ~sel_i[3];
  assign N196 = ~sel_i[1];
  assign N276 = sel_i[5] & N197 & (sel_i[2] & N198) & sel_i[1];
  assign N197 = ~sel_i[3];
  assign N198 = ~sel_i[0];
  assign N278 = sel_i[5] & N199 & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N199 = ~sel_i[3];
  assign N280 = sel_i[5] & sel_i[3] & (N200 & N201) & N202;
  assign N200 = ~sel_i[2];
  assign N201 = ~sel_i[0];
  assign N202 = ~sel_i[1];
  assign N282 = sel_i[5] & sel_i[3] & (N203 & sel_i[0]) & N204;
  assign N203 = ~sel_i[2];
  assign N204 = ~sel_i[1];
  assign N284 = sel_i[5] & sel_i[3] & (N205 & N206) & sel_i[1];
  assign N205 = ~sel_i[2];
  assign N206 = ~sel_i[0];
  assign N286 = sel_i[5] & sel_i[3] & (N207 & sel_i[0]) & sel_i[1];
  assign N207 = ~sel_i[2];
  assign N288 = sel_i[5] & sel_i[3] & (sel_i[2] & N208) & N209;
  assign N208 = ~sel_i[0];
  assign N209 = ~sel_i[1];
  assign N290 = sel_i[5] & sel_i[3] & (sel_i[2] & sel_i[0]) & N210;
  assign N210 = ~sel_i[1];
  assign N292 = sel_i[5] & sel_i[3] & (sel_i[2] & N211) & sel_i[1];
  assign N211 = ~sel_i[0];
  assign N294 = sel_i[5] & sel_i[3] & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N296 = sel_i[5] & sel_i[4] & N212;
  assign N212 = ~sel_i[0];
  assign N298 = sel_i[5] & sel_i[4] & sel_i[0];
  assign data_o[31] = (N213)? data_i[31] : 
                      (N214)? data_i[63] : 
                      (N215)? data_i[95] : 
                      (N216)? data_i[127] : 
                      (N217)? data_i[159] : 
                      (N218)? data_i[191] : 
                      (N219)? data_i[223] : 
                      (N220)? data_i[255] : 
                      (N221)? data_i[287] : 
                      (N222)? data_i[319] : 
                      (N223)? data_i[351] : 
                      (N224)? data_i[383] : 
                      (N225)? data_i[415] : 
                      (N226)? data_i[447] : 
                      (N227)? data_i[479] : 
                      (N228)? data_i[511] : 
                      (N229)? data_i[543] : 
                      (N230)? data_i[575] : 
                      (N231)? data_i[607] : 
                      (N232)? data_i[639] : 
                      (N233)? data_i[671] : 
                      (N234)? data_i[703] : 
                      (N235)? data_i[735] : 
                      (N236)? data_i[767] : 
                      (N237)? data_i[799] : 
                      (N238)? data_i[831] : 
                      (N239)? data_i[863] : 
                      (N240)? data_i[895] : 
                      (N241)? data_i[927] : 
                      (N242)? data_i[959] : 
                      (N243)? data_i[991] : 
                      (N244)? data_i[1023] : 
                      (N245)? data_i[1055] : 
                      (N246)? data_i[1087] : 
                      (N247)? data_i[1119] : 
                      (N248)? data_i[1151] : 
                      (N249)? data_i[1183] : 
                      (N250)? data_i[1215] : 
                      (N251)? data_i[1247] : 
                      (N252)? data_i[1279] : 
                      (N253)? data_i[1311] : 
                      (N254)? data_i[1343] : 
                      (N255)? data_i[1375] : 
                      (N256)? data_i[1407] : 
                      (N257)? data_i[1439] : 
                      (N258)? data_i[1471] : 
                      (N259)? data_i[1503] : 
                      (N260)? data_i[1535] : 
                      (N261)? data_i[1567] : 
                      (N262)? data_i[1599] : 1'b0;
  assign N213 = N263;
  assign N214 = N265;
  assign N215 = N267;
  assign N216 = N269;
  assign N217 = N271;
  assign N218 = N273;
  assign N219 = N275;
  assign N220 = N277;
  assign N221 = N279;
  assign N222 = N281;
  assign N223 = N283;
  assign N224 = N285;
  assign N225 = N287;
  assign N226 = N289;
  assign N227 = N291;
  assign N228 = N293;
  assign N229 = N295;
  assign N230 = N297;
  assign N231 = N299;
  assign N232 = N300;
  assign N233 = N301;
  assign N234 = N302;
  assign N235 = N303;
  assign N236 = N304;
  assign N237 = N305;
  assign N238 = N306;
  assign N239 = N307;
  assign N240 = N308;
  assign N241 = N309;
  assign N242 = N310;
  assign N243 = N311;
  assign N244 = N312;
  assign N245 = N264;
  assign N246 = N266;
  assign N247 = N268;
  assign N248 = N270;
  assign N249 = N272;
  assign N250 = N274;
  assign N251 = N276;
  assign N252 = N278;
  assign N253 = N280;
  assign N254 = N282;
  assign N255 = N284;
  assign N256 = N286;
  assign N257 = N288;
  assign N258 = N290;
  assign N259 = N292;
  assign N260 = N294;
  assign N261 = N296;
  assign N262 = N298;
  assign data_o[30] = (N213)? data_i[30] : 
                      (N214)? data_i[62] : 
                      (N215)? data_i[94] : 
                      (N216)? data_i[126] : 
                      (N217)? data_i[158] : 
                      (N218)? data_i[190] : 
                      (N219)? data_i[222] : 
                      (N220)? data_i[254] : 
                      (N221)? data_i[286] : 
                      (N222)? data_i[318] : 
                      (N223)? data_i[350] : 
                      (N224)? data_i[382] : 
                      (N225)? data_i[414] : 
                      (N226)? data_i[446] : 
                      (N227)? data_i[478] : 
                      (N228)? data_i[510] : 
                      (N229)? data_i[542] : 
                      (N230)? data_i[574] : 
                      (N231)? data_i[606] : 
                      (N232)? data_i[638] : 
                      (N233)? data_i[670] : 
                      (N234)? data_i[702] : 
                      (N235)? data_i[734] : 
                      (N236)? data_i[766] : 
                      (N237)? data_i[798] : 
                      (N238)? data_i[830] : 
                      (N239)? data_i[862] : 
                      (N240)? data_i[894] : 
                      (N241)? data_i[926] : 
                      (N242)? data_i[958] : 
                      (N243)? data_i[990] : 
                      (N244)? data_i[1022] : 
                      (N245)? data_i[1054] : 
                      (N246)? data_i[1086] : 
                      (N247)? data_i[1118] : 
                      (N248)? data_i[1150] : 
                      (N249)? data_i[1182] : 
                      (N250)? data_i[1214] : 
                      (N251)? data_i[1246] : 
                      (N252)? data_i[1278] : 
                      (N253)? data_i[1310] : 
                      (N254)? data_i[1342] : 
                      (N255)? data_i[1374] : 
                      (N256)? data_i[1406] : 
                      (N257)? data_i[1438] : 
                      (N258)? data_i[1470] : 
                      (N259)? data_i[1502] : 
                      (N260)? data_i[1534] : 
                      (N261)? data_i[1566] : 
                      (N262)? data_i[1598] : 1'b0;
  assign data_o[29] = (N213)? data_i[29] : 
                      (N214)? data_i[61] : 
                      (N215)? data_i[93] : 
                      (N216)? data_i[125] : 
                      (N217)? data_i[157] : 
                      (N218)? data_i[189] : 
                      (N219)? data_i[221] : 
                      (N220)? data_i[253] : 
                      (N221)? data_i[285] : 
                      (N222)? data_i[317] : 
                      (N223)? data_i[349] : 
                      (N224)? data_i[381] : 
                      (N225)? data_i[413] : 
                      (N226)? data_i[445] : 
                      (N227)? data_i[477] : 
                      (N228)? data_i[509] : 
                      (N229)? data_i[541] : 
                      (N230)? data_i[573] : 
                      (N231)? data_i[605] : 
                      (N232)? data_i[637] : 
                      (N233)? data_i[669] : 
                      (N234)? data_i[701] : 
                      (N235)? data_i[733] : 
                      (N236)? data_i[765] : 
                      (N237)? data_i[797] : 
                      (N238)? data_i[829] : 
                      (N239)? data_i[861] : 
                      (N240)? data_i[893] : 
                      (N241)? data_i[925] : 
                      (N242)? data_i[957] : 
                      (N243)? data_i[989] : 
                      (N244)? data_i[1021] : 
                      (N245)? data_i[1053] : 
                      (N246)? data_i[1085] : 
                      (N247)? data_i[1117] : 
                      (N248)? data_i[1149] : 
                      (N249)? data_i[1181] : 
                      (N250)? data_i[1213] : 
                      (N251)? data_i[1245] : 
                      (N252)? data_i[1277] : 
                      (N253)? data_i[1309] : 
                      (N254)? data_i[1341] : 
                      (N255)? data_i[1373] : 
                      (N256)? data_i[1405] : 
                      (N257)? data_i[1437] : 
                      (N258)? data_i[1469] : 
                      (N259)? data_i[1501] : 
                      (N260)? data_i[1533] : 
                      (N261)? data_i[1565] : 
                      (N262)? data_i[1597] : 1'b0;
  assign data_o[28] = (N213)? data_i[28] : 
                      (N214)? data_i[60] : 
                      (N215)? data_i[92] : 
                      (N216)? data_i[124] : 
                      (N217)? data_i[156] : 
                      (N218)? data_i[188] : 
                      (N219)? data_i[220] : 
                      (N220)? data_i[252] : 
                      (N221)? data_i[284] : 
                      (N222)? data_i[316] : 
                      (N223)? data_i[348] : 
                      (N224)? data_i[380] : 
                      (N225)? data_i[412] : 
                      (N226)? data_i[444] : 
                      (N227)? data_i[476] : 
                      (N228)? data_i[508] : 
                      (N229)? data_i[540] : 
                      (N230)? data_i[572] : 
                      (N231)? data_i[604] : 
                      (N232)? data_i[636] : 
                      (N233)? data_i[668] : 
                      (N234)? data_i[700] : 
                      (N235)? data_i[732] : 
                      (N236)? data_i[764] : 
                      (N237)? data_i[796] : 
                      (N238)? data_i[828] : 
                      (N239)? data_i[860] : 
                      (N240)? data_i[892] : 
                      (N241)? data_i[924] : 
                      (N242)? data_i[956] : 
                      (N243)? data_i[988] : 
                      (N244)? data_i[1020] : 
                      (N245)? data_i[1052] : 
                      (N246)? data_i[1084] : 
                      (N247)? data_i[1116] : 
                      (N248)? data_i[1148] : 
                      (N249)? data_i[1180] : 
                      (N250)? data_i[1212] : 
                      (N251)? data_i[1244] : 
                      (N252)? data_i[1276] : 
                      (N253)? data_i[1308] : 
                      (N254)? data_i[1340] : 
                      (N255)? data_i[1372] : 
                      (N256)? data_i[1404] : 
                      (N257)? data_i[1436] : 
                      (N258)? data_i[1468] : 
                      (N259)? data_i[1500] : 
                      (N260)? data_i[1532] : 
                      (N261)? data_i[1564] : 
                      (N262)? data_i[1596] : 1'b0;
  assign data_o[27] = (N213)? data_i[27] : 
                      (N214)? data_i[59] : 
                      (N215)? data_i[91] : 
                      (N216)? data_i[123] : 
                      (N217)? data_i[155] : 
                      (N218)? data_i[187] : 
                      (N219)? data_i[219] : 
                      (N220)? data_i[251] : 
                      (N221)? data_i[283] : 
                      (N222)? data_i[315] : 
                      (N223)? data_i[347] : 
                      (N224)? data_i[379] : 
                      (N225)? data_i[411] : 
                      (N226)? data_i[443] : 
                      (N227)? data_i[475] : 
                      (N228)? data_i[507] : 
                      (N229)? data_i[539] : 
                      (N230)? data_i[571] : 
                      (N231)? data_i[603] : 
                      (N232)? data_i[635] : 
                      (N233)? data_i[667] : 
                      (N234)? data_i[699] : 
                      (N235)? data_i[731] : 
                      (N236)? data_i[763] : 
                      (N237)? data_i[795] : 
                      (N238)? data_i[827] : 
                      (N239)? data_i[859] : 
                      (N240)? data_i[891] : 
                      (N241)? data_i[923] : 
                      (N242)? data_i[955] : 
                      (N243)? data_i[987] : 
                      (N244)? data_i[1019] : 
                      (N245)? data_i[1051] : 
                      (N246)? data_i[1083] : 
                      (N247)? data_i[1115] : 
                      (N248)? data_i[1147] : 
                      (N249)? data_i[1179] : 
                      (N250)? data_i[1211] : 
                      (N251)? data_i[1243] : 
                      (N252)? data_i[1275] : 
                      (N253)? data_i[1307] : 
                      (N254)? data_i[1339] : 
                      (N255)? data_i[1371] : 
                      (N256)? data_i[1403] : 
                      (N257)? data_i[1435] : 
                      (N258)? data_i[1467] : 
                      (N259)? data_i[1499] : 
                      (N260)? data_i[1531] : 
                      (N261)? data_i[1563] : 
                      (N262)? data_i[1595] : 1'b0;
  assign data_o[26] = (N213)? data_i[26] : 
                      (N214)? data_i[58] : 
                      (N215)? data_i[90] : 
                      (N216)? data_i[122] : 
                      (N217)? data_i[154] : 
                      (N218)? data_i[186] : 
                      (N219)? data_i[218] : 
                      (N220)? data_i[250] : 
                      (N221)? data_i[282] : 
                      (N222)? data_i[314] : 
                      (N223)? data_i[346] : 
                      (N224)? data_i[378] : 
                      (N225)? data_i[410] : 
                      (N226)? data_i[442] : 
                      (N227)? data_i[474] : 
                      (N228)? data_i[506] : 
                      (N229)? data_i[538] : 
                      (N230)? data_i[570] : 
                      (N231)? data_i[602] : 
                      (N232)? data_i[634] : 
                      (N233)? data_i[666] : 
                      (N234)? data_i[698] : 
                      (N235)? data_i[730] : 
                      (N236)? data_i[762] : 
                      (N237)? data_i[794] : 
                      (N238)? data_i[826] : 
                      (N239)? data_i[858] : 
                      (N240)? data_i[890] : 
                      (N241)? data_i[922] : 
                      (N242)? data_i[954] : 
                      (N243)? data_i[986] : 
                      (N244)? data_i[1018] : 
                      (N245)? data_i[1050] : 
                      (N246)? data_i[1082] : 
                      (N247)? data_i[1114] : 
                      (N248)? data_i[1146] : 
                      (N249)? data_i[1178] : 
                      (N250)? data_i[1210] : 
                      (N251)? data_i[1242] : 
                      (N252)? data_i[1274] : 
                      (N253)? data_i[1306] : 
                      (N254)? data_i[1338] : 
                      (N255)? data_i[1370] : 
                      (N256)? data_i[1402] : 
                      (N257)? data_i[1434] : 
                      (N258)? data_i[1466] : 
                      (N259)? data_i[1498] : 
                      (N260)? data_i[1530] : 
                      (N261)? data_i[1562] : 
                      (N262)? data_i[1594] : 1'b0;
  assign data_o[25] = (N213)? data_i[25] : 
                      (N214)? data_i[57] : 
                      (N215)? data_i[89] : 
                      (N216)? data_i[121] : 
                      (N217)? data_i[153] : 
                      (N218)? data_i[185] : 
                      (N219)? data_i[217] : 
                      (N220)? data_i[249] : 
                      (N221)? data_i[281] : 
                      (N222)? data_i[313] : 
                      (N223)? data_i[345] : 
                      (N224)? data_i[377] : 
                      (N225)? data_i[409] : 
                      (N226)? data_i[441] : 
                      (N227)? data_i[473] : 
                      (N228)? data_i[505] : 
                      (N229)? data_i[537] : 
                      (N230)? data_i[569] : 
                      (N231)? data_i[601] : 
                      (N232)? data_i[633] : 
                      (N233)? data_i[665] : 
                      (N234)? data_i[697] : 
                      (N235)? data_i[729] : 
                      (N236)? data_i[761] : 
                      (N237)? data_i[793] : 
                      (N238)? data_i[825] : 
                      (N239)? data_i[857] : 
                      (N240)? data_i[889] : 
                      (N241)? data_i[921] : 
                      (N242)? data_i[953] : 
                      (N243)? data_i[985] : 
                      (N244)? data_i[1017] : 
                      (N245)? data_i[1049] : 
                      (N246)? data_i[1081] : 
                      (N247)? data_i[1113] : 
                      (N248)? data_i[1145] : 
                      (N249)? data_i[1177] : 
                      (N250)? data_i[1209] : 
                      (N251)? data_i[1241] : 
                      (N252)? data_i[1273] : 
                      (N253)? data_i[1305] : 
                      (N254)? data_i[1337] : 
                      (N255)? data_i[1369] : 
                      (N256)? data_i[1401] : 
                      (N257)? data_i[1433] : 
                      (N258)? data_i[1465] : 
                      (N259)? data_i[1497] : 
                      (N260)? data_i[1529] : 
                      (N261)? data_i[1561] : 
                      (N262)? data_i[1593] : 1'b0;
  assign data_o[24] = (N213)? data_i[24] : 
                      (N214)? data_i[56] : 
                      (N215)? data_i[88] : 
                      (N216)? data_i[120] : 
                      (N217)? data_i[152] : 
                      (N218)? data_i[184] : 
                      (N219)? data_i[216] : 
                      (N220)? data_i[248] : 
                      (N221)? data_i[280] : 
                      (N222)? data_i[312] : 
                      (N223)? data_i[344] : 
                      (N224)? data_i[376] : 
                      (N225)? data_i[408] : 
                      (N226)? data_i[440] : 
                      (N227)? data_i[472] : 
                      (N228)? data_i[504] : 
                      (N229)? data_i[536] : 
                      (N230)? data_i[568] : 
                      (N231)? data_i[600] : 
                      (N232)? data_i[632] : 
                      (N233)? data_i[664] : 
                      (N234)? data_i[696] : 
                      (N235)? data_i[728] : 
                      (N236)? data_i[760] : 
                      (N237)? data_i[792] : 
                      (N238)? data_i[824] : 
                      (N239)? data_i[856] : 
                      (N240)? data_i[888] : 
                      (N241)? data_i[920] : 
                      (N242)? data_i[952] : 
                      (N243)? data_i[984] : 
                      (N244)? data_i[1016] : 
                      (N245)? data_i[1048] : 
                      (N246)? data_i[1080] : 
                      (N247)? data_i[1112] : 
                      (N248)? data_i[1144] : 
                      (N249)? data_i[1176] : 
                      (N250)? data_i[1208] : 
                      (N251)? data_i[1240] : 
                      (N252)? data_i[1272] : 
                      (N253)? data_i[1304] : 
                      (N254)? data_i[1336] : 
                      (N255)? data_i[1368] : 
                      (N256)? data_i[1400] : 
                      (N257)? data_i[1432] : 
                      (N258)? data_i[1464] : 
                      (N259)? data_i[1496] : 
                      (N260)? data_i[1528] : 
                      (N261)? data_i[1560] : 
                      (N262)? data_i[1592] : 1'b0;
  assign data_o[23] = (N213)? data_i[23] : 
                      (N214)? data_i[55] : 
                      (N215)? data_i[87] : 
                      (N216)? data_i[119] : 
                      (N217)? data_i[151] : 
                      (N218)? data_i[183] : 
                      (N219)? data_i[215] : 
                      (N220)? data_i[247] : 
                      (N221)? data_i[279] : 
                      (N222)? data_i[311] : 
                      (N223)? data_i[343] : 
                      (N224)? data_i[375] : 
                      (N225)? data_i[407] : 
                      (N226)? data_i[439] : 
                      (N227)? data_i[471] : 
                      (N228)? data_i[503] : 
                      (N229)? data_i[535] : 
                      (N230)? data_i[567] : 
                      (N231)? data_i[599] : 
                      (N232)? data_i[631] : 
                      (N233)? data_i[663] : 
                      (N234)? data_i[695] : 
                      (N235)? data_i[727] : 
                      (N236)? data_i[759] : 
                      (N237)? data_i[791] : 
                      (N238)? data_i[823] : 
                      (N239)? data_i[855] : 
                      (N240)? data_i[887] : 
                      (N241)? data_i[919] : 
                      (N242)? data_i[951] : 
                      (N243)? data_i[983] : 
                      (N244)? data_i[1015] : 
                      (N245)? data_i[1047] : 
                      (N246)? data_i[1079] : 
                      (N247)? data_i[1111] : 
                      (N248)? data_i[1143] : 
                      (N249)? data_i[1175] : 
                      (N250)? data_i[1207] : 
                      (N251)? data_i[1239] : 
                      (N252)? data_i[1271] : 
                      (N253)? data_i[1303] : 
                      (N254)? data_i[1335] : 
                      (N255)? data_i[1367] : 
                      (N256)? data_i[1399] : 
                      (N257)? data_i[1431] : 
                      (N258)? data_i[1463] : 
                      (N259)? data_i[1495] : 
                      (N260)? data_i[1527] : 
                      (N261)? data_i[1559] : 
                      (N262)? data_i[1591] : 1'b0;
  assign data_o[22] = (N213)? data_i[22] : 
                      (N214)? data_i[54] : 
                      (N215)? data_i[86] : 
                      (N216)? data_i[118] : 
                      (N217)? data_i[150] : 
                      (N218)? data_i[182] : 
                      (N219)? data_i[214] : 
                      (N220)? data_i[246] : 
                      (N221)? data_i[278] : 
                      (N222)? data_i[310] : 
                      (N223)? data_i[342] : 
                      (N224)? data_i[374] : 
                      (N225)? data_i[406] : 
                      (N226)? data_i[438] : 
                      (N227)? data_i[470] : 
                      (N228)? data_i[502] : 
                      (N229)? data_i[534] : 
                      (N230)? data_i[566] : 
                      (N231)? data_i[598] : 
                      (N232)? data_i[630] : 
                      (N233)? data_i[662] : 
                      (N234)? data_i[694] : 
                      (N235)? data_i[726] : 
                      (N236)? data_i[758] : 
                      (N237)? data_i[790] : 
                      (N238)? data_i[822] : 
                      (N239)? data_i[854] : 
                      (N240)? data_i[886] : 
                      (N241)? data_i[918] : 
                      (N242)? data_i[950] : 
                      (N243)? data_i[982] : 
                      (N244)? data_i[1014] : 
                      (N245)? data_i[1046] : 
                      (N246)? data_i[1078] : 
                      (N247)? data_i[1110] : 
                      (N248)? data_i[1142] : 
                      (N249)? data_i[1174] : 
                      (N250)? data_i[1206] : 
                      (N251)? data_i[1238] : 
                      (N252)? data_i[1270] : 
                      (N253)? data_i[1302] : 
                      (N254)? data_i[1334] : 
                      (N255)? data_i[1366] : 
                      (N256)? data_i[1398] : 
                      (N257)? data_i[1430] : 
                      (N258)? data_i[1462] : 
                      (N259)? data_i[1494] : 
                      (N260)? data_i[1526] : 
                      (N261)? data_i[1558] : 
                      (N262)? data_i[1590] : 1'b0;
  assign data_o[21] = (N213)? data_i[21] : 
                      (N214)? data_i[53] : 
                      (N215)? data_i[85] : 
                      (N216)? data_i[117] : 
                      (N217)? data_i[149] : 
                      (N218)? data_i[181] : 
                      (N219)? data_i[213] : 
                      (N220)? data_i[245] : 
                      (N221)? data_i[277] : 
                      (N222)? data_i[309] : 
                      (N223)? data_i[341] : 
                      (N224)? data_i[373] : 
                      (N225)? data_i[405] : 
                      (N226)? data_i[437] : 
                      (N227)? data_i[469] : 
                      (N228)? data_i[501] : 
                      (N229)? data_i[533] : 
                      (N230)? data_i[565] : 
                      (N231)? data_i[597] : 
                      (N232)? data_i[629] : 
                      (N233)? data_i[661] : 
                      (N234)? data_i[693] : 
                      (N235)? data_i[725] : 
                      (N236)? data_i[757] : 
                      (N237)? data_i[789] : 
                      (N238)? data_i[821] : 
                      (N239)? data_i[853] : 
                      (N240)? data_i[885] : 
                      (N241)? data_i[917] : 
                      (N242)? data_i[949] : 
                      (N243)? data_i[981] : 
                      (N244)? data_i[1013] : 
                      (N245)? data_i[1045] : 
                      (N246)? data_i[1077] : 
                      (N247)? data_i[1109] : 
                      (N248)? data_i[1141] : 
                      (N249)? data_i[1173] : 
                      (N250)? data_i[1205] : 
                      (N251)? data_i[1237] : 
                      (N252)? data_i[1269] : 
                      (N253)? data_i[1301] : 
                      (N254)? data_i[1333] : 
                      (N255)? data_i[1365] : 
                      (N256)? data_i[1397] : 
                      (N257)? data_i[1429] : 
                      (N258)? data_i[1461] : 
                      (N259)? data_i[1493] : 
                      (N260)? data_i[1525] : 
                      (N261)? data_i[1557] : 
                      (N262)? data_i[1589] : 1'b0;
  assign data_o[20] = (N213)? data_i[20] : 
                      (N214)? data_i[52] : 
                      (N215)? data_i[84] : 
                      (N216)? data_i[116] : 
                      (N217)? data_i[148] : 
                      (N218)? data_i[180] : 
                      (N219)? data_i[212] : 
                      (N220)? data_i[244] : 
                      (N221)? data_i[276] : 
                      (N222)? data_i[308] : 
                      (N223)? data_i[340] : 
                      (N224)? data_i[372] : 
                      (N225)? data_i[404] : 
                      (N226)? data_i[436] : 
                      (N227)? data_i[468] : 
                      (N228)? data_i[500] : 
                      (N229)? data_i[532] : 
                      (N230)? data_i[564] : 
                      (N231)? data_i[596] : 
                      (N232)? data_i[628] : 
                      (N233)? data_i[660] : 
                      (N234)? data_i[692] : 
                      (N235)? data_i[724] : 
                      (N236)? data_i[756] : 
                      (N237)? data_i[788] : 
                      (N238)? data_i[820] : 
                      (N239)? data_i[852] : 
                      (N240)? data_i[884] : 
                      (N241)? data_i[916] : 
                      (N242)? data_i[948] : 
                      (N243)? data_i[980] : 
                      (N244)? data_i[1012] : 
                      (N245)? data_i[1044] : 
                      (N246)? data_i[1076] : 
                      (N247)? data_i[1108] : 
                      (N248)? data_i[1140] : 
                      (N249)? data_i[1172] : 
                      (N250)? data_i[1204] : 
                      (N251)? data_i[1236] : 
                      (N252)? data_i[1268] : 
                      (N253)? data_i[1300] : 
                      (N254)? data_i[1332] : 
                      (N255)? data_i[1364] : 
                      (N256)? data_i[1396] : 
                      (N257)? data_i[1428] : 
                      (N258)? data_i[1460] : 
                      (N259)? data_i[1492] : 
                      (N260)? data_i[1524] : 
                      (N261)? data_i[1556] : 
                      (N262)? data_i[1588] : 1'b0;
  assign data_o[19] = (N213)? data_i[19] : 
                      (N214)? data_i[51] : 
                      (N215)? data_i[83] : 
                      (N216)? data_i[115] : 
                      (N217)? data_i[147] : 
                      (N218)? data_i[179] : 
                      (N219)? data_i[211] : 
                      (N220)? data_i[243] : 
                      (N221)? data_i[275] : 
                      (N222)? data_i[307] : 
                      (N223)? data_i[339] : 
                      (N224)? data_i[371] : 
                      (N225)? data_i[403] : 
                      (N226)? data_i[435] : 
                      (N227)? data_i[467] : 
                      (N228)? data_i[499] : 
                      (N229)? data_i[531] : 
                      (N230)? data_i[563] : 
                      (N231)? data_i[595] : 
                      (N232)? data_i[627] : 
                      (N233)? data_i[659] : 
                      (N234)? data_i[691] : 
                      (N235)? data_i[723] : 
                      (N236)? data_i[755] : 
                      (N237)? data_i[787] : 
                      (N238)? data_i[819] : 
                      (N239)? data_i[851] : 
                      (N240)? data_i[883] : 
                      (N241)? data_i[915] : 
                      (N242)? data_i[947] : 
                      (N243)? data_i[979] : 
                      (N244)? data_i[1011] : 
                      (N245)? data_i[1043] : 
                      (N246)? data_i[1075] : 
                      (N247)? data_i[1107] : 
                      (N248)? data_i[1139] : 
                      (N249)? data_i[1171] : 
                      (N250)? data_i[1203] : 
                      (N251)? data_i[1235] : 
                      (N252)? data_i[1267] : 
                      (N253)? data_i[1299] : 
                      (N254)? data_i[1331] : 
                      (N255)? data_i[1363] : 
                      (N256)? data_i[1395] : 
                      (N257)? data_i[1427] : 
                      (N258)? data_i[1459] : 
                      (N259)? data_i[1491] : 
                      (N260)? data_i[1523] : 
                      (N261)? data_i[1555] : 
                      (N262)? data_i[1587] : 1'b0;
  assign data_o[18] = (N213)? data_i[18] : 
                      (N214)? data_i[50] : 
                      (N215)? data_i[82] : 
                      (N216)? data_i[114] : 
                      (N217)? data_i[146] : 
                      (N218)? data_i[178] : 
                      (N219)? data_i[210] : 
                      (N220)? data_i[242] : 
                      (N221)? data_i[274] : 
                      (N222)? data_i[306] : 
                      (N223)? data_i[338] : 
                      (N224)? data_i[370] : 
                      (N225)? data_i[402] : 
                      (N226)? data_i[434] : 
                      (N227)? data_i[466] : 
                      (N228)? data_i[498] : 
                      (N229)? data_i[530] : 
                      (N230)? data_i[562] : 
                      (N231)? data_i[594] : 
                      (N232)? data_i[626] : 
                      (N233)? data_i[658] : 
                      (N234)? data_i[690] : 
                      (N235)? data_i[722] : 
                      (N236)? data_i[754] : 
                      (N237)? data_i[786] : 
                      (N238)? data_i[818] : 
                      (N239)? data_i[850] : 
                      (N240)? data_i[882] : 
                      (N241)? data_i[914] : 
                      (N242)? data_i[946] : 
                      (N243)? data_i[978] : 
                      (N244)? data_i[1010] : 
                      (N245)? data_i[1042] : 
                      (N246)? data_i[1074] : 
                      (N247)? data_i[1106] : 
                      (N248)? data_i[1138] : 
                      (N249)? data_i[1170] : 
                      (N250)? data_i[1202] : 
                      (N251)? data_i[1234] : 
                      (N252)? data_i[1266] : 
                      (N253)? data_i[1298] : 
                      (N254)? data_i[1330] : 
                      (N255)? data_i[1362] : 
                      (N256)? data_i[1394] : 
                      (N257)? data_i[1426] : 
                      (N258)? data_i[1458] : 
                      (N259)? data_i[1490] : 
                      (N260)? data_i[1522] : 
                      (N261)? data_i[1554] : 
                      (N262)? data_i[1586] : 1'b0;
  assign data_o[17] = (N213)? data_i[17] : 
                      (N214)? data_i[49] : 
                      (N215)? data_i[81] : 
                      (N216)? data_i[113] : 
                      (N217)? data_i[145] : 
                      (N218)? data_i[177] : 
                      (N219)? data_i[209] : 
                      (N220)? data_i[241] : 
                      (N221)? data_i[273] : 
                      (N222)? data_i[305] : 
                      (N223)? data_i[337] : 
                      (N224)? data_i[369] : 
                      (N225)? data_i[401] : 
                      (N226)? data_i[433] : 
                      (N227)? data_i[465] : 
                      (N228)? data_i[497] : 
                      (N229)? data_i[529] : 
                      (N230)? data_i[561] : 
                      (N231)? data_i[593] : 
                      (N232)? data_i[625] : 
                      (N233)? data_i[657] : 
                      (N234)? data_i[689] : 
                      (N235)? data_i[721] : 
                      (N236)? data_i[753] : 
                      (N237)? data_i[785] : 
                      (N238)? data_i[817] : 
                      (N239)? data_i[849] : 
                      (N240)? data_i[881] : 
                      (N241)? data_i[913] : 
                      (N242)? data_i[945] : 
                      (N243)? data_i[977] : 
                      (N244)? data_i[1009] : 
                      (N245)? data_i[1041] : 
                      (N246)? data_i[1073] : 
                      (N247)? data_i[1105] : 
                      (N248)? data_i[1137] : 
                      (N249)? data_i[1169] : 
                      (N250)? data_i[1201] : 
                      (N251)? data_i[1233] : 
                      (N252)? data_i[1265] : 
                      (N253)? data_i[1297] : 
                      (N254)? data_i[1329] : 
                      (N255)? data_i[1361] : 
                      (N256)? data_i[1393] : 
                      (N257)? data_i[1425] : 
                      (N258)? data_i[1457] : 
                      (N259)? data_i[1489] : 
                      (N260)? data_i[1521] : 
                      (N261)? data_i[1553] : 
                      (N262)? data_i[1585] : 1'b0;
  assign data_o[16] = (N213)? data_i[16] : 
                      (N214)? data_i[48] : 
                      (N215)? data_i[80] : 
                      (N216)? data_i[112] : 
                      (N217)? data_i[144] : 
                      (N218)? data_i[176] : 
                      (N219)? data_i[208] : 
                      (N220)? data_i[240] : 
                      (N221)? data_i[272] : 
                      (N222)? data_i[304] : 
                      (N223)? data_i[336] : 
                      (N224)? data_i[368] : 
                      (N225)? data_i[400] : 
                      (N226)? data_i[432] : 
                      (N227)? data_i[464] : 
                      (N228)? data_i[496] : 
                      (N229)? data_i[528] : 
                      (N230)? data_i[560] : 
                      (N231)? data_i[592] : 
                      (N232)? data_i[624] : 
                      (N233)? data_i[656] : 
                      (N234)? data_i[688] : 
                      (N235)? data_i[720] : 
                      (N236)? data_i[752] : 
                      (N237)? data_i[784] : 
                      (N238)? data_i[816] : 
                      (N239)? data_i[848] : 
                      (N240)? data_i[880] : 
                      (N241)? data_i[912] : 
                      (N242)? data_i[944] : 
                      (N243)? data_i[976] : 
                      (N244)? data_i[1008] : 
                      (N245)? data_i[1040] : 
                      (N246)? data_i[1072] : 
                      (N247)? data_i[1104] : 
                      (N248)? data_i[1136] : 
                      (N249)? data_i[1168] : 
                      (N250)? data_i[1200] : 
                      (N251)? data_i[1232] : 
                      (N252)? data_i[1264] : 
                      (N253)? data_i[1296] : 
                      (N254)? data_i[1328] : 
                      (N255)? data_i[1360] : 
                      (N256)? data_i[1392] : 
                      (N257)? data_i[1424] : 
                      (N258)? data_i[1456] : 
                      (N259)? data_i[1488] : 
                      (N260)? data_i[1520] : 
                      (N261)? data_i[1552] : 
                      (N262)? data_i[1584] : 1'b0;
  assign data_o[15] = (N213)? data_i[15] : 
                      (N214)? data_i[47] : 
                      (N215)? data_i[79] : 
                      (N216)? data_i[111] : 
                      (N217)? data_i[143] : 
                      (N218)? data_i[175] : 
                      (N219)? data_i[207] : 
                      (N220)? data_i[239] : 
                      (N221)? data_i[271] : 
                      (N222)? data_i[303] : 
                      (N223)? data_i[335] : 
                      (N224)? data_i[367] : 
                      (N225)? data_i[399] : 
                      (N226)? data_i[431] : 
                      (N227)? data_i[463] : 
                      (N228)? data_i[495] : 
                      (N229)? data_i[527] : 
                      (N230)? data_i[559] : 
                      (N231)? data_i[591] : 
                      (N232)? data_i[623] : 
                      (N233)? data_i[655] : 
                      (N234)? data_i[687] : 
                      (N235)? data_i[719] : 
                      (N236)? data_i[751] : 
                      (N237)? data_i[783] : 
                      (N238)? data_i[815] : 
                      (N239)? data_i[847] : 
                      (N240)? data_i[879] : 
                      (N241)? data_i[911] : 
                      (N242)? data_i[943] : 
                      (N243)? data_i[975] : 
                      (N244)? data_i[1007] : 
                      (N245)? data_i[1039] : 
                      (N246)? data_i[1071] : 
                      (N247)? data_i[1103] : 
                      (N248)? data_i[1135] : 
                      (N249)? data_i[1167] : 
                      (N250)? data_i[1199] : 
                      (N251)? data_i[1231] : 
                      (N252)? data_i[1263] : 
                      (N253)? data_i[1295] : 
                      (N254)? data_i[1327] : 
                      (N255)? data_i[1359] : 
                      (N256)? data_i[1391] : 
                      (N257)? data_i[1423] : 
                      (N258)? data_i[1455] : 
                      (N259)? data_i[1487] : 
                      (N260)? data_i[1519] : 
                      (N261)? data_i[1551] : 
                      (N262)? data_i[1583] : 1'b0;
  assign data_o[14] = (N213)? data_i[14] : 
                      (N214)? data_i[46] : 
                      (N215)? data_i[78] : 
                      (N216)? data_i[110] : 
                      (N217)? data_i[142] : 
                      (N218)? data_i[174] : 
                      (N219)? data_i[206] : 
                      (N220)? data_i[238] : 
                      (N221)? data_i[270] : 
                      (N222)? data_i[302] : 
                      (N223)? data_i[334] : 
                      (N224)? data_i[366] : 
                      (N225)? data_i[398] : 
                      (N226)? data_i[430] : 
                      (N227)? data_i[462] : 
                      (N228)? data_i[494] : 
                      (N229)? data_i[526] : 
                      (N230)? data_i[558] : 
                      (N231)? data_i[590] : 
                      (N232)? data_i[622] : 
                      (N233)? data_i[654] : 
                      (N234)? data_i[686] : 
                      (N235)? data_i[718] : 
                      (N236)? data_i[750] : 
                      (N237)? data_i[782] : 
                      (N238)? data_i[814] : 
                      (N239)? data_i[846] : 
                      (N240)? data_i[878] : 
                      (N241)? data_i[910] : 
                      (N242)? data_i[942] : 
                      (N243)? data_i[974] : 
                      (N244)? data_i[1006] : 
                      (N245)? data_i[1038] : 
                      (N246)? data_i[1070] : 
                      (N247)? data_i[1102] : 
                      (N248)? data_i[1134] : 
                      (N249)? data_i[1166] : 
                      (N250)? data_i[1198] : 
                      (N251)? data_i[1230] : 
                      (N252)? data_i[1262] : 
                      (N253)? data_i[1294] : 
                      (N254)? data_i[1326] : 
                      (N255)? data_i[1358] : 
                      (N256)? data_i[1390] : 
                      (N257)? data_i[1422] : 
                      (N258)? data_i[1454] : 
                      (N259)? data_i[1486] : 
                      (N260)? data_i[1518] : 
                      (N261)? data_i[1550] : 
                      (N262)? data_i[1582] : 1'b0;
  assign data_o[13] = (N213)? data_i[13] : 
                      (N214)? data_i[45] : 
                      (N215)? data_i[77] : 
                      (N216)? data_i[109] : 
                      (N217)? data_i[141] : 
                      (N218)? data_i[173] : 
                      (N219)? data_i[205] : 
                      (N220)? data_i[237] : 
                      (N221)? data_i[269] : 
                      (N222)? data_i[301] : 
                      (N223)? data_i[333] : 
                      (N224)? data_i[365] : 
                      (N225)? data_i[397] : 
                      (N226)? data_i[429] : 
                      (N227)? data_i[461] : 
                      (N228)? data_i[493] : 
                      (N229)? data_i[525] : 
                      (N230)? data_i[557] : 
                      (N231)? data_i[589] : 
                      (N232)? data_i[621] : 
                      (N233)? data_i[653] : 
                      (N234)? data_i[685] : 
                      (N235)? data_i[717] : 
                      (N236)? data_i[749] : 
                      (N237)? data_i[781] : 
                      (N238)? data_i[813] : 
                      (N239)? data_i[845] : 
                      (N240)? data_i[877] : 
                      (N241)? data_i[909] : 
                      (N242)? data_i[941] : 
                      (N243)? data_i[973] : 
                      (N244)? data_i[1005] : 
                      (N245)? data_i[1037] : 
                      (N246)? data_i[1069] : 
                      (N247)? data_i[1101] : 
                      (N248)? data_i[1133] : 
                      (N249)? data_i[1165] : 
                      (N250)? data_i[1197] : 
                      (N251)? data_i[1229] : 
                      (N252)? data_i[1261] : 
                      (N253)? data_i[1293] : 
                      (N254)? data_i[1325] : 
                      (N255)? data_i[1357] : 
                      (N256)? data_i[1389] : 
                      (N257)? data_i[1421] : 
                      (N258)? data_i[1453] : 
                      (N259)? data_i[1485] : 
                      (N260)? data_i[1517] : 
                      (N261)? data_i[1549] : 
                      (N262)? data_i[1581] : 1'b0;
  assign data_o[12] = (N213)? data_i[12] : 
                      (N214)? data_i[44] : 
                      (N215)? data_i[76] : 
                      (N216)? data_i[108] : 
                      (N217)? data_i[140] : 
                      (N218)? data_i[172] : 
                      (N219)? data_i[204] : 
                      (N220)? data_i[236] : 
                      (N221)? data_i[268] : 
                      (N222)? data_i[300] : 
                      (N223)? data_i[332] : 
                      (N224)? data_i[364] : 
                      (N225)? data_i[396] : 
                      (N226)? data_i[428] : 
                      (N227)? data_i[460] : 
                      (N228)? data_i[492] : 
                      (N229)? data_i[524] : 
                      (N230)? data_i[556] : 
                      (N231)? data_i[588] : 
                      (N232)? data_i[620] : 
                      (N233)? data_i[652] : 
                      (N234)? data_i[684] : 
                      (N235)? data_i[716] : 
                      (N236)? data_i[748] : 
                      (N237)? data_i[780] : 
                      (N238)? data_i[812] : 
                      (N239)? data_i[844] : 
                      (N240)? data_i[876] : 
                      (N241)? data_i[908] : 
                      (N242)? data_i[940] : 
                      (N243)? data_i[972] : 
                      (N244)? data_i[1004] : 
                      (N245)? data_i[1036] : 
                      (N246)? data_i[1068] : 
                      (N247)? data_i[1100] : 
                      (N248)? data_i[1132] : 
                      (N249)? data_i[1164] : 
                      (N250)? data_i[1196] : 
                      (N251)? data_i[1228] : 
                      (N252)? data_i[1260] : 
                      (N253)? data_i[1292] : 
                      (N254)? data_i[1324] : 
                      (N255)? data_i[1356] : 
                      (N256)? data_i[1388] : 
                      (N257)? data_i[1420] : 
                      (N258)? data_i[1452] : 
                      (N259)? data_i[1484] : 
                      (N260)? data_i[1516] : 
                      (N261)? data_i[1548] : 
                      (N262)? data_i[1580] : 1'b0;
  assign data_o[11] = (N213)? data_i[11] : 
                      (N214)? data_i[43] : 
                      (N215)? data_i[75] : 
                      (N216)? data_i[107] : 
                      (N217)? data_i[139] : 
                      (N218)? data_i[171] : 
                      (N219)? data_i[203] : 
                      (N220)? data_i[235] : 
                      (N221)? data_i[267] : 
                      (N222)? data_i[299] : 
                      (N223)? data_i[331] : 
                      (N224)? data_i[363] : 
                      (N225)? data_i[395] : 
                      (N226)? data_i[427] : 
                      (N227)? data_i[459] : 
                      (N228)? data_i[491] : 
                      (N229)? data_i[523] : 
                      (N230)? data_i[555] : 
                      (N231)? data_i[587] : 
                      (N232)? data_i[619] : 
                      (N233)? data_i[651] : 
                      (N234)? data_i[683] : 
                      (N235)? data_i[715] : 
                      (N236)? data_i[747] : 
                      (N237)? data_i[779] : 
                      (N238)? data_i[811] : 
                      (N239)? data_i[843] : 
                      (N240)? data_i[875] : 
                      (N241)? data_i[907] : 
                      (N242)? data_i[939] : 
                      (N243)? data_i[971] : 
                      (N244)? data_i[1003] : 
                      (N245)? data_i[1035] : 
                      (N246)? data_i[1067] : 
                      (N247)? data_i[1099] : 
                      (N248)? data_i[1131] : 
                      (N249)? data_i[1163] : 
                      (N250)? data_i[1195] : 
                      (N251)? data_i[1227] : 
                      (N252)? data_i[1259] : 
                      (N253)? data_i[1291] : 
                      (N254)? data_i[1323] : 
                      (N255)? data_i[1355] : 
                      (N256)? data_i[1387] : 
                      (N257)? data_i[1419] : 
                      (N258)? data_i[1451] : 
                      (N259)? data_i[1483] : 
                      (N260)? data_i[1515] : 
                      (N261)? data_i[1547] : 
                      (N262)? data_i[1579] : 1'b0;
  assign data_o[10] = (N213)? data_i[10] : 
                      (N214)? data_i[42] : 
                      (N215)? data_i[74] : 
                      (N216)? data_i[106] : 
                      (N217)? data_i[138] : 
                      (N218)? data_i[170] : 
                      (N219)? data_i[202] : 
                      (N220)? data_i[234] : 
                      (N221)? data_i[266] : 
                      (N222)? data_i[298] : 
                      (N223)? data_i[330] : 
                      (N224)? data_i[362] : 
                      (N225)? data_i[394] : 
                      (N226)? data_i[426] : 
                      (N227)? data_i[458] : 
                      (N228)? data_i[490] : 
                      (N229)? data_i[522] : 
                      (N230)? data_i[554] : 
                      (N231)? data_i[586] : 
                      (N232)? data_i[618] : 
                      (N233)? data_i[650] : 
                      (N234)? data_i[682] : 
                      (N235)? data_i[714] : 
                      (N236)? data_i[746] : 
                      (N237)? data_i[778] : 
                      (N238)? data_i[810] : 
                      (N239)? data_i[842] : 
                      (N240)? data_i[874] : 
                      (N241)? data_i[906] : 
                      (N242)? data_i[938] : 
                      (N243)? data_i[970] : 
                      (N244)? data_i[1002] : 
                      (N245)? data_i[1034] : 
                      (N246)? data_i[1066] : 
                      (N247)? data_i[1098] : 
                      (N248)? data_i[1130] : 
                      (N249)? data_i[1162] : 
                      (N250)? data_i[1194] : 
                      (N251)? data_i[1226] : 
                      (N252)? data_i[1258] : 
                      (N253)? data_i[1290] : 
                      (N254)? data_i[1322] : 
                      (N255)? data_i[1354] : 
                      (N256)? data_i[1386] : 
                      (N257)? data_i[1418] : 
                      (N258)? data_i[1450] : 
                      (N259)? data_i[1482] : 
                      (N260)? data_i[1514] : 
                      (N261)? data_i[1546] : 
                      (N262)? data_i[1578] : 1'b0;
  assign data_o[9] = (N213)? data_i[9] : 
                     (N214)? data_i[41] : 
                     (N215)? data_i[73] : 
                     (N216)? data_i[105] : 
                     (N217)? data_i[137] : 
                     (N218)? data_i[169] : 
                     (N219)? data_i[201] : 
                     (N220)? data_i[233] : 
                     (N221)? data_i[265] : 
                     (N222)? data_i[297] : 
                     (N223)? data_i[329] : 
                     (N224)? data_i[361] : 
                     (N225)? data_i[393] : 
                     (N226)? data_i[425] : 
                     (N227)? data_i[457] : 
                     (N228)? data_i[489] : 
                     (N229)? data_i[521] : 
                     (N230)? data_i[553] : 
                     (N231)? data_i[585] : 
                     (N232)? data_i[617] : 
                     (N233)? data_i[649] : 
                     (N234)? data_i[681] : 
                     (N235)? data_i[713] : 
                     (N236)? data_i[745] : 
                     (N237)? data_i[777] : 
                     (N238)? data_i[809] : 
                     (N239)? data_i[841] : 
                     (N240)? data_i[873] : 
                     (N241)? data_i[905] : 
                     (N242)? data_i[937] : 
                     (N243)? data_i[969] : 
                     (N244)? data_i[1001] : 
                     (N245)? data_i[1033] : 
                     (N246)? data_i[1065] : 
                     (N247)? data_i[1097] : 
                     (N248)? data_i[1129] : 
                     (N249)? data_i[1161] : 
                     (N250)? data_i[1193] : 
                     (N251)? data_i[1225] : 
                     (N252)? data_i[1257] : 
                     (N253)? data_i[1289] : 
                     (N254)? data_i[1321] : 
                     (N255)? data_i[1353] : 
                     (N256)? data_i[1385] : 
                     (N257)? data_i[1417] : 
                     (N258)? data_i[1449] : 
                     (N259)? data_i[1481] : 
                     (N260)? data_i[1513] : 
                     (N261)? data_i[1545] : 
                     (N262)? data_i[1577] : 1'b0;
  assign data_o[8] = (N213)? data_i[8] : 
                     (N214)? data_i[40] : 
                     (N215)? data_i[72] : 
                     (N216)? data_i[104] : 
                     (N217)? data_i[136] : 
                     (N218)? data_i[168] : 
                     (N219)? data_i[200] : 
                     (N220)? data_i[232] : 
                     (N221)? data_i[264] : 
                     (N222)? data_i[296] : 
                     (N223)? data_i[328] : 
                     (N224)? data_i[360] : 
                     (N225)? data_i[392] : 
                     (N226)? data_i[424] : 
                     (N227)? data_i[456] : 
                     (N228)? data_i[488] : 
                     (N229)? data_i[520] : 
                     (N230)? data_i[552] : 
                     (N231)? data_i[584] : 
                     (N232)? data_i[616] : 
                     (N233)? data_i[648] : 
                     (N234)? data_i[680] : 
                     (N235)? data_i[712] : 
                     (N236)? data_i[744] : 
                     (N237)? data_i[776] : 
                     (N238)? data_i[808] : 
                     (N239)? data_i[840] : 
                     (N240)? data_i[872] : 
                     (N241)? data_i[904] : 
                     (N242)? data_i[936] : 
                     (N243)? data_i[968] : 
                     (N244)? data_i[1000] : 
                     (N245)? data_i[1032] : 
                     (N246)? data_i[1064] : 
                     (N247)? data_i[1096] : 
                     (N248)? data_i[1128] : 
                     (N249)? data_i[1160] : 
                     (N250)? data_i[1192] : 
                     (N251)? data_i[1224] : 
                     (N252)? data_i[1256] : 
                     (N253)? data_i[1288] : 
                     (N254)? data_i[1320] : 
                     (N255)? data_i[1352] : 
                     (N256)? data_i[1384] : 
                     (N257)? data_i[1416] : 
                     (N258)? data_i[1448] : 
                     (N259)? data_i[1480] : 
                     (N260)? data_i[1512] : 
                     (N261)? data_i[1544] : 
                     (N262)? data_i[1576] : 1'b0;
  assign data_o[7] = (N213)? data_i[7] : 
                     (N214)? data_i[39] : 
                     (N215)? data_i[71] : 
                     (N216)? data_i[103] : 
                     (N217)? data_i[135] : 
                     (N218)? data_i[167] : 
                     (N219)? data_i[199] : 
                     (N220)? data_i[231] : 
                     (N221)? data_i[263] : 
                     (N222)? data_i[295] : 
                     (N223)? data_i[327] : 
                     (N224)? data_i[359] : 
                     (N225)? data_i[391] : 
                     (N226)? data_i[423] : 
                     (N227)? data_i[455] : 
                     (N228)? data_i[487] : 
                     (N229)? data_i[519] : 
                     (N230)? data_i[551] : 
                     (N231)? data_i[583] : 
                     (N232)? data_i[615] : 
                     (N233)? data_i[647] : 
                     (N234)? data_i[679] : 
                     (N235)? data_i[711] : 
                     (N236)? data_i[743] : 
                     (N237)? data_i[775] : 
                     (N238)? data_i[807] : 
                     (N239)? data_i[839] : 
                     (N240)? data_i[871] : 
                     (N241)? data_i[903] : 
                     (N242)? data_i[935] : 
                     (N243)? data_i[967] : 
                     (N244)? data_i[999] : 
                     (N245)? data_i[1031] : 
                     (N246)? data_i[1063] : 
                     (N247)? data_i[1095] : 
                     (N248)? data_i[1127] : 
                     (N249)? data_i[1159] : 
                     (N250)? data_i[1191] : 
                     (N251)? data_i[1223] : 
                     (N252)? data_i[1255] : 
                     (N253)? data_i[1287] : 
                     (N254)? data_i[1319] : 
                     (N255)? data_i[1351] : 
                     (N256)? data_i[1383] : 
                     (N257)? data_i[1415] : 
                     (N258)? data_i[1447] : 
                     (N259)? data_i[1479] : 
                     (N260)? data_i[1511] : 
                     (N261)? data_i[1543] : 
                     (N262)? data_i[1575] : 1'b0;
  assign data_o[6] = (N213)? data_i[6] : 
                     (N214)? data_i[38] : 
                     (N215)? data_i[70] : 
                     (N216)? data_i[102] : 
                     (N217)? data_i[134] : 
                     (N218)? data_i[166] : 
                     (N219)? data_i[198] : 
                     (N220)? data_i[230] : 
                     (N221)? data_i[262] : 
                     (N222)? data_i[294] : 
                     (N223)? data_i[326] : 
                     (N224)? data_i[358] : 
                     (N225)? data_i[390] : 
                     (N226)? data_i[422] : 
                     (N227)? data_i[454] : 
                     (N228)? data_i[486] : 
                     (N229)? data_i[518] : 
                     (N230)? data_i[550] : 
                     (N231)? data_i[582] : 
                     (N232)? data_i[614] : 
                     (N233)? data_i[646] : 
                     (N234)? data_i[678] : 
                     (N235)? data_i[710] : 
                     (N236)? data_i[742] : 
                     (N237)? data_i[774] : 
                     (N238)? data_i[806] : 
                     (N239)? data_i[838] : 
                     (N240)? data_i[870] : 
                     (N241)? data_i[902] : 
                     (N242)? data_i[934] : 
                     (N243)? data_i[966] : 
                     (N244)? data_i[998] : 
                     (N245)? data_i[1030] : 
                     (N246)? data_i[1062] : 
                     (N247)? data_i[1094] : 
                     (N248)? data_i[1126] : 
                     (N249)? data_i[1158] : 
                     (N250)? data_i[1190] : 
                     (N251)? data_i[1222] : 
                     (N252)? data_i[1254] : 
                     (N253)? data_i[1286] : 
                     (N254)? data_i[1318] : 
                     (N255)? data_i[1350] : 
                     (N256)? data_i[1382] : 
                     (N257)? data_i[1414] : 
                     (N258)? data_i[1446] : 
                     (N259)? data_i[1478] : 
                     (N260)? data_i[1510] : 
                     (N261)? data_i[1542] : 
                     (N262)? data_i[1574] : 1'b0;
  assign data_o[5] = (N213)? data_i[5] : 
                     (N214)? data_i[37] : 
                     (N215)? data_i[69] : 
                     (N216)? data_i[101] : 
                     (N217)? data_i[133] : 
                     (N218)? data_i[165] : 
                     (N219)? data_i[197] : 
                     (N220)? data_i[229] : 
                     (N221)? data_i[261] : 
                     (N222)? data_i[293] : 
                     (N223)? data_i[325] : 
                     (N224)? data_i[357] : 
                     (N225)? data_i[389] : 
                     (N226)? data_i[421] : 
                     (N227)? data_i[453] : 
                     (N228)? data_i[485] : 
                     (N229)? data_i[517] : 
                     (N230)? data_i[549] : 
                     (N231)? data_i[581] : 
                     (N232)? data_i[613] : 
                     (N233)? data_i[645] : 
                     (N234)? data_i[677] : 
                     (N235)? data_i[709] : 
                     (N236)? data_i[741] : 
                     (N237)? data_i[773] : 
                     (N238)? data_i[805] : 
                     (N239)? data_i[837] : 
                     (N240)? data_i[869] : 
                     (N241)? data_i[901] : 
                     (N242)? data_i[933] : 
                     (N243)? data_i[965] : 
                     (N244)? data_i[997] : 
                     (N245)? data_i[1029] : 
                     (N246)? data_i[1061] : 
                     (N247)? data_i[1093] : 
                     (N248)? data_i[1125] : 
                     (N249)? data_i[1157] : 
                     (N250)? data_i[1189] : 
                     (N251)? data_i[1221] : 
                     (N252)? data_i[1253] : 
                     (N253)? data_i[1285] : 
                     (N254)? data_i[1317] : 
                     (N255)? data_i[1349] : 
                     (N256)? data_i[1381] : 
                     (N257)? data_i[1413] : 
                     (N258)? data_i[1445] : 
                     (N259)? data_i[1477] : 
                     (N260)? data_i[1509] : 
                     (N261)? data_i[1541] : 
                     (N262)? data_i[1573] : 1'b0;
  assign data_o[4] = (N213)? data_i[4] : 
                     (N214)? data_i[36] : 
                     (N215)? data_i[68] : 
                     (N216)? data_i[100] : 
                     (N217)? data_i[132] : 
                     (N218)? data_i[164] : 
                     (N219)? data_i[196] : 
                     (N220)? data_i[228] : 
                     (N221)? data_i[260] : 
                     (N222)? data_i[292] : 
                     (N223)? data_i[324] : 
                     (N224)? data_i[356] : 
                     (N225)? data_i[388] : 
                     (N226)? data_i[420] : 
                     (N227)? data_i[452] : 
                     (N228)? data_i[484] : 
                     (N229)? data_i[516] : 
                     (N230)? data_i[548] : 
                     (N231)? data_i[580] : 
                     (N232)? data_i[612] : 
                     (N233)? data_i[644] : 
                     (N234)? data_i[676] : 
                     (N235)? data_i[708] : 
                     (N236)? data_i[740] : 
                     (N237)? data_i[772] : 
                     (N238)? data_i[804] : 
                     (N239)? data_i[836] : 
                     (N240)? data_i[868] : 
                     (N241)? data_i[900] : 
                     (N242)? data_i[932] : 
                     (N243)? data_i[964] : 
                     (N244)? data_i[996] : 
                     (N245)? data_i[1028] : 
                     (N246)? data_i[1060] : 
                     (N247)? data_i[1092] : 
                     (N248)? data_i[1124] : 
                     (N249)? data_i[1156] : 
                     (N250)? data_i[1188] : 
                     (N251)? data_i[1220] : 
                     (N252)? data_i[1252] : 
                     (N253)? data_i[1284] : 
                     (N254)? data_i[1316] : 
                     (N255)? data_i[1348] : 
                     (N256)? data_i[1380] : 
                     (N257)? data_i[1412] : 
                     (N258)? data_i[1444] : 
                     (N259)? data_i[1476] : 
                     (N260)? data_i[1508] : 
                     (N261)? data_i[1540] : 
                     (N262)? data_i[1572] : 1'b0;
  assign data_o[3] = (N213)? data_i[3] : 
                     (N214)? data_i[35] : 
                     (N215)? data_i[67] : 
                     (N216)? data_i[99] : 
                     (N217)? data_i[131] : 
                     (N218)? data_i[163] : 
                     (N219)? data_i[195] : 
                     (N220)? data_i[227] : 
                     (N221)? data_i[259] : 
                     (N222)? data_i[291] : 
                     (N223)? data_i[323] : 
                     (N224)? data_i[355] : 
                     (N225)? data_i[387] : 
                     (N226)? data_i[419] : 
                     (N227)? data_i[451] : 
                     (N228)? data_i[483] : 
                     (N229)? data_i[515] : 
                     (N230)? data_i[547] : 
                     (N231)? data_i[579] : 
                     (N232)? data_i[611] : 
                     (N233)? data_i[643] : 
                     (N234)? data_i[675] : 
                     (N235)? data_i[707] : 
                     (N236)? data_i[739] : 
                     (N237)? data_i[771] : 
                     (N238)? data_i[803] : 
                     (N239)? data_i[835] : 
                     (N240)? data_i[867] : 
                     (N241)? data_i[899] : 
                     (N242)? data_i[931] : 
                     (N243)? data_i[963] : 
                     (N244)? data_i[995] : 
                     (N245)? data_i[1027] : 
                     (N246)? data_i[1059] : 
                     (N247)? data_i[1091] : 
                     (N248)? data_i[1123] : 
                     (N249)? data_i[1155] : 
                     (N250)? data_i[1187] : 
                     (N251)? data_i[1219] : 
                     (N252)? data_i[1251] : 
                     (N253)? data_i[1283] : 
                     (N254)? data_i[1315] : 
                     (N255)? data_i[1347] : 
                     (N256)? data_i[1379] : 
                     (N257)? data_i[1411] : 
                     (N258)? data_i[1443] : 
                     (N259)? data_i[1475] : 
                     (N260)? data_i[1507] : 
                     (N261)? data_i[1539] : 
                     (N262)? data_i[1571] : 1'b0;
  assign data_o[2] = (N213)? data_i[2] : 
                     (N214)? data_i[34] : 
                     (N215)? data_i[66] : 
                     (N216)? data_i[98] : 
                     (N217)? data_i[130] : 
                     (N218)? data_i[162] : 
                     (N219)? data_i[194] : 
                     (N220)? data_i[226] : 
                     (N221)? data_i[258] : 
                     (N222)? data_i[290] : 
                     (N223)? data_i[322] : 
                     (N224)? data_i[354] : 
                     (N225)? data_i[386] : 
                     (N226)? data_i[418] : 
                     (N227)? data_i[450] : 
                     (N228)? data_i[482] : 
                     (N229)? data_i[514] : 
                     (N230)? data_i[546] : 
                     (N231)? data_i[578] : 
                     (N232)? data_i[610] : 
                     (N233)? data_i[642] : 
                     (N234)? data_i[674] : 
                     (N235)? data_i[706] : 
                     (N236)? data_i[738] : 
                     (N237)? data_i[770] : 
                     (N238)? data_i[802] : 
                     (N239)? data_i[834] : 
                     (N240)? data_i[866] : 
                     (N241)? data_i[898] : 
                     (N242)? data_i[930] : 
                     (N243)? data_i[962] : 
                     (N244)? data_i[994] : 
                     (N245)? data_i[1026] : 
                     (N246)? data_i[1058] : 
                     (N247)? data_i[1090] : 
                     (N248)? data_i[1122] : 
                     (N249)? data_i[1154] : 
                     (N250)? data_i[1186] : 
                     (N251)? data_i[1218] : 
                     (N252)? data_i[1250] : 
                     (N253)? data_i[1282] : 
                     (N254)? data_i[1314] : 
                     (N255)? data_i[1346] : 
                     (N256)? data_i[1378] : 
                     (N257)? data_i[1410] : 
                     (N258)? data_i[1442] : 
                     (N259)? data_i[1474] : 
                     (N260)? data_i[1506] : 
                     (N261)? data_i[1538] : 
                     (N262)? data_i[1570] : 1'b0;
  assign data_o[1] = (N213)? data_i[1] : 
                     (N214)? data_i[33] : 
                     (N215)? data_i[65] : 
                     (N216)? data_i[97] : 
                     (N217)? data_i[129] : 
                     (N218)? data_i[161] : 
                     (N219)? data_i[193] : 
                     (N220)? data_i[225] : 
                     (N221)? data_i[257] : 
                     (N222)? data_i[289] : 
                     (N223)? data_i[321] : 
                     (N224)? data_i[353] : 
                     (N225)? data_i[385] : 
                     (N226)? data_i[417] : 
                     (N227)? data_i[449] : 
                     (N228)? data_i[481] : 
                     (N229)? data_i[513] : 
                     (N230)? data_i[545] : 
                     (N231)? data_i[577] : 
                     (N232)? data_i[609] : 
                     (N233)? data_i[641] : 
                     (N234)? data_i[673] : 
                     (N235)? data_i[705] : 
                     (N236)? data_i[737] : 
                     (N237)? data_i[769] : 
                     (N238)? data_i[801] : 
                     (N239)? data_i[833] : 
                     (N240)? data_i[865] : 
                     (N241)? data_i[897] : 
                     (N242)? data_i[929] : 
                     (N243)? data_i[961] : 
                     (N244)? data_i[993] : 
                     (N245)? data_i[1025] : 
                     (N246)? data_i[1057] : 
                     (N247)? data_i[1089] : 
                     (N248)? data_i[1121] : 
                     (N249)? data_i[1153] : 
                     (N250)? data_i[1185] : 
                     (N251)? data_i[1217] : 
                     (N252)? data_i[1249] : 
                     (N253)? data_i[1281] : 
                     (N254)? data_i[1313] : 
                     (N255)? data_i[1345] : 
                     (N256)? data_i[1377] : 
                     (N257)? data_i[1409] : 
                     (N258)? data_i[1441] : 
                     (N259)? data_i[1473] : 
                     (N260)? data_i[1505] : 
                     (N261)? data_i[1537] : 
                     (N262)? data_i[1569] : 1'b0;
  assign data_o[0] = (N213)? data_i[0] : 
                     (N214)? data_i[32] : 
                     (N215)? data_i[64] : 
                     (N216)? data_i[96] : 
                     (N217)? data_i[128] : 
                     (N218)? data_i[160] : 
                     (N219)? data_i[192] : 
                     (N220)? data_i[224] : 
                     (N221)? data_i[256] : 
                     (N222)? data_i[288] : 
                     (N223)? data_i[320] : 
                     (N224)? data_i[352] : 
                     (N225)? data_i[384] : 
                     (N226)? data_i[416] : 
                     (N227)? data_i[448] : 
                     (N228)? data_i[480] : 
                     (N229)? data_i[512] : 
                     (N230)? data_i[544] : 
                     (N231)? data_i[576] : 
                     (N232)? data_i[608] : 
                     (N233)? data_i[640] : 
                     (N234)? data_i[672] : 
                     (N235)? data_i[704] : 
                     (N236)? data_i[736] : 
                     (N237)? data_i[768] : 
                     (N238)? data_i[800] : 
                     (N239)? data_i[832] : 
                     (N240)? data_i[864] : 
                     (N241)? data_i[896] : 
                     (N242)? data_i[928] : 
                     (N243)? data_i[960] : 
                     (N244)? data_i[992] : 
                     (N245)? data_i[1024] : 
                     (N246)? data_i[1056] : 
                     (N247)? data_i[1088] : 
                     (N248)? data_i[1120] : 
                     (N249)? data_i[1152] : 
                     (N250)? data_i[1184] : 
                     (N251)? data_i[1216] : 
                     (N252)? data_i[1248] : 
                     (N253)? data_i[1280] : 
                     (N254)? data_i[1312] : 
                     (N255)? data_i[1344] : 
                     (N256)? data_i[1376] : 
                     (N257)? data_i[1408] : 
                     (N258)? data_i[1440] : 
                     (N259)? data_i[1472] : 
                     (N260)? data_i[1504] : 
                     (N261)? data_i[1536] : 
                     (N262)? data_i[1568] : 1'b0;

endmodule



module bsg_parallel_in_serial_out_dynamic
(
  clk_i,
  reset_i,
  v_i,
  len_i,
  data_i,
  ready_o,
  v_o,
  len_v_o,
  data_o,
  yumi_i
);

  input [5:0] len_i;
  input [1599:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output len_v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,len_v_o,count_r_is_last,up_li,clear_li,N0,N1,N2,N3,N4,N6;
  wire [5:0] len_lo,count_lo;
  wire [1599:0] fifo_data_lo;

  bsg_two_fifo_width_p6
  go_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o),
    .data_i(len_i),
    .v_i(v_i),
    .v_o(v_o),
    .data_o(len_lo),
    .yumi_i(clear_li)
  );


  bsg_two_fifo_width_p1600
  data_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(v_i),
    .data_o(fifo_data_lo),
    .yumi_i(clear_li)
  );

  assign count_r_is_last = count_lo == len_lo;

  bsg_counter_clear_up_max_val_p49_init_val_p0
  ctr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(clear_li),
    .up_i(up_li),
    .count_o(count_lo)
  );


  bsg_mux_width_p32_els_p50
  data_mux
  (
    .data_i(fifo_data_lo),
    .sel_i(count_lo),
    .data_o(data_o)
  );

  assign N0 = count_lo[4] | count_lo[5];
  assign N1 = count_lo[3] | N0;
  assign N2 = count_lo[2] | N1;
  assign N3 = count_lo[1] | N2;
  assign N4 = count_lo[0] | N3;
  assign len_v_o = ~N4;
  assign up_li = yumi_i & N6;
  assign N6 = ~count_r_is_last;
  assign clear_li = yumi_i & count_r_is_last;

endmodule

