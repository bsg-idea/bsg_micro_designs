

module top
(
  i,
  shamt_i,
  sticky_o
);

  input [127:0] i;
  input [7:0] shamt_i;
  output sticky_o;

  bsg_fpu_sticky
  wrapper
  (
    .i(i),
    .shamt_i(shamt_i),
    .sticky_o(sticky_o)
  );


endmodule



module bsg_scan_width_p128_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [127:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire t_3__127_,t_3__126_,t_3__125_,t_3__124_,t_3__123_,t_3__122_,t_3__121_,t_3__120_,
  t_3__119_,t_3__118_,t_3__117_,t_3__116_,t_3__115_,t_3__114_,t_3__113_,t_3__112_,
  t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,t_3__106_,t_3__105_,t_3__104_,
  t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,t_3__98_,t_3__97_,t_3__96_,
  t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,t_3__89_,t_3__88_,t_3__87_,
  t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,t_3__81_,t_3__80_,t_3__79_,t_3__78_,
  t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,t_3__72_,t_3__71_,t_3__70_,t_3__69_,
  t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,t_3__63_,t_3__62_,t_3__61_,t_3__60_,
  t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,t_3__54_,t_3__53_,t_3__52_,
  t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,
  t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,
  t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,
  t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,
  t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,
  t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__127_,t_2__126_,t_2__125_,
  t_2__124_,t_2__123_,t_2__122_,t_2__121_,t_2__120_,t_2__119_,t_2__118_,t_2__117_,
  t_2__116_,t_2__115_,t_2__114_,t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,
  t_2__108_,t_2__107_,t_2__106_,t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,
  t_2__100_,t_2__99_,t_2__98_,t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,
  t_2__92_,t_2__91_,t_2__90_,t_2__89_,t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,
  t_2__83_,t_2__82_,t_2__81_,t_2__80_,t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,
  t_2__74_,t_2__73_,t_2__72_,t_2__71_,t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,
  t_2__65_,t_2__64_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,
  t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,
  t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,
  t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,
  t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_1__127_,t_1__126_,t_1__125_,t_1__124_,t_1__123_,t_1__122_,
  t_1__121_,t_1__120_,t_1__119_,t_1__118_,t_1__117_,t_1__116_,t_1__115_,t_1__114_,
  t_1__113_,t_1__112_,t_1__111_,t_1__110_,t_1__109_,t_1__108_,t_1__107_,t_1__106_,
  t_1__105_,t_1__104_,t_1__103_,t_1__102_,t_1__101_,t_1__100_,t_1__99_,t_1__98_,
  t_1__97_,t_1__96_,t_1__95_,t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,t_1__89_,
  t_1__88_,t_1__87_,t_1__86_,t_1__85_,t_1__84_,t_1__83_,t_1__82_,t_1__81_,t_1__80_,
  t_1__79_,t_1__78_,t_1__77_,t_1__76_,t_1__75_,t_1__74_,t_1__73_,t_1__72_,
  t_1__71_,t_1__70_,t_1__69_,t_1__68_,t_1__67_,t_1__66_,t_1__65_,t_1__64_,t_1__63_,
  t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,t_1__57_,t_1__56_,t_1__55_,t_1__54_,
  t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,
  t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,
  t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,
  t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,
  t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,
  t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_,t_6__127_,
  t_6__126_,t_6__125_,t_6__124_,t_6__123_,t_6__122_,t_6__121_,t_6__120_,t_6__119_,
  t_6__118_,t_6__117_,t_6__116_,t_6__115_,t_6__114_,t_6__113_,t_6__112_,t_6__111_,
  t_6__110_,t_6__109_,t_6__108_,t_6__107_,t_6__106_,t_6__105_,t_6__104_,t_6__103_,
  t_6__102_,t_6__101_,t_6__100_,t_6__99_,t_6__98_,t_6__97_,t_6__96_,t_6__95_,
  t_6__94_,t_6__93_,t_6__92_,t_6__91_,t_6__90_,t_6__89_,t_6__88_,t_6__87_,t_6__86_,
  t_6__85_,t_6__84_,t_6__83_,t_6__82_,t_6__81_,t_6__80_,t_6__79_,t_6__78_,t_6__77_,
  t_6__76_,t_6__75_,t_6__74_,t_6__73_,t_6__72_,t_6__71_,t_6__70_,t_6__69_,t_6__68_,
  t_6__67_,t_6__66_,t_6__65_,t_6__64_,t_6__63_,t_6__62_,t_6__61_,t_6__60_,t_6__59_,
  t_6__58_,t_6__57_,t_6__56_,t_6__55_,t_6__54_,t_6__53_,t_6__52_,t_6__51_,t_6__50_,
  t_6__49_,t_6__48_,t_6__47_,t_6__46_,t_6__45_,t_6__44_,t_6__43_,t_6__42_,
  t_6__41_,t_6__40_,t_6__39_,t_6__38_,t_6__37_,t_6__36_,t_6__35_,t_6__34_,t_6__33_,
  t_6__32_,t_6__31_,t_6__30_,t_6__29_,t_6__28_,t_6__27_,t_6__26_,t_6__25_,t_6__24_,
  t_6__23_,t_6__22_,t_6__21_,t_6__20_,t_6__19_,t_6__18_,t_6__17_,t_6__16_,t_6__15_,
  t_6__14_,t_6__13_,t_6__12_,t_6__11_,t_6__10_,t_6__9_,t_6__8_,t_6__7_,t_6__6_,t_6__5_,
  t_6__4_,t_6__3_,t_6__2_,t_6__1_,t_6__0_,t_5__127_,t_5__126_,t_5__125_,t_5__124_,
  t_5__123_,t_5__122_,t_5__121_,t_5__120_,t_5__119_,t_5__118_,t_5__117_,t_5__116_,
  t_5__115_,t_5__114_,t_5__113_,t_5__112_,t_5__111_,t_5__110_,t_5__109_,t_5__108_,
  t_5__107_,t_5__106_,t_5__105_,t_5__104_,t_5__103_,t_5__102_,t_5__101_,t_5__100_,
  t_5__99_,t_5__98_,t_5__97_,t_5__96_,t_5__95_,t_5__94_,t_5__93_,t_5__92_,
  t_5__91_,t_5__90_,t_5__89_,t_5__88_,t_5__87_,t_5__86_,t_5__85_,t_5__84_,t_5__83_,
  t_5__82_,t_5__81_,t_5__80_,t_5__79_,t_5__78_,t_5__77_,t_5__76_,t_5__75_,t_5__74_,
  t_5__73_,t_5__72_,t_5__71_,t_5__70_,t_5__69_,t_5__68_,t_5__67_,t_5__66_,t_5__65_,
  t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,
  t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,
  t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,
  t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,
  t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,
  t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,
  t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,
  t_5__1_,t_5__0_,t_4__127_,t_4__126_,t_4__125_,t_4__124_,t_4__123_,t_4__122_,t_4__121_,
  t_4__120_,t_4__119_,t_4__118_,t_4__117_,t_4__116_,t_4__115_,t_4__114_,t_4__113_,
  t_4__112_,t_4__111_,t_4__110_,t_4__109_,t_4__108_,t_4__107_,t_4__106_,t_4__105_,
  t_4__104_,t_4__103_,t_4__102_,t_4__101_,t_4__100_,t_4__99_,t_4__98_,t_4__97_,
  t_4__96_,t_4__95_,t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,t_4__89_,t_4__88_,
  t_4__87_,t_4__86_,t_4__85_,t_4__84_,t_4__83_,t_4__82_,t_4__81_,t_4__80_,t_4__79_,
  t_4__78_,t_4__77_,t_4__76_,t_4__75_,t_4__74_,t_4__73_,t_4__72_,t_4__71_,t_4__70_,
  t_4__69_,t_4__68_,t_4__67_,t_4__66_,t_4__65_,t_4__64_,t_4__63_,t_4__62_,
  t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,
  t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,
  t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,
  t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,
  t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,
  t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,
  t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_;
  assign t_1__127_ = i[0] | 1'b0;
  assign t_1__126_ = i[1] | i[0];
  assign t_1__125_ = i[2] | i[1];
  assign t_1__124_ = i[3] | i[2];
  assign t_1__123_ = i[4] | i[3];
  assign t_1__122_ = i[5] | i[4];
  assign t_1__121_ = i[6] | i[5];
  assign t_1__120_ = i[7] | i[6];
  assign t_1__119_ = i[8] | i[7];
  assign t_1__118_ = i[9] | i[8];
  assign t_1__117_ = i[10] | i[9];
  assign t_1__116_ = i[11] | i[10];
  assign t_1__115_ = i[12] | i[11];
  assign t_1__114_ = i[13] | i[12];
  assign t_1__113_ = i[14] | i[13];
  assign t_1__112_ = i[15] | i[14];
  assign t_1__111_ = i[16] | i[15];
  assign t_1__110_ = i[17] | i[16];
  assign t_1__109_ = i[18] | i[17];
  assign t_1__108_ = i[19] | i[18];
  assign t_1__107_ = i[20] | i[19];
  assign t_1__106_ = i[21] | i[20];
  assign t_1__105_ = i[22] | i[21];
  assign t_1__104_ = i[23] | i[22];
  assign t_1__103_ = i[24] | i[23];
  assign t_1__102_ = i[25] | i[24];
  assign t_1__101_ = i[26] | i[25];
  assign t_1__100_ = i[27] | i[26];
  assign t_1__99_ = i[28] | i[27];
  assign t_1__98_ = i[29] | i[28];
  assign t_1__97_ = i[30] | i[29];
  assign t_1__96_ = i[31] | i[30];
  assign t_1__95_ = i[32] | i[31];
  assign t_1__94_ = i[33] | i[32];
  assign t_1__93_ = i[34] | i[33];
  assign t_1__92_ = i[35] | i[34];
  assign t_1__91_ = i[36] | i[35];
  assign t_1__90_ = i[37] | i[36];
  assign t_1__89_ = i[38] | i[37];
  assign t_1__88_ = i[39] | i[38];
  assign t_1__87_ = i[40] | i[39];
  assign t_1__86_ = i[41] | i[40];
  assign t_1__85_ = i[42] | i[41];
  assign t_1__84_ = i[43] | i[42];
  assign t_1__83_ = i[44] | i[43];
  assign t_1__82_ = i[45] | i[44];
  assign t_1__81_ = i[46] | i[45];
  assign t_1__80_ = i[47] | i[46];
  assign t_1__79_ = i[48] | i[47];
  assign t_1__78_ = i[49] | i[48];
  assign t_1__77_ = i[50] | i[49];
  assign t_1__76_ = i[51] | i[50];
  assign t_1__75_ = i[52] | i[51];
  assign t_1__74_ = i[53] | i[52];
  assign t_1__73_ = i[54] | i[53];
  assign t_1__72_ = i[55] | i[54];
  assign t_1__71_ = i[56] | i[55];
  assign t_1__70_ = i[57] | i[56];
  assign t_1__69_ = i[58] | i[57];
  assign t_1__68_ = i[59] | i[58];
  assign t_1__67_ = i[60] | i[59];
  assign t_1__66_ = i[61] | i[60];
  assign t_1__65_ = i[62] | i[61];
  assign t_1__64_ = i[63] | i[62];
  assign t_1__63_ = i[64] | i[63];
  assign t_1__62_ = i[65] | i[64];
  assign t_1__61_ = i[66] | i[65];
  assign t_1__60_ = i[67] | i[66];
  assign t_1__59_ = i[68] | i[67];
  assign t_1__58_ = i[69] | i[68];
  assign t_1__57_ = i[70] | i[69];
  assign t_1__56_ = i[71] | i[70];
  assign t_1__55_ = i[72] | i[71];
  assign t_1__54_ = i[73] | i[72];
  assign t_1__53_ = i[74] | i[73];
  assign t_1__52_ = i[75] | i[74];
  assign t_1__51_ = i[76] | i[75];
  assign t_1__50_ = i[77] | i[76];
  assign t_1__49_ = i[78] | i[77];
  assign t_1__48_ = i[79] | i[78];
  assign t_1__47_ = i[80] | i[79];
  assign t_1__46_ = i[81] | i[80];
  assign t_1__45_ = i[82] | i[81];
  assign t_1__44_ = i[83] | i[82];
  assign t_1__43_ = i[84] | i[83];
  assign t_1__42_ = i[85] | i[84];
  assign t_1__41_ = i[86] | i[85];
  assign t_1__40_ = i[87] | i[86];
  assign t_1__39_ = i[88] | i[87];
  assign t_1__38_ = i[89] | i[88];
  assign t_1__37_ = i[90] | i[89];
  assign t_1__36_ = i[91] | i[90];
  assign t_1__35_ = i[92] | i[91];
  assign t_1__34_ = i[93] | i[92];
  assign t_1__33_ = i[94] | i[93];
  assign t_1__32_ = i[95] | i[94];
  assign t_1__31_ = i[96] | i[95];
  assign t_1__30_ = i[97] | i[96];
  assign t_1__29_ = i[98] | i[97];
  assign t_1__28_ = i[99] | i[98];
  assign t_1__27_ = i[100] | i[99];
  assign t_1__26_ = i[101] | i[100];
  assign t_1__25_ = i[102] | i[101];
  assign t_1__24_ = i[103] | i[102];
  assign t_1__23_ = i[104] | i[103];
  assign t_1__22_ = i[105] | i[104];
  assign t_1__21_ = i[106] | i[105];
  assign t_1__20_ = i[107] | i[106];
  assign t_1__19_ = i[108] | i[107];
  assign t_1__18_ = i[109] | i[108];
  assign t_1__17_ = i[110] | i[109];
  assign t_1__16_ = i[111] | i[110];
  assign t_1__15_ = i[112] | i[111];
  assign t_1__14_ = i[113] | i[112];
  assign t_1__13_ = i[114] | i[113];
  assign t_1__12_ = i[115] | i[114];
  assign t_1__11_ = i[116] | i[115];
  assign t_1__10_ = i[117] | i[116];
  assign t_1__9_ = i[118] | i[117];
  assign t_1__8_ = i[119] | i[118];
  assign t_1__7_ = i[120] | i[119];
  assign t_1__6_ = i[121] | i[120];
  assign t_1__5_ = i[122] | i[121];
  assign t_1__4_ = i[123] | i[122];
  assign t_1__3_ = i[124] | i[123];
  assign t_1__2_ = i[125] | i[124];
  assign t_1__1_ = i[126] | i[125];
  assign t_1__0_ = i[127] | i[126];
  assign t_2__127_ = t_1__127_ | 1'b0;
  assign t_2__126_ = t_1__126_ | 1'b0;
  assign t_2__125_ = t_1__125_ | t_1__127_;
  assign t_2__124_ = t_1__124_ | t_1__126_;
  assign t_2__123_ = t_1__123_ | t_1__125_;
  assign t_2__122_ = t_1__122_ | t_1__124_;
  assign t_2__121_ = t_1__121_ | t_1__123_;
  assign t_2__120_ = t_1__120_ | t_1__122_;
  assign t_2__119_ = t_1__119_ | t_1__121_;
  assign t_2__118_ = t_1__118_ | t_1__120_;
  assign t_2__117_ = t_1__117_ | t_1__119_;
  assign t_2__116_ = t_1__116_ | t_1__118_;
  assign t_2__115_ = t_1__115_ | t_1__117_;
  assign t_2__114_ = t_1__114_ | t_1__116_;
  assign t_2__113_ = t_1__113_ | t_1__115_;
  assign t_2__112_ = t_1__112_ | t_1__114_;
  assign t_2__111_ = t_1__111_ | t_1__113_;
  assign t_2__110_ = t_1__110_ | t_1__112_;
  assign t_2__109_ = t_1__109_ | t_1__111_;
  assign t_2__108_ = t_1__108_ | t_1__110_;
  assign t_2__107_ = t_1__107_ | t_1__109_;
  assign t_2__106_ = t_1__106_ | t_1__108_;
  assign t_2__105_ = t_1__105_ | t_1__107_;
  assign t_2__104_ = t_1__104_ | t_1__106_;
  assign t_2__103_ = t_1__103_ | t_1__105_;
  assign t_2__102_ = t_1__102_ | t_1__104_;
  assign t_2__101_ = t_1__101_ | t_1__103_;
  assign t_2__100_ = t_1__100_ | t_1__102_;
  assign t_2__99_ = t_1__99_ | t_1__101_;
  assign t_2__98_ = t_1__98_ | t_1__100_;
  assign t_2__97_ = t_1__97_ | t_1__99_;
  assign t_2__96_ = t_1__96_ | t_1__98_;
  assign t_2__95_ = t_1__95_ | t_1__97_;
  assign t_2__94_ = t_1__94_ | t_1__96_;
  assign t_2__93_ = t_1__93_ | t_1__95_;
  assign t_2__92_ = t_1__92_ | t_1__94_;
  assign t_2__91_ = t_1__91_ | t_1__93_;
  assign t_2__90_ = t_1__90_ | t_1__92_;
  assign t_2__89_ = t_1__89_ | t_1__91_;
  assign t_2__88_ = t_1__88_ | t_1__90_;
  assign t_2__87_ = t_1__87_ | t_1__89_;
  assign t_2__86_ = t_1__86_ | t_1__88_;
  assign t_2__85_ = t_1__85_ | t_1__87_;
  assign t_2__84_ = t_1__84_ | t_1__86_;
  assign t_2__83_ = t_1__83_ | t_1__85_;
  assign t_2__82_ = t_1__82_ | t_1__84_;
  assign t_2__81_ = t_1__81_ | t_1__83_;
  assign t_2__80_ = t_1__80_ | t_1__82_;
  assign t_2__79_ = t_1__79_ | t_1__81_;
  assign t_2__78_ = t_1__78_ | t_1__80_;
  assign t_2__77_ = t_1__77_ | t_1__79_;
  assign t_2__76_ = t_1__76_ | t_1__78_;
  assign t_2__75_ = t_1__75_ | t_1__77_;
  assign t_2__74_ = t_1__74_ | t_1__76_;
  assign t_2__73_ = t_1__73_ | t_1__75_;
  assign t_2__72_ = t_1__72_ | t_1__74_;
  assign t_2__71_ = t_1__71_ | t_1__73_;
  assign t_2__70_ = t_1__70_ | t_1__72_;
  assign t_2__69_ = t_1__69_ | t_1__71_;
  assign t_2__68_ = t_1__68_ | t_1__70_;
  assign t_2__67_ = t_1__67_ | t_1__69_;
  assign t_2__66_ = t_1__66_ | t_1__68_;
  assign t_2__65_ = t_1__65_ | t_1__67_;
  assign t_2__64_ = t_1__64_ | t_1__66_;
  assign t_2__63_ = t_1__63_ | t_1__65_;
  assign t_2__62_ = t_1__62_ | t_1__64_;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__127_ = t_2__127_ | 1'b0;
  assign t_3__126_ = t_2__126_ | 1'b0;
  assign t_3__125_ = t_2__125_ | 1'b0;
  assign t_3__124_ = t_2__124_ | 1'b0;
  assign t_3__123_ = t_2__123_ | t_2__127_;
  assign t_3__122_ = t_2__122_ | t_2__126_;
  assign t_3__121_ = t_2__121_ | t_2__125_;
  assign t_3__120_ = t_2__120_ | t_2__124_;
  assign t_3__119_ = t_2__119_ | t_2__123_;
  assign t_3__118_ = t_2__118_ | t_2__122_;
  assign t_3__117_ = t_2__117_ | t_2__121_;
  assign t_3__116_ = t_2__116_ | t_2__120_;
  assign t_3__115_ = t_2__115_ | t_2__119_;
  assign t_3__114_ = t_2__114_ | t_2__118_;
  assign t_3__113_ = t_2__113_ | t_2__117_;
  assign t_3__112_ = t_2__112_ | t_2__116_;
  assign t_3__111_ = t_2__111_ | t_2__115_;
  assign t_3__110_ = t_2__110_ | t_2__114_;
  assign t_3__109_ = t_2__109_ | t_2__113_;
  assign t_3__108_ = t_2__108_ | t_2__112_;
  assign t_3__107_ = t_2__107_ | t_2__111_;
  assign t_3__106_ = t_2__106_ | t_2__110_;
  assign t_3__105_ = t_2__105_ | t_2__109_;
  assign t_3__104_ = t_2__104_ | t_2__108_;
  assign t_3__103_ = t_2__103_ | t_2__107_;
  assign t_3__102_ = t_2__102_ | t_2__106_;
  assign t_3__101_ = t_2__101_ | t_2__105_;
  assign t_3__100_ = t_2__100_ | t_2__104_;
  assign t_3__99_ = t_2__99_ | t_2__103_;
  assign t_3__98_ = t_2__98_ | t_2__102_;
  assign t_3__97_ = t_2__97_ | t_2__101_;
  assign t_3__96_ = t_2__96_ | t_2__100_;
  assign t_3__95_ = t_2__95_ | t_2__99_;
  assign t_3__94_ = t_2__94_ | t_2__98_;
  assign t_3__93_ = t_2__93_ | t_2__97_;
  assign t_3__92_ = t_2__92_ | t_2__96_;
  assign t_3__91_ = t_2__91_ | t_2__95_;
  assign t_3__90_ = t_2__90_ | t_2__94_;
  assign t_3__89_ = t_2__89_ | t_2__93_;
  assign t_3__88_ = t_2__88_ | t_2__92_;
  assign t_3__87_ = t_2__87_ | t_2__91_;
  assign t_3__86_ = t_2__86_ | t_2__90_;
  assign t_3__85_ = t_2__85_ | t_2__89_;
  assign t_3__84_ = t_2__84_ | t_2__88_;
  assign t_3__83_ = t_2__83_ | t_2__87_;
  assign t_3__82_ = t_2__82_ | t_2__86_;
  assign t_3__81_ = t_2__81_ | t_2__85_;
  assign t_3__80_ = t_2__80_ | t_2__84_;
  assign t_3__79_ = t_2__79_ | t_2__83_;
  assign t_3__78_ = t_2__78_ | t_2__82_;
  assign t_3__77_ = t_2__77_ | t_2__81_;
  assign t_3__76_ = t_2__76_ | t_2__80_;
  assign t_3__75_ = t_2__75_ | t_2__79_;
  assign t_3__74_ = t_2__74_ | t_2__78_;
  assign t_3__73_ = t_2__73_ | t_2__77_;
  assign t_3__72_ = t_2__72_ | t_2__76_;
  assign t_3__71_ = t_2__71_ | t_2__75_;
  assign t_3__70_ = t_2__70_ | t_2__74_;
  assign t_3__69_ = t_2__69_ | t_2__73_;
  assign t_3__68_ = t_2__68_ | t_2__72_;
  assign t_3__67_ = t_2__67_ | t_2__71_;
  assign t_3__66_ = t_2__66_ | t_2__70_;
  assign t_3__65_ = t_2__65_ | t_2__69_;
  assign t_3__64_ = t_2__64_ | t_2__68_;
  assign t_3__63_ = t_2__63_ | t_2__67_;
  assign t_3__62_ = t_2__62_ | t_2__66_;
  assign t_3__61_ = t_2__61_ | t_2__65_;
  assign t_3__60_ = t_2__60_ | t_2__64_;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__127_ = t_3__127_ | 1'b0;
  assign t_4__126_ = t_3__126_ | 1'b0;
  assign t_4__125_ = t_3__125_ | 1'b0;
  assign t_4__124_ = t_3__124_ | 1'b0;
  assign t_4__123_ = t_3__123_ | 1'b0;
  assign t_4__122_ = t_3__122_ | 1'b0;
  assign t_4__121_ = t_3__121_ | 1'b0;
  assign t_4__120_ = t_3__120_ | 1'b0;
  assign t_4__119_ = t_3__119_ | t_3__127_;
  assign t_4__118_ = t_3__118_ | t_3__126_;
  assign t_4__117_ = t_3__117_ | t_3__125_;
  assign t_4__116_ = t_3__116_ | t_3__124_;
  assign t_4__115_ = t_3__115_ | t_3__123_;
  assign t_4__114_ = t_3__114_ | t_3__122_;
  assign t_4__113_ = t_3__113_ | t_3__121_;
  assign t_4__112_ = t_3__112_ | t_3__120_;
  assign t_4__111_ = t_3__111_ | t_3__119_;
  assign t_4__110_ = t_3__110_ | t_3__118_;
  assign t_4__109_ = t_3__109_ | t_3__117_;
  assign t_4__108_ = t_3__108_ | t_3__116_;
  assign t_4__107_ = t_3__107_ | t_3__115_;
  assign t_4__106_ = t_3__106_ | t_3__114_;
  assign t_4__105_ = t_3__105_ | t_3__113_;
  assign t_4__104_ = t_3__104_ | t_3__112_;
  assign t_4__103_ = t_3__103_ | t_3__111_;
  assign t_4__102_ = t_3__102_ | t_3__110_;
  assign t_4__101_ = t_3__101_ | t_3__109_;
  assign t_4__100_ = t_3__100_ | t_3__108_;
  assign t_4__99_ = t_3__99_ | t_3__107_;
  assign t_4__98_ = t_3__98_ | t_3__106_;
  assign t_4__97_ = t_3__97_ | t_3__105_;
  assign t_4__96_ = t_3__96_ | t_3__104_;
  assign t_4__95_ = t_3__95_ | t_3__103_;
  assign t_4__94_ = t_3__94_ | t_3__102_;
  assign t_4__93_ = t_3__93_ | t_3__101_;
  assign t_4__92_ = t_3__92_ | t_3__100_;
  assign t_4__91_ = t_3__91_ | t_3__99_;
  assign t_4__90_ = t_3__90_ | t_3__98_;
  assign t_4__89_ = t_3__89_ | t_3__97_;
  assign t_4__88_ = t_3__88_ | t_3__96_;
  assign t_4__87_ = t_3__87_ | t_3__95_;
  assign t_4__86_ = t_3__86_ | t_3__94_;
  assign t_4__85_ = t_3__85_ | t_3__93_;
  assign t_4__84_ = t_3__84_ | t_3__92_;
  assign t_4__83_ = t_3__83_ | t_3__91_;
  assign t_4__82_ = t_3__82_ | t_3__90_;
  assign t_4__81_ = t_3__81_ | t_3__89_;
  assign t_4__80_ = t_3__80_ | t_3__88_;
  assign t_4__79_ = t_3__79_ | t_3__87_;
  assign t_4__78_ = t_3__78_ | t_3__86_;
  assign t_4__77_ = t_3__77_ | t_3__85_;
  assign t_4__76_ = t_3__76_ | t_3__84_;
  assign t_4__75_ = t_3__75_ | t_3__83_;
  assign t_4__74_ = t_3__74_ | t_3__82_;
  assign t_4__73_ = t_3__73_ | t_3__81_;
  assign t_4__72_ = t_3__72_ | t_3__80_;
  assign t_4__71_ = t_3__71_ | t_3__79_;
  assign t_4__70_ = t_3__70_ | t_3__78_;
  assign t_4__69_ = t_3__69_ | t_3__77_;
  assign t_4__68_ = t_3__68_ | t_3__76_;
  assign t_4__67_ = t_3__67_ | t_3__75_;
  assign t_4__66_ = t_3__66_ | t_3__74_;
  assign t_4__65_ = t_3__65_ | t_3__73_;
  assign t_4__64_ = t_3__64_ | t_3__72_;
  assign t_4__63_ = t_3__63_ | t_3__71_;
  assign t_4__62_ = t_3__62_ | t_3__70_;
  assign t_4__61_ = t_3__61_ | t_3__69_;
  assign t_4__60_ = t_3__60_ | t_3__68_;
  assign t_4__59_ = t_3__59_ | t_3__67_;
  assign t_4__58_ = t_3__58_ | t_3__66_;
  assign t_4__57_ = t_3__57_ | t_3__65_;
  assign t_4__56_ = t_3__56_ | t_3__64_;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__127_ = t_4__127_ | 1'b0;
  assign t_5__126_ = t_4__126_ | 1'b0;
  assign t_5__125_ = t_4__125_ | 1'b0;
  assign t_5__124_ = t_4__124_ | 1'b0;
  assign t_5__123_ = t_4__123_ | 1'b0;
  assign t_5__122_ = t_4__122_ | 1'b0;
  assign t_5__121_ = t_4__121_ | 1'b0;
  assign t_5__120_ = t_4__120_ | 1'b0;
  assign t_5__119_ = t_4__119_ | 1'b0;
  assign t_5__118_ = t_4__118_ | 1'b0;
  assign t_5__117_ = t_4__117_ | 1'b0;
  assign t_5__116_ = t_4__116_ | 1'b0;
  assign t_5__115_ = t_4__115_ | 1'b0;
  assign t_5__114_ = t_4__114_ | 1'b0;
  assign t_5__113_ = t_4__113_ | 1'b0;
  assign t_5__112_ = t_4__112_ | 1'b0;
  assign t_5__111_ = t_4__111_ | t_4__127_;
  assign t_5__110_ = t_4__110_ | t_4__126_;
  assign t_5__109_ = t_4__109_ | t_4__125_;
  assign t_5__108_ = t_4__108_ | t_4__124_;
  assign t_5__107_ = t_4__107_ | t_4__123_;
  assign t_5__106_ = t_4__106_ | t_4__122_;
  assign t_5__105_ = t_4__105_ | t_4__121_;
  assign t_5__104_ = t_4__104_ | t_4__120_;
  assign t_5__103_ = t_4__103_ | t_4__119_;
  assign t_5__102_ = t_4__102_ | t_4__118_;
  assign t_5__101_ = t_4__101_ | t_4__117_;
  assign t_5__100_ = t_4__100_ | t_4__116_;
  assign t_5__99_ = t_4__99_ | t_4__115_;
  assign t_5__98_ = t_4__98_ | t_4__114_;
  assign t_5__97_ = t_4__97_ | t_4__113_;
  assign t_5__96_ = t_4__96_ | t_4__112_;
  assign t_5__95_ = t_4__95_ | t_4__111_;
  assign t_5__94_ = t_4__94_ | t_4__110_;
  assign t_5__93_ = t_4__93_ | t_4__109_;
  assign t_5__92_ = t_4__92_ | t_4__108_;
  assign t_5__91_ = t_4__91_ | t_4__107_;
  assign t_5__90_ = t_4__90_ | t_4__106_;
  assign t_5__89_ = t_4__89_ | t_4__105_;
  assign t_5__88_ = t_4__88_ | t_4__104_;
  assign t_5__87_ = t_4__87_ | t_4__103_;
  assign t_5__86_ = t_4__86_ | t_4__102_;
  assign t_5__85_ = t_4__85_ | t_4__101_;
  assign t_5__84_ = t_4__84_ | t_4__100_;
  assign t_5__83_ = t_4__83_ | t_4__99_;
  assign t_5__82_ = t_4__82_ | t_4__98_;
  assign t_5__81_ = t_4__81_ | t_4__97_;
  assign t_5__80_ = t_4__80_ | t_4__96_;
  assign t_5__79_ = t_4__79_ | t_4__95_;
  assign t_5__78_ = t_4__78_ | t_4__94_;
  assign t_5__77_ = t_4__77_ | t_4__93_;
  assign t_5__76_ = t_4__76_ | t_4__92_;
  assign t_5__75_ = t_4__75_ | t_4__91_;
  assign t_5__74_ = t_4__74_ | t_4__90_;
  assign t_5__73_ = t_4__73_ | t_4__89_;
  assign t_5__72_ = t_4__72_ | t_4__88_;
  assign t_5__71_ = t_4__71_ | t_4__87_;
  assign t_5__70_ = t_4__70_ | t_4__86_;
  assign t_5__69_ = t_4__69_ | t_4__85_;
  assign t_5__68_ = t_4__68_ | t_4__84_;
  assign t_5__67_ = t_4__67_ | t_4__83_;
  assign t_5__66_ = t_4__66_ | t_4__82_;
  assign t_5__65_ = t_4__65_ | t_4__81_;
  assign t_5__64_ = t_4__64_ | t_4__80_;
  assign t_5__63_ = t_4__63_ | t_4__79_;
  assign t_5__62_ = t_4__62_ | t_4__78_;
  assign t_5__61_ = t_4__61_ | t_4__77_;
  assign t_5__60_ = t_4__60_ | t_4__76_;
  assign t_5__59_ = t_4__59_ | t_4__75_;
  assign t_5__58_ = t_4__58_ | t_4__74_;
  assign t_5__57_ = t_4__57_ | t_4__73_;
  assign t_5__56_ = t_4__56_ | t_4__72_;
  assign t_5__55_ = t_4__55_ | t_4__71_;
  assign t_5__54_ = t_4__54_ | t_4__70_;
  assign t_5__53_ = t_4__53_ | t_4__69_;
  assign t_5__52_ = t_4__52_ | t_4__68_;
  assign t_5__51_ = t_4__51_ | t_4__67_;
  assign t_5__50_ = t_4__50_ | t_4__66_;
  assign t_5__49_ = t_4__49_ | t_4__65_;
  assign t_5__48_ = t_4__48_ | t_4__64_;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign t_6__127_ = t_5__127_ | 1'b0;
  assign t_6__126_ = t_5__126_ | 1'b0;
  assign t_6__125_ = t_5__125_ | 1'b0;
  assign t_6__124_ = t_5__124_ | 1'b0;
  assign t_6__123_ = t_5__123_ | 1'b0;
  assign t_6__122_ = t_5__122_ | 1'b0;
  assign t_6__121_ = t_5__121_ | 1'b0;
  assign t_6__120_ = t_5__120_ | 1'b0;
  assign t_6__119_ = t_5__119_ | 1'b0;
  assign t_6__118_ = t_5__118_ | 1'b0;
  assign t_6__117_ = t_5__117_ | 1'b0;
  assign t_6__116_ = t_5__116_ | 1'b0;
  assign t_6__115_ = t_5__115_ | 1'b0;
  assign t_6__114_ = t_5__114_ | 1'b0;
  assign t_6__113_ = t_5__113_ | 1'b0;
  assign t_6__112_ = t_5__112_ | 1'b0;
  assign t_6__111_ = t_5__111_ | 1'b0;
  assign t_6__110_ = t_5__110_ | 1'b0;
  assign t_6__109_ = t_5__109_ | 1'b0;
  assign t_6__108_ = t_5__108_ | 1'b0;
  assign t_6__107_ = t_5__107_ | 1'b0;
  assign t_6__106_ = t_5__106_ | 1'b0;
  assign t_6__105_ = t_5__105_ | 1'b0;
  assign t_6__104_ = t_5__104_ | 1'b0;
  assign t_6__103_ = t_5__103_ | 1'b0;
  assign t_6__102_ = t_5__102_ | 1'b0;
  assign t_6__101_ = t_5__101_ | 1'b0;
  assign t_6__100_ = t_5__100_ | 1'b0;
  assign t_6__99_ = t_5__99_ | 1'b0;
  assign t_6__98_ = t_5__98_ | 1'b0;
  assign t_6__97_ = t_5__97_ | 1'b0;
  assign t_6__96_ = t_5__96_ | 1'b0;
  assign t_6__95_ = t_5__95_ | t_5__127_;
  assign t_6__94_ = t_5__94_ | t_5__126_;
  assign t_6__93_ = t_5__93_ | t_5__125_;
  assign t_6__92_ = t_5__92_ | t_5__124_;
  assign t_6__91_ = t_5__91_ | t_5__123_;
  assign t_6__90_ = t_5__90_ | t_5__122_;
  assign t_6__89_ = t_5__89_ | t_5__121_;
  assign t_6__88_ = t_5__88_ | t_5__120_;
  assign t_6__87_ = t_5__87_ | t_5__119_;
  assign t_6__86_ = t_5__86_ | t_5__118_;
  assign t_6__85_ = t_5__85_ | t_5__117_;
  assign t_6__84_ = t_5__84_ | t_5__116_;
  assign t_6__83_ = t_5__83_ | t_5__115_;
  assign t_6__82_ = t_5__82_ | t_5__114_;
  assign t_6__81_ = t_5__81_ | t_5__113_;
  assign t_6__80_ = t_5__80_ | t_5__112_;
  assign t_6__79_ = t_5__79_ | t_5__111_;
  assign t_6__78_ = t_5__78_ | t_5__110_;
  assign t_6__77_ = t_5__77_ | t_5__109_;
  assign t_6__76_ = t_5__76_ | t_5__108_;
  assign t_6__75_ = t_5__75_ | t_5__107_;
  assign t_6__74_ = t_5__74_ | t_5__106_;
  assign t_6__73_ = t_5__73_ | t_5__105_;
  assign t_6__72_ = t_5__72_ | t_5__104_;
  assign t_6__71_ = t_5__71_ | t_5__103_;
  assign t_6__70_ = t_5__70_ | t_5__102_;
  assign t_6__69_ = t_5__69_ | t_5__101_;
  assign t_6__68_ = t_5__68_ | t_5__100_;
  assign t_6__67_ = t_5__67_ | t_5__99_;
  assign t_6__66_ = t_5__66_ | t_5__98_;
  assign t_6__65_ = t_5__65_ | t_5__97_;
  assign t_6__64_ = t_5__64_ | t_5__96_;
  assign t_6__63_ = t_5__63_ | t_5__95_;
  assign t_6__62_ = t_5__62_ | t_5__94_;
  assign t_6__61_ = t_5__61_ | t_5__93_;
  assign t_6__60_ = t_5__60_ | t_5__92_;
  assign t_6__59_ = t_5__59_ | t_5__91_;
  assign t_6__58_ = t_5__58_ | t_5__90_;
  assign t_6__57_ = t_5__57_ | t_5__89_;
  assign t_6__56_ = t_5__56_ | t_5__88_;
  assign t_6__55_ = t_5__55_ | t_5__87_;
  assign t_6__54_ = t_5__54_ | t_5__86_;
  assign t_6__53_ = t_5__53_ | t_5__85_;
  assign t_6__52_ = t_5__52_ | t_5__84_;
  assign t_6__51_ = t_5__51_ | t_5__83_;
  assign t_6__50_ = t_5__50_ | t_5__82_;
  assign t_6__49_ = t_5__49_ | t_5__81_;
  assign t_6__48_ = t_5__48_ | t_5__80_;
  assign t_6__47_ = t_5__47_ | t_5__79_;
  assign t_6__46_ = t_5__46_ | t_5__78_;
  assign t_6__45_ = t_5__45_ | t_5__77_;
  assign t_6__44_ = t_5__44_ | t_5__76_;
  assign t_6__43_ = t_5__43_ | t_5__75_;
  assign t_6__42_ = t_5__42_ | t_5__74_;
  assign t_6__41_ = t_5__41_ | t_5__73_;
  assign t_6__40_ = t_5__40_ | t_5__72_;
  assign t_6__39_ = t_5__39_ | t_5__71_;
  assign t_6__38_ = t_5__38_ | t_5__70_;
  assign t_6__37_ = t_5__37_ | t_5__69_;
  assign t_6__36_ = t_5__36_ | t_5__68_;
  assign t_6__35_ = t_5__35_ | t_5__67_;
  assign t_6__34_ = t_5__34_ | t_5__66_;
  assign t_6__33_ = t_5__33_ | t_5__65_;
  assign t_6__32_ = t_5__32_ | t_5__64_;
  assign t_6__31_ = t_5__31_ | t_5__63_;
  assign t_6__30_ = t_5__30_ | t_5__62_;
  assign t_6__29_ = t_5__29_ | t_5__61_;
  assign t_6__28_ = t_5__28_ | t_5__60_;
  assign t_6__27_ = t_5__27_ | t_5__59_;
  assign t_6__26_ = t_5__26_ | t_5__58_;
  assign t_6__25_ = t_5__25_ | t_5__57_;
  assign t_6__24_ = t_5__24_ | t_5__56_;
  assign t_6__23_ = t_5__23_ | t_5__55_;
  assign t_6__22_ = t_5__22_ | t_5__54_;
  assign t_6__21_ = t_5__21_ | t_5__53_;
  assign t_6__20_ = t_5__20_ | t_5__52_;
  assign t_6__19_ = t_5__19_ | t_5__51_;
  assign t_6__18_ = t_5__18_ | t_5__50_;
  assign t_6__17_ = t_5__17_ | t_5__49_;
  assign t_6__16_ = t_5__16_ | t_5__48_;
  assign t_6__15_ = t_5__15_ | t_5__47_;
  assign t_6__14_ = t_5__14_ | t_5__46_;
  assign t_6__13_ = t_5__13_ | t_5__45_;
  assign t_6__12_ = t_5__12_ | t_5__44_;
  assign t_6__11_ = t_5__11_ | t_5__43_;
  assign t_6__10_ = t_5__10_ | t_5__42_;
  assign t_6__9_ = t_5__9_ | t_5__41_;
  assign t_6__8_ = t_5__8_ | t_5__40_;
  assign t_6__7_ = t_5__7_ | t_5__39_;
  assign t_6__6_ = t_5__6_ | t_5__38_;
  assign t_6__5_ = t_5__5_ | t_5__37_;
  assign t_6__4_ = t_5__4_ | t_5__36_;
  assign t_6__3_ = t_5__3_ | t_5__35_;
  assign t_6__2_ = t_5__2_ | t_5__34_;
  assign t_6__1_ = t_5__1_ | t_5__33_;
  assign t_6__0_ = t_5__0_ | t_5__32_;
  assign o[0] = t_6__127_ | 1'b0;
  assign o[1] = t_6__126_ | 1'b0;
  assign o[2] = t_6__125_ | 1'b0;
  assign o[3] = t_6__124_ | 1'b0;
  assign o[4] = t_6__123_ | 1'b0;
  assign o[5] = t_6__122_ | 1'b0;
  assign o[6] = t_6__121_ | 1'b0;
  assign o[7] = t_6__120_ | 1'b0;
  assign o[8] = t_6__119_ | 1'b0;
  assign o[9] = t_6__118_ | 1'b0;
  assign o[10] = t_6__117_ | 1'b0;
  assign o[11] = t_6__116_ | 1'b0;
  assign o[12] = t_6__115_ | 1'b0;
  assign o[13] = t_6__114_ | 1'b0;
  assign o[14] = t_6__113_ | 1'b0;
  assign o[15] = t_6__112_ | 1'b0;
  assign o[16] = t_6__111_ | 1'b0;
  assign o[17] = t_6__110_ | 1'b0;
  assign o[18] = t_6__109_ | 1'b0;
  assign o[19] = t_6__108_ | 1'b0;
  assign o[20] = t_6__107_ | 1'b0;
  assign o[21] = t_6__106_ | 1'b0;
  assign o[22] = t_6__105_ | 1'b0;
  assign o[23] = t_6__104_ | 1'b0;
  assign o[24] = t_6__103_ | 1'b0;
  assign o[25] = t_6__102_ | 1'b0;
  assign o[26] = t_6__101_ | 1'b0;
  assign o[27] = t_6__100_ | 1'b0;
  assign o[28] = t_6__99_ | 1'b0;
  assign o[29] = t_6__98_ | 1'b0;
  assign o[30] = t_6__97_ | 1'b0;
  assign o[31] = t_6__96_ | 1'b0;
  assign o[32] = t_6__95_ | 1'b0;
  assign o[33] = t_6__94_ | 1'b0;
  assign o[34] = t_6__93_ | 1'b0;
  assign o[35] = t_6__92_ | 1'b0;
  assign o[36] = t_6__91_ | 1'b0;
  assign o[37] = t_6__90_ | 1'b0;
  assign o[38] = t_6__89_ | 1'b0;
  assign o[39] = t_6__88_ | 1'b0;
  assign o[40] = t_6__87_ | 1'b0;
  assign o[41] = t_6__86_ | 1'b0;
  assign o[42] = t_6__85_ | 1'b0;
  assign o[43] = t_6__84_ | 1'b0;
  assign o[44] = t_6__83_ | 1'b0;
  assign o[45] = t_6__82_ | 1'b0;
  assign o[46] = t_6__81_ | 1'b0;
  assign o[47] = t_6__80_ | 1'b0;
  assign o[48] = t_6__79_ | 1'b0;
  assign o[49] = t_6__78_ | 1'b0;
  assign o[50] = t_6__77_ | 1'b0;
  assign o[51] = t_6__76_ | 1'b0;
  assign o[52] = t_6__75_ | 1'b0;
  assign o[53] = t_6__74_ | 1'b0;
  assign o[54] = t_6__73_ | 1'b0;
  assign o[55] = t_6__72_ | 1'b0;
  assign o[56] = t_6__71_ | 1'b0;
  assign o[57] = t_6__70_ | 1'b0;
  assign o[58] = t_6__69_ | 1'b0;
  assign o[59] = t_6__68_ | 1'b0;
  assign o[60] = t_6__67_ | 1'b0;
  assign o[61] = t_6__66_ | 1'b0;
  assign o[62] = t_6__65_ | 1'b0;
  assign o[63] = t_6__64_ | 1'b0;
  assign o[64] = t_6__63_ | t_6__127_;
  assign o[65] = t_6__62_ | t_6__126_;
  assign o[66] = t_6__61_ | t_6__125_;
  assign o[67] = t_6__60_ | t_6__124_;
  assign o[68] = t_6__59_ | t_6__123_;
  assign o[69] = t_6__58_ | t_6__122_;
  assign o[70] = t_6__57_ | t_6__121_;
  assign o[71] = t_6__56_ | t_6__120_;
  assign o[72] = t_6__55_ | t_6__119_;
  assign o[73] = t_6__54_ | t_6__118_;
  assign o[74] = t_6__53_ | t_6__117_;
  assign o[75] = t_6__52_ | t_6__116_;
  assign o[76] = t_6__51_ | t_6__115_;
  assign o[77] = t_6__50_ | t_6__114_;
  assign o[78] = t_6__49_ | t_6__113_;
  assign o[79] = t_6__48_ | t_6__112_;
  assign o[80] = t_6__47_ | t_6__111_;
  assign o[81] = t_6__46_ | t_6__110_;
  assign o[82] = t_6__45_ | t_6__109_;
  assign o[83] = t_6__44_ | t_6__108_;
  assign o[84] = t_6__43_ | t_6__107_;
  assign o[85] = t_6__42_ | t_6__106_;
  assign o[86] = t_6__41_ | t_6__105_;
  assign o[87] = t_6__40_ | t_6__104_;
  assign o[88] = t_6__39_ | t_6__103_;
  assign o[89] = t_6__38_ | t_6__102_;
  assign o[90] = t_6__37_ | t_6__101_;
  assign o[91] = t_6__36_ | t_6__100_;
  assign o[92] = t_6__35_ | t_6__99_;
  assign o[93] = t_6__34_ | t_6__98_;
  assign o[94] = t_6__33_ | t_6__97_;
  assign o[95] = t_6__32_ | t_6__96_;
  assign o[96] = t_6__31_ | t_6__95_;
  assign o[97] = t_6__30_ | t_6__94_;
  assign o[98] = t_6__29_ | t_6__93_;
  assign o[99] = t_6__28_ | t_6__92_;
  assign o[100] = t_6__27_ | t_6__91_;
  assign o[101] = t_6__26_ | t_6__90_;
  assign o[102] = t_6__25_ | t_6__89_;
  assign o[103] = t_6__24_ | t_6__88_;
  assign o[104] = t_6__23_ | t_6__87_;
  assign o[105] = t_6__22_ | t_6__86_;
  assign o[106] = t_6__21_ | t_6__85_;
  assign o[107] = t_6__20_ | t_6__84_;
  assign o[108] = t_6__19_ | t_6__83_;
  assign o[109] = t_6__18_ | t_6__82_;
  assign o[110] = t_6__17_ | t_6__81_;
  assign o[111] = t_6__16_ | t_6__80_;
  assign o[112] = t_6__15_ | t_6__79_;
  assign o[113] = t_6__14_ | t_6__78_;
  assign o[114] = t_6__13_ | t_6__77_;
  assign o[115] = t_6__12_ | t_6__76_;
  assign o[116] = t_6__11_ | t_6__75_;
  assign o[117] = t_6__10_ | t_6__74_;
  assign o[118] = t_6__9_ | t_6__73_;
  assign o[119] = t_6__8_ | t_6__72_;
  assign o[120] = t_6__7_ | t_6__71_;
  assign o[121] = t_6__6_ | t_6__70_;
  assign o[122] = t_6__5_ | t_6__69_;
  assign o[123] = t_6__4_ | t_6__68_;
  assign o[124] = t_6__3_ | t_6__67_;
  assign o[125] = t_6__2_ | t_6__66_;
  assign o[126] = t_6__1_ | t_6__65_;
  assign o[127] = t_6__0_ | t_6__64_;

endmodule



module bsg_fpu_sticky
(
  i,
  shamt_i,
  sticky_o
);

  input [127:0] i;
  input [7:0] shamt_i;
  output sticky_o;
  wire sticky_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,
  N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
  N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,
  N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,
  N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,
  N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,
  N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,
  N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
  N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,
  N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,
  N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
  N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,
  N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,
  N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,
  N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,
  N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,
  N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,
  N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,
  N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,
  N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,
  N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,
  N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,
  N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,
  N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,
  N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,
  N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,
  N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,
  N1343,N1344;
  wire [127:0] scan_out;

  bsg_scan_width_p128_or_p1_lo_to_hi_p1
  scan0
  (
    .i(i),
    .o(scan_out)
  );

  assign N1214 = shamt_i > { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign N1216 = N0 & N1 & (N2 & N3) & (N4 & N5 & (N6 & N7));
  assign N0 = ~shamt_i[7];
  assign N1 = ~shamt_i[6];
  assign N2 = ~shamt_i[5];
  assign N3 = ~shamt_i[4];
  assign N4 = ~shamt_i[3];
  assign N5 = ~shamt_i[2];
  assign N6 = ~shamt_i[0];
  assign N7 = ~shamt_i[1];
  assign N8 = N13 & N14;
  assign N9 = N8 & N15;
  assign N10 = N9 & N16;
  assign N11 = N10 & N17;
  assign N12 = N11 & shamt_i[0];
  assign N1217 = N12 & N18;
  assign N13 = ~shamt_i[6];
  assign N14 = ~shamt_i[5];
  assign N15 = ~shamt_i[4];
  assign N16 = ~shamt_i[3];
  assign N17 = ~shamt_i[2];
  assign N18 = ~shamt_i[1];
  assign N19 = N24 & N25;
  assign N20 = N19 & N26;
  assign N21 = N20 & N27;
  assign N22 = N21 & N28;
  assign N23 = N22 & N29;
  assign N1218 = N23 & shamt_i[1];
  assign N24 = ~shamt_i[6];
  assign N25 = ~shamt_i[5];
  assign N26 = ~shamt_i[4];
  assign N27 = ~shamt_i[3];
  assign N28 = ~shamt_i[2];
  assign N29 = ~shamt_i[0];
  assign N30 = N35 & N36;
  assign N31 = N30 & N37;
  assign N32 = N31 & N38;
  assign N33 = N32 & N39;
  assign N34 = N33 & shamt_i[0];
  assign N1219 = N34 & shamt_i[1];
  assign N35 = ~shamt_i[6];
  assign N36 = ~shamt_i[5];
  assign N37 = ~shamt_i[4];
  assign N38 = ~shamt_i[3];
  assign N39 = ~shamt_i[2];
  assign N40 = N45 & N46;
  assign N41 = N40 & N47;
  assign N42 = N41 & N48;
  assign N43 = N42 & shamt_i[2];
  assign N44 = N43 & N49;
  assign N1220 = N44 & N50;
  assign N45 = ~shamt_i[6];
  assign N46 = ~shamt_i[5];
  assign N47 = ~shamt_i[4];
  assign N48 = ~shamt_i[3];
  assign N49 = ~shamt_i[0];
  assign N50 = ~shamt_i[1];
  assign N51 = N56 & N57;
  assign N52 = N51 & N58;
  assign N53 = N52 & N59;
  assign N54 = N53 & shamt_i[2];
  assign N55 = N54 & shamt_i[0];
  assign N1221 = N55 & N60;
  assign N56 = ~shamt_i[6];
  assign N57 = ~shamt_i[5];
  assign N58 = ~shamt_i[4];
  assign N59 = ~shamt_i[3];
  assign N60 = ~shamt_i[1];
  assign N61 = N66 & N67;
  assign N62 = N61 & N68;
  assign N63 = N62 & N69;
  assign N64 = N63 & shamt_i[2];
  assign N65 = N64 & N70;
  assign N1222 = N65 & shamt_i[1];
  assign N66 = ~shamt_i[6];
  assign N67 = ~shamt_i[5];
  assign N68 = ~shamt_i[4];
  assign N69 = ~shamt_i[3];
  assign N70 = ~shamt_i[0];
  assign N71 = N76 & N77;
  assign N72 = N71 & N78;
  assign N73 = N72 & N79;
  assign N74 = N73 & shamt_i[2];
  assign N75 = N74 & shamt_i[0];
  assign N1223 = N75 & shamt_i[1];
  assign N76 = ~shamt_i[6];
  assign N77 = ~shamt_i[5];
  assign N78 = ~shamt_i[4];
  assign N79 = ~shamt_i[3];
  assign N80 = N85 & N86;
  assign N81 = N80 & N87;
  assign N82 = N81 & shamt_i[3];
  assign N83 = N82 & N88;
  assign N84 = N83 & N89;
  assign N1224 = N84 & N90;
  assign N85 = ~shamt_i[6];
  assign N86 = ~shamt_i[5];
  assign N87 = ~shamt_i[4];
  assign N88 = ~shamt_i[2];
  assign N89 = ~shamt_i[0];
  assign N90 = ~shamt_i[1];
  assign N91 = N96 & N97;
  assign N92 = N91 & N98;
  assign N93 = N92 & shamt_i[3];
  assign N94 = N93 & N99;
  assign N95 = N94 & shamt_i[0];
  assign N1225 = N95 & N100;
  assign N96 = ~shamt_i[6];
  assign N97 = ~shamt_i[5];
  assign N98 = ~shamt_i[4];
  assign N99 = ~shamt_i[2];
  assign N100 = ~shamt_i[1];
  assign N101 = N106 & N107;
  assign N102 = N101 & N108;
  assign N103 = N102 & shamt_i[3];
  assign N104 = N103 & N109;
  assign N105 = N104 & N110;
  assign N1226 = N105 & shamt_i[1];
  assign N106 = ~shamt_i[6];
  assign N107 = ~shamt_i[5];
  assign N108 = ~shamt_i[4];
  assign N109 = ~shamt_i[2];
  assign N110 = ~shamt_i[0];
  assign N111 = N116 & N117;
  assign N112 = N111 & N118;
  assign N113 = N112 & shamt_i[3];
  assign N114 = N113 & N119;
  assign N115 = N114 & shamt_i[0];
  assign N1227 = N115 & shamt_i[1];
  assign N116 = ~shamt_i[6];
  assign N117 = ~shamt_i[5];
  assign N118 = ~shamt_i[4];
  assign N119 = ~shamt_i[2];
  assign N120 = N125 & N126;
  assign N121 = N120 & N127;
  assign N122 = N121 & shamt_i[3];
  assign N123 = N122 & shamt_i[2];
  assign N124 = N123 & N128;
  assign N1228 = N124 & N129;
  assign N125 = ~shamt_i[6];
  assign N126 = ~shamt_i[5];
  assign N127 = ~shamt_i[4];
  assign N128 = ~shamt_i[0];
  assign N129 = ~shamt_i[1];
  assign N130 = N135 & N136;
  assign N131 = N130 & N137;
  assign N132 = N131 & shamt_i[3];
  assign N133 = N132 & shamt_i[2];
  assign N134 = N133 & shamt_i[0];
  assign N1229 = N134 & N138;
  assign N135 = ~shamt_i[6];
  assign N136 = ~shamt_i[5];
  assign N137 = ~shamt_i[4];
  assign N138 = ~shamt_i[1];
  assign N139 = N144 & N145;
  assign N140 = N139 & N146;
  assign N141 = N140 & shamt_i[3];
  assign N142 = N141 & shamt_i[2];
  assign N143 = N142 & N147;
  assign N1230 = N143 & shamt_i[1];
  assign N144 = ~shamt_i[6];
  assign N145 = ~shamt_i[5];
  assign N146 = ~shamt_i[4];
  assign N147 = ~shamt_i[0];
  assign N148 = N153 & N154;
  assign N149 = N148 & N155;
  assign N150 = N149 & shamt_i[3];
  assign N151 = N150 & shamt_i[2];
  assign N152 = N151 & shamt_i[0];
  assign N1231 = N152 & shamt_i[1];
  assign N153 = ~shamt_i[6];
  assign N154 = ~shamt_i[5];
  assign N155 = ~shamt_i[4];
  assign N156 = N161 & N162;
  assign N157 = N156 & shamt_i[4];
  assign N158 = N157 & N163;
  assign N159 = N158 & N164;
  assign N160 = N159 & N165;
  assign N1232 = N160 & N166;
  assign N161 = ~shamt_i[6];
  assign N162 = ~shamt_i[5];
  assign N163 = ~shamt_i[3];
  assign N164 = ~shamt_i[2];
  assign N165 = ~shamt_i[0];
  assign N166 = ~shamt_i[1];
  assign N167 = N172 & N173;
  assign N168 = N167 & shamt_i[4];
  assign N169 = N168 & N174;
  assign N170 = N169 & N175;
  assign N171 = N170 & shamt_i[0];
  assign N1233 = N171 & N176;
  assign N172 = ~shamt_i[6];
  assign N173 = ~shamt_i[5];
  assign N174 = ~shamt_i[3];
  assign N175 = ~shamt_i[2];
  assign N176 = ~shamt_i[1];
  assign N177 = N182 & N183;
  assign N178 = N177 & shamt_i[4];
  assign N179 = N178 & N184;
  assign N180 = N179 & N185;
  assign N181 = N180 & N186;
  assign N1234 = N181 & shamt_i[1];
  assign N182 = ~shamt_i[6];
  assign N183 = ~shamt_i[5];
  assign N184 = ~shamt_i[3];
  assign N185 = ~shamt_i[2];
  assign N186 = ~shamt_i[0];
  assign N187 = N192 & N193;
  assign N188 = N187 & shamt_i[4];
  assign N189 = N188 & N194;
  assign N190 = N189 & N195;
  assign N191 = N190 & shamt_i[0];
  assign N1235 = N191 & shamt_i[1];
  assign N192 = ~shamt_i[6];
  assign N193 = ~shamt_i[5];
  assign N194 = ~shamt_i[3];
  assign N195 = ~shamt_i[2];
  assign N196 = N201 & N202;
  assign N197 = N196 & shamt_i[4];
  assign N198 = N197 & N203;
  assign N199 = N198 & shamt_i[2];
  assign N200 = N199 & N204;
  assign N1236 = N200 & N205;
  assign N201 = ~shamt_i[6];
  assign N202 = ~shamt_i[5];
  assign N203 = ~shamt_i[3];
  assign N204 = ~shamt_i[0];
  assign N205 = ~shamt_i[1];
  assign N206 = N211 & N212;
  assign N207 = N206 & shamt_i[4];
  assign N208 = N207 & N213;
  assign N209 = N208 & shamt_i[2];
  assign N210 = N209 & shamt_i[0];
  assign N1237 = N210 & N214;
  assign N211 = ~shamt_i[6];
  assign N212 = ~shamt_i[5];
  assign N213 = ~shamt_i[3];
  assign N214 = ~shamt_i[1];
  assign N215 = N220 & N221;
  assign N216 = N215 & shamt_i[4];
  assign N217 = N216 & N222;
  assign N218 = N217 & shamt_i[2];
  assign N219 = N218 & N223;
  assign N1238 = N219 & shamt_i[1];
  assign N220 = ~shamt_i[6];
  assign N221 = ~shamt_i[5];
  assign N222 = ~shamt_i[3];
  assign N223 = ~shamt_i[0];
  assign N224 = N229 & N230;
  assign N225 = N224 & shamt_i[4];
  assign N226 = N225 & N231;
  assign N227 = N226 & shamt_i[2];
  assign N228 = N227 & shamt_i[0];
  assign N1239 = N228 & shamt_i[1];
  assign N229 = ~shamt_i[6];
  assign N230 = ~shamt_i[5];
  assign N231 = ~shamt_i[3];
  assign N232 = N237 & N238;
  assign N233 = N232 & shamt_i[4];
  assign N234 = N233 & shamt_i[3];
  assign N235 = N234 & N239;
  assign N236 = N235 & N240;
  assign N1240 = N236 & N241;
  assign N237 = ~shamt_i[6];
  assign N238 = ~shamt_i[5];
  assign N239 = ~shamt_i[2];
  assign N240 = ~shamt_i[0];
  assign N241 = ~shamt_i[1];
  assign N242 = N247 & N248;
  assign N243 = N242 & shamt_i[4];
  assign N244 = N243 & shamt_i[3];
  assign N245 = N244 & N249;
  assign N246 = N245 & shamt_i[0];
  assign N1241 = N246 & N250;
  assign N247 = ~shamt_i[6];
  assign N248 = ~shamt_i[5];
  assign N249 = ~shamt_i[2];
  assign N250 = ~shamt_i[1];
  assign N251 = N256 & N257;
  assign N252 = N251 & shamt_i[4];
  assign N253 = N252 & shamt_i[3];
  assign N254 = N253 & N258;
  assign N255 = N254 & N259;
  assign N1242 = N255 & shamt_i[1];
  assign N256 = ~shamt_i[6];
  assign N257 = ~shamt_i[5];
  assign N258 = ~shamt_i[2];
  assign N259 = ~shamt_i[0];
  assign N260 = N265 & N266;
  assign N261 = N260 & shamt_i[4];
  assign N262 = N261 & shamt_i[3];
  assign N263 = N262 & N267;
  assign N264 = N263 & shamt_i[0];
  assign N1243 = N264 & shamt_i[1];
  assign N265 = ~shamt_i[6];
  assign N266 = ~shamt_i[5];
  assign N267 = ~shamt_i[2];
  assign N268 = N273 & N274;
  assign N269 = N268 & shamt_i[4];
  assign N270 = N269 & shamt_i[3];
  assign N271 = N270 & shamt_i[2];
  assign N272 = N271 & N275;
  assign N1244 = N272 & N276;
  assign N273 = ~shamt_i[6];
  assign N274 = ~shamt_i[5];
  assign N275 = ~shamt_i[0];
  assign N276 = ~shamt_i[1];
  assign N277 = N282 & N283;
  assign N278 = N277 & shamt_i[4];
  assign N279 = N278 & shamt_i[3];
  assign N280 = N279 & shamt_i[2];
  assign N281 = N280 & shamt_i[0];
  assign N1245 = N281 & N284;
  assign N282 = ~shamt_i[6];
  assign N283 = ~shamt_i[5];
  assign N284 = ~shamt_i[1];
  assign N285 = N290 & N291;
  assign N286 = N285 & shamt_i[4];
  assign N287 = N286 & shamt_i[3];
  assign N288 = N287 & shamt_i[2];
  assign N289 = N288 & N292;
  assign N1246 = N289 & shamt_i[1];
  assign N290 = ~shamt_i[6];
  assign N291 = ~shamt_i[5];
  assign N292 = ~shamt_i[0];
  assign N293 = N298 & N299;
  assign N294 = N293 & shamt_i[4];
  assign N295 = N294 & shamt_i[3];
  assign N296 = N295 & shamt_i[2];
  assign N297 = N296 & shamt_i[0];
  assign N1247 = N297 & shamt_i[1];
  assign N298 = ~shamt_i[6];
  assign N299 = ~shamt_i[5];
  assign N300 = N305 & shamt_i[5];
  assign N301 = N300 & N306;
  assign N302 = N301 & N307;
  assign N303 = N302 & N308;
  assign N304 = N303 & N309;
  assign N1248 = N304 & N310;
  assign N305 = ~shamt_i[6];
  assign N306 = ~shamt_i[4];
  assign N307 = ~shamt_i[3];
  assign N308 = ~shamt_i[2];
  assign N309 = ~shamt_i[0];
  assign N310 = ~shamt_i[1];
  assign N311 = N316 & shamt_i[5];
  assign N312 = N311 & N317;
  assign N313 = N312 & N318;
  assign N314 = N313 & N319;
  assign N315 = N314 & shamt_i[0];
  assign N1249 = N315 & N320;
  assign N316 = ~shamt_i[6];
  assign N317 = ~shamt_i[4];
  assign N318 = ~shamt_i[3];
  assign N319 = ~shamt_i[2];
  assign N320 = ~shamt_i[1];
  assign N321 = N326 & shamt_i[5];
  assign N322 = N321 & N327;
  assign N323 = N322 & N328;
  assign N324 = N323 & N329;
  assign N325 = N324 & N330;
  assign N1250 = N325 & shamt_i[1];
  assign N326 = ~shamt_i[6];
  assign N327 = ~shamt_i[4];
  assign N328 = ~shamt_i[3];
  assign N329 = ~shamt_i[2];
  assign N330 = ~shamt_i[0];
  assign N331 = N336 & shamt_i[5];
  assign N332 = N331 & N337;
  assign N333 = N332 & N338;
  assign N334 = N333 & N339;
  assign N335 = N334 & shamt_i[0];
  assign N1251 = N335 & shamt_i[1];
  assign N336 = ~shamt_i[6];
  assign N337 = ~shamt_i[4];
  assign N338 = ~shamt_i[3];
  assign N339 = ~shamt_i[2];
  assign N340 = N345 & shamt_i[5];
  assign N341 = N340 & N346;
  assign N342 = N341 & N347;
  assign N343 = N342 & shamt_i[2];
  assign N344 = N343 & N348;
  assign N1252 = N344 & N349;
  assign N345 = ~shamt_i[6];
  assign N346 = ~shamt_i[4];
  assign N347 = ~shamt_i[3];
  assign N348 = ~shamt_i[0];
  assign N349 = ~shamt_i[1];
  assign N350 = N355 & shamt_i[5];
  assign N351 = N350 & N356;
  assign N352 = N351 & N357;
  assign N353 = N352 & shamt_i[2];
  assign N354 = N353 & shamt_i[0];
  assign N1253 = N354 & N358;
  assign N355 = ~shamt_i[6];
  assign N356 = ~shamt_i[4];
  assign N357 = ~shamt_i[3];
  assign N358 = ~shamt_i[1];
  assign N359 = N364 & shamt_i[5];
  assign N360 = N359 & N365;
  assign N361 = N360 & N366;
  assign N362 = N361 & shamt_i[2];
  assign N363 = N362 & N367;
  assign N1254 = N363 & shamt_i[1];
  assign N364 = ~shamt_i[6];
  assign N365 = ~shamt_i[4];
  assign N366 = ~shamt_i[3];
  assign N367 = ~shamt_i[0];
  assign N368 = N373 & shamt_i[5];
  assign N369 = N368 & N374;
  assign N370 = N369 & N375;
  assign N371 = N370 & shamt_i[2];
  assign N372 = N371 & shamt_i[0];
  assign N1255 = N372 & shamt_i[1];
  assign N373 = ~shamt_i[6];
  assign N374 = ~shamt_i[4];
  assign N375 = ~shamt_i[3];
  assign N376 = N381 & shamt_i[5];
  assign N377 = N376 & N382;
  assign N378 = N377 & shamt_i[3];
  assign N379 = N378 & N383;
  assign N380 = N379 & N384;
  assign N1256 = N380 & N385;
  assign N381 = ~shamt_i[6];
  assign N382 = ~shamt_i[4];
  assign N383 = ~shamt_i[2];
  assign N384 = ~shamt_i[0];
  assign N385 = ~shamt_i[1];
  assign N386 = N391 & shamt_i[5];
  assign N387 = N386 & N392;
  assign N388 = N387 & shamt_i[3];
  assign N389 = N388 & N393;
  assign N390 = N389 & shamt_i[0];
  assign N1257 = N390 & N394;
  assign N391 = ~shamt_i[6];
  assign N392 = ~shamt_i[4];
  assign N393 = ~shamt_i[2];
  assign N394 = ~shamt_i[1];
  assign N395 = N400 & shamt_i[5];
  assign N396 = N395 & N401;
  assign N397 = N396 & shamt_i[3];
  assign N398 = N397 & N402;
  assign N399 = N398 & N403;
  assign N1258 = N399 & shamt_i[1];
  assign N400 = ~shamt_i[6];
  assign N401 = ~shamt_i[4];
  assign N402 = ~shamt_i[2];
  assign N403 = ~shamt_i[0];
  assign N404 = N409 & shamt_i[5];
  assign N405 = N404 & N410;
  assign N406 = N405 & shamt_i[3];
  assign N407 = N406 & N411;
  assign N408 = N407 & shamt_i[0];
  assign N1259 = N408 & shamt_i[1];
  assign N409 = ~shamt_i[6];
  assign N410 = ~shamt_i[4];
  assign N411 = ~shamt_i[2];
  assign N412 = N417 & shamt_i[5];
  assign N413 = N412 & N418;
  assign N414 = N413 & shamt_i[3];
  assign N415 = N414 & shamt_i[2];
  assign N416 = N415 & N419;
  assign N1260 = N416 & N420;
  assign N417 = ~shamt_i[6];
  assign N418 = ~shamt_i[4];
  assign N419 = ~shamt_i[0];
  assign N420 = ~shamt_i[1];
  assign N421 = N426 & shamt_i[5];
  assign N422 = N421 & N427;
  assign N423 = N422 & shamt_i[3];
  assign N424 = N423 & shamt_i[2];
  assign N425 = N424 & shamt_i[0];
  assign N1261 = N425 & N428;
  assign N426 = ~shamt_i[6];
  assign N427 = ~shamt_i[4];
  assign N428 = ~shamt_i[1];
  assign N429 = N434 & shamt_i[5];
  assign N430 = N429 & N435;
  assign N431 = N430 & shamt_i[3];
  assign N432 = N431 & shamt_i[2];
  assign N433 = N432 & N436;
  assign N1262 = N433 & shamt_i[1];
  assign N434 = ~shamt_i[6];
  assign N435 = ~shamt_i[4];
  assign N436 = ~shamt_i[0];
  assign N437 = N442 & shamt_i[5];
  assign N438 = N437 & N443;
  assign N439 = N438 & shamt_i[3];
  assign N440 = N439 & shamt_i[2];
  assign N441 = N440 & shamt_i[0];
  assign N1263 = N441 & shamt_i[1];
  assign N442 = ~shamt_i[6];
  assign N443 = ~shamt_i[4];
  assign N444 = N449 & shamt_i[5];
  assign N445 = N444 & shamt_i[4];
  assign N446 = N445 & N450;
  assign N447 = N446 & N451;
  assign N448 = N447 & N452;
  assign N1264 = N448 & N453;
  assign N449 = ~shamt_i[6];
  assign N450 = ~shamt_i[3];
  assign N451 = ~shamt_i[2];
  assign N452 = ~shamt_i[0];
  assign N453 = ~shamt_i[1];
  assign N454 = N459 & shamt_i[5];
  assign N455 = N454 & shamt_i[4];
  assign N456 = N455 & N460;
  assign N457 = N456 & N461;
  assign N458 = N457 & shamt_i[0];
  assign N1265 = N458 & N462;
  assign N459 = ~shamt_i[6];
  assign N460 = ~shamt_i[3];
  assign N461 = ~shamt_i[2];
  assign N462 = ~shamt_i[1];
  assign N463 = N468 & shamt_i[5];
  assign N464 = N463 & shamt_i[4];
  assign N465 = N464 & N469;
  assign N466 = N465 & N470;
  assign N467 = N466 & N471;
  assign N1266 = N467 & shamt_i[1];
  assign N468 = ~shamt_i[6];
  assign N469 = ~shamt_i[3];
  assign N470 = ~shamt_i[2];
  assign N471 = ~shamt_i[0];
  assign N472 = N477 & shamt_i[5];
  assign N473 = N472 & shamt_i[4];
  assign N474 = N473 & N478;
  assign N475 = N474 & N479;
  assign N476 = N475 & shamt_i[0];
  assign N1267 = N476 & shamt_i[1];
  assign N477 = ~shamt_i[6];
  assign N478 = ~shamt_i[3];
  assign N479 = ~shamt_i[2];
  assign N480 = N485 & shamt_i[5];
  assign N481 = N480 & shamt_i[4];
  assign N482 = N481 & N486;
  assign N483 = N482 & shamt_i[2];
  assign N484 = N483 & N487;
  assign N1268 = N484 & N488;
  assign N485 = ~shamt_i[6];
  assign N486 = ~shamt_i[3];
  assign N487 = ~shamt_i[0];
  assign N488 = ~shamt_i[1];
  assign N489 = N494 & shamt_i[5];
  assign N490 = N489 & shamt_i[4];
  assign N491 = N490 & N495;
  assign N492 = N491 & shamt_i[2];
  assign N493 = N492 & shamt_i[0];
  assign N1269 = N493 & N496;
  assign N494 = ~shamt_i[6];
  assign N495 = ~shamt_i[3];
  assign N496 = ~shamt_i[1];
  assign N497 = N502 & shamt_i[5];
  assign N498 = N497 & shamt_i[4];
  assign N499 = N498 & N503;
  assign N500 = N499 & shamt_i[2];
  assign N501 = N500 & N504;
  assign N1270 = N501 & shamt_i[1];
  assign N502 = ~shamt_i[6];
  assign N503 = ~shamt_i[3];
  assign N504 = ~shamt_i[0];
  assign N505 = N510 & shamt_i[5];
  assign N506 = N505 & shamt_i[4];
  assign N507 = N506 & N511;
  assign N508 = N507 & shamt_i[2];
  assign N509 = N508 & shamt_i[0];
  assign N1271 = N509 & shamt_i[1];
  assign N510 = ~shamt_i[6];
  assign N511 = ~shamt_i[3];
  assign N512 = N517 & shamt_i[5];
  assign N513 = N512 & shamt_i[4];
  assign N514 = N513 & shamt_i[3];
  assign N515 = N514 & N518;
  assign N516 = N515 & N519;
  assign N1272 = N516 & N520;
  assign N517 = ~shamt_i[6];
  assign N518 = ~shamt_i[2];
  assign N519 = ~shamt_i[0];
  assign N520 = ~shamt_i[1];
  assign N521 = N526 & shamt_i[5];
  assign N522 = N521 & shamt_i[4];
  assign N523 = N522 & shamt_i[3];
  assign N524 = N523 & N527;
  assign N525 = N524 & shamt_i[0];
  assign N1273 = N525 & N528;
  assign N526 = ~shamt_i[6];
  assign N527 = ~shamt_i[2];
  assign N528 = ~shamt_i[1];
  assign N529 = N534 & shamt_i[5];
  assign N530 = N529 & shamt_i[4];
  assign N531 = N530 & shamt_i[3];
  assign N532 = N531 & N535;
  assign N533 = N532 & N536;
  assign N1274 = N533 & shamt_i[1];
  assign N534 = ~shamt_i[6];
  assign N535 = ~shamt_i[2];
  assign N536 = ~shamt_i[0];
  assign N537 = N542 & shamt_i[5];
  assign N538 = N537 & shamt_i[4];
  assign N539 = N538 & shamt_i[3];
  assign N540 = N539 & N543;
  assign N541 = N540 & shamt_i[0];
  assign N1275 = N541 & shamt_i[1];
  assign N542 = ~shamt_i[6];
  assign N543 = ~shamt_i[2];
  assign N544 = N549 & shamt_i[5];
  assign N545 = N544 & shamt_i[4];
  assign N546 = N545 & shamt_i[3];
  assign N547 = N546 & shamt_i[2];
  assign N548 = N547 & N550;
  assign N1276 = N548 & N551;
  assign N549 = ~shamt_i[6];
  assign N550 = ~shamt_i[0];
  assign N551 = ~shamt_i[1];
  assign N552 = N557 & shamt_i[5];
  assign N553 = N552 & shamt_i[4];
  assign N554 = N553 & shamt_i[3];
  assign N555 = N554 & shamt_i[2];
  assign N556 = N555 & shamt_i[0];
  assign N1277 = N556 & N558;
  assign N557 = ~shamt_i[6];
  assign N558 = ~shamt_i[1];
  assign N559 = N564 & shamt_i[5];
  assign N560 = N559 & shamt_i[4];
  assign N561 = N560 & shamt_i[3];
  assign N562 = N561 & shamt_i[2];
  assign N563 = N562 & N565;
  assign N1278 = N563 & shamt_i[1];
  assign N564 = ~shamt_i[6];
  assign N565 = ~shamt_i[0];
  assign N566 = N571 & shamt_i[5];
  assign N567 = N566 & shamt_i[4];
  assign N568 = N567 & shamt_i[3];
  assign N569 = N568 & shamt_i[2];
  assign N570 = N569 & shamt_i[0];
  assign N1279 = N570 & shamt_i[1];
  assign N571 = ~shamt_i[6];
  assign N572 = shamt_i[6] & N577;
  assign N573 = N572 & N578;
  assign N574 = N573 & N579;
  assign N575 = N574 & N580;
  assign N576 = N575 & N581;
  assign N1280 = N576 & N582;
  assign N577 = ~shamt_i[5];
  assign N578 = ~shamt_i[4];
  assign N579 = ~shamt_i[3];
  assign N580 = ~shamt_i[2];
  assign N581 = ~shamt_i[0];
  assign N582 = ~shamt_i[1];
  assign N583 = shamt_i[6] & N588;
  assign N584 = N583 & N589;
  assign N585 = N584 & N590;
  assign N586 = N585 & N591;
  assign N587 = N586 & shamt_i[0];
  assign N1281 = N587 & N592;
  assign N588 = ~shamt_i[5];
  assign N589 = ~shamt_i[4];
  assign N590 = ~shamt_i[3];
  assign N591 = ~shamt_i[2];
  assign N592 = ~shamt_i[1];
  assign N593 = shamt_i[6] & N598;
  assign N594 = N593 & N599;
  assign N595 = N594 & N600;
  assign N596 = N595 & N601;
  assign N597 = N596 & N602;
  assign N1282 = N597 & shamt_i[1];
  assign N598 = ~shamt_i[5];
  assign N599 = ~shamt_i[4];
  assign N600 = ~shamt_i[3];
  assign N601 = ~shamt_i[2];
  assign N602 = ~shamt_i[0];
  assign N603 = shamt_i[6] & N608;
  assign N604 = N603 & N609;
  assign N605 = N604 & N610;
  assign N606 = N605 & N611;
  assign N607 = N606 & shamt_i[0];
  assign N1283 = N607 & shamt_i[1];
  assign N608 = ~shamt_i[5];
  assign N609 = ~shamt_i[4];
  assign N610 = ~shamt_i[3];
  assign N611 = ~shamt_i[2];
  assign N612 = shamt_i[6] & N617;
  assign N613 = N612 & N618;
  assign N614 = N613 & N619;
  assign N615 = N614 & shamt_i[2];
  assign N616 = N615 & N620;
  assign N1284 = N616 & N621;
  assign N617 = ~shamt_i[5];
  assign N618 = ~shamt_i[4];
  assign N619 = ~shamt_i[3];
  assign N620 = ~shamt_i[0];
  assign N621 = ~shamt_i[1];
  assign N622 = shamt_i[6] & N627;
  assign N623 = N622 & N628;
  assign N624 = N623 & N629;
  assign N625 = N624 & shamt_i[2];
  assign N626 = N625 & shamt_i[0];
  assign N1285 = N626 & N630;
  assign N627 = ~shamt_i[5];
  assign N628 = ~shamt_i[4];
  assign N629 = ~shamt_i[3];
  assign N630 = ~shamt_i[1];
  assign N631 = shamt_i[6] & N636;
  assign N632 = N631 & N637;
  assign N633 = N632 & N638;
  assign N634 = N633 & shamt_i[2];
  assign N635 = N634 & N639;
  assign N1286 = N635 & shamt_i[1];
  assign N636 = ~shamt_i[5];
  assign N637 = ~shamt_i[4];
  assign N638 = ~shamt_i[3];
  assign N639 = ~shamt_i[0];
  assign N640 = shamt_i[6] & N645;
  assign N641 = N640 & N646;
  assign N642 = N641 & N647;
  assign N643 = N642 & shamt_i[2];
  assign N644 = N643 & shamt_i[0];
  assign N1287 = N644 & shamt_i[1];
  assign N645 = ~shamt_i[5];
  assign N646 = ~shamt_i[4];
  assign N647 = ~shamt_i[3];
  assign N648 = shamt_i[6] & N653;
  assign N649 = N648 & N654;
  assign N650 = N649 & shamt_i[3];
  assign N651 = N650 & N655;
  assign N652 = N651 & N656;
  assign N1288 = N652 & N657;
  assign N653 = ~shamt_i[5];
  assign N654 = ~shamt_i[4];
  assign N655 = ~shamt_i[2];
  assign N656 = ~shamt_i[0];
  assign N657 = ~shamt_i[1];
  assign N658 = shamt_i[6] & N663;
  assign N659 = N658 & N664;
  assign N660 = N659 & shamt_i[3];
  assign N661 = N660 & N665;
  assign N662 = N661 & shamt_i[0];
  assign N1289 = N662 & N666;
  assign N663 = ~shamt_i[5];
  assign N664 = ~shamt_i[4];
  assign N665 = ~shamt_i[2];
  assign N666 = ~shamt_i[1];
  assign N667 = shamt_i[6] & N672;
  assign N668 = N667 & N673;
  assign N669 = N668 & shamt_i[3];
  assign N670 = N669 & N674;
  assign N671 = N670 & N675;
  assign N1290 = N671 & shamt_i[1];
  assign N672 = ~shamt_i[5];
  assign N673 = ~shamt_i[4];
  assign N674 = ~shamt_i[2];
  assign N675 = ~shamt_i[0];
  assign N676 = shamt_i[6] & N681;
  assign N677 = N676 & N682;
  assign N678 = N677 & shamt_i[3];
  assign N679 = N678 & N683;
  assign N680 = N679 & shamt_i[0];
  assign N1291 = N680 & shamt_i[1];
  assign N681 = ~shamt_i[5];
  assign N682 = ~shamt_i[4];
  assign N683 = ~shamt_i[2];
  assign N684 = shamt_i[6] & N689;
  assign N685 = N684 & N690;
  assign N686 = N685 & shamt_i[3];
  assign N687 = N686 & shamt_i[2];
  assign N688 = N687 & N691;
  assign N1292 = N688 & N692;
  assign N689 = ~shamt_i[5];
  assign N690 = ~shamt_i[4];
  assign N691 = ~shamt_i[0];
  assign N692 = ~shamt_i[1];
  assign N693 = shamt_i[6] & N698;
  assign N694 = N693 & N699;
  assign N695 = N694 & shamt_i[3];
  assign N696 = N695 & shamt_i[2];
  assign N697 = N696 & shamt_i[0];
  assign N1293 = N697 & N700;
  assign N698 = ~shamt_i[5];
  assign N699 = ~shamt_i[4];
  assign N700 = ~shamt_i[1];
  assign N701 = shamt_i[6] & N706;
  assign N702 = N701 & N707;
  assign N703 = N702 & shamt_i[3];
  assign N704 = N703 & shamt_i[2];
  assign N705 = N704 & N708;
  assign N1294 = N705 & shamt_i[1];
  assign N706 = ~shamt_i[5];
  assign N707 = ~shamt_i[4];
  assign N708 = ~shamt_i[0];
  assign N709 = shamt_i[6] & N714;
  assign N710 = N709 & N715;
  assign N711 = N710 & shamt_i[3];
  assign N712 = N711 & shamt_i[2];
  assign N713 = N712 & shamt_i[0];
  assign N1295 = N713 & shamt_i[1];
  assign N714 = ~shamt_i[5];
  assign N715 = ~shamt_i[4];
  assign N716 = shamt_i[6] & N721;
  assign N717 = N716 & shamt_i[4];
  assign N718 = N717 & N722;
  assign N719 = N718 & N723;
  assign N720 = N719 & N724;
  assign N1296 = N720 & N725;
  assign N721 = ~shamt_i[5];
  assign N722 = ~shamt_i[3];
  assign N723 = ~shamt_i[2];
  assign N724 = ~shamt_i[0];
  assign N725 = ~shamt_i[1];
  assign N726 = shamt_i[6] & N731;
  assign N727 = N726 & shamt_i[4];
  assign N728 = N727 & N732;
  assign N729 = N728 & N733;
  assign N730 = N729 & shamt_i[0];
  assign N1297 = N730 & N734;
  assign N731 = ~shamt_i[5];
  assign N732 = ~shamt_i[3];
  assign N733 = ~shamt_i[2];
  assign N734 = ~shamt_i[1];
  assign N735 = shamt_i[6] & N740;
  assign N736 = N735 & shamt_i[4];
  assign N737 = N736 & N741;
  assign N738 = N737 & N742;
  assign N739 = N738 & N743;
  assign N1298 = N739 & shamt_i[1];
  assign N740 = ~shamt_i[5];
  assign N741 = ~shamt_i[3];
  assign N742 = ~shamt_i[2];
  assign N743 = ~shamt_i[0];
  assign N744 = shamt_i[6] & N749;
  assign N745 = N744 & shamt_i[4];
  assign N746 = N745 & N750;
  assign N747 = N746 & N751;
  assign N748 = N747 & shamt_i[0];
  assign N1299 = N748 & shamt_i[1];
  assign N749 = ~shamt_i[5];
  assign N750 = ~shamt_i[3];
  assign N751 = ~shamt_i[2];
  assign N752 = shamt_i[6] & N757;
  assign N753 = N752 & shamt_i[4];
  assign N754 = N753 & N758;
  assign N755 = N754 & shamt_i[2];
  assign N756 = N755 & N759;
  assign N1300 = N756 & N760;
  assign N757 = ~shamt_i[5];
  assign N758 = ~shamt_i[3];
  assign N759 = ~shamt_i[0];
  assign N760 = ~shamt_i[1];
  assign N761 = shamt_i[6] & N766;
  assign N762 = N761 & shamt_i[4];
  assign N763 = N762 & N767;
  assign N764 = N763 & shamt_i[2];
  assign N765 = N764 & shamt_i[0];
  assign N1301 = N765 & N768;
  assign N766 = ~shamt_i[5];
  assign N767 = ~shamt_i[3];
  assign N768 = ~shamt_i[1];
  assign N769 = shamt_i[6] & N774;
  assign N770 = N769 & shamt_i[4];
  assign N771 = N770 & N775;
  assign N772 = N771 & shamt_i[2];
  assign N773 = N772 & N776;
  assign N1302 = N773 & shamt_i[1];
  assign N774 = ~shamt_i[5];
  assign N775 = ~shamt_i[3];
  assign N776 = ~shamt_i[0];
  assign N777 = shamt_i[6] & N782;
  assign N778 = N777 & shamt_i[4];
  assign N779 = N778 & N783;
  assign N780 = N779 & shamt_i[2];
  assign N781 = N780 & shamt_i[0];
  assign N1303 = N781 & shamt_i[1];
  assign N782 = ~shamt_i[5];
  assign N783 = ~shamt_i[3];
  assign N784 = shamt_i[6] & N789;
  assign N785 = N784 & shamt_i[4];
  assign N786 = N785 & shamt_i[3];
  assign N787 = N786 & N790;
  assign N788 = N787 & N791;
  assign N1304 = N788 & N792;
  assign N789 = ~shamt_i[5];
  assign N790 = ~shamt_i[2];
  assign N791 = ~shamt_i[0];
  assign N792 = ~shamt_i[1];
  assign N793 = shamt_i[6] & N798;
  assign N794 = N793 & shamt_i[4];
  assign N795 = N794 & shamt_i[3];
  assign N796 = N795 & N799;
  assign N797 = N796 & shamt_i[0];
  assign N1305 = N797 & N800;
  assign N798 = ~shamt_i[5];
  assign N799 = ~shamt_i[2];
  assign N800 = ~shamt_i[1];
  assign N801 = shamt_i[6] & N806;
  assign N802 = N801 & shamt_i[4];
  assign N803 = N802 & shamt_i[3];
  assign N804 = N803 & N807;
  assign N805 = N804 & N808;
  assign N1306 = N805 & shamt_i[1];
  assign N806 = ~shamt_i[5];
  assign N807 = ~shamt_i[2];
  assign N808 = ~shamt_i[0];
  assign N809 = shamt_i[6] & N814;
  assign N810 = N809 & shamt_i[4];
  assign N811 = N810 & shamt_i[3];
  assign N812 = N811 & N815;
  assign N813 = N812 & shamt_i[0];
  assign N1307 = N813 & shamt_i[1];
  assign N814 = ~shamt_i[5];
  assign N815 = ~shamt_i[2];
  assign N816 = shamt_i[6] & N821;
  assign N817 = N816 & shamt_i[4];
  assign N818 = N817 & shamt_i[3];
  assign N819 = N818 & shamt_i[2];
  assign N820 = N819 & N822;
  assign N1308 = N820 & N823;
  assign N821 = ~shamt_i[5];
  assign N822 = ~shamt_i[0];
  assign N823 = ~shamt_i[1];
  assign N824 = shamt_i[6] & N829;
  assign N825 = N824 & shamt_i[4];
  assign N826 = N825 & shamt_i[3];
  assign N827 = N826 & shamt_i[2];
  assign N828 = N827 & shamt_i[0];
  assign N1309 = N828 & N830;
  assign N829 = ~shamt_i[5];
  assign N830 = ~shamt_i[1];
  assign N831 = shamt_i[6] & N836;
  assign N832 = N831 & shamt_i[4];
  assign N833 = N832 & shamt_i[3];
  assign N834 = N833 & shamt_i[2];
  assign N835 = N834 & N837;
  assign N1310 = N835 & shamt_i[1];
  assign N836 = ~shamt_i[5];
  assign N837 = ~shamt_i[0];
  assign N838 = shamt_i[6] & N843;
  assign N839 = N838 & shamt_i[4];
  assign N840 = N839 & shamt_i[3];
  assign N841 = N840 & shamt_i[2];
  assign N842 = N841 & shamt_i[0];
  assign N1311 = N842 & shamt_i[1];
  assign N843 = ~shamt_i[5];
  assign N844 = shamt_i[6] & shamt_i[5];
  assign N845 = N844 & N849;
  assign N846 = N845 & N850;
  assign N847 = N846 & N851;
  assign N848 = N847 & N852;
  assign N1312 = N848 & N853;
  assign N849 = ~shamt_i[4];
  assign N850 = ~shamt_i[3];
  assign N851 = ~shamt_i[2];
  assign N852 = ~shamt_i[0];
  assign N853 = ~shamt_i[1];
  assign N854 = shamt_i[6] & shamt_i[5];
  assign N855 = N854 & N859;
  assign N856 = N855 & N860;
  assign N857 = N856 & N861;
  assign N858 = N857 & shamt_i[0];
  assign N1313 = N858 & N862;
  assign N859 = ~shamt_i[4];
  assign N860 = ~shamt_i[3];
  assign N861 = ~shamt_i[2];
  assign N862 = ~shamt_i[1];
  assign N863 = shamt_i[6] & shamt_i[5];
  assign N864 = N863 & N868;
  assign N865 = N864 & N869;
  assign N866 = N865 & N870;
  assign N867 = N866 & N871;
  assign N1314 = N867 & shamt_i[1];
  assign N868 = ~shamt_i[4];
  assign N869 = ~shamt_i[3];
  assign N870 = ~shamt_i[2];
  assign N871 = ~shamt_i[0];
  assign N872 = shamt_i[6] & shamt_i[5];
  assign N873 = N872 & N877;
  assign N874 = N873 & N878;
  assign N875 = N874 & N879;
  assign N876 = N875 & shamt_i[0];
  assign N1315 = N876 & shamt_i[1];
  assign N877 = ~shamt_i[4];
  assign N878 = ~shamt_i[3];
  assign N879 = ~shamt_i[2];
  assign N880 = shamt_i[6] & shamt_i[5];
  assign N881 = N880 & N885;
  assign N882 = N881 & N886;
  assign N883 = N882 & shamt_i[2];
  assign N884 = N883 & N887;
  assign N1316 = N884 & N888;
  assign N885 = ~shamt_i[4];
  assign N886 = ~shamt_i[3];
  assign N887 = ~shamt_i[0];
  assign N888 = ~shamt_i[1];
  assign N889 = shamt_i[6] & shamt_i[5];
  assign N890 = N889 & N894;
  assign N891 = N890 & N895;
  assign N892 = N891 & shamt_i[2];
  assign N893 = N892 & shamt_i[0];
  assign N1317 = N893 & N896;
  assign N894 = ~shamt_i[4];
  assign N895 = ~shamt_i[3];
  assign N896 = ~shamt_i[1];
  assign N897 = shamt_i[6] & shamt_i[5];
  assign N898 = N897 & N902;
  assign N899 = N898 & N903;
  assign N900 = N899 & shamt_i[2];
  assign N901 = N900 & N904;
  assign N1318 = N901 & shamt_i[1];
  assign N902 = ~shamt_i[4];
  assign N903 = ~shamt_i[3];
  assign N904 = ~shamt_i[0];
  assign N905 = shamt_i[6] & shamt_i[5];
  assign N906 = N905 & N910;
  assign N907 = N906 & N911;
  assign N908 = N907 & shamt_i[2];
  assign N909 = N908 & shamt_i[0];
  assign N1319 = N909 & shamt_i[1];
  assign N910 = ~shamt_i[4];
  assign N911 = ~shamt_i[3];
  assign N912 = shamt_i[6] & shamt_i[5];
  assign N913 = N912 & N917;
  assign N914 = N913 & shamt_i[3];
  assign N915 = N914 & N918;
  assign N916 = N915 & N919;
  assign N1320 = N916 & N920;
  assign N917 = ~shamt_i[4];
  assign N918 = ~shamt_i[2];
  assign N919 = ~shamt_i[0];
  assign N920 = ~shamt_i[1];
  assign N921 = shamt_i[6] & shamt_i[5];
  assign N922 = N921 & N926;
  assign N923 = N922 & shamt_i[3];
  assign N924 = N923 & N927;
  assign N925 = N924 & shamt_i[0];
  assign N1321 = N925 & N928;
  assign N926 = ~shamt_i[4];
  assign N927 = ~shamt_i[2];
  assign N928 = ~shamt_i[1];
  assign N929 = shamt_i[6] & shamt_i[5];
  assign N930 = N929 & N934;
  assign N931 = N930 & shamt_i[3];
  assign N932 = N931 & N935;
  assign N933 = N932 & N936;
  assign N1322 = N933 & shamt_i[1];
  assign N934 = ~shamt_i[4];
  assign N935 = ~shamt_i[2];
  assign N936 = ~shamt_i[0];
  assign N937 = shamt_i[6] & shamt_i[5];
  assign N938 = N937 & N942;
  assign N939 = N938 & shamt_i[3];
  assign N940 = N939 & N943;
  assign N941 = N940 & shamt_i[0];
  assign N1323 = N941 & shamt_i[1];
  assign N942 = ~shamt_i[4];
  assign N943 = ~shamt_i[2];
  assign N944 = shamt_i[6] & shamt_i[5];
  assign N945 = N944 & N949;
  assign N946 = N945 & shamt_i[3];
  assign N947 = N946 & shamt_i[2];
  assign N948 = N947 & N950;
  assign N1324 = N948 & N951;
  assign N949 = ~shamt_i[4];
  assign N950 = ~shamt_i[0];
  assign N951 = ~shamt_i[1];
  assign N952 = shamt_i[6] & shamt_i[5];
  assign N953 = N952 & N957;
  assign N954 = N953 & shamt_i[3];
  assign N955 = N954 & shamt_i[2];
  assign N956 = N955 & shamt_i[0];
  assign N1325 = N956 & N958;
  assign N957 = ~shamt_i[4];
  assign N958 = ~shamt_i[1];
  assign N959 = shamt_i[6] & shamt_i[5];
  assign N960 = N959 & N964;
  assign N961 = N960 & shamt_i[3];
  assign N962 = N961 & shamt_i[2];
  assign N963 = N962 & N965;
  assign N1326 = N963 & shamt_i[1];
  assign N964 = ~shamt_i[4];
  assign N965 = ~shamt_i[0];
  assign N966 = shamt_i[6] & shamt_i[5];
  assign N967 = N966 & N971;
  assign N968 = N967 & shamt_i[3];
  assign N969 = N968 & shamt_i[2];
  assign N970 = N969 & shamt_i[0];
  assign N1327 = N970 & shamt_i[1];
  assign N971 = ~shamt_i[4];
  assign N972 = shamt_i[6] & shamt_i[5];
  assign N973 = N972 & shamt_i[4];
  assign N974 = N973 & N977;
  assign N975 = N974 & N978;
  assign N976 = N975 & N979;
  assign N1328 = N976 & N980;
  assign N977 = ~shamt_i[3];
  assign N978 = ~shamt_i[2];
  assign N979 = ~shamt_i[0];
  assign N980 = ~shamt_i[1];
  assign N981 = shamt_i[6] & shamt_i[5];
  assign N982 = N981 & shamt_i[4];
  assign N983 = N982 & N986;
  assign N984 = N983 & N987;
  assign N985 = N984 & shamt_i[0];
  assign N1329 = N985 & N988;
  assign N986 = ~shamt_i[3];
  assign N987 = ~shamt_i[2];
  assign N988 = ~shamt_i[1];
  assign N989 = shamt_i[6] & shamt_i[5];
  assign N990 = N989 & shamt_i[4];
  assign N991 = N990 & N994;
  assign N992 = N991 & N995;
  assign N993 = N992 & N996;
  assign N1330 = N993 & shamt_i[1];
  assign N994 = ~shamt_i[3];
  assign N995 = ~shamt_i[2];
  assign N996 = ~shamt_i[0];
  assign N997 = shamt_i[6] & shamt_i[5];
  assign N998 = N997 & shamt_i[4];
  assign N999 = N998 & N1002;
  assign N1000 = N999 & N1003;
  assign N1001 = N1000 & shamt_i[0];
  assign N1331 = N1001 & shamt_i[1];
  assign N1002 = ~shamt_i[3];
  assign N1003 = ~shamt_i[2];
  assign N1004 = shamt_i[6] & shamt_i[5];
  assign N1005 = N1004 & shamt_i[4];
  assign N1006 = N1005 & N1009;
  assign N1007 = N1006 & shamt_i[2];
  assign N1008 = N1007 & N1010;
  assign N1332 = N1008 & N1011;
  assign N1009 = ~shamt_i[3];
  assign N1010 = ~shamt_i[0];
  assign N1011 = ~shamt_i[1];
  assign N1012 = shamt_i[6] & shamt_i[5];
  assign N1013 = N1012 & shamt_i[4];
  assign N1014 = N1013 & N1017;
  assign N1015 = N1014 & shamt_i[2];
  assign N1016 = N1015 & shamt_i[0];
  assign N1333 = N1016 & N1018;
  assign N1017 = ~shamt_i[3];
  assign N1018 = ~shamt_i[1];
  assign N1019 = shamt_i[6] & shamt_i[5];
  assign N1020 = N1019 & shamt_i[4];
  assign N1021 = N1020 & N1024;
  assign N1022 = N1021 & shamt_i[2];
  assign N1023 = N1022 & N1025;
  assign N1334 = N1023 & shamt_i[1];
  assign N1024 = ~shamt_i[3];
  assign N1025 = ~shamt_i[0];
  assign N1026 = shamt_i[6] & shamt_i[5];
  assign N1027 = N1026 & shamt_i[4];
  assign N1028 = N1027 & N1031;
  assign N1029 = N1028 & shamt_i[2];
  assign N1030 = N1029 & shamt_i[0];
  assign N1335 = N1030 & shamt_i[1];
  assign N1031 = ~shamt_i[3];
  assign N1032 = shamt_i[6] & shamt_i[5];
  assign N1033 = N1032 & shamt_i[4];
  assign N1034 = N1033 & shamt_i[3];
  assign N1035 = N1034 & N1037;
  assign N1036 = N1035 & N1038;
  assign N1336 = N1036 & N1039;
  assign N1037 = ~shamt_i[2];
  assign N1038 = ~shamt_i[0];
  assign N1039 = ~shamt_i[1];
  assign N1040 = shamt_i[6] & shamt_i[5];
  assign N1041 = N1040 & shamt_i[4];
  assign N1042 = N1041 & shamt_i[3];
  assign N1043 = N1042 & N1045;
  assign N1044 = N1043 & shamt_i[0];
  assign N1337 = N1044 & N1046;
  assign N1045 = ~shamt_i[2];
  assign N1046 = ~shamt_i[1];
  assign N1047 = shamt_i[6] & shamt_i[5];
  assign N1048 = N1047 & shamt_i[4];
  assign N1049 = N1048 & shamt_i[3];
  assign N1050 = N1049 & N1052;
  assign N1051 = N1050 & N1053;
  assign N1338 = N1051 & shamt_i[1];
  assign N1052 = ~shamt_i[2];
  assign N1053 = ~shamt_i[0];
  assign N1054 = shamt_i[6] & shamt_i[5];
  assign N1055 = N1054 & shamt_i[4];
  assign N1056 = N1055 & shamt_i[3];
  assign N1057 = N1056 & N1059;
  assign N1058 = N1057 & shamt_i[0];
  assign N1339 = N1058 & shamt_i[1];
  assign N1059 = ~shamt_i[2];
  assign N1060 = shamt_i[6] & shamt_i[5];
  assign N1061 = N1060 & shamt_i[4];
  assign N1062 = N1061 & shamt_i[3];
  assign N1063 = N1062 & shamt_i[2];
  assign N1064 = N1063 & N1065;
  assign N1340 = N1064 & N1066;
  assign N1065 = ~shamt_i[0];
  assign N1066 = ~shamt_i[1];
  assign N1067 = shamt_i[6] & shamt_i[5];
  assign N1068 = N1067 & shamt_i[4];
  assign N1069 = N1068 & shamt_i[3];
  assign N1070 = N1069 & shamt_i[2];
  assign N1071 = N1070 & shamt_i[0];
  assign N1341 = N1071 & N1072;
  assign N1072 = ~shamt_i[1];
  assign N1073 = shamt_i[6] & shamt_i[5];
  assign N1074 = N1073 & shamt_i[4];
  assign N1075 = N1074 & shamt_i[3];
  assign N1076 = N1075 & shamt_i[2];
  assign N1077 = N1076 & N1078;
  assign N1342 = N1077 & shamt_i[1];
  assign N1078 = ~shamt_i[0];
  assign N1079 = shamt_i[6] & shamt_i[5];
  assign N1080 = N1079 & shamt_i[4];
  assign N1081 = N1080 & shamt_i[3];
  assign N1082 = N1081 & shamt_i[2];
  assign N1083 = N1082 & shamt_i[0];
  assign N1343 = N1083 & shamt_i[1];
  assign sticky_o = (N1084)? scan_out[127] : 
                    (N1215)? N1344 : 1'b0;
  assign N1084 = N1214;
  assign N1344 = (N1085)? 1'b0 : 
                 (N1086)? scan_out[0] : 
                 (N1087)? scan_out[1] : 
                 (N1088)? scan_out[2] : 
                 (N1089)? scan_out[3] : 
                 (N1090)? scan_out[4] : 
                 (N1091)? scan_out[5] : 
                 (N1092)? scan_out[6] : 
                 (N1093)? scan_out[7] : 
                 (N1094)? scan_out[8] : 
                 (N1095)? scan_out[9] : 
                 (N1096)? scan_out[10] : 
                 (N1097)? scan_out[11] : 
                 (N1098)? scan_out[12] : 
                 (N1099)? scan_out[13] : 
                 (N1100)? scan_out[14] : 
                 (N1101)? scan_out[15] : 
                 (N1102)? scan_out[16] : 
                 (N1103)? scan_out[17] : 
                 (N1104)? scan_out[18] : 
                 (N1105)? scan_out[19] : 
                 (N1106)? scan_out[20] : 
                 (N1107)? scan_out[21] : 
                 (N1108)? scan_out[22] : 
                 (N1109)? scan_out[23] : 
                 (N1110)? scan_out[24] : 
                 (N1111)? scan_out[25] : 
                 (N1112)? scan_out[26] : 
                 (N1113)? scan_out[27] : 
                 (N1114)? scan_out[28] : 
                 (N1115)? scan_out[29] : 
                 (N1116)? scan_out[30] : 
                 (N1117)? scan_out[31] : 
                 (N1118)? scan_out[32] : 
                 (N1119)? scan_out[33] : 
                 (N1120)? scan_out[34] : 
                 (N1121)? scan_out[35] : 
                 (N1122)? scan_out[36] : 
                 (N1123)? scan_out[37] : 
                 (N1124)? scan_out[38] : 
                 (N1125)? scan_out[39] : 
                 (N1126)? scan_out[40] : 
                 (N1127)? scan_out[41] : 
                 (N1128)? scan_out[42] : 
                 (N1129)? scan_out[43] : 
                 (N1130)? scan_out[44] : 
                 (N1131)? scan_out[45] : 
                 (N1132)? scan_out[46] : 
                 (N1133)? scan_out[47] : 
                 (N1134)? scan_out[48] : 
                 (N1135)? scan_out[49] : 
                 (N1136)? scan_out[50] : 
                 (N1137)? scan_out[51] : 
                 (N1138)? scan_out[52] : 
                 (N1139)? scan_out[53] : 
                 (N1140)? scan_out[54] : 
                 (N1141)? scan_out[55] : 
                 (N1142)? scan_out[56] : 
                 (N1143)? scan_out[57] : 
                 (N1144)? scan_out[58] : 
                 (N1145)? scan_out[59] : 
                 (N1146)? scan_out[60] : 
                 (N1147)? scan_out[61] : 
                 (N1148)? scan_out[62] : 
                 (N1149)? scan_out[63] : 
                 (N1150)? scan_out[64] : 
                 (N1151)? scan_out[65] : 
                 (N1152)? scan_out[66] : 
                 (N1153)? scan_out[67] : 
                 (N1154)? scan_out[68] : 
                 (N1155)? scan_out[69] : 
                 (N1156)? scan_out[70] : 
                 (N1157)? scan_out[71] : 
                 (N1158)? scan_out[72] : 
                 (N1159)? scan_out[73] : 
                 (N1160)? scan_out[74] : 
                 (N1161)? scan_out[75] : 
                 (N1162)? scan_out[76] : 
                 (N1163)? scan_out[77] : 
                 (N1164)? scan_out[78] : 
                 (N1165)? scan_out[79] : 
                 (N1166)? scan_out[80] : 
                 (N1167)? scan_out[81] : 
                 (N1168)? scan_out[82] : 
                 (N1169)? scan_out[83] : 
                 (N1170)? scan_out[84] : 
                 (N1171)? scan_out[85] : 
                 (N1172)? scan_out[86] : 
                 (N1173)? scan_out[87] : 
                 (N1174)? scan_out[88] : 
                 (N1175)? scan_out[89] : 
                 (N1176)? scan_out[90] : 
                 (N1177)? scan_out[91] : 
                 (N1178)? scan_out[92] : 
                 (N1179)? scan_out[93] : 
                 (N1180)? scan_out[94] : 
                 (N1181)? scan_out[95] : 
                 (N1182)? scan_out[96] : 
                 (N1183)? scan_out[97] : 
                 (N1184)? scan_out[98] : 
                 (N1185)? scan_out[99] : 
                 (N1186)? scan_out[100] : 
                 (N1187)? scan_out[101] : 
                 (N1188)? scan_out[102] : 
                 (N1189)? scan_out[103] : 
                 (N1190)? scan_out[104] : 
                 (N1191)? scan_out[105] : 
                 (N1192)? scan_out[106] : 
                 (N1193)? scan_out[107] : 
                 (N1194)? scan_out[108] : 
                 (N1195)? scan_out[109] : 
                 (N1196)? scan_out[110] : 
                 (N1197)? scan_out[111] : 
                 (N1198)? scan_out[112] : 
                 (N1199)? scan_out[113] : 
                 (N1200)? scan_out[114] : 
                 (N1201)? scan_out[115] : 
                 (N1202)? scan_out[116] : 
                 (N1203)? scan_out[117] : 
                 (N1204)? scan_out[118] : 
                 (N1205)? scan_out[119] : 
                 (N1206)? scan_out[120] : 
                 (N1207)? scan_out[121] : 
                 (N1208)? scan_out[122] : 
                 (N1209)? scan_out[123] : 
                 (N1210)? scan_out[124] : 
                 (N1211)? scan_out[125] : 
                 (N1212)? scan_out[126] : 
                 (N1213)? scan_out[127] : 1'b0;
  assign N1085 = N1216;
  assign N1086 = N1217;
  assign N1087 = N1218;
  assign N1088 = N1219;
  assign N1089 = N1220;
  assign N1090 = N1221;
  assign N1091 = N1222;
  assign N1092 = N1223;
  assign N1093 = N1224;
  assign N1094 = N1225;
  assign N1095 = N1226;
  assign N1096 = N1227;
  assign N1097 = N1228;
  assign N1098 = N1229;
  assign N1099 = N1230;
  assign N1100 = N1231;
  assign N1101 = N1232;
  assign N1102 = N1233;
  assign N1103 = N1234;
  assign N1104 = N1235;
  assign N1105 = N1236;
  assign N1106 = N1237;
  assign N1107 = N1238;
  assign N1108 = N1239;
  assign N1109 = N1240;
  assign N1110 = N1241;
  assign N1111 = N1242;
  assign N1112 = N1243;
  assign N1113 = N1244;
  assign N1114 = N1245;
  assign N1115 = N1246;
  assign N1116 = N1247;
  assign N1117 = N1248;
  assign N1118 = N1249;
  assign N1119 = N1250;
  assign N1120 = N1251;
  assign N1121 = N1252;
  assign N1122 = N1253;
  assign N1123 = N1254;
  assign N1124 = N1255;
  assign N1125 = N1256;
  assign N1126 = N1257;
  assign N1127 = N1258;
  assign N1128 = N1259;
  assign N1129 = N1260;
  assign N1130 = N1261;
  assign N1131 = N1262;
  assign N1132 = N1263;
  assign N1133 = N1264;
  assign N1134 = N1265;
  assign N1135 = N1266;
  assign N1136 = N1267;
  assign N1137 = N1268;
  assign N1138 = N1269;
  assign N1139 = N1270;
  assign N1140 = N1271;
  assign N1141 = N1272;
  assign N1142 = N1273;
  assign N1143 = N1274;
  assign N1144 = N1275;
  assign N1145 = N1276;
  assign N1146 = N1277;
  assign N1147 = N1278;
  assign N1148 = N1279;
  assign N1149 = N1280;
  assign N1150 = N1281;
  assign N1151 = N1282;
  assign N1152 = N1283;
  assign N1153 = N1284;
  assign N1154 = N1285;
  assign N1155 = N1286;
  assign N1156 = N1287;
  assign N1157 = N1288;
  assign N1158 = N1289;
  assign N1159 = N1290;
  assign N1160 = N1291;
  assign N1161 = N1292;
  assign N1162 = N1293;
  assign N1163 = N1294;
  assign N1164 = N1295;
  assign N1165 = N1296;
  assign N1166 = N1297;
  assign N1167 = N1298;
  assign N1168 = N1299;
  assign N1169 = N1300;
  assign N1170 = N1301;
  assign N1171 = N1302;
  assign N1172 = N1303;
  assign N1173 = N1304;
  assign N1174 = N1305;
  assign N1175 = N1306;
  assign N1176 = N1307;
  assign N1177 = N1308;
  assign N1178 = N1309;
  assign N1179 = N1310;
  assign N1180 = N1311;
  assign N1181 = N1312;
  assign N1182 = N1313;
  assign N1183 = N1314;
  assign N1184 = N1315;
  assign N1185 = N1316;
  assign N1186 = N1317;
  assign N1187 = N1318;
  assign N1188 = N1319;
  assign N1189 = N1320;
  assign N1190 = N1321;
  assign N1191 = N1322;
  assign N1192 = N1323;
  assign N1193 = N1324;
  assign N1194 = N1325;
  assign N1195 = N1326;
  assign N1196 = N1327;
  assign N1197 = N1328;
  assign N1198 = N1329;
  assign N1199 = N1330;
  assign N1200 = N1331;
  assign N1201 = N1332;
  assign N1202 = N1333;
  assign N1203 = N1334;
  assign N1204 = N1335;
  assign N1205 = N1336;
  assign N1206 = N1337;
  assign N1207 = N1338;
  assign N1208 = N1339;
  assign N1209 = N1340;
  assign N1210 = N1341;
  assign N1211 = N1342;
  assign N1212 = N1343;
  assign N1213 = shamt_i[7];
  assign N1215 = ~N1214;

endmodule

