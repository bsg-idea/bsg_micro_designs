

module top
(
  i,
  o
);

  input [63:0] i;
  output [16383:0] o;

  bsg_expand_bitmask
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_expand_bitmask
(
  i,
  o
);

  input [63:0] i;
  output [16383:0] o;
  wire [16383:0] o;
  assign o[16128] = i[63];
  assign o[16129] = i[63];
  assign o[16130] = i[63];
  assign o[16131] = i[63];
  assign o[16132] = i[63];
  assign o[16133] = i[63];
  assign o[16134] = i[63];
  assign o[16135] = i[63];
  assign o[16136] = i[63];
  assign o[16137] = i[63];
  assign o[16138] = i[63];
  assign o[16139] = i[63];
  assign o[16140] = i[63];
  assign o[16141] = i[63];
  assign o[16142] = i[63];
  assign o[16143] = i[63];
  assign o[16144] = i[63];
  assign o[16145] = i[63];
  assign o[16146] = i[63];
  assign o[16147] = i[63];
  assign o[16148] = i[63];
  assign o[16149] = i[63];
  assign o[16150] = i[63];
  assign o[16151] = i[63];
  assign o[16152] = i[63];
  assign o[16153] = i[63];
  assign o[16154] = i[63];
  assign o[16155] = i[63];
  assign o[16156] = i[63];
  assign o[16157] = i[63];
  assign o[16158] = i[63];
  assign o[16159] = i[63];
  assign o[16160] = i[63];
  assign o[16161] = i[63];
  assign o[16162] = i[63];
  assign o[16163] = i[63];
  assign o[16164] = i[63];
  assign o[16165] = i[63];
  assign o[16166] = i[63];
  assign o[16167] = i[63];
  assign o[16168] = i[63];
  assign o[16169] = i[63];
  assign o[16170] = i[63];
  assign o[16171] = i[63];
  assign o[16172] = i[63];
  assign o[16173] = i[63];
  assign o[16174] = i[63];
  assign o[16175] = i[63];
  assign o[16176] = i[63];
  assign o[16177] = i[63];
  assign o[16178] = i[63];
  assign o[16179] = i[63];
  assign o[16180] = i[63];
  assign o[16181] = i[63];
  assign o[16182] = i[63];
  assign o[16183] = i[63];
  assign o[16184] = i[63];
  assign o[16185] = i[63];
  assign o[16186] = i[63];
  assign o[16187] = i[63];
  assign o[16188] = i[63];
  assign o[16189] = i[63];
  assign o[16190] = i[63];
  assign o[16191] = i[63];
  assign o[16192] = i[63];
  assign o[16193] = i[63];
  assign o[16194] = i[63];
  assign o[16195] = i[63];
  assign o[16196] = i[63];
  assign o[16197] = i[63];
  assign o[16198] = i[63];
  assign o[16199] = i[63];
  assign o[16200] = i[63];
  assign o[16201] = i[63];
  assign o[16202] = i[63];
  assign o[16203] = i[63];
  assign o[16204] = i[63];
  assign o[16205] = i[63];
  assign o[16206] = i[63];
  assign o[16207] = i[63];
  assign o[16208] = i[63];
  assign o[16209] = i[63];
  assign o[16210] = i[63];
  assign o[16211] = i[63];
  assign o[16212] = i[63];
  assign o[16213] = i[63];
  assign o[16214] = i[63];
  assign o[16215] = i[63];
  assign o[16216] = i[63];
  assign o[16217] = i[63];
  assign o[16218] = i[63];
  assign o[16219] = i[63];
  assign o[16220] = i[63];
  assign o[16221] = i[63];
  assign o[16222] = i[63];
  assign o[16223] = i[63];
  assign o[16224] = i[63];
  assign o[16225] = i[63];
  assign o[16226] = i[63];
  assign o[16227] = i[63];
  assign o[16228] = i[63];
  assign o[16229] = i[63];
  assign o[16230] = i[63];
  assign o[16231] = i[63];
  assign o[16232] = i[63];
  assign o[16233] = i[63];
  assign o[16234] = i[63];
  assign o[16235] = i[63];
  assign o[16236] = i[63];
  assign o[16237] = i[63];
  assign o[16238] = i[63];
  assign o[16239] = i[63];
  assign o[16240] = i[63];
  assign o[16241] = i[63];
  assign o[16242] = i[63];
  assign o[16243] = i[63];
  assign o[16244] = i[63];
  assign o[16245] = i[63];
  assign o[16246] = i[63];
  assign o[16247] = i[63];
  assign o[16248] = i[63];
  assign o[16249] = i[63];
  assign o[16250] = i[63];
  assign o[16251] = i[63];
  assign o[16252] = i[63];
  assign o[16253] = i[63];
  assign o[16254] = i[63];
  assign o[16255] = i[63];
  assign o[16256] = i[63];
  assign o[16257] = i[63];
  assign o[16258] = i[63];
  assign o[16259] = i[63];
  assign o[16260] = i[63];
  assign o[16261] = i[63];
  assign o[16262] = i[63];
  assign o[16263] = i[63];
  assign o[16264] = i[63];
  assign o[16265] = i[63];
  assign o[16266] = i[63];
  assign o[16267] = i[63];
  assign o[16268] = i[63];
  assign o[16269] = i[63];
  assign o[16270] = i[63];
  assign o[16271] = i[63];
  assign o[16272] = i[63];
  assign o[16273] = i[63];
  assign o[16274] = i[63];
  assign o[16275] = i[63];
  assign o[16276] = i[63];
  assign o[16277] = i[63];
  assign o[16278] = i[63];
  assign o[16279] = i[63];
  assign o[16280] = i[63];
  assign o[16281] = i[63];
  assign o[16282] = i[63];
  assign o[16283] = i[63];
  assign o[16284] = i[63];
  assign o[16285] = i[63];
  assign o[16286] = i[63];
  assign o[16287] = i[63];
  assign o[16288] = i[63];
  assign o[16289] = i[63];
  assign o[16290] = i[63];
  assign o[16291] = i[63];
  assign o[16292] = i[63];
  assign o[16293] = i[63];
  assign o[16294] = i[63];
  assign o[16295] = i[63];
  assign o[16296] = i[63];
  assign o[16297] = i[63];
  assign o[16298] = i[63];
  assign o[16299] = i[63];
  assign o[16300] = i[63];
  assign o[16301] = i[63];
  assign o[16302] = i[63];
  assign o[16303] = i[63];
  assign o[16304] = i[63];
  assign o[16305] = i[63];
  assign o[16306] = i[63];
  assign o[16307] = i[63];
  assign o[16308] = i[63];
  assign o[16309] = i[63];
  assign o[16310] = i[63];
  assign o[16311] = i[63];
  assign o[16312] = i[63];
  assign o[16313] = i[63];
  assign o[16314] = i[63];
  assign o[16315] = i[63];
  assign o[16316] = i[63];
  assign o[16317] = i[63];
  assign o[16318] = i[63];
  assign o[16319] = i[63];
  assign o[16320] = i[63];
  assign o[16321] = i[63];
  assign o[16322] = i[63];
  assign o[16323] = i[63];
  assign o[16324] = i[63];
  assign o[16325] = i[63];
  assign o[16326] = i[63];
  assign o[16327] = i[63];
  assign o[16328] = i[63];
  assign o[16329] = i[63];
  assign o[16330] = i[63];
  assign o[16331] = i[63];
  assign o[16332] = i[63];
  assign o[16333] = i[63];
  assign o[16334] = i[63];
  assign o[16335] = i[63];
  assign o[16336] = i[63];
  assign o[16337] = i[63];
  assign o[16338] = i[63];
  assign o[16339] = i[63];
  assign o[16340] = i[63];
  assign o[16341] = i[63];
  assign o[16342] = i[63];
  assign o[16343] = i[63];
  assign o[16344] = i[63];
  assign o[16345] = i[63];
  assign o[16346] = i[63];
  assign o[16347] = i[63];
  assign o[16348] = i[63];
  assign o[16349] = i[63];
  assign o[16350] = i[63];
  assign o[16351] = i[63];
  assign o[16352] = i[63];
  assign o[16353] = i[63];
  assign o[16354] = i[63];
  assign o[16355] = i[63];
  assign o[16356] = i[63];
  assign o[16357] = i[63];
  assign o[16358] = i[63];
  assign o[16359] = i[63];
  assign o[16360] = i[63];
  assign o[16361] = i[63];
  assign o[16362] = i[63];
  assign o[16363] = i[63];
  assign o[16364] = i[63];
  assign o[16365] = i[63];
  assign o[16366] = i[63];
  assign o[16367] = i[63];
  assign o[16368] = i[63];
  assign o[16369] = i[63];
  assign o[16370] = i[63];
  assign o[16371] = i[63];
  assign o[16372] = i[63];
  assign o[16373] = i[63];
  assign o[16374] = i[63];
  assign o[16375] = i[63];
  assign o[16376] = i[63];
  assign o[16377] = i[63];
  assign o[16378] = i[63];
  assign o[16379] = i[63];
  assign o[16380] = i[63];
  assign o[16381] = i[63];
  assign o[16382] = i[63];
  assign o[16383] = i[63];
  assign o[15872] = i[62];
  assign o[15873] = i[62];
  assign o[15874] = i[62];
  assign o[15875] = i[62];
  assign o[15876] = i[62];
  assign o[15877] = i[62];
  assign o[15878] = i[62];
  assign o[15879] = i[62];
  assign o[15880] = i[62];
  assign o[15881] = i[62];
  assign o[15882] = i[62];
  assign o[15883] = i[62];
  assign o[15884] = i[62];
  assign o[15885] = i[62];
  assign o[15886] = i[62];
  assign o[15887] = i[62];
  assign o[15888] = i[62];
  assign o[15889] = i[62];
  assign o[15890] = i[62];
  assign o[15891] = i[62];
  assign o[15892] = i[62];
  assign o[15893] = i[62];
  assign o[15894] = i[62];
  assign o[15895] = i[62];
  assign o[15896] = i[62];
  assign o[15897] = i[62];
  assign o[15898] = i[62];
  assign o[15899] = i[62];
  assign o[15900] = i[62];
  assign o[15901] = i[62];
  assign o[15902] = i[62];
  assign o[15903] = i[62];
  assign o[15904] = i[62];
  assign o[15905] = i[62];
  assign o[15906] = i[62];
  assign o[15907] = i[62];
  assign o[15908] = i[62];
  assign o[15909] = i[62];
  assign o[15910] = i[62];
  assign o[15911] = i[62];
  assign o[15912] = i[62];
  assign o[15913] = i[62];
  assign o[15914] = i[62];
  assign o[15915] = i[62];
  assign o[15916] = i[62];
  assign o[15917] = i[62];
  assign o[15918] = i[62];
  assign o[15919] = i[62];
  assign o[15920] = i[62];
  assign o[15921] = i[62];
  assign o[15922] = i[62];
  assign o[15923] = i[62];
  assign o[15924] = i[62];
  assign o[15925] = i[62];
  assign o[15926] = i[62];
  assign o[15927] = i[62];
  assign o[15928] = i[62];
  assign o[15929] = i[62];
  assign o[15930] = i[62];
  assign o[15931] = i[62];
  assign o[15932] = i[62];
  assign o[15933] = i[62];
  assign o[15934] = i[62];
  assign o[15935] = i[62];
  assign o[15936] = i[62];
  assign o[15937] = i[62];
  assign o[15938] = i[62];
  assign o[15939] = i[62];
  assign o[15940] = i[62];
  assign o[15941] = i[62];
  assign o[15942] = i[62];
  assign o[15943] = i[62];
  assign o[15944] = i[62];
  assign o[15945] = i[62];
  assign o[15946] = i[62];
  assign o[15947] = i[62];
  assign o[15948] = i[62];
  assign o[15949] = i[62];
  assign o[15950] = i[62];
  assign o[15951] = i[62];
  assign o[15952] = i[62];
  assign o[15953] = i[62];
  assign o[15954] = i[62];
  assign o[15955] = i[62];
  assign o[15956] = i[62];
  assign o[15957] = i[62];
  assign o[15958] = i[62];
  assign o[15959] = i[62];
  assign o[15960] = i[62];
  assign o[15961] = i[62];
  assign o[15962] = i[62];
  assign o[15963] = i[62];
  assign o[15964] = i[62];
  assign o[15965] = i[62];
  assign o[15966] = i[62];
  assign o[15967] = i[62];
  assign o[15968] = i[62];
  assign o[15969] = i[62];
  assign o[15970] = i[62];
  assign o[15971] = i[62];
  assign o[15972] = i[62];
  assign o[15973] = i[62];
  assign o[15974] = i[62];
  assign o[15975] = i[62];
  assign o[15976] = i[62];
  assign o[15977] = i[62];
  assign o[15978] = i[62];
  assign o[15979] = i[62];
  assign o[15980] = i[62];
  assign o[15981] = i[62];
  assign o[15982] = i[62];
  assign o[15983] = i[62];
  assign o[15984] = i[62];
  assign o[15985] = i[62];
  assign o[15986] = i[62];
  assign o[15987] = i[62];
  assign o[15988] = i[62];
  assign o[15989] = i[62];
  assign o[15990] = i[62];
  assign o[15991] = i[62];
  assign o[15992] = i[62];
  assign o[15993] = i[62];
  assign o[15994] = i[62];
  assign o[15995] = i[62];
  assign o[15996] = i[62];
  assign o[15997] = i[62];
  assign o[15998] = i[62];
  assign o[15999] = i[62];
  assign o[16000] = i[62];
  assign o[16001] = i[62];
  assign o[16002] = i[62];
  assign o[16003] = i[62];
  assign o[16004] = i[62];
  assign o[16005] = i[62];
  assign o[16006] = i[62];
  assign o[16007] = i[62];
  assign o[16008] = i[62];
  assign o[16009] = i[62];
  assign o[16010] = i[62];
  assign o[16011] = i[62];
  assign o[16012] = i[62];
  assign o[16013] = i[62];
  assign o[16014] = i[62];
  assign o[16015] = i[62];
  assign o[16016] = i[62];
  assign o[16017] = i[62];
  assign o[16018] = i[62];
  assign o[16019] = i[62];
  assign o[16020] = i[62];
  assign o[16021] = i[62];
  assign o[16022] = i[62];
  assign o[16023] = i[62];
  assign o[16024] = i[62];
  assign o[16025] = i[62];
  assign o[16026] = i[62];
  assign o[16027] = i[62];
  assign o[16028] = i[62];
  assign o[16029] = i[62];
  assign o[16030] = i[62];
  assign o[16031] = i[62];
  assign o[16032] = i[62];
  assign o[16033] = i[62];
  assign o[16034] = i[62];
  assign o[16035] = i[62];
  assign o[16036] = i[62];
  assign o[16037] = i[62];
  assign o[16038] = i[62];
  assign o[16039] = i[62];
  assign o[16040] = i[62];
  assign o[16041] = i[62];
  assign o[16042] = i[62];
  assign o[16043] = i[62];
  assign o[16044] = i[62];
  assign o[16045] = i[62];
  assign o[16046] = i[62];
  assign o[16047] = i[62];
  assign o[16048] = i[62];
  assign o[16049] = i[62];
  assign o[16050] = i[62];
  assign o[16051] = i[62];
  assign o[16052] = i[62];
  assign o[16053] = i[62];
  assign o[16054] = i[62];
  assign o[16055] = i[62];
  assign o[16056] = i[62];
  assign o[16057] = i[62];
  assign o[16058] = i[62];
  assign o[16059] = i[62];
  assign o[16060] = i[62];
  assign o[16061] = i[62];
  assign o[16062] = i[62];
  assign o[16063] = i[62];
  assign o[16064] = i[62];
  assign o[16065] = i[62];
  assign o[16066] = i[62];
  assign o[16067] = i[62];
  assign o[16068] = i[62];
  assign o[16069] = i[62];
  assign o[16070] = i[62];
  assign o[16071] = i[62];
  assign o[16072] = i[62];
  assign o[16073] = i[62];
  assign o[16074] = i[62];
  assign o[16075] = i[62];
  assign o[16076] = i[62];
  assign o[16077] = i[62];
  assign o[16078] = i[62];
  assign o[16079] = i[62];
  assign o[16080] = i[62];
  assign o[16081] = i[62];
  assign o[16082] = i[62];
  assign o[16083] = i[62];
  assign o[16084] = i[62];
  assign o[16085] = i[62];
  assign o[16086] = i[62];
  assign o[16087] = i[62];
  assign o[16088] = i[62];
  assign o[16089] = i[62];
  assign o[16090] = i[62];
  assign o[16091] = i[62];
  assign o[16092] = i[62];
  assign o[16093] = i[62];
  assign o[16094] = i[62];
  assign o[16095] = i[62];
  assign o[16096] = i[62];
  assign o[16097] = i[62];
  assign o[16098] = i[62];
  assign o[16099] = i[62];
  assign o[16100] = i[62];
  assign o[16101] = i[62];
  assign o[16102] = i[62];
  assign o[16103] = i[62];
  assign o[16104] = i[62];
  assign o[16105] = i[62];
  assign o[16106] = i[62];
  assign o[16107] = i[62];
  assign o[16108] = i[62];
  assign o[16109] = i[62];
  assign o[16110] = i[62];
  assign o[16111] = i[62];
  assign o[16112] = i[62];
  assign o[16113] = i[62];
  assign o[16114] = i[62];
  assign o[16115] = i[62];
  assign o[16116] = i[62];
  assign o[16117] = i[62];
  assign o[16118] = i[62];
  assign o[16119] = i[62];
  assign o[16120] = i[62];
  assign o[16121] = i[62];
  assign o[16122] = i[62];
  assign o[16123] = i[62];
  assign o[16124] = i[62];
  assign o[16125] = i[62];
  assign o[16126] = i[62];
  assign o[16127] = i[62];
  assign o[15616] = i[61];
  assign o[15617] = i[61];
  assign o[15618] = i[61];
  assign o[15619] = i[61];
  assign o[15620] = i[61];
  assign o[15621] = i[61];
  assign o[15622] = i[61];
  assign o[15623] = i[61];
  assign o[15624] = i[61];
  assign o[15625] = i[61];
  assign o[15626] = i[61];
  assign o[15627] = i[61];
  assign o[15628] = i[61];
  assign o[15629] = i[61];
  assign o[15630] = i[61];
  assign o[15631] = i[61];
  assign o[15632] = i[61];
  assign o[15633] = i[61];
  assign o[15634] = i[61];
  assign o[15635] = i[61];
  assign o[15636] = i[61];
  assign o[15637] = i[61];
  assign o[15638] = i[61];
  assign o[15639] = i[61];
  assign o[15640] = i[61];
  assign o[15641] = i[61];
  assign o[15642] = i[61];
  assign o[15643] = i[61];
  assign o[15644] = i[61];
  assign o[15645] = i[61];
  assign o[15646] = i[61];
  assign o[15647] = i[61];
  assign o[15648] = i[61];
  assign o[15649] = i[61];
  assign o[15650] = i[61];
  assign o[15651] = i[61];
  assign o[15652] = i[61];
  assign o[15653] = i[61];
  assign o[15654] = i[61];
  assign o[15655] = i[61];
  assign o[15656] = i[61];
  assign o[15657] = i[61];
  assign o[15658] = i[61];
  assign o[15659] = i[61];
  assign o[15660] = i[61];
  assign o[15661] = i[61];
  assign o[15662] = i[61];
  assign o[15663] = i[61];
  assign o[15664] = i[61];
  assign o[15665] = i[61];
  assign o[15666] = i[61];
  assign o[15667] = i[61];
  assign o[15668] = i[61];
  assign o[15669] = i[61];
  assign o[15670] = i[61];
  assign o[15671] = i[61];
  assign o[15672] = i[61];
  assign o[15673] = i[61];
  assign o[15674] = i[61];
  assign o[15675] = i[61];
  assign o[15676] = i[61];
  assign o[15677] = i[61];
  assign o[15678] = i[61];
  assign o[15679] = i[61];
  assign o[15680] = i[61];
  assign o[15681] = i[61];
  assign o[15682] = i[61];
  assign o[15683] = i[61];
  assign o[15684] = i[61];
  assign o[15685] = i[61];
  assign o[15686] = i[61];
  assign o[15687] = i[61];
  assign o[15688] = i[61];
  assign o[15689] = i[61];
  assign o[15690] = i[61];
  assign o[15691] = i[61];
  assign o[15692] = i[61];
  assign o[15693] = i[61];
  assign o[15694] = i[61];
  assign o[15695] = i[61];
  assign o[15696] = i[61];
  assign o[15697] = i[61];
  assign o[15698] = i[61];
  assign o[15699] = i[61];
  assign o[15700] = i[61];
  assign o[15701] = i[61];
  assign o[15702] = i[61];
  assign o[15703] = i[61];
  assign o[15704] = i[61];
  assign o[15705] = i[61];
  assign o[15706] = i[61];
  assign o[15707] = i[61];
  assign o[15708] = i[61];
  assign o[15709] = i[61];
  assign o[15710] = i[61];
  assign o[15711] = i[61];
  assign o[15712] = i[61];
  assign o[15713] = i[61];
  assign o[15714] = i[61];
  assign o[15715] = i[61];
  assign o[15716] = i[61];
  assign o[15717] = i[61];
  assign o[15718] = i[61];
  assign o[15719] = i[61];
  assign o[15720] = i[61];
  assign o[15721] = i[61];
  assign o[15722] = i[61];
  assign o[15723] = i[61];
  assign o[15724] = i[61];
  assign o[15725] = i[61];
  assign o[15726] = i[61];
  assign o[15727] = i[61];
  assign o[15728] = i[61];
  assign o[15729] = i[61];
  assign o[15730] = i[61];
  assign o[15731] = i[61];
  assign o[15732] = i[61];
  assign o[15733] = i[61];
  assign o[15734] = i[61];
  assign o[15735] = i[61];
  assign o[15736] = i[61];
  assign o[15737] = i[61];
  assign o[15738] = i[61];
  assign o[15739] = i[61];
  assign o[15740] = i[61];
  assign o[15741] = i[61];
  assign o[15742] = i[61];
  assign o[15743] = i[61];
  assign o[15744] = i[61];
  assign o[15745] = i[61];
  assign o[15746] = i[61];
  assign o[15747] = i[61];
  assign o[15748] = i[61];
  assign o[15749] = i[61];
  assign o[15750] = i[61];
  assign o[15751] = i[61];
  assign o[15752] = i[61];
  assign o[15753] = i[61];
  assign o[15754] = i[61];
  assign o[15755] = i[61];
  assign o[15756] = i[61];
  assign o[15757] = i[61];
  assign o[15758] = i[61];
  assign o[15759] = i[61];
  assign o[15760] = i[61];
  assign o[15761] = i[61];
  assign o[15762] = i[61];
  assign o[15763] = i[61];
  assign o[15764] = i[61];
  assign o[15765] = i[61];
  assign o[15766] = i[61];
  assign o[15767] = i[61];
  assign o[15768] = i[61];
  assign o[15769] = i[61];
  assign o[15770] = i[61];
  assign o[15771] = i[61];
  assign o[15772] = i[61];
  assign o[15773] = i[61];
  assign o[15774] = i[61];
  assign o[15775] = i[61];
  assign o[15776] = i[61];
  assign o[15777] = i[61];
  assign o[15778] = i[61];
  assign o[15779] = i[61];
  assign o[15780] = i[61];
  assign o[15781] = i[61];
  assign o[15782] = i[61];
  assign o[15783] = i[61];
  assign o[15784] = i[61];
  assign o[15785] = i[61];
  assign o[15786] = i[61];
  assign o[15787] = i[61];
  assign o[15788] = i[61];
  assign o[15789] = i[61];
  assign o[15790] = i[61];
  assign o[15791] = i[61];
  assign o[15792] = i[61];
  assign o[15793] = i[61];
  assign o[15794] = i[61];
  assign o[15795] = i[61];
  assign o[15796] = i[61];
  assign o[15797] = i[61];
  assign o[15798] = i[61];
  assign o[15799] = i[61];
  assign o[15800] = i[61];
  assign o[15801] = i[61];
  assign o[15802] = i[61];
  assign o[15803] = i[61];
  assign o[15804] = i[61];
  assign o[15805] = i[61];
  assign o[15806] = i[61];
  assign o[15807] = i[61];
  assign o[15808] = i[61];
  assign o[15809] = i[61];
  assign o[15810] = i[61];
  assign o[15811] = i[61];
  assign o[15812] = i[61];
  assign o[15813] = i[61];
  assign o[15814] = i[61];
  assign o[15815] = i[61];
  assign o[15816] = i[61];
  assign o[15817] = i[61];
  assign o[15818] = i[61];
  assign o[15819] = i[61];
  assign o[15820] = i[61];
  assign o[15821] = i[61];
  assign o[15822] = i[61];
  assign o[15823] = i[61];
  assign o[15824] = i[61];
  assign o[15825] = i[61];
  assign o[15826] = i[61];
  assign o[15827] = i[61];
  assign o[15828] = i[61];
  assign o[15829] = i[61];
  assign o[15830] = i[61];
  assign o[15831] = i[61];
  assign o[15832] = i[61];
  assign o[15833] = i[61];
  assign o[15834] = i[61];
  assign o[15835] = i[61];
  assign o[15836] = i[61];
  assign o[15837] = i[61];
  assign o[15838] = i[61];
  assign o[15839] = i[61];
  assign o[15840] = i[61];
  assign o[15841] = i[61];
  assign o[15842] = i[61];
  assign o[15843] = i[61];
  assign o[15844] = i[61];
  assign o[15845] = i[61];
  assign o[15846] = i[61];
  assign o[15847] = i[61];
  assign o[15848] = i[61];
  assign o[15849] = i[61];
  assign o[15850] = i[61];
  assign o[15851] = i[61];
  assign o[15852] = i[61];
  assign o[15853] = i[61];
  assign o[15854] = i[61];
  assign o[15855] = i[61];
  assign o[15856] = i[61];
  assign o[15857] = i[61];
  assign o[15858] = i[61];
  assign o[15859] = i[61];
  assign o[15860] = i[61];
  assign o[15861] = i[61];
  assign o[15862] = i[61];
  assign o[15863] = i[61];
  assign o[15864] = i[61];
  assign o[15865] = i[61];
  assign o[15866] = i[61];
  assign o[15867] = i[61];
  assign o[15868] = i[61];
  assign o[15869] = i[61];
  assign o[15870] = i[61];
  assign o[15871] = i[61];
  assign o[15360] = i[60];
  assign o[15361] = i[60];
  assign o[15362] = i[60];
  assign o[15363] = i[60];
  assign o[15364] = i[60];
  assign o[15365] = i[60];
  assign o[15366] = i[60];
  assign o[15367] = i[60];
  assign o[15368] = i[60];
  assign o[15369] = i[60];
  assign o[15370] = i[60];
  assign o[15371] = i[60];
  assign o[15372] = i[60];
  assign o[15373] = i[60];
  assign o[15374] = i[60];
  assign o[15375] = i[60];
  assign o[15376] = i[60];
  assign o[15377] = i[60];
  assign o[15378] = i[60];
  assign o[15379] = i[60];
  assign o[15380] = i[60];
  assign o[15381] = i[60];
  assign o[15382] = i[60];
  assign o[15383] = i[60];
  assign o[15384] = i[60];
  assign o[15385] = i[60];
  assign o[15386] = i[60];
  assign o[15387] = i[60];
  assign o[15388] = i[60];
  assign o[15389] = i[60];
  assign o[15390] = i[60];
  assign o[15391] = i[60];
  assign o[15392] = i[60];
  assign o[15393] = i[60];
  assign o[15394] = i[60];
  assign o[15395] = i[60];
  assign o[15396] = i[60];
  assign o[15397] = i[60];
  assign o[15398] = i[60];
  assign o[15399] = i[60];
  assign o[15400] = i[60];
  assign o[15401] = i[60];
  assign o[15402] = i[60];
  assign o[15403] = i[60];
  assign o[15404] = i[60];
  assign o[15405] = i[60];
  assign o[15406] = i[60];
  assign o[15407] = i[60];
  assign o[15408] = i[60];
  assign o[15409] = i[60];
  assign o[15410] = i[60];
  assign o[15411] = i[60];
  assign o[15412] = i[60];
  assign o[15413] = i[60];
  assign o[15414] = i[60];
  assign o[15415] = i[60];
  assign o[15416] = i[60];
  assign o[15417] = i[60];
  assign o[15418] = i[60];
  assign o[15419] = i[60];
  assign o[15420] = i[60];
  assign o[15421] = i[60];
  assign o[15422] = i[60];
  assign o[15423] = i[60];
  assign o[15424] = i[60];
  assign o[15425] = i[60];
  assign o[15426] = i[60];
  assign o[15427] = i[60];
  assign o[15428] = i[60];
  assign o[15429] = i[60];
  assign o[15430] = i[60];
  assign o[15431] = i[60];
  assign o[15432] = i[60];
  assign o[15433] = i[60];
  assign o[15434] = i[60];
  assign o[15435] = i[60];
  assign o[15436] = i[60];
  assign o[15437] = i[60];
  assign o[15438] = i[60];
  assign o[15439] = i[60];
  assign o[15440] = i[60];
  assign o[15441] = i[60];
  assign o[15442] = i[60];
  assign o[15443] = i[60];
  assign o[15444] = i[60];
  assign o[15445] = i[60];
  assign o[15446] = i[60];
  assign o[15447] = i[60];
  assign o[15448] = i[60];
  assign o[15449] = i[60];
  assign o[15450] = i[60];
  assign o[15451] = i[60];
  assign o[15452] = i[60];
  assign o[15453] = i[60];
  assign o[15454] = i[60];
  assign o[15455] = i[60];
  assign o[15456] = i[60];
  assign o[15457] = i[60];
  assign o[15458] = i[60];
  assign o[15459] = i[60];
  assign o[15460] = i[60];
  assign o[15461] = i[60];
  assign o[15462] = i[60];
  assign o[15463] = i[60];
  assign o[15464] = i[60];
  assign o[15465] = i[60];
  assign o[15466] = i[60];
  assign o[15467] = i[60];
  assign o[15468] = i[60];
  assign o[15469] = i[60];
  assign o[15470] = i[60];
  assign o[15471] = i[60];
  assign o[15472] = i[60];
  assign o[15473] = i[60];
  assign o[15474] = i[60];
  assign o[15475] = i[60];
  assign o[15476] = i[60];
  assign o[15477] = i[60];
  assign o[15478] = i[60];
  assign o[15479] = i[60];
  assign o[15480] = i[60];
  assign o[15481] = i[60];
  assign o[15482] = i[60];
  assign o[15483] = i[60];
  assign o[15484] = i[60];
  assign o[15485] = i[60];
  assign o[15486] = i[60];
  assign o[15487] = i[60];
  assign o[15488] = i[60];
  assign o[15489] = i[60];
  assign o[15490] = i[60];
  assign o[15491] = i[60];
  assign o[15492] = i[60];
  assign o[15493] = i[60];
  assign o[15494] = i[60];
  assign o[15495] = i[60];
  assign o[15496] = i[60];
  assign o[15497] = i[60];
  assign o[15498] = i[60];
  assign o[15499] = i[60];
  assign o[15500] = i[60];
  assign o[15501] = i[60];
  assign o[15502] = i[60];
  assign o[15503] = i[60];
  assign o[15504] = i[60];
  assign o[15505] = i[60];
  assign o[15506] = i[60];
  assign o[15507] = i[60];
  assign o[15508] = i[60];
  assign o[15509] = i[60];
  assign o[15510] = i[60];
  assign o[15511] = i[60];
  assign o[15512] = i[60];
  assign o[15513] = i[60];
  assign o[15514] = i[60];
  assign o[15515] = i[60];
  assign o[15516] = i[60];
  assign o[15517] = i[60];
  assign o[15518] = i[60];
  assign o[15519] = i[60];
  assign o[15520] = i[60];
  assign o[15521] = i[60];
  assign o[15522] = i[60];
  assign o[15523] = i[60];
  assign o[15524] = i[60];
  assign o[15525] = i[60];
  assign o[15526] = i[60];
  assign o[15527] = i[60];
  assign o[15528] = i[60];
  assign o[15529] = i[60];
  assign o[15530] = i[60];
  assign o[15531] = i[60];
  assign o[15532] = i[60];
  assign o[15533] = i[60];
  assign o[15534] = i[60];
  assign o[15535] = i[60];
  assign o[15536] = i[60];
  assign o[15537] = i[60];
  assign o[15538] = i[60];
  assign o[15539] = i[60];
  assign o[15540] = i[60];
  assign o[15541] = i[60];
  assign o[15542] = i[60];
  assign o[15543] = i[60];
  assign o[15544] = i[60];
  assign o[15545] = i[60];
  assign o[15546] = i[60];
  assign o[15547] = i[60];
  assign o[15548] = i[60];
  assign o[15549] = i[60];
  assign o[15550] = i[60];
  assign o[15551] = i[60];
  assign o[15552] = i[60];
  assign o[15553] = i[60];
  assign o[15554] = i[60];
  assign o[15555] = i[60];
  assign o[15556] = i[60];
  assign o[15557] = i[60];
  assign o[15558] = i[60];
  assign o[15559] = i[60];
  assign o[15560] = i[60];
  assign o[15561] = i[60];
  assign o[15562] = i[60];
  assign o[15563] = i[60];
  assign o[15564] = i[60];
  assign o[15565] = i[60];
  assign o[15566] = i[60];
  assign o[15567] = i[60];
  assign o[15568] = i[60];
  assign o[15569] = i[60];
  assign o[15570] = i[60];
  assign o[15571] = i[60];
  assign o[15572] = i[60];
  assign o[15573] = i[60];
  assign o[15574] = i[60];
  assign o[15575] = i[60];
  assign o[15576] = i[60];
  assign o[15577] = i[60];
  assign o[15578] = i[60];
  assign o[15579] = i[60];
  assign o[15580] = i[60];
  assign o[15581] = i[60];
  assign o[15582] = i[60];
  assign o[15583] = i[60];
  assign o[15584] = i[60];
  assign o[15585] = i[60];
  assign o[15586] = i[60];
  assign o[15587] = i[60];
  assign o[15588] = i[60];
  assign o[15589] = i[60];
  assign o[15590] = i[60];
  assign o[15591] = i[60];
  assign o[15592] = i[60];
  assign o[15593] = i[60];
  assign o[15594] = i[60];
  assign o[15595] = i[60];
  assign o[15596] = i[60];
  assign o[15597] = i[60];
  assign o[15598] = i[60];
  assign o[15599] = i[60];
  assign o[15600] = i[60];
  assign o[15601] = i[60];
  assign o[15602] = i[60];
  assign o[15603] = i[60];
  assign o[15604] = i[60];
  assign o[15605] = i[60];
  assign o[15606] = i[60];
  assign o[15607] = i[60];
  assign o[15608] = i[60];
  assign o[15609] = i[60];
  assign o[15610] = i[60];
  assign o[15611] = i[60];
  assign o[15612] = i[60];
  assign o[15613] = i[60];
  assign o[15614] = i[60];
  assign o[15615] = i[60];
  assign o[15104] = i[59];
  assign o[15105] = i[59];
  assign o[15106] = i[59];
  assign o[15107] = i[59];
  assign o[15108] = i[59];
  assign o[15109] = i[59];
  assign o[15110] = i[59];
  assign o[15111] = i[59];
  assign o[15112] = i[59];
  assign o[15113] = i[59];
  assign o[15114] = i[59];
  assign o[15115] = i[59];
  assign o[15116] = i[59];
  assign o[15117] = i[59];
  assign o[15118] = i[59];
  assign o[15119] = i[59];
  assign o[15120] = i[59];
  assign o[15121] = i[59];
  assign o[15122] = i[59];
  assign o[15123] = i[59];
  assign o[15124] = i[59];
  assign o[15125] = i[59];
  assign o[15126] = i[59];
  assign o[15127] = i[59];
  assign o[15128] = i[59];
  assign o[15129] = i[59];
  assign o[15130] = i[59];
  assign o[15131] = i[59];
  assign o[15132] = i[59];
  assign o[15133] = i[59];
  assign o[15134] = i[59];
  assign o[15135] = i[59];
  assign o[15136] = i[59];
  assign o[15137] = i[59];
  assign o[15138] = i[59];
  assign o[15139] = i[59];
  assign o[15140] = i[59];
  assign o[15141] = i[59];
  assign o[15142] = i[59];
  assign o[15143] = i[59];
  assign o[15144] = i[59];
  assign o[15145] = i[59];
  assign o[15146] = i[59];
  assign o[15147] = i[59];
  assign o[15148] = i[59];
  assign o[15149] = i[59];
  assign o[15150] = i[59];
  assign o[15151] = i[59];
  assign o[15152] = i[59];
  assign o[15153] = i[59];
  assign o[15154] = i[59];
  assign o[15155] = i[59];
  assign o[15156] = i[59];
  assign o[15157] = i[59];
  assign o[15158] = i[59];
  assign o[15159] = i[59];
  assign o[15160] = i[59];
  assign o[15161] = i[59];
  assign o[15162] = i[59];
  assign o[15163] = i[59];
  assign o[15164] = i[59];
  assign o[15165] = i[59];
  assign o[15166] = i[59];
  assign o[15167] = i[59];
  assign o[15168] = i[59];
  assign o[15169] = i[59];
  assign o[15170] = i[59];
  assign o[15171] = i[59];
  assign o[15172] = i[59];
  assign o[15173] = i[59];
  assign o[15174] = i[59];
  assign o[15175] = i[59];
  assign o[15176] = i[59];
  assign o[15177] = i[59];
  assign o[15178] = i[59];
  assign o[15179] = i[59];
  assign o[15180] = i[59];
  assign o[15181] = i[59];
  assign o[15182] = i[59];
  assign o[15183] = i[59];
  assign o[15184] = i[59];
  assign o[15185] = i[59];
  assign o[15186] = i[59];
  assign o[15187] = i[59];
  assign o[15188] = i[59];
  assign o[15189] = i[59];
  assign o[15190] = i[59];
  assign o[15191] = i[59];
  assign o[15192] = i[59];
  assign o[15193] = i[59];
  assign o[15194] = i[59];
  assign o[15195] = i[59];
  assign o[15196] = i[59];
  assign o[15197] = i[59];
  assign o[15198] = i[59];
  assign o[15199] = i[59];
  assign o[15200] = i[59];
  assign o[15201] = i[59];
  assign o[15202] = i[59];
  assign o[15203] = i[59];
  assign o[15204] = i[59];
  assign o[15205] = i[59];
  assign o[15206] = i[59];
  assign o[15207] = i[59];
  assign o[15208] = i[59];
  assign o[15209] = i[59];
  assign o[15210] = i[59];
  assign o[15211] = i[59];
  assign o[15212] = i[59];
  assign o[15213] = i[59];
  assign o[15214] = i[59];
  assign o[15215] = i[59];
  assign o[15216] = i[59];
  assign o[15217] = i[59];
  assign o[15218] = i[59];
  assign o[15219] = i[59];
  assign o[15220] = i[59];
  assign o[15221] = i[59];
  assign o[15222] = i[59];
  assign o[15223] = i[59];
  assign o[15224] = i[59];
  assign o[15225] = i[59];
  assign o[15226] = i[59];
  assign o[15227] = i[59];
  assign o[15228] = i[59];
  assign o[15229] = i[59];
  assign o[15230] = i[59];
  assign o[15231] = i[59];
  assign o[15232] = i[59];
  assign o[15233] = i[59];
  assign o[15234] = i[59];
  assign o[15235] = i[59];
  assign o[15236] = i[59];
  assign o[15237] = i[59];
  assign o[15238] = i[59];
  assign o[15239] = i[59];
  assign o[15240] = i[59];
  assign o[15241] = i[59];
  assign o[15242] = i[59];
  assign o[15243] = i[59];
  assign o[15244] = i[59];
  assign o[15245] = i[59];
  assign o[15246] = i[59];
  assign o[15247] = i[59];
  assign o[15248] = i[59];
  assign o[15249] = i[59];
  assign o[15250] = i[59];
  assign o[15251] = i[59];
  assign o[15252] = i[59];
  assign o[15253] = i[59];
  assign o[15254] = i[59];
  assign o[15255] = i[59];
  assign o[15256] = i[59];
  assign o[15257] = i[59];
  assign o[15258] = i[59];
  assign o[15259] = i[59];
  assign o[15260] = i[59];
  assign o[15261] = i[59];
  assign o[15262] = i[59];
  assign o[15263] = i[59];
  assign o[15264] = i[59];
  assign o[15265] = i[59];
  assign o[15266] = i[59];
  assign o[15267] = i[59];
  assign o[15268] = i[59];
  assign o[15269] = i[59];
  assign o[15270] = i[59];
  assign o[15271] = i[59];
  assign o[15272] = i[59];
  assign o[15273] = i[59];
  assign o[15274] = i[59];
  assign o[15275] = i[59];
  assign o[15276] = i[59];
  assign o[15277] = i[59];
  assign o[15278] = i[59];
  assign o[15279] = i[59];
  assign o[15280] = i[59];
  assign o[15281] = i[59];
  assign o[15282] = i[59];
  assign o[15283] = i[59];
  assign o[15284] = i[59];
  assign o[15285] = i[59];
  assign o[15286] = i[59];
  assign o[15287] = i[59];
  assign o[15288] = i[59];
  assign o[15289] = i[59];
  assign o[15290] = i[59];
  assign o[15291] = i[59];
  assign o[15292] = i[59];
  assign o[15293] = i[59];
  assign o[15294] = i[59];
  assign o[15295] = i[59];
  assign o[15296] = i[59];
  assign o[15297] = i[59];
  assign o[15298] = i[59];
  assign o[15299] = i[59];
  assign o[15300] = i[59];
  assign o[15301] = i[59];
  assign o[15302] = i[59];
  assign o[15303] = i[59];
  assign o[15304] = i[59];
  assign o[15305] = i[59];
  assign o[15306] = i[59];
  assign o[15307] = i[59];
  assign o[15308] = i[59];
  assign o[15309] = i[59];
  assign o[15310] = i[59];
  assign o[15311] = i[59];
  assign o[15312] = i[59];
  assign o[15313] = i[59];
  assign o[15314] = i[59];
  assign o[15315] = i[59];
  assign o[15316] = i[59];
  assign o[15317] = i[59];
  assign o[15318] = i[59];
  assign o[15319] = i[59];
  assign o[15320] = i[59];
  assign o[15321] = i[59];
  assign o[15322] = i[59];
  assign o[15323] = i[59];
  assign o[15324] = i[59];
  assign o[15325] = i[59];
  assign o[15326] = i[59];
  assign o[15327] = i[59];
  assign o[15328] = i[59];
  assign o[15329] = i[59];
  assign o[15330] = i[59];
  assign o[15331] = i[59];
  assign o[15332] = i[59];
  assign o[15333] = i[59];
  assign o[15334] = i[59];
  assign o[15335] = i[59];
  assign o[15336] = i[59];
  assign o[15337] = i[59];
  assign o[15338] = i[59];
  assign o[15339] = i[59];
  assign o[15340] = i[59];
  assign o[15341] = i[59];
  assign o[15342] = i[59];
  assign o[15343] = i[59];
  assign o[15344] = i[59];
  assign o[15345] = i[59];
  assign o[15346] = i[59];
  assign o[15347] = i[59];
  assign o[15348] = i[59];
  assign o[15349] = i[59];
  assign o[15350] = i[59];
  assign o[15351] = i[59];
  assign o[15352] = i[59];
  assign o[15353] = i[59];
  assign o[15354] = i[59];
  assign o[15355] = i[59];
  assign o[15356] = i[59];
  assign o[15357] = i[59];
  assign o[15358] = i[59];
  assign o[15359] = i[59];
  assign o[14848] = i[58];
  assign o[14849] = i[58];
  assign o[14850] = i[58];
  assign o[14851] = i[58];
  assign o[14852] = i[58];
  assign o[14853] = i[58];
  assign o[14854] = i[58];
  assign o[14855] = i[58];
  assign o[14856] = i[58];
  assign o[14857] = i[58];
  assign o[14858] = i[58];
  assign o[14859] = i[58];
  assign o[14860] = i[58];
  assign o[14861] = i[58];
  assign o[14862] = i[58];
  assign o[14863] = i[58];
  assign o[14864] = i[58];
  assign o[14865] = i[58];
  assign o[14866] = i[58];
  assign o[14867] = i[58];
  assign o[14868] = i[58];
  assign o[14869] = i[58];
  assign o[14870] = i[58];
  assign o[14871] = i[58];
  assign o[14872] = i[58];
  assign o[14873] = i[58];
  assign o[14874] = i[58];
  assign o[14875] = i[58];
  assign o[14876] = i[58];
  assign o[14877] = i[58];
  assign o[14878] = i[58];
  assign o[14879] = i[58];
  assign o[14880] = i[58];
  assign o[14881] = i[58];
  assign o[14882] = i[58];
  assign o[14883] = i[58];
  assign o[14884] = i[58];
  assign o[14885] = i[58];
  assign o[14886] = i[58];
  assign o[14887] = i[58];
  assign o[14888] = i[58];
  assign o[14889] = i[58];
  assign o[14890] = i[58];
  assign o[14891] = i[58];
  assign o[14892] = i[58];
  assign o[14893] = i[58];
  assign o[14894] = i[58];
  assign o[14895] = i[58];
  assign o[14896] = i[58];
  assign o[14897] = i[58];
  assign o[14898] = i[58];
  assign o[14899] = i[58];
  assign o[14900] = i[58];
  assign o[14901] = i[58];
  assign o[14902] = i[58];
  assign o[14903] = i[58];
  assign o[14904] = i[58];
  assign o[14905] = i[58];
  assign o[14906] = i[58];
  assign o[14907] = i[58];
  assign o[14908] = i[58];
  assign o[14909] = i[58];
  assign o[14910] = i[58];
  assign o[14911] = i[58];
  assign o[14912] = i[58];
  assign o[14913] = i[58];
  assign o[14914] = i[58];
  assign o[14915] = i[58];
  assign o[14916] = i[58];
  assign o[14917] = i[58];
  assign o[14918] = i[58];
  assign o[14919] = i[58];
  assign o[14920] = i[58];
  assign o[14921] = i[58];
  assign o[14922] = i[58];
  assign o[14923] = i[58];
  assign o[14924] = i[58];
  assign o[14925] = i[58];
  assign o[14926] = i[58];
  assign o[14927] = i[58];
  assign o[14928] = i[58];
  assign o[14929] = i[58];
  assign o[14930] = i[58];
  assign o[14931] = i[58];
  assign o[14932] = i[58];
  assign o[14933] = i[58];
  assign o[14934] = i[58];
  assign o[14935] = i[58];
  assign o[14936] = i[58];
  assign o[14937] = i[58];
  assign o[14938] = i[58];
  assign o[14939] = i[58];
  assign o[14940] = i[58];
  assign o[14941] = i[58];
  assign o[14942] = i[58];
  assign o[14943] = i[58];
  assign o[14944] = i[58];
  assign o[14945] = i[58];
  assign o[14946] = i[58];
  assign o[14947] = i[58];
  assign o[14948] = i[58];
  assign o[14949] = i[58];
  assign o[14950] = i[58];
  assign o[14951] = i[58];
  assign o[14952] = i[58];
  assign o[14953] = i[58];
  assign o[14954] = i[58];
  assign o[14955] = i[58];
  assign o[14956] = i[58];
  assign o[14957] = i[58];
  assign o[14958] = i[58];
  assign o[14959] = i[58];
  assign o[14960] = i[58];
  assign o[14961] = i[58];
  assign o[14962] = i[58];
  assign o[14963] = i[58];
  assign o[14964] = i[58];
  assign o[14965] = i[58];
  assign o[14966] = i[58];
  assign o[14967] = i[58];
  assign o[14968] = i[58];
  assign o[14969] = i[58];
  assign o[14970] = i[58];
  assign o[14971] = i[58];
  assign o[14972] = i[58];
  assign o[14973] = i[58];
  assign o[14974] = i[58];
  assign o[14975] = i[58];
  assign o[14976] = i[58];
  assign o[14977] = i[58];
  assign o[14978] = i[58];
  assign o[14979] = i[58];
  assign o[14980] = i[58];
  assign o[14981] = i[58];
  assign o[14982] = i[58];
  assign o[14983] = i[58];
  assign o[14984] = i[58];
  assign o[14985] = i[58];
  assign o[14986] = i[58];
  assign o[14987] = i[58];
  assign o[14988] = i[58];
  assign o[14989] = i[58];
  assign o[14990] = i[58];
  assign o[14991] = i[58];
  assign o[14992] = i[58];
  assign o[14993] = i[58];
  assign o[14994] = i[58];
  assign o[14995] = i[58];
  assign o[14996] = i[58];
  assign o[14997] = i[58];
  assign o[14998] = i[58];
  assign o[14999] = i[58];
  assign o[15000] = i[58];
  assign o[15001] = i[58];
  assign o[15002] = i[58];
  assign o[15003] = i[58];
  assign o[15004] = i[58];
  assign o[15005] = i[58];
  assign o[15006] = i[58];
  assign o[15007] = i[58];
  assign o[15008] = i[58];
  assign o[15009] = i[58];
  assign o[15010] = i[58];
  assign o[15011] = i[58];
  assign o[15012] = i[58];
  assign o[15013] = i[58];
  assign o[15014] = i[58];
  assign o[15015] = i[58];
  assign o[15016] = i[58];
  assign o[15017] = i[58];
  assign o[15018] = i[58];
  assign o[15019] = i[58];
  assign o[15020] = i[58];
  assign o[15021] = i[58];
  assign o[15022] = i[58];
  assign o[15023] = i[58];
  assign o[15024] = i[58];
  assign o[15025] = i[58];
  assign o[15026] = i[58];
  assign o[15027] = i[58];
  assign o[15028] = i[58];
  assign o[15029] = i[58];
  assign o[15030] = i[58];
  assign o[15031] = i[58];
  assign o[15032] = i[58];
  assign o[15033] = i[58];
  assign o[15034] = i[58];
  assign o[15035] = i[58];
  assign o[15036] = i[58];
  assign o[15037] = i[58];
  assign o[15038] = i[58];
  assign o[15039] = i[58];
  assign o[15040] = i[58];
  assign o[15041] = i[58];
  assign o[15042] = i[58];
  assign o[15043] = i[58];
  assign o[15044] = i[58];
  assign o[15045] = i[58];
  assign o[15046] = i[58];
  assign o[15047] = i[58];
  assign o[15048] = i[58];
  assign o[15049] = i[58];
  assign o[15050] = i[58];
  assign o[15051] = i[58];
  assign o[15052] = i[58];
  assign o[15053] = i[58];
  assign o[15054] = i[58];
  assign o[15055] = i[58];
  assign o[15056] = i[58];
  assign o[15057] = i[58];
  assign o[15058] = i[58];
  assign o[15059] = i[58];
  assign o[15060] = i[58];
  assign o[15061] = i[58];
  assign o[15062] = i[58];
  assign o[15063] = i[58];
  assign o[15064] = i[58];
  assign o[15065] = i[58];
  assign o[15066] = i[58];
  assign o[15067] = i[58];
  assign o[15068] = i[58];
  assign o[15069] = i[58];
  assign o[15070] = i[58];
  assign o[15071] = i[58];
  assign o[15072] = i[58];
  assign o[15073] = i[58];
  assign o[15074] = i[58];
  assign o[15075] = i[58];
  assign o[15076] = i[58];
  assign o[15077] = i[58];
  assign o[15078] = i[58];
  assign o[15079] = i[58];
  assign o[15080] = i[58];
  assign o[15081] = i[58];
  assign o[15082] = i[58];
  assign o[15083] = i[58];
  assign o[15084] = i[58];
  assign o[15085] = i[58];
  assign o[15086] = i[58];
  assign o[15087] = i[58];
  assign o[15088] = i[58];
  assign o[15089] = i[58];
  assign o[15090] = i[58];
  assign o[15091] = i[58];
  assign o[15092] = i[58];
  assign o[15093] = i[58];
  assign o[15094] = i[58];
  assign o[15095] = i[58];
  assign o[15096] = i[58];
  assign o[15097] = i[58];
  assign o[15098] = i[58];
  assign o[15099] = i[58];
  assign o[15100] = i[58];
  assign o[15101] = i[58];
  assign o[15102] = i[58];
  assign o[15103] = i[58];
  assign o[14592] = i[57];
  assign o[14593] = i[57];
  assign o[14594] = i[57];
  assign o[14595] = i[57];
  assign o[14596] = i[57];
  assign o[14597] = i[57];
  assign o[14598] = i[57];
  assign o[14599] = i[57];
  assign o[14600] = i[57];
  assign o[14601] = i[57];
  assign o[14602] = i[57];
  assign o[14603] = i[57];
  assign o[14604] = i[57];
  assign o[14605] = i[57];
  assign o[14606] = i[57];
  assign o[14607] = i[57];
  assign o[14608] = i[57];
  assign o[14609] = i[57];
  assign o[14610] = i[57];
  assign o[14611] = i[57];
  assign o[14612] = i[57];
  assign o[14613] = i[57];
  assign o[14614] = i[57];
  assign o[14615] = i[57];
  assign o[14616] = i[57];
  assign o[14617] = i[57];
  assign o[14618] = i[57];
  assign o[14619] = i[57];
  assign o[14620] = i[57];
  assign o[14621] = i[57];
  assign o[14622] = i[57];
  assign o[14623] = i[57];
  assign o[14624] = i[57];
  assign o[14625] = i[57];
  assign o[14626] = i[57];
  assign o[14627] = i[57];
  assign o[14628] = i[57];
  assign o[14629] = i[57];
  assign o[14630] = i[57];
  assign o[14631] = i[57];
  assign o[14632] = i[57];
  assign o[14633] = i[57];
  assign o[14634] = i[57];
  assign o[14635] = i[57];
  assign o[14636] = i[57];
  assign o[14637] = i[57];
  assign o[14638] = i[57];
  assign o[14639] = i[57];
  assign o[14640] = i[57];
  assign o[14641] = i[57];
  assign o[14642] = i[57];
  assign o[14643] = i[57];
  assign o[14644] = i[57];
  assign o[14645] = i[57];
  assign o[14646] = i[57];
  assign o[14647] = i[57];
  assign o[14648] = i[57];
  assign o[14649] = i[57];
  assign o[14650] = i[57];
  assign o[14651] = i[57];
  assign o[14652] = i[57];
  assign o[14653] = i[57];
  assign o[14654] = i[57];
  assign o[14655] = i[57];
  assign o[14656] = i[57];
  assign o[14657] = i[57];
  assign o[14658] = i[57];
  assign o[14659] = i[57];
  assign o[14660] = i[57];
  assign o[14661] = i[57];
  assign o[14662] = i[57];
  assign o[14663] = i[57];
  assign o[14664] = i[57];
  assign o[14665] = i[57];
  assign o[14666] = i[57];
  assign o[14667] = i[57];
  assign o[14668] = i[57];
  assign o[14669] = i[57];
  assign o[14670] = i[57];
  assign o[14671] = i[57];
  assign o[14672] = i[57];
  assign o[14673] = i[57];
  assign o[14674] = i[57];
  assign o[14675] = i[57];
  assign o[14676] = i[57];
  assign o[14677] = i[57];
  assign o[14678] = i[57];
  assign o[14679] = i[57];
  assign o[14680] = i[57];
  assign o[14681] = i[57];
  assign o[14682] = i[57];
  assign o[14683] = i[57];
  assign o[14684] = i[57];
  assign o[14685] = i[57];
  assign o[14686] = i[57];
  assign o[14687] = i[57];
  assign o[14688] = i[57];
  assign o[14689] = i[57];
  assign o[14690] = i[57];
  assign o[14691] = i[57];
  assign o[14692] = i[57];
  assign o[14693] = i[57];
  assign o[14694] = i[57];
  assign o[14695] = i[57];
  assign o[14696] = i[57];
  assign o[14697] = i[57];
  assign o[14698] = i[57];
  assign o[14699] = i[57];
  assign o[14700] = i[57];
  assign o[14701] = i[57];
  assign o[14702] = i[57];
  assign o[14703] = i[57];
  assign o[14704] = i[57];
  assign o[14705] = i[57];
  assign o[14706] = i[57];
  assign o[14707] = i[57];
  assign o[14708] = i[57];
  assign o[14709] = i[57];
  assign o[14710] = i[57];
  assign o[14711] = i[57];
  assign o[14712] = i[57];
  assign o[14713] = i[57];
  assign o[14714] = i[57];
  assign o[14715] = i[57];
  assign o[14716] = i[57];
  assign o[14717] = i[57];
  assign o[14718] = i[57];
  assign o[14719] = i[57];
  assign o[14720] = i[57];
  assign o[14721] = i[57];
  assign o[14722] = i[57];
  assign o[14723] = i[57];
  assign o[14724] = i[57];
  assign o[14725] = i[57];
  assign o[14726] = i[57];
  assign o[14727] = i[57];
  assign o[14728] = i[57];
  assign o[14729] = i[57];
  assign o[14730] = i[57];
  assign o[14731] = i[57];
  assign o[14732] = i[57];
  assign o[14733] = i[57];
  assign o[14734] = i[57];
  assign o[14735] = i[57];
  assign o[14736] = i[57];
  assign o[14737] = i[57];
  assign o[14738] = i[57];
  assign o[14739] = i[57];
  assign o[14740] = i[57];
  assign o[14741] = i[57];
  assign o[14742] = i[57];
  assign o[14743] = i[57];
  assign o[14744] = i[57];
  assign o[14745] = i[57];
  assign o[14746] = i[57];
  assign o[14747] = i[57];
  assign o[14748] = i[57];
  assign o[14749] = i[57];
  assign o[14750] = i[57];
  assign o[14751] = i[57];
  assign o[14752] = i[57];
  assign o[14753] = i[57];
  assign o[14754] = i[57];
  assign o[14755] = i[57];
  assign o[14756] = i[57];
  assign o[14757] = i[57];
  assign o[14758] = i[57];
  assign o[14759] = i[57];
  assign o[14760] = i[57];
  assign o[14761] = i[57];
  assign o[14762] = i[57];
  assign o[14763] = i[57];
  assign o[14764] = i[57];
  assign o[14765] = i[57];
  assign o[14766] = i[57];
  assign o[14767] = i[57];
  assign o[14768] = i[57];
  assign o[14769] = i[57];
  assign o[14770] = i[57];
  assign o[14771] = i[57];
  assign o[14772] = i[57];
  assign o[14773] = i[57];
  assign o[14774] = i[57];
  assign o[14775] = i[57];
  assign o[14776] = i[57];
  assign o[14777] = i[57];
  assign o[14778] = i[57];
  assign o[14779] = i[57];
  assign o[14780] = i[57];
  assign o[14781] = i[57];
  assign o[14782] = i[57];
  assign o[14783] = i[57];
  assign o[14784] = i[57];
  assign o[14785] = i[57];
  assign o[14786] = i[57];
  assign o[14787] = i[57];
  assign o[14788] = i[57];
  assign o[14789] = i[57];
  assign o[14790] = i[57];
  assign o[14791] = i[57];
  assign o[14792] = i[57];
  assign o[14793] = i[57];
  assign o[14794] = i[57];
  assign o[14795] = i[57];
  assign o[14796] = i[57];
  assign o[14797] = i[57];
  assign o[14798] = i[57];
  assign o[14799] = i[57];
  assign o[14800] = i[57];
  assign o[14801] = i[57];
  assign o[14802] = i[57];
  assign o[14803] = i[57];
  assign o[14804] = i[57];
  assign o[14805] = i[57];
  assign o[14806] = i[57];
  assign o[14807] = i[57];
  assign o[14808] = i[57];
  assign o[14809] = i[57];
  assign o[14810] = i[57];
  assign o[14811] = i[57];
  assign o[14812] = i[57];
  assign o[14813] = i[57];
  assign o[14814] = i[57];
  assign o[14815] = i[57];
  assign o[14816] = i[57];
  assign o[14817] = i[57];
  assign o[14818] = i[57];
  assign o[14819] = i[57];
  assign o[14820] = i[57];
  assign o[14821] = i[57];
  assign o[14822] = i[57];
  assign o[14823] = i[57];
  assign o[14824] = i[57];
  assign o[14825] = i[57];
  assign o[14826] = i[57];
  assign o[14827] = i[57];
  assign o[14828] = i[57];
  assign o[14829] = i[57];
  assign o[14830] = i[57];
  assign o[14831] = i[57];
  assign o[14832] = i[57];
  assign o[14833] = i[57];
  assign o[14834] = i[57];
  assign o[14835] = i[57];
  assign o[14836] = i[57];
  assign o[14837] = i[57];
  assign o[14838] = i[57];
  assign o[14839] = i[57];
  assign o[14840] = i[57];
  assign o[14841] = i[57];
  assign o[14842] = i[57];
  assign o[14843] = i[57];
  assign o[14844] = i[57];
  assign o[14845] = i[57];
  assign o[14846] = i[57];
  assign o[14847] = i[57];
  assign o[14336] = i[56];
  assign o[14337] = i[56];
  assign o[14338] = i[56];
  assign o[14339] = i[56];
  assign o[14340] = i[56];
  assign o[14341] = i[56];
  assign o[14342] = i[56];
  assign o[14343] = i[56];
  assign o[14344] = i[56];
  assign o[14345] = i[56];
  assign o[14346] = i[56];
  assign o[14347] = i[56];
  assign o[14348] = i[56];
  assign o[14349] = i[56];
  assign o[14350] = i[56];
  assign o[14351] = i[56];
  assign o[14352] = i[56];
  assign o[14353] = i[56];
  assign o[14354] = i[56];
  assign o[14355] = i[56];
  assign o[14356] = i[56];
  assign o[14357] = i[56];
  assign o[14358] = i[56];
  assign o[14359] = i[56];
  assign o[14360] = i[56];
  assign o[14361] = i[56];
  assign o[14362] = i[56];
  assign o[14363] = i[56];
  assign o[14364] = i[56];
  assign o[14365] = i[56];
  assign o[14366] = i[56];
  assign o[14367] = i[56];
  assign o[14368] = i[56];
  assign o[14369] = i[56];
  assign o[14370] = i[56];
  assign o[14371] = i[56];
  assign o[14372] = i[56];
  assign o[14373] = i[56];
  assign o[14374] = i[56];
  assign o[14375] = i[56];
  assign o[14376] = i[56];
  assign o[14377] = i[56];
  assign o[14378] = i[56];
  assign o[14379] = i[56];
  assign o[14380] = i[56];
  assign o[14381] = i[56];
  assign o[14382] = i[56];
  assign o[14383] = i[56];
  assign o[14384] = i[56];
  assign o[14385] = i[56];
  assign o[14386] = i[56];
  assign o[14387] = i[56];
  assign o[14388] = i[56];
  assign o[14389] = i[56];
  assign o[14390] = i[56];
  assign o[14391] = i[56];
  assign o[14392] = i[56];
  assign o[14393] = i[56];
  assign o[14394] = i[56];
  assign o[14395] = i[56];
  assign o[14396] = i[56];
  assign o[14397] = i[56];
  assign o[14398] = i[56];
  assign o[14399] = i[56];
  assign o[14400] = i[56];
  assign o[14401] = i[56];
  assign o[14402] = i[56];
  assign o[14403] = i[56];
  assign o[14404] = i[56];
  assign o[14405] = i[56];
  assign o[14406] = i[56];
  assign o[14407] = i[56];
  assign o[14408] = i[56];
  assign o[14409] = i[56];
  assign o[14410] = i[56];
  assign o[14411] = i[56];
  assign o[14412] = i[56];
  assign o[14413] = i[56];
  assign o[14414] = i[56];
  assign o[14415] = i[56];
  assign o[14416] = i[56];
  assign o[14417] = i[56];
  assign o[14418] = i[56];
  assign o[14419] = i[56];
  assign o[14420] = i[56];
  assign o[14421] = i[56];
  assign o[14422] = i[56];
  assign o[14423] = i[56];
  assign o[14424] = i[56];
  assign o[14425] = i[56];
  assign o[14426] = i[56];
  assign o[14427] = i[56];
  assign o[14428] = i[56];
  assign o[14429] = i[56];
  assign o[14430] = i[56];
  assign o[14431] = i[56];
  assign o[14432] = i[56];
  assign o[14433] = i[56];
  assign o[14434] = i[56];
  assign o[14435] = i[56];
  assign o[14436] = i[56];
  assign o[14437] = i[56];
  assign o[14438] = i[56];
  assign o[14439] = i[56];
  assign o[14440] = i[56];
  assign o[14441] = i[56];
  assign o[14442] = i[56];
  assign o[14443] = i[56];
  assign o[14444] = i[56];
  assign o[14445] = i[56];
  assign o[14446] = i[56];
  assign o[14447] = i[56];
  assign o[14448] = i[56];
  assign o[14449] = i[56];
  assign o[14450] = i[56];
  assign o[14451] = i[56];
  assign o[14452] = i[56];
  assign o[14453] = i[56];
  assign o[14454] = i[56];
  assign o[14455] = i[56];
  assign o[14456] = i[56];
  assign o[14457] = i[56];
  assign o[14458] = i[56];
  assign o[14459] = i[56];
  assign o[14460] = i[56];
  assign o[14461] = i[56];
  assign o[14462] = i[56];
  assign o[14463] = i[56];
  assign o[14464] = i[56];
  assign o[14465] = i[56];
  assign o[14466] = i[56];
  assign o[14467] = i[56];
  assign o[14468] = i[56];
  assign o[14469] = i[56];
  assign o[14470] = i[56];
  assign o[14471] = i[56];
  assign o[14472] = i[56];
  assign o[14473] = i[56];
  assign o[14474] = i[56];
  assign o[14475] = i[56];
  assign o[14476] = i[56];
  assign o[14477] = i[56];
  assign o[14478] = i[56];
  assign o[14479] = i[56];
  assign o[14480] = i[56];
  assign o[14481] = i[56];
  assign o[14482] = i[56];
  assign o[14483] = i[56];
  assign o[14484] = i[56];
  assign o[14485] = i[56];
  assign o[14486] = i[56];
  assign o[14487] = i[56];
  assign o[14488] = i[56];
  assign o[14489] = i[56];
  assign o[14490] = i[56];
  assign o[14491] = i[56];
  assign o[14492] = i[56];
  assign o[14493] = i[56];
  assign o[14494] = i[56];
  assign o[14495] = i[56];
  assign o[14496] = i[56];
  assign o[14497] = i[56];
  assign o[14498] = i[56];
  assign o[14499] = i[56];
  assign o[14500] = i[56];
  assign o[14501] = i[56];
  assign o[14502] = i[56];
  assign o[14503] = i[56];
  assign o[14504] = i[56];
  assign o[14505] = i[56];
  assign o[14506] = i[56];
  assign o[14507] = i[56];
  assign o[14508] = i[56];
  assign o[14509] = i[56];
  assign o[14510] = i[56];
  assign o[14511] = i[56];
  assign o[14512] = i[56];
  assign o[14513] = i[56];
  assign o[14514] = i[56];
  assign o[14515] = i[56];
  assign o[14516] = i[56];
  assign o[14517] = i[56];
  assign o[14518] = i[56];
  assign o[14519] = i[56];
  assign o[14520] = i[56];
  assign o[14521] = i[56];
  assign o[14522] = i[56];
  assign o[14523] = i[56];
  assign o[14524] = i[56];
  assign o[14525] = i[56];
  assign o[14526] = i[56];
  assign o[14527] = i[56];
  assign o[14528] = i[56];
  assign o[14529] = i[56];
  assign o[14530] = i[56];
  assign o[14531] = i[56];
  assign o[14532] = i[56];
  assign o[14533] = i[56];
  assign o[14534] = i[56];
  assign o[14535] = i[56];
  assign o[14536] = i[56];
  assign o[14537] = i[56];
  assign o[14538] = i[56];
  assign o[14539] = i[56];
  assign o[14540] = i[56];
  assign o[14541] = i[56];
  assign o[14542] = i[56];
  assign o[14543] = i[56];
  assign o[14544] = i[56];
  assign o[14545] = i[56];
  assign o[14546] = i[56];
  assign o[14547] = i[56];
  assign o[14548] = i[56];
  assign o[14549] = i[56];
  assign o[14550] = i[56];
  assign o[14551] = i[56];
  assign o[14552] = i[56];
  assign o[14553] = i[56];
  assign o[14554] = i[56];
  assign o[14555] = i[56];
  assign o[14556] = i[56];
  assign o[14557] = i[56];
  assign o[14558] = i[56];
  assign o[14559] = i[56];
  assign o[14560] = i[56];
  assign o[14561] = i[56];
  assign o[14562] = i[56];
  assign o[14563] = i[56];
  assign o[14564] = i[56];
  assign o[14565] = i[56];
  assign o[14566] = i[56];
  assign o[14567] = i[56];
  assign o[14568] = i[56];
  assign o[14569] = i[56];
  assign o[14570] = i[56];
  assign o[14571] = i[56];
  assign o[14572] = i[56];
  assign o[14573] = i[56];
  assign o[14574] = i[56];
  assign o[14575] = i[56];
  assign o[14576] = i[56];
  assign o[14577] = i[56];
  assign o[14578] = i[56];
  assign o[14579] = i[56];
  assign o[14580] = i[56];
  assign o[14581] = i[56];
  assign o[14582] = i[56];
  assign o[14583] = i[56];
  assign o[14584] = i[56];
  assign o[14585] = i[56];
  assign o[14586] = i[56];
  assign o[14587] = i[56];
  assign o[14588] = i[56];
  assign o[14589] = i[56];
  assign o[14590] = i[56];
  assign o[14591] = i[56];
  assign o[14080] = i[55];
  assign o[14081] = i[55];
  assign o[14082] = i[55];
  assign o[14083] = i[55];
  assign o[14084] = i[55];
  assign o[14085] = i[55];
  assign o[14086] = i[55];
  assign o[14087] = i[55];
  assign o[14088] = i[55];
  assign o[14089] = i[55];
  assign o[14090] = i[55];
  assign o[14091] = i[55];
  assign o[14092] = i[55];
  assign o[14093] = i[55];
  assign o[14094] = i[55];
  assign o[14095] = i[55];
  assign o[14096] = i[55];
  assign o[14097] = i[55];
  assign o[14098] = i[55];
  assign o[14099] = i[55];
  assign o[14100] = i[55];
  assign o[14101] = i[55];
  assign o[14102] = i[55];
  assign o[14103] = i[55];
  assign o[14104] = i[55];
  assign o[14105] = i[55];
  assign o[14106] = i[55];
  assign o[14107] = i[55];
  assign o[14108] = i[55];
  assign o[14109] = i[55];
  assign o[14110] = i[55];
  assign o[14111] = i[55];
  assign o[14112] = i[55];
  assign o[14113] = i[55];
  assign o[14114] = i[55];
  assign o[14115] = i[55];
  assign o[14116] = i[55];
  assign o[14117] = i[55];
  assign o[14118] = i[55];
  assign o[14119] = i[55];
  assign o[14120] = i[55];
  assign o[14121] = i[55];
  assign o[14122] = i[55];
  assign o[14123] = i[55];
  assign o[14124] = i[55];
  assign o[14125] = i[55];
  assign o[14126] = i[55];
  assign o[14127] = i[55];
  assign o[14128] = i[55];
  assign o[14129] = i[55];
  assign o[14130] = i[55];
  assign o[14131] = i[55];
  assign o[14132] = i[55];
  assign o[14133] = i[55];
  assign o[14134] = i[55];
  assign o[14135] = i[55];
  assign o[14136] = i[55];
  assign o[14137] = i[55];
  assign o[14138] = i[55];
  assign o[14139] = i[55];
  assign o[14140] = i[55];
  assign o[14141] = i[55];
  assign o[14142] = i[55];
  assign o[14143] = i[55];
  assign o[14144] = i[55];
  assign o[14145] = i[55];
  assign o[14146] = i[55];
  assign o[14147] = i[55];
  assign o[14148] = i[55];
  assign o[14149] = i[55];
  assign o[14150] = i[55];
  assign o[14151] = i[55];
  assign o[14152] = i[55];
  assign o[14153] = i[55];
  assign o[14154] = i[55];
  assign o[14155] = i[55];
  assign o[14156] = i[55];
  assign o[14157] = i[55];
  assign o[14158] = i[55];
  assign o[14159] = i[55];
  assign o[14160] = i[55];
  assign o[14161] = i[55];
  assign o[14162] = i[55];
  assign o[14163] = i[55];
  assign o[14164] = i[55];
  assign o[14165] = i[55];
  assign o[14166] = i[55];
  assign o[14167] = i[55];
  assign o[14168] = i[55];
  assign o[14169] = i[55];
  assign o[14170] = i[55];
  assign o[14171] = i[55];
  assign o[14172] = i[55];
  assign o[14173] = i[55];
  assign o[14174] = i[55];
  assign o[14175] = i[55];
  assign o[14176] = i[55];
  assign o[14177] = i[55];
  assign o[14178] = i[55];
  assign o[14179] = i[55];
  assign o[14180] = i[55];
  assign o[14181] = i[55];
  assign o[14182] = i[55];
  assign o[14183] = i[55];
  assign o[14184] = i[55];
  assign o[14185] = i[55];
  assign o[14186] = i[55];
  assign o[14187] = i[55];
  assign o[14188] = i[55];
  assign o[14189] = i[55];
  assign o[14190] = i[55];
  assign o[14191] = i[55];
  assign o[14192] = i[55];
  assign o[14193] = i[55];
  assign o[14194] = i[55];
  assign o[14195] = i[55];
  assign o[14196] = i[55];
  assign o[14197] = i[55];
  assign o[14198] = i[55];
  assign o[14199] = i[55];
  assign o[14200] = i[55];
  assign o[14201] = i[55];
  assign o[14202] = i[55];
  assign o[14203] = i[55];
  assign o[14204] = i[55];
  assign o[14205] = i[55];
  assign o[14206] = i[55];
  assign o[14207] = i[55];
  assign o[14208] = i[55];
  assign o[14209] = i[55];
  assign o[14210] = i[55];
  assign o[14211] = i[55];
  assign o[14212] = i[55];
  assign o[14213] = i[55];
  assign o[14214] = i[55];
  assign o[14215] = i[55];
  assign o[14216] = i[55];
  assign o[14217] = i[55];
  assign o[14218] = i[55];
  assign o[14219] = i[55];
  assign o[14220] = i[55];
  assign o[14221] = i[55];
  assign o[14222] = i[55];
  assign o[14223] = i[55];
  assign o[14224] = i[55];
  assign o[14225] = i[55];
  assign o[14226] = i[55];
  assign o[14227] = i[55];
  assign o[14228] = i[55];
  assign o[14229] = i[55];
  assign o[14230] = i[55];
  assign o[14231] = i[55];
  assign o[14232] = i[55];
  assign o[14233] = i[55];
  assign o[14234] = i[55];
  assign o[14235] = i[55];
  assign o[14236] = i[55];
  assign o[14237] = i[55];
  assign o[14238] = i[55];
  assign o[14239] = i[55];
  assign o[14240] = i[55];
  assign o[14241] = i[55];
  assign o[14242] = i[55];
  assign o[14243] = i[55];
  assign o[14244] = i[55];
  assign o[14245] = i[55];
  assign o[14246] = i[55];
  assign o[14247] = i[55];
  assign o[14248] = i[55];
  assign o[14249] = i[55];
  assign o[14250] = i[55];
  assign o[14251] = i[55];
  assign o[14252] = i[55];
  assign o[14253] = i[55];
  assign o[14254] = i[55];
  assign o[14255] = i[55];
  assign o[14256] = i[55];
  assign o[14257] = i[55];
  assign o[14258] = i[55];
  assign o[14259] = i[55];
  assign o[14260] = i[55];
  assign o[14261] = i[55];
  assign o[14262] = i[55];
  assign o[14263] = i[55];
  assign o[14264] = i[55];
  assign o[14265] = i[55];
  assign o[14266] = i[55];
  assign o[14267] = i[55];
  assign o[14268] = i[55];
  assign o[14269] = i[55];
  assign o[14270] = i[55];
  assign o[14271] = i[55];
  assign o[14272] = i[55];
  assign o[14273] = i[55];
  assign o[14274] = i[55];
  assign o[14275] = i[55];
  assign o[14276] = i[55];
  assign o[14277] = i[55];
  assign o[14278] = i[55];
  assign o[14279] = i[55];
  assign o[14280] = i[55];
  assign o[14281] = i[55];
  assign o[14282] = i[55];
  assign o[14283] = i[55];
  assign o[14284] = i[55];
  assign o[14285] = i[55];
  assign o[14286] = i[55];
  assign o[14287] = i[55];
  assign o[14288] = i[55];
  assign o[14289] = i[55];
  assign o[14290] = i[55];
  assign o[14291] = i[55];
  assign o[14292] = i[55];
  assign o[14293] = i[55];
  assign o[14294] = i[55];
  assign o[14295] = i[55];
  assign o[14296] = i[55];
  assign o[14297] = i[55];
  assign o[14298] = i[55];
  assign o[14299] = i[55];
  assign o[14300] = i[55];
  assign o[14301] = i[55];
  assign o[14302] = i[55];
  assign o[14303] = i[55];
  assign o[14304] = i[55];
  assign o[14305] = i[55];
  assign o[14306] = i[55];
  assign o[14307] = i[55];
  assign o[14308] = i[55];
  assign o[14309] = i[55];
  assign o[14310] = i[55];
  assign o[14311] = i[55];
  assign o[14312] = i[55];
  assign o[14313] = i[55];
  assign o[14314] = i[55];
  assign o[14315] = i[55];
  assign o[14316] = i[55];
  assign o[14317] = i[55];
  assign o[14318] = i[55];
  assign o[14319] = i[55];
  assign o[14320] = i[55];
  assign o[14321] = i[55];
  assign o[14322] = i[55];
  assign o[14323] = i[55];
  assign o[14324] = i[55];
  assign o[14325] = i[55];
  assign o[14326] = i[55];
  assign o[14327] = i[55];
  assign o[14328] = i[55];
  assign o[14329] = i[55];
  assign o[14330] = i[55];
  assign o[14331] = i[55];
  assign o[14332] = i[55];
  assign o[14333] = i[55];
  assign o[14334] = i[55];
  assign o[14335] = i[55];
  assign o[13824] = i[54];
  assign o[13825] = i[54];
  assign o[13826] = i[54];
  assign o[13827] = i[54];
  assign o[13828] = i[54];
  assign o[13829] = i[54];
  assign o[13830] = i[54];
  assign o[13831] = i[54];
  assign o[13832] = i[54];
  assign o[13833] = i[54];
  assign o[13834] = i[54];
  assign o[13835] = i[54];
  assign o[13836] = i[54];
  assign o[13837] = i[54];
  assign o[13838] = i[54];
  assign o[13839] = i[54];
  assign o[13840] = i[54];
  assign o[13841] = i[54];
  assign o[13842] = i[54];
  assign o[13843] = i[54];
  assign o[13844] = i[54];
  assign o[13845] = i[54];
  assign o[13846] = i[54];
  assign o[13847] = i[54];
  assign o[13848] = i[54];
  assign o[13849] = i[54];
  assign o[13850] = i[54];
  assign o[13851] = i[54];
  assign o[13852] = i[54];
  assign o[13853] = i[54];
  assign o[13854] = i[54];
  assign o[13855] = i[54];
  assign o[13856] = i[54];
  assign o[13857] = i[54];
  assign o[13858] = i[54];
  assign o[13859] = i[54];
  assign o[13860] = i[54];
  assign o[13861] = i[54];
  assign o[13862] = i[54];
  assign o[13863] = i[54];
  assign o[13864] = i[54];
  assign o[13865] = i[54];
  assign o[13866] = i[54];
  assign o[13867] = i[54];
  assign o[13868] = i[54];
  assign o[13869] = i[54];
  assign o[13870] = i[54];
  assign o[13871] = i[54];
  assign o[13872] = i[54];
  assign o[13873] = i[54];
  assign o[13874] = i[54];
  assign o[13875] = i[54];
  assign o[13876] = i[54];
  assign o[13877] = i[54];
  assign o[13878] = i[54];
  assign o[13879] = i[54];
  assign o[13880] = i[54];
  assign o[13881] = i[54];
  assign o[13882] = i[54];
  assign o[13883] = i[54];
  assign o[13884] = i[54];
  assign o[13885] = i[54];
  assign o[13886] = i[54];
  assign o[13887] = i[54];
  assign o[13888] = i[54];
  assign o[13889] = i[54];
  assign o[13890] = i[54];
  assign o[13891] = i[54];
  assign o[13892] = i[54];
  assign o[13893] = i[54];
  assign o[13894] = i[54];
  assign o[13895] = i[54];
  assign o[13896] = i[54];
  assign o[13897] = i[54];
  assign o[13898] = i[54];
  assign o[13899] = i[54];
  assign o[13900] = i[54];
  assign o[13901] = i[54];
  assign o[13902] = i[54];
  assign o[13903] = i[54];
  assign o[13904] = i[54];
  assign o[13905] = i[54];
  assign o[13906] = i[54];
  assign o[13907] = i[54];
  assign o[13908] = i[54];
  assign o[13909] = i[54];
  assign o[13910] = i[54];
  assign o[13911] = i[54];
  assign o[13912] = i[54];
  assign o[13913] = i[54];
  assign o[13914] = i[54];
  assign o[13915] = i[54];
  assign o[13916] = i[54];
  assign o[13917] = i[54];
  assign o[13918] = i[54];
  assign o[13919] = i[54];
  assign o[13920] = i[54];
  assign o[13921] = i[54];
  assign o[13922] = i[54];
  assign o[13923] = i[54];
  assign o[13924] = i[54];
  assign o[13925] = i[54];
  assign o[13926] = i[54];
  assign o[13927] = i[54];
  assign o[13928] = i[54];
  assign o[13929] = i[54];
  assign o[13930] = i[54];
  assign o[13931] = i[54];
  assign o[13932] = i[54];
  assign o[13933] = i[54];
  assign o[13934] = i[54];
  assign o[13935] = i[54];
  assign o[13936] = i[54];
  assign o[13937] = i[54];
  assign o[13938] = i[54];
  assign o[13939] = i[54];
  assign o[13940] = i[54];
  assign o[13941] = i[54];
  assign o[13942] = i[54];
  assign o[13943] = i[54];
  assign o[13944] = i[54];
  assign o[13945] = i[54];
  assign o[13946] = i[54];
  assign o[13947] = i[54];
  assign o[13948] = i[54];
  assign o[13949] = i[54];
  assign o[13950] = i[54];
  assign o[13951] = i[54];
  assign o[13952] = i[54];
  assign o[13953] = i[54];
  assign o[13954] = i[54];
  assign o[13955] = i[54];
  assign o[13956] = i[54];
  assign o[13957] = i[54];
  assign o[13958] = i[54];
  assign o[13959] = i[54];
  assign o[13960] = i[54];
  assign o[13961] = i[54];
  assign o[13962] = i[54];
  assign o[13963] = i[54];
  assign o[13964] = i[54];
  assign o[13965] = i[54];
  assign o[13966] = i[54];
  assign o[13967] = i[54];
  assign o[13968] = i[54];
  assign o[13969] = i[54];
  assign o[13970] = i[54];
  assign o[13971] = i[54];
  assign o[13972] = i[54];
  assign o[13973] = i[54];
  assign o[13974] = i[54];
  assign o[13975] = i[54];
  assign o[13976] = i[54];
  assign o[13977] = i[54];
  assign o[13978] = i[54];
  assign o[13979] = i[54];
  assign o[13980] = i[54];
  assign o[13981] = i[54];
  assign o[13982] = i[54];
  assign o[13983] = i[54];
  assign o[13984] = i[54];
  assign o[13985] = i[54];
  assign o[13986] = i[54];
  assign o[13987] = i[54];
  assign o[13988] = i[54];
  assign o[13989] = i[54];
  assign o[13990] = i[54];
  assign o[13991] = i[54];
  assign o[13992] = i[54];
  assign o[13993] = i[54];
  assign o[13994] = i[54];
  assign o[13995] = i[54];
  assign o[13996] = i[54];
  assign o[13997] = i[54];
  assign o[13998] = i[54];
  assign o[13999] = i[54];
  assign o[14000] = i[54];
  assign o[14001] = i[54];
  assign o[14002] = i[54];
  assign o[14003] = i[54];
  assign o[14004] = i[54];
  assign o[14005] = i[54];
  assign o[14006] = i[54];
  assign o[14007] = i[54];
  assign o[14008] = i[54];
  assign o[14009] = i[54];
  assign o[14010] = i[54];
  assign o[14011] = i[54];
  assign o[14012] = i[54];
  assign o[14013] = i[54];
  assign o[14014] = i[54];
  assign o[14015] = i[54];
  assign o[14016] = i[54];
  assign o[14017] = i[54];
  assign o[14018] = i[54];
  assign o[14019] = i[54];
  assign o[14020] = i[54];
  assign o[14021] = i[54];
  assign o[14022] = i[54];
  assign o[14023] = i[54];
  assign o[14024] = i[54];
  assign o[14025] = i[54];
  assign o[14026] = i[54];
  assign o[14027] = i[54];
  assign o[14028] = i[54];
  assign o[14029] = i[54];
  assign o[14030] = i[54];
  assign o[14031] = i[54];
  assign o[14032] = i[54];
  assign o[14033] = i[54];
  assign o[14034] = i[54];
  assign o[14035] = i[54];
  assign o[14036] = i[54];
  assign o[14037] = i[54];
  assign o[14038] = i[54];
  assign o[14039] = i[54];
  assign o[14040] = i[54];
  assign o[14041] = i[54];
  assign o[14042] = i[54];
  assign o[14043] = i[54];
  assign o[14044] = i[54];
  assign o[14045] = i[54];
  assign o[14046] = i[54];
  assign o[14047] = i[54];
  assign o[14048] = i[54];
  assign o[14049] = i[54];
  assign o[14050] = i[54];
  assign o[14051] = i[54];
  assign o[14052] = i[54];
  assign o[14053] = i[54];
  assign o[14054] = i[54];
  assign o[14055] = i[54];
  assign o[14056] = i[54];
  assign o[14057] = i[54];
  assign o[14058] = i[54];
  assign o[14059] = i[54];
  assign o[14060] = i[54];
  assign o[14061] = i[54];
  assign o[14062] = i[54];
  assign o[14063] = i[54];
  assign o[14064] = i[54];
  assign o[14065] = i[54];
  assign o[14066] = i[54];
  assign o[14067] = i[54];
  assign o[14068] = i[54];
  assign o[14069] = i[54];
  assign o[14070] = i[54];
  assign o[14071] = i[54];
  assign o[14072] = i[54];
  assign o[14073] = i[54];
  assign o[14074] = i[54];
  assign o[14075] = i[54];
  assign o[14076] = i[54];
  assign o[14077] = i[54];
  assign o[14078] = i[54];
  assign o[14079] = i[54];
  assign o[13568] = i[53];
  assign o[13569] = i[53];
  assign o[13570] = i[53];
  assign o[13571] = i[53];
  assign o[13572] = i[53];
  assign o[13573] = i[53];
  assign o[13574] = i[53];
  assign o[13575] = i[53];
  assign o[13576] = i[53];
  assign o[13577] = i[53];
  assign o[13578] = i[53];
  assign o[13579] = i[53];
  assign o[13580] = i[53];
  assign o[13581] = i[53];
  assign o[13582] = i[53];
  assign o[13583] = i[53];
  assign o[13584] = i[53];
  assign o[13585] = i[53];
  assign o[13586] = i[53];
  assign o[13587] = i[53];
  assign o[13588] = i[53];
  assign o[13589] = i[53];
  assign o[13590] = i[53];
  assign o[13591] = i[53];
  assign o[13592] = i[53];
  assign o[13593] = i[53];
  assign o[13594] = i[53];
  assign o[13595] = i[53];
  assign o[13596] = i[53];
  assign o[13597] = i[53];
  assign o[13598] = i[53];
  assign o[13599] = i[53];
  assign o[13600] = i[53];
  assign o[13601] = i[53];
  assign o[13602] = i[53];
  assign o[13603] = i[53];
  assign o[13604] = i[53];
  assign o[13605] = i[53];
  assign o[13606] = i[53];
  assign o[13607] = i[53];
  assign o[13608] = i[53];
  assign o[13609] = i[53];
  assign o[13610] = i[53];
  assign o[13611] = i[53];
  assign o[13612] = i[53];
  assign o[13613] = i[53];
  assign o[13614] = i[53];
  assign o[13615] = i[53];
  assign o[13616] = i[53];
  assign o[13617] = i[53];
  assign o[13618] = i[53];
  assign o[13619] = i[53];
  assign o[13620] = i[53];
  assign o[13621] = i[53];
  assign o[13622] = i[53];
  assign o[13623] = i[53];
  assign o[13624] = i[53];
  assign o[13625] = i[53];
  assign o[13626] = i[53];
  assign o[13627] = i[53];
  assign o[13628] = i[53];
  assign o[13629] = i[53];
  assign o[13630] = i[53];
  assign o[13631] = i[53];
  assign o[13632] = i[53];
  assign o[13633] = i[53];
  assign o[13634] = i[53];
  assign o[13635] = i[53];
  assign o[13636] = i[53];
  assign o[13637] = i[53];
  assign o[13638] = i[53];
  assign o[13639] = i[53];
  assign o[13640] = i[53];
  assign o[13641] = i[53];
  assign o[13642] = i[53];
  assign o[13643] = i[53];
  assign o[13644] = i[53];
  assign o[13645] = i[53];
  assign o[13646] = i[53];
  assign o[13647] = i[53];
  assign o[13648] = i[53];
  assign o[13649] = i[53];
  assign o[13650] = i[53];
  assign o[13651] = i[53];
  assign o[13652] = i[53];
  assign o[13653] = i[53];
  assign o[13654] = i[53];
  assign o[13655] = i[53];
  assign o[13656] = i[53];
  assign o[13657] = i[53];
  assign o[13658] = i[53];
  assign o[13659] = i[53];
  assign o[13660] = i[53];
  assign o[13661] = i[53];
  assign o[13662] = i[53];
  assign o[13663] = i[53];
  assign o[13664] = i[53];
  assign o[13665] = i[53];
  assign o[13666] = i[53];
  assign o[13667] = i[53];
  assign o[13668] = i[53];
  assign o[13669] = i[53];
  assign o[13670] = i[53];
  assign o[13671] = i[53];
  assign o[13672] = i[53];
  assign o[13673] = i[53];
  assign o[13674] = i[53];
  assign o[13675] = i[53];
  assign o[13676] = i[53];
  assign o[13677] = i[53];
  assign o[13678] = i[53];
  assign o[13679] = i[53];
  assign o[13680] = i[53];
  assign o[13681] = i[53];
  assign o[13682] = i[53];
  assign o[13683] = i[53];
  assign o[13684] = i[53];
  assign o[13685] = i[53];
  assign o[13686] = i[53];
  assign o[13687] = i[53];
  assign o[13688] = i[53];
  assign o[13689] = i[53];
  assign o[13690] = i[53];
  assign o[13691] = i[53];
  assign o[13692] = i[53];
  assign o[13693] = i[53];
  assign o[13694] = i[53];
  assign o[13695] = i[53];
  assign o[13696] = i[53];
  assign o[13697] = i[53];
  assign o[13698] = i[53];
  assign o[13699] = i[53];
  assign o[13700] = i[53];
  assign o[13701] = i[53];
  assign o[13702] = i[53];
  assign o[13703] = i[53];
  assign o[13704] = i[53];
  assign o[13705] = i[53];
  assign o[13706] = i[53];
  assign o[13707] = i[53];
  assign o[13708] = i[53];
  assign o[13709] = i[53];
  assign o[13710] = i[53];
  assign o[13711] = i[53];
  assign o[13712] = i[53];
  assign o[13713] = i[53];
  assign o[13714] = i[53];
  assign o[13715] = i[53];
  assign o[13716] = i[53];
  assign o[13717] = i[53];
  assign o[13718] = i[53];
  assign o[13719] = i[53];
  assign o[13720] = i[53];
  assign o[13721] = i[53];
  assign o[13722] = i[53];
  assign o[13723] = i[53];
  assign o[13724] = i[53];
  assign o[13725] = i[53];
  assign o[13726] = i[53];
  assign o[13727] = i[53];
  assign o[13728] = i[53];
  assign o[13729] = i[53];
  assign o[13730] = i[53];
  assign o[13731] = i[53];
  assign o[13732] = i[53];
  assign o[13733] = i[53];
  assign o[13734] = i[53];
  assign o[13735] = i[53];
  assign o[13736] = i[53];
  assign o[13737] = i[53];
  assign o[13738] = i[53];
  assign o[13739] = i[53];
  assign o[13740] = i[53];
  assign o[13741] = i[53];
  assign o[13742] = i[53];
  assign o[13743] = i[53];
  assign o[13744] = i[53];
  assign o[13745] = i[53];
  assign o[13746] = i[53];
  assign o[13747] = i[53];
  assign o[13748] = i[53];
  assign o[13749] = i[53];
  assign o[13750] = i[53];
  assign o[13751] = i[53];
  assign o[13752] = i[53];
  assign o[13753] = i[53];
  assign o[13754] = i[53];
  assign o[13755] = i[53];
  assign o[13756] = i[53];
  assign o[13757] = i[53];
  assign o[13758] = i[53];
  assign o[13759] = i[53];
  assign o[13760] = i[53];
  assign o[13761] = i[53];
  assign o[13762] = i[53];
  assign o[13763] = i[53];
  assign o[13764] = i[53];
  assign o[13765] = i[53];
  assign o[13766] = i[53];
  assign o[13767] = i[53];
  assign o[13768] = i[53];
  assign o[13769] = i[53];
  assign o[13770] = i[53];
  assign o[13771] = i[53];
  assign o[13772] = i[53];
  assign o[13773] = i[53];
  assign o[13774] = i[53];
  assign o[13775] = i[53];
  assign o[13776] = i[53];
  assign o[13777] = i[53];
  assign o[13778] = i[53];
  assign o[13779] = i[53];
  assign o[13780] = i[53];
  assign o[13781] = i[53];
  assign o[13782] = i[53];
  assign o[13783] = i[53];
  assign o[13784] = i[53];
  assign o[13785] = i[53];
  assign o[13786] = i[53];
  assign o[13787] = i[53];
  assign o[13788] = i[53];
  assign o[13789] = i[53];
  assign o[13790] = i[53];
  assign o[13791] = i[53];
  assign o[13792] = i[53];
  assign o[13793] = i[53];
  assign o[13794] = i[53];
  assign o[13795] = i[53];
  assign o[13796] = i[53];
  assign o[13797] = i[53];
  assign o[13798] = i[53];
  assign o[13799] = i[53];
  assign o[13800] = i[53];
  assign o[13801] = i[53];
  assign o[13802] = i[53];
  assign o[13803] = i[53];
  assign o[13804] = i[53];
  assign o[13805] = i[53];
  assign o[13806] = i[53];
  assign o[13807] = i[53];
  assign o[13808] = i[53];
  assign o[13809] = i[53];
  assign o[13810] = i[53];
  assign o[13811] = i[53];
  assign o[13812] = i[53];
  assign o[13813] = i[53];
  assign o[13814] = i[53];
  assign o[13815] = i[53];
  assign o[13816] = i[53];
  assign o[13817] = i[53];
  assign o[13818] = i[53];
  assign o[13819] = i[53];
  assign o[13820] = i[53];
  assign o[13821] = i[53];
  assign o[13822] = i[53];
  assign o[13823] = i[53];
  assign o[13312] = i[52];
  assign o[13313] = i[52];
  assign o[13314] = i[52];
  assign o[13315] = i[52];
  assign o[13316] = i[52];
  assign o[13317] = i[52];
  assign o[13318] = i[52];
  assign o[13319] = i[52];
  assign o[13320] = i[52];
  assign o[13321] = i[52];
  assign o[13322] = i[52];
  assign o[13323] = i[52];
  assign o[13324] = i[52];
  assign o[13325] = i[52];
  assign o[13326] = i[52];
  assign o[13327] = i[52];
  assign o[13328] = i[52];
  assign o[13329] = i[52];
  assign o[13330] = i[52];
  assign o[13331] = i[52];
  assign o[13332] = i[52];
  assign o[13333] = i[52];
  assign o[13334] = i[52];
  assign o[13335] = i[52];
  assign o[13336] = i[52];
  assign o[13337] = i[52];
  assign o[13338] = i[52];
  assign o[13339] = i[52];
  assign o[13340] = i[52];
  assign o[13341] = i[52];
  assign o[13342] = i[52];
  assign o[13343] = i[52];
  assign o[13344] = i[52];
  assign o[13345] = i[52];
  assign o[13346] = i[52];
  assign o[13347] = i[52];
  assign o[13348] = i[52];
  assign o[13349] = i[52];
  assign o[13350] = i[52];
  assign o[13351] = i[52];
  assign o[13352] = i[52];
  assign o[13353] = i[52];
  assign o[13354] = i[52];
  assign o[13355] = i[52];
  assign o[13356] = i[52];
  assign o[13357] = i[52];
  assign o[13358] = i[52];
  assign o[13359] = i[52];
  assign o[13360] = i[52];
  assign o[13361] = i[52];
  assign o[13362] = i[52];
  assign o[13363] = i[52];
  assign o[13364] = i[52];
  assign o[13365] = i[52];
  assign o[13366] = i[52];
  assign o[13367] = i[52];
  assign o[13368] = i[52];
  assign o[13369] = i[52];
  assign o[13370] = i[52];
  assign o[13371] = i[52];
  assign o[13372] = i[52];
  assign o[13373] = i[52];
  assign o[13374] = i[52];
  assign o[13375] = i[52];
  assign o[13376] = i[52];
  assign o[13377] = i[52];
  assign o[13378] = i[52];
  assign o[13379] = i[52];
  assign o[13380] = i[52];
  assign o[13381] = i[52];
  assign o[13382] = i[52];
  assign o[13383] = i[52];
  assign o[13384] = i[52];
  assign o[13385] = i[52];
  assign o[13386] = i[52];
  assign o[13387] = i[52];
  assign o[13388] = i[52];
  assign o[13389] = i[52];
  assign o[13390] = i[52];
  assign o[13391] = i[52];
  assign o[13392] = i[52];
  assign o[13393] = i[52];
  assign o[13394] = i[52];
  assign o[13395] = i[52];
  assign o[13396] = i[52];
  assign o[13397] = i[52];
  assign o[13398] = i[52];
  assign o[13399] = i[52];
  assign o[13400] = i[52];
  assign o[13401] = i[52];
  assign o[13402] = i[52];
  assign o[13403] = i[52];
  assign o[13404] = i[52];
  assign o[13405] = i[52];
  assign o[13406] = i[52];
  assign o[13407] = i[52];
  assign o[13408] = i[52];
  assign o[13409] = i[52];
  assign o[13410] = i[52];
  assign o[13411] = i[52];
  assign o[13412] = i[52];
  assign o[13413] = i[52];
  assign o[13414] = i[52];
  assign o[13415] = i[52];
  assign o[13416] = i[52];
  assign o[13417] = i[52];
  assign o[13418] = i[52];
  assign o[13419] = i[52];
  assign o[13420] = i[52];
  assign o[13421] = i[52];
  assign o[13422] = i[52];
  assign o[13423] = i[52];
  assign o[13424] = i[52];
  assign o[13425] = i[52];
  assign o[13426] = i[52];
  assign o[13427] = i[52];
  assign o[13428] = i[52];
  assign o[13429] = i[52];
  assign o[13430] = i[52];
  assign o[13431] = i[52];
  assign o[13432] = i[52];
  assign o[13433] = i[52];
  assign o[13434] = i[52];
  assign o[13435] = i[52];
  assign o[13436] = i[52];
  assign o[13437] = i[52];
  assign o[13438] = i[52];
  assign o[13439] = i[52];
  assign o[13440] = i[52];
  assign o[13441] = i[52];
  assign o[13442] = i[52];
  assign o[13443] = i[52];
  assign o[13444] = i[52];
  assign o[13445] = i[52];
  assign o[13446] = i[52];
  assign o[13447] = i[52];
  assign o[13448] = i[52];
  assign o[13449] = i[52];
  assign o[13450] = i[52];
  assign o[13451] = i[52];
  assign o[13452] = i[52];
  assign o[13453] = i[52];
  assign o[13454] = i[52];
  assign o[13455] = i[52];
  assign o[13456] = i[52];
  assign o[13457] = i[52];
  assign o[13458] = i[52];
  assign o[13459] = i[52];
  assign o[13460] = i[52];
  assign o[13461] = i[52];
  assign o[13462] = i[52];
  assign o[13463] = i[52];
  assign o[13464] = i[52];
  assign o[13465] = i[52];
  assign o[13466] = i[52];
  assign o[13467] = i[52];
  assign o[13468] = i[52];
  assign o[13469] = i[52];
  assign o[13470] = i[52];
  assign o[13471] = i[52];
  assign o[13472] = i[52];
  assign o[13473] = i[52];
  assign o[13474] = i[52];
  assign o[13475] = i[52];
  assign o[13476] = i[52];
  assign o[13477] = i[52];
  assign o[13478] = i[52];
  assign o[13479] = i[52];
  assign o[13480] = i[52];
  assign o[13481] = i[52];
  assign o[13482] = i[52];
  assign o[13483] = i[52];
  assign o[13484] = i[52];
  assign o[13485] = i[52];
  assign o[13486] = i[52];
  assign o[13487] = i[52];
  assign o[13488] = i[52];
  assign o[13489] = i[52];
  assign o[13490] = i[52];
  assign o[13491] = i[52];
  assign o[13492] = i[52];
  assign o[13493] = i[52];
  assign o[13494] = i[52];
  assign o[13495] = i[52];
  assign o[13496] = i[52];
  assign o[13497] = i[52];
  assign o[13498] = i[52];
  assign o[13499] = i[52];
  assign o[13500] = i[52];
  assign o[13501] = i[52];
  assign o[13502] = i[52];
  assign o[13503] = i[52];
  assign o[13504] = i[52];
  assign o[13505] = i[52];
  assign o[13506] = i[52];
  assign o[13507] = i[52];
  assign o[13508] = i[52];
  assign o[13509] = i[52];
  assign o[13510] = i[52];
  assign o[13511] = i[52];
  assign o[13512] = i[52];
  assign o[13513] = i[52];
  assign o[13514] = i[52];
  assign o[13515] = i[52];
  assign o[13516] = i[52];
  assign o[13517] = i[52];
  assign o[13518] = i[52];
  assign o[13519] = i[52];
  assign o[13520] = i[52];
  assign o[13521] = i[52];
  assign o[13522] = i[52];
  assign o[13523] = i[52];
  assign o[13524] = i[52];
  assign o[13525] = i[52];
  assign o[13526] = i[52];
  assign o[13527] = i[52];
  assign o[13528] = i[52];
  assign o[13529] = i[52];
  assign o[13530] = i[52];
  assign o[13531] = i[52];
  assign o[13532] = i[52];
  assign o[13533] = i[52];
  assign o[13534] = i[52];
  assign o[13535] = i[52];
  assign o[13536] = i[52];
  assign o[13537] = i[52];
  assign o[13538] = i[52];
  assign o[13539] = i[52];
  assign o[13540] = i[52];
  assign o[13541] = i[52];
  assign o[13542] = i[52];
  assign o[13543] = i[52];
  assign o[13544] = i[52];
  assign o[13545] = i[52];
  assign o[13546] = i[52];
  assign o[13547] = i[52];
  assign o[13548] = i[52];
  assign o[13549] = i[52];
  assign o[13550] = i[52];
  assign o[13551] = i[52];
  assign o[13552] = i[52];
  assign o[13553] = i[52];
  assign o[13554] = i[52];
  assign o[13555] = i[52];
  assign o[13556] = i[52];
  assign o[13557] = i[52];
  assign o[13558] = i[52];
  assign o[13559] = i[52];
  assign o[13560] = i[52];
  assign o[13561] = i[52];
  assign o[13562] = i[52];
  assign o[13563] = i[52];
  assign o[13564] = i[52];
  assign o[13565] = i[52];
  assign o[13566] = i[52];
  assign o[13567] = i[52];
  assign o[13056] = i[51];
  assign o[13057] = i[51];
  assign o[13058] = i[51];
  assign o[13059] = i[51];
  assign o[13060] = i[51];
  assign o[13061] = i[51];
  assign o[13062] = i[51];
  assign o[13063] = i[51];
  assign o[13064] = i[51];
  assign o[13065] = i[51];
  assign o[13066] = i[51];
  assign o[13067] = i[51];
  assign o[13068] = i[51];
  assign o[13069] = i[51];
  assign o[13070] = i[51];
  assign o[13071] = i[51];
  assign o[13072] = i[51];
  assign o[13073] = i[51];
  assign o[13074] = i[51];
  assign o[13075] = i[51];
  assign o[13076] = i[51];
  assign o[13077] = i[51];
  assign o[13078] = i[51];
  assign o[13079] = i[51];
  assign o[13080] = i[51];
  assign o[13081] = i[51];
  assign o[13082] = i[51];
  assign o[13083] = i[51];
  assign o[13084] = i[51];
  assign o[13085] = i[51];
  assign o[13086] = i[51];
  assign o[13087] = i[51];
  assign o[13088] = i[51];
  assign o[13089] = i[51];
  assign o[13090] = i[51];
  assign o[13091] = i[51];
  assign o[13092] = i[51];
  assign o[13093] = i[51];
  assign o[13094] = i[51];
  assign o[13095] = i[51];
  assign o[13096] = i[51];
  assign o[13097] = i[51];
  assign o[13098] = i[51];
  assign o[13099] = i[51];
  assign o[13100] = i[51];
  assign o[13101] = i[51];
  assign o[13102] = i[51];
  assign o[13103] = i[51];
  assign o[13104] = i[51];
  assign o[13105] = i[51];
  assign o[13106] = i[51];
  assign o[13107] = i[51];
  assign o[13108] = i[51];
  assign o[13109] = i[51];
  assign o[13110] = i[51];
  assign o[13111] = i[51];
  assign o[13112] = i[51];
  assign o[13113] = i[51];
  assign o[13114] = i[51];
  assign o[13115] = i[51];
  assign o[13116] = i[51];
  assign o[13117] = i[51];
  assign o[13118] = i[51];
  assign o[13119] = i[51];
  assign o[13120] = i[51];
  assign o[13121] = i[51];
  assign o[13122] = i[51];
  assign o[13123] = i[51];
  assign o[13124] = i[51];
  assign o[13125] = i[51];
  assign o[13126] = i[51];
  assign o[13127] = i[51];
  assign o[13128] = i[51];
  assign o[13129] = i[51];
  assign o[13130] = i[51];
  assign o[13131] = i[51];
  assign o[13132] = i[51];
  assign o[13133] = i[51];
  assign o[13134] = i[51];
  assign o[13135] = i[51];
  assign o[13136] = i[51];
  assign o[13137] = i[51];
  assign o[13138] = i[51];
  assign o[13139] = i[51];
  assign o[13140] = i[51];
  assign o[13141] = i[51];
  assign o[13142] = i[51];
  assign o[13143] = i[51];
  assign o[13144] = i[51];
  assign o[13145] = i[51];
  assign o[13146] = i[51];
  assign o[13147] = i[51];
  assign o[13148] = i[51];
  assign o[13149] = i[51];
  assign o[13150] = i[51];
  assign o[13151] = i[51];
  assign o[13152] = i[51];
  assign o[13153] = i[51];
  assign o[13154] = i[51];
  assign o[13155] = i[51];
  assign o[13156] = i[51];
  assign o[13157] = i[51];
  assign o[13158] = i[51];
  assign o[13159] = i[51];
  assign o[13160] = i[51];
  assign o[13161] = i[51];
  assign o[13162] = i[51];
  assign o[13163] = i[51];
  assign o[13164] = i[51];
  assign o[13165] = i[51];
  assign o[13166] = i[51];
  assign o[13167] = i[51];
  assign o[13168] = i[51];
  assign o[13169] = i[51];
  assign o[13170] = i[51];
  assign o[13171] = i[51];
  assign o[13172] = i[51];
  assign o[13173] = i[51];
  assign o[13174] = i[51];
  assign o[13175] = i[51];
  assign o[13176] = i[51];
  assign o[13177] = i[51];
  assign o[13178] = i[51];
  assign o[13179] = i[51];
  assign o[13180] = i[51];
  assign o[13181] = i[51];
  assign o[13182] = i[51];
  assign o[13183] = i[51];
  assign o[13184] = i[51];
  assign o[13185] = i[51];
  assign o[13186] = i[51];
  assign o[13187] = i[51];
  assign o[13188] = i[51];
  assign o[13189] = i[51];
  assign o[13190] = i[51];
  assign o[13191] = i[51];
  assign o[13192] = i[51];
  assign o[13193] = i[51];
  assign o[13194] = i[51];
  assign o[13195] = i[51];
  assign o[13196] = i[51];
  assign o[13197] = i[51];
  assign o[13198] = i[51];
  assign o[13199] = i[51];
  assign o[13200] = i[51];
  assign o[13201] = i[51];
  assign o[13202] = i[51];
  assign o[13203] = i[51];
  assign o[13204] = i[51];
  assign o[13205] = i[51];
  assign o[13206] = i[51];
  assign o[13207] = i[51];
  assign o[13208] = i[51];
  assign o[13209] = i[51];
  assign o[13210] = i[51];
  assign o[13211] = i[51];
  assign o[13212] = i[51];
  assign o[13213] = i[51];
  assign o[13214] = i[51];
  assign o[13215] = i[51];
  assign o[13216] = i[51];
  assign o[13217] = i[51];
  assign o[13218] = i[51];
  assign o[13219] = i[51];
  assign o[13220] = i[51];
  assign o[13221] = i[51];
  assign o[13222] = i[51];
  assign o[13223] = i[51];
  assign o[13224] = i[51];
  assign o[13225] = i[51];
  assign o[13226] = i[51];
  assign o[13227] = i[51];
  assign o[13228] = i[51];
  assign o[13229] = i[51];
  assign o[13230] = i[51];
  assign o[13231] = i[51];
  assign o[13232] = i[51];
  assign o[13233] = i[51];
  assign o[13234] = i[51];
  assign o[13235] = i[51];
  assign o[13236] = i[51];
  assign o[13237] = i[51];
  assign o[13238] = i[51];
  assign o[13239] = i[51];
  assign o[13240] = i[51];
  assign o[13241] = i[51];
  assign o[13242] = i[51];
  assign o[13243] = i[51];
  assign o[13244] = i[51];
  assign o[13245] = i[51];
  assign o[13246] = i[51];
  assign o[13247] = i[51];
  assign o[13248] = i[51];
  assign o[13249] = i[51];
  assign o[13250] = i[51];
  assign o[13251] = i[51];
  assign o[13252] = i[51];
  assign o[13253] = i[51];
  assign o[13254] = i[51];
  assign o[13255] = i[51];
  assign o[13256] = i[51];
  assign o[13257] = i[51];
  assign o[13258] = i[51];
  assign o[13259] = i[51];
  assign o[13260] = i[51];
  assign o[13261] = i[51];
  assign o[13262] = i[51];
  assign o[13263] = i[51];
  assign o[13264] = i[51];
  assign o[13265] = i[51];
  assign o[13266] = i[51];
  assign o[13267] = i[51];
  assign o[13268] = i[51];
  assign o[13269] = i[51];
  assign o[13270] = i[51];
  assign o[13271] = i[51];
  assign o[13272] = i[51];
  assign o[13273] = i[51];
  assign o[13274] = i[51];
  assign o[13275] = i[51];
  assign o[13276] = i[51];
  assign o[13277] = i[51];
  assign o[13278] = i[51];
  assign o[13279] = i[51];
  assign o[13280] = i[51];
  assign o[13281] = i[51];
  assign o[13282] = i[51];
  assign o[13283] = i[51];
  assign o[13284] = i[51];
  assign o[13285] = i[51];
  assign o[13286] = i[51];
  assign o[13287] = i[51];
  assign o[13288] = i[51];
  assign o[13289] = i[51];
  assign o[13290] = i[51];
  assign o[13291] = i[51];
  assign o[13292] = i[51];
  assign o[13293] = i[51];
  assign o[13294] = i[51];
  assign o[13295] = i[51];
  assign o[13296] = i[51];
  assign o[13297] = i[51];
  assign o[13298] = i[51];
  assign o[13299] = i[51];
  assign o[13300] = i[51];
  assign o[13301] = i[51];
  assign o[13302] = i[51];
  assign o[13303] = i[51];
  assign o[13304] = i[51];
  assign o[13305] = i[51];
  assign o[13306] = i[51];
  assign o[13307] = i[51];
  assign o[13308] = i[51];
  assign o[13309] = i[51];
  assign o[13310] = i[51];
  assign o[13311] = i[51];
  assign o[12800] = i[50];
  assign o[12801] = i[50];
  assign o[12802] = i[50];
  assign o[12803] = i[50];
  assign o[12804] = i[50];
  assign o[12805] = i[50];
  assign o[12806] = i[50];
  assign o[12807] = i[50];
  assign o[12808] = i[50];
  assign o[12809] = i[50];
  assign o[12810] = i[50];
  assign o[12811] = i[50];
  assign o[12812] = i[50];
  assign o[12813] = i[50];
  assign o[12814] = i[50];
  assign o[12815] = i[50];
  assign o[12816] = i[50];
  assign o[12817] = i[50];
  assign o[12818] = i[50];
  assign o[12819] = i[50];
  assign o[12820] = i[50];
  assign o[12821] = i[50];
  assign o[12822] = i[50];
  assign o[12823] = i[50];
  assign o[12824] = i[50];
  assign o[12825] = i[50];
  assign o[12826] = i[50];
  assign o[12827] = i[50];
  assign o[12828] = i[50];
  assign o[12829] = i[50];
  assign o[12830] = i[50];
  assign o[12831] = i[50];
  assign o[12832] = i[50];
  assign o[12833] = i[50];
  assign o[12834] = i[50];
  assign o[12835] = i[50];
  assign o[12836] = i[50];
  assign o[12837] = i[50];
  assign o[12838] = i[50];
  assign o[12839] = i[50];
  assign o[12840] = i[50];
  assign o[12841] = i[50];
  assign o[12842] = i[50];
  assign o[12843] = i[50];
  assign o[12844] = i[50];
  assign o[12845] = i[50];
  assign o[12846] = i[50];
  assign o[12847] = i[50];
  assign o[12848] = i[50];
  assign o[12849] = i[50];
  assign o[12850] = i[50];
  assign o[12851] = i[50];
  assign o[12852] = i[50];
  assign o[12853] = i[50];
  assign o[12854] = i[50];
  assign o[12855] = i[50];
  assign o[12856] = i[50];
  assign o[12857] = i[50];
  assign o[12858] = i[50];
  assign o[12859] = i[50];
  assign o[12860] = i[50];
  assign o[12861] = i[50];
  assign o[12862] = i[50];
  assign o[12863] = i[50];
  assign o[12864] = i[50];
  assign o[12865] = i[50];
  assign o[12866] = i[50];
  assign o[12867] = i[50];
  assign o[12868] = i[50];
  assign o[12869] = i[50];
  assign o[12870] = i[50];
  assign o[12871] = i[50];
  assign o[12872] = i[50];
  assign o[12873] = i[50];
  assign o[12874] = i[50];
  assign o[12875] = i[50];
  assign o[12876] = i[50];
  assign o[12877] = i[50];
  assign o[12878] = i[50];
  assign o[12879] = i[50];
  assign o[12880] = i[50];
  assign o[12881] = i[50];
  assign o[12882] = i[50];
  assign o[12883] = i[50];
  assign o[12884] = i[50];
  assign o[12885] = i[50];
  assign o[12886] = i[50];
  assign o[12887] = i[50];
  assign o[12888] = i[50];
  assign o[12889] = i[50];
  assign o[12890] = i[50];
  assign o[12891] = i[50];
  assign o[12892] = i[50];
  assign o[12893] = i[50];
  assign o[12894] = i[50];
  assign o[12895] = i[50];
  assign o[12896] = i[50];
  assign o[12897] = i[50];
  assign o[12898] = i[50];
  assign o[12899] = i[50];
  assign o[12900] = i[50];
  assign o[12901] = i[50];
  assign o[12902] = i[50];
  assign o[12903] = i[50];
  assign o[12904] = i[50];
  assign o[12905] = i[50];
  assign o[12906] = i[50];
  assign o[12907] = i[50];
  assign o[12908] = i[50];
  assign o[12909] = i[50];
  assign o[12910] = i[50];
  assign o[12911] = i[50];
  assign o[12912] = i[50];
  assign o[12913] = i[50];
  assign o[12914] = i[50];
  assign o[12915] = i[50];
  assign o[12916] = i[50];
  assign o[12917] = i[50];
  assign o[12918] = i[50];
  assign o[12919] = i[50];
  assign o[12920] = i[50];
  assign o[12921] = i[50];
  assign o[12922] = i[50];
  assign o[12923] = i[50];
  assign o[12924] = i[50];
  assign o[12925] = i[50];
  assign o[12926] = i[50];
  assign o[12927] = i[50];
  assign o[12928] = i[50];
  assign o[12929] = i[50];
  assign o[12930] = i[50];
  assign o[12931] = i[50];
  assign o[12932] = i[50];
  assign o[12933] = i[50];
  assign o[12934] = i[50];
  assign o[12935] = i[50];
  assign o[12936] = i[50];
  assign o[12937] = i[50];
  assign o[12938] = i[50];
  assign o[12939] = i[50];
  assign o[12940] = i[50];
  assign o[12941] = i[50];
  assign o[12942] = i[50];
  assign o[12943] = i[50];
  assign o[12944] = i[50];
  assign o[12945] = i[50];
  assign o[12946] = i[50];
  assign o[12947] = i[50];
  assign o[12948] = i[50];
  assign o[12949] = i[50];
  assign o[12950] = i[50];
  assign o[12951] = i[50];
  assign o[12952] = i[50];
  assign o[12953] = i[50];
  assign o[12954] = i[50];
  assign o[12955] = i[50];
  assign o[12956] = i[50];
  assign o[12957] = i[50];
  assign o[12958] = i[50];
  assign o[12959] = i[50];
  assign o[12960] = i[50];
  assign o[12961] = i[50];
  assign o[12962] = i[50];
  assign o[12963] = i[50];
  assign o[12964] = i[50];
  assign o[12965] = i[50];
  assign o[12966] = i[50];
  assign o[12967] = i[50];
  assign o[12968] = i[50];
  assign o[12969] = i[50];
  assign o[12970] = i[50];
  assign o[12971] = i[50];
  assign o[12972] = i[50];
  assign o[12973] = i[50];
  assign o[12974] = i[50];
  assign o[12975] = i[50];
  assign o[12976] = i[50];
  assign o[12977] = i[50];
  assign o[12978] = i[50];
  assign o[12979] = i[50];
  assign o[12980] = i[50];
  assign o[12981] = i[50];
  assign o[12982] = i[50];
  assign o[12983] = i[50];
  assign o[12984] = i[50];
  assign o[12985] = i[50];
  assign o[12986] = i[50];
  assign o[12987] = i[50];
  assign o[12988] = i[50];
  assign o[12989] = i[50];
  assign o[12990] = i[50];
  assign o[12991] = i[50];
  assign o[12992] = i[50];
  assign o[12993] = i[50];
  assign o[12994] = i[50];
  assign o[12995] = i[50];
  assign o[12996] = i[50];
  assign o[12997] = i[50];
  assign o[12998] = i[50];
  assign o[12999] = i[50];
  assign o[13000] = i[50];
  assign o[13001] = i[50];
  assign o[13002] = i[50];
  assign o[13003] = i[50];
  assign o[13004] = i[50];
  assign o[13005] = i[50];
  assign o[13006] = i[50];
  assign o[13007] = i[50];
  assign o[13008] = i[50];
  assign o[13009] = i[50];
  assign o[13010] = i[50];
  assign o[13011] = i[50];
  assign o[13012] = i[50];
  assign o[13013] = i[50];
  assign o[13014] = i[50];
  assign o[13015] = i[50];
  assign o[13016] = i[50];
  assign o[13017] = i[50];
  assign o[13018] = i[50];
  assign o[13019] = i[50];
  assign o[13020] = i[50];
  assign o[13021] = i[50];
  assign o[13022] = i[50];
  assign o[13023] = i[50];
  assign o[13024] = i[50];
  assign o[13025] = i[50];
  assign o[13026] = i[50];
  assign o[13027] = i[50];
  assign o[13028] = i[50];
  assign o[13029] = i[50];
  assign o[13030] = i[50];
  assign o[13031] = i[50];
  assign o[13032] = i[50];
  assign o[13033] = i[50];
  assign o[13034] = i[50];
  assign o[13035] = i[50];
  assign o[13036] = i[50];
  assign o[13037] = i[50];
  assign o[13038] = i[50];
  assign o[13039] = i[50];
  assign o[13040] = i[50];
  assign o[13041] = i[50];
  assign o[13042] = i[50];
  assign o[13043] = i[50];
  assign o[13044] = i[50];
  assign o[13045] = i[50];
  assign o[13046] = i[50];
  assign o[13047] = i[50];
  assign o[13048] = i[50];
  assign o[13049] = i[50];
  assign o[13050] = i[50];
  assign o[13051] = i[50];
  assign o[13052] = i[50];
  assign o[13053] = i[50];
  assign o[13054] = i[50];
  assign o[13055] = i[50];
  assign o[12544] = i[49];
  assign o[12545] = i[49];
  assign o[12546] = i[49];
  assign o[12547] = i[49];
  assign o[12548] = i[49];
  assign o[12549] = i[49];
  assign o[12550] = i[49];
  assign o[12551] = i[49];
  assign o[12552] = i[49];
  assign o[12553] = i[49];
  assign o[12554] = i[49];
  assign o[12555] = i[49];
  assign o[12556] = i[49];
  assign o[12557] = i[49];
  assign o[12558] = i[49];
  assign o[12559] = i[49];
  assign o[12560] = i[49];
  assign o[12561] = i[49];
  assign o[12562] = i[49];
  assign o[12563] = i[49];
  assign o[12564] = i[49];
  assign o[12565] = i[49];
  assign o[12566] = i[49];
  assign o[12567] = i[49];
  assign o[12568] = i[49];
  assign o[12569] = i[49];
  assign o[12570] = i[49];
  assign o[12571] = i[49];
  assign o[12572] = i[49];
  assign o[12573] = i[49];
  assign o[12574] = i[49];
  assign o[12575] = i[49];
  assign o[12576] = i[49];
  assign o[12577] = i[49];
  assign o[12578] = i[49];
  assign o[12579] = i[49];
  assign o[12580] = i[49];
  assign o[12581] = i[49];
  assign o[12582] = i[49];
  assign o[12583] = i[49];
  assign o[12584] = i[49];
  assign o[12585] = i[49];
  assign o[12586] = i[49];
  assign o[12587] = i[49];
  assign o[12588] = i[49];
  assign o[12589] = i[49];
  assign o[12590] = i[49];
  assign o[12591] = i[49];
  assign o[12592] = i[49];
  assign o[12593] = i[49];
  assign o[12594] = i[49];
  assign o[12595] = i[49];
  assign o[12596] = i[49];
  assign o[12597] = i[49];
  assign o[12598] = i[49];
  assign o[12599] = i[49];
  assign o[12600] = i[49];
  assign o[12601] = i[49];
  assign o[12602] = i[49];
  assign o[12603] = i[49];
  assign o[12604] = i[49];
  assign o[12605] = i[49];
  assign o[12606] = i[49];
  assign o[12607] = i[49];
  assign o[12608] = i[49];
  assign o[12609] = i[49];
  assign o[12610] = i[49];
  assign o[12611] = i[49];
  assign o[12612] = i[49];
  assign o[12613] = i[49];
  assign o[12614] = i[49];
  assign o[12615] = i[49];
  assign o[12616] = i[49];
  assign o[12617] = i[49];
  assign o[12618] = i[49];
  assign o[12619] = i[49];
  assign o[12620] = i[49];
  assign o[12621] = i[49];
  assign o[12622] = i[49];
  assign o[12623] = i[49];
  assign o[12624] = i[49];
  assign o[12625] = i[49];
  assign o[12626] = i[49];
  assign o[12627] = i[49];
  assign o[12628] = i[49];
  assign o[12629] = i[49];
  assign o[12630] = i[49];
  assign o[12631] = i[49];
  assign o[12632] = i[49];
  assign o[12633] = i[49];
  assign o[12634] = i[49];
  assign o[12635] = i[49];
  assign o[12636] = i[49];
  assign o[12637] = i[49];
  assign o[12638] = i[49];
  assign o[12639] = i[49];
  assign o[12640] = i[49];
  assign o[12641] = i[49];
  assign o[12642] = i[49];
  assign o[12643] = i[49];
  assign o[12644] = i[49];
  assign o[12645] = i[49];
  assign o[12646] = i[49];
  assign o[12647] = i[49];
  assign o[12648] = i[49];
  assign o[12649] = i[49];
  assign o[12650] = i[49];
  assign o[12651] = i[49];
  assign o[12652] = i[49];
  assign o[12653] = i[49];
  assign o[12654] = i[49];
  assign o[12655] = i[49];
  assign o[12656] = i[49];
  assign o[12657] = i[49];
  assign o[12658] = i[49];
  assign o[12659] = i[49];
  assign o[12660] = i[49];
  assign o[12661] = i[49];
  assign o[12662] = i[49];
  assign o[12663] = i[49];
  assign o[12664] = i[49];
  assign o[12665] = i[49];
  assign o[12666] = i[49];
  assign o[12667] = i[49];
  assign o[12668] = i[49];
  assign o[12669] = i[49];
  assign o[12670] = i[49];
  assign o[12671] = i[49];
  assign o[12672] = i[49];
  assign o[12673] = i[49];
  assign o[12674] = i[49];
  assign o[12675] = i[49];
  assign o[12676] = i[49];
  assign o[12677] = i[49];
  assign o[12678] = i[49];
  assign o[12679] = i[49];
  assign o[12680] = i[49];
  assign o[12681] = i[49];
  assign o[12682] = i[49];
  assign o[12683] = i[49];
  assign o[12684] = i[49];
  assign o[12685] = i[49];
  assign o[12686] = i[49];
  assign o[12687] = i[49];
  assign o[12688] = i[49];
  assign o[12689] = i[49];
  assign o[12690] = i[49];
  assign o[12691] = i[49];
  assign o[12692] = i[49];
  assign o[12693] = i[49];
  assign o[12694] = i[49];
  assign o[12695] = i[49];
  assign o[12696] = i[49];
  assign o[12697] = i[49];
  assign o[12698] = i[49];
  assign o[12699] = i[49];
  assign o[12700] = i[49];
  assign o[12701] = i[49];
  assign o[12702] = i[49];
  assign o[12703] = i[49];
  assign o[12704] = i[49];
  assign o[12705] = i[49];
  assign o[12706] = i[49];
  assign o[12707] = i[49];
  assign o[12708] = i[49];
  assign o[12709] = i[49];
  assign o[12710] = i[49];
  assign o[12711] = i[49];
  assign o[12712] = i[49];
  assign o[12713] = i[49];
  assign o[12714] = i[49];
  assign o[12715] = i[49];
  assign o[12716] = i[49];
  assign o[12717] = i[49];
  assign o[12718] = i[49];
  assign o[12719] = i[49];
  assign o[12720] = i[49];
  assign o[12721] = i[49];
  assign o[12722] = i[49];
  assign o[12723] = i[49];
  assign o[12724] = i[49];
  assign o[12725] = i[49];
  assign o[12726] = i[49];
  assign o[12727] = i[49];
  assign o[12728] = i[49];
  assign o[12729] = i[49];
  assign o[12730] = i[49];
  assign o[12731] = i[49];
  assign o[12732] = i[49];
  assign o[12733] = i[49];
  assign o[12734] = i[49];
  assign o[12735] = i[49];
  assign o[12736] = i[49];
  assign o[12737] = i[49];
  assign o[12738] = i[49];
  assign o[12739] = i[49];
  assign o[12740] = i[49];
  assign o[12741] = i[49];
  assign o[12742] = i[49];
  assign o[12743] = i[49];
  assign o[12744] = i[49];
  assign o[12745] = i[49];
  assign o[12746] = i[49];
  assign o[12747] = i[49];
  assign o[12748] = i[49];
  assign o[12749] = i[49];
  assign o[12750] = i[49];
  assign o[12751] = i[49];
  assign o[12752] = i[49];
  assign o[12753] = i[49];
  assign o[12754] = i[49];
  assign o[12755] = i[49];
  assign o[12756] = i[49];
  assign o[12757] = i[49];
  assign o[12758] = i[49];
  assign o[12759] = i[49];
  assign o[12760] = i[49];
  assign o[12761] = i[49];
  assign o[12762] = i[49];
  assign o[12763] = i[49];
  assign o[12764] = i[49];
  assign o[12765] = i[49];
  assign o[12766] = i[49];
  assign o[12767] = i[49];
  assign o[12768] = i[49];
  assign o[12769] = i[49];
  assign o[12770] = i[49];
  assign o[12771] = i[49];
  assign o[12772] = i[49];
  assign o[12773] = i[49];
  assign o[12774] = i[49];
  assign o[12775] = i[49];
  assign o[12776] = i[49];
  assign o[12777] = i[49];
  assign o[12778] = i[49];
  assign o[12779] = i[49];
  assign o[12780] = i[49];
  assign o[12781] = i[49];
  assign o[12782] = i[49];
  assign o[12783] = i[49];
  assign o[12784] = i[49];
  assign o[12785] = i[49];
  assign o[12786] = i[49];
  assign o[12787] = i[49];
  assign o[12788] = i[49];
  assign o[12789] = i[49];
  assign o[12790] = i[49];
  assign o[12791] = i[49];
  assign o[12792] = i[49];
  assign o[12793] = i[49];
  assign o[12794] = i[49];
  assign o[12795] = i[49];
  assign o[12796] = i[49];
  assign o[12797] = i[49];
  assign o[12798] = i[49];
  assign o[12799] = i[49];
  assign o[12288] = i[48];
  assign o[12289] = i[48];
  assign o[12290] = i[48];
  assign o[12291] = i[48];
  assign o[12292] = i[48];
  assign o[12293] = i[48];
  assign o[12294] = i[48];
  assign o[12295] = i[48];
  assign o[12296] = i[48];
  assign o[12297] = i[48];
  assign o[12298] = i[48];
  assign o[12299] = i[48];
  assign o[12300] = i[48];
  assign o[12301] = i[48];
  assign o[12302] = i[48];
  assign o[12303] = i[48];
  assign o[12304] = i[48];
  assign o[12305] = i[48];
  assign o[12306] = i[48];
  assign o[12307] = i[48];
  assign o[12308] = i[48];
  assign o[12309] = i[48];
  assign o[12310] = i[48];
  assign o[12311] = i[48];
  assign o[12312] = i[48];
  assign o[12313] = i[48];
  assign o[12314] = i[48];
  assign o[12315] = i[48];
  assign o[12316] = i[48];
  assign o[12317] = i[48];
  assign o[12318] = i[48];
  assign o[12319] = i[48];
  assign o[12320] = i[48];
  assign o[12321] = i[48];
  assign o[12322] = i[48];
  assign o[12323] = i[48];
  assign o[12324] = i[48];
  assign o[12325] = i[48];
  assign o[12326] = i[48];
  assign o[12327] = i[48];
  assign o[12328] = i[48];
  assign o[12329] = i[48];
  assign o[12330] = i[48];
  assign o[12331] = i[48];
  assign o[12332] = i[48];
  assign o[12333] = i[48];
  assign o[12334] = i[48];
  assign o[12335] = i[48];
  assign o[12336] = i[48];
  assign o[12337] = i[48];
  assign o[12338] = i[48];
  assign o[12339] = i[48];
  assign o[12340] = i[48];
  assign o[12341] = i[48];
  assign o[12342] = i[48];
  assign o[12343] = i[48];
  assign o[12344] = i[48];
  assign o[12345] = i[48];
  assign o[12346] = i[48];
  assign o[12347] = i[48];
  assign o[12348] = i[48];
  assign o[12349] = i[48];
  assign o[12350] = i[48];
  assign o[12351] = i[48];
  assign o[12352] = i[48];
  assign o[12353] = i[48];
  assign o[12354] = i[48];
  assign o[12355] = i[48];
  assign o[12356] = i[48];
  assign o[12357] = i[48];
  assign o[12358] = i[48];
  assign o[12359] = i[48];
  assign o[12360] = i[48];
  assign o[12361] = i[48];
  assign o[12362] = i[48];
  assign o[12363] = i[48];
  assign o[12364] = i[48];
  assign o[12365] = i[48];
  assign o[12366] = i[48];
  assign o[12367] = i[48];
  assign o[12368] = i[48];
  assign o[12369] = i[48];
  assign o[12370] = i[48];
  assign o[12371] = i[48];
  assign o[12372] = i[48];
  assign o[12373] = i[48];
  assign o[12374] = i[48];
  assign o[12375] = i[48];
  assign o[12376] = i[48];
  assign o[12377] = i[48];
  assign o[12378] = i[48];
  assign o[12379] = i[48];
  assign o[12380] = i[48];
  assign o[12381] = i[48];
  assign o[12382] = i[48];
  assign o[12383] = i[48];
  assign o[12384] = i[48];
  assign o[12385] = i[48];
  assign o[12386] = i[48];
  assign o[12387] = i[48];
  assign o[12388] = i[48];
  assign o[12389] = i[48];
  assign o[12390] = i[48];
  assign o[12391] = i[48];
  assign o[12392] = i[48];
  assign o[12393] = i[48];
  assign o[12394] = i[48];
  assign o[12395] = i[48];
  assign o[12396] = i[48];
  assign o[12397] = i[48];
  assign o[12398] = i[48];
  assign o[12399] = i[48];
  assign o[12400] = i[48];
  assign o[12401] = i[48];
  assign o[12402] = i[48];
  assign o[12403] = i[48];
  assign o[12404] = i[48];
  assign o[12405] = i[48];
  assign o[12406] = i[48];
  assign o[12407] = i[48];
  assign o[12408] = i[48];
  assign o[12409] = i[48];
  assign o[12410] = i[48];
  assign o[12411] = i[48];
  assign o[12412] = i[48];
  assign o[12413] = i[48];
  assign o[12414] = i[48];
  assign o[12415] = i[48];
  assign o[12416] = i[48];
  assign o[12417] = i[48];
  assign o[12418] = i[48];
  assign o[12419] = i[48];
  assign o[12420] = i[48];
  assign o[12421] = i[48];
  assign o[12422] = i[48];
  assign o[12423] = i[48];
  assign o[12424] = i[48];
  assign o[12425] = i[48];
  assign o[12426] = i[48];
  assign o[12427] = i[48];
  assign o[12428] = i[48];
  assign o[12429] = i[48];
  assign o[12430] = i[48];
  assign o[12431] = i[48];
  assign o[12432] = i[48];
  assign o[12433] = i[48];
  assign o[12434] = i[48];
  assign o[12435] = i[48];
  assign o[12436] = i[48];
  assign o[12437] = i[48];
  assign o[12438] = i[48];
  assign o[12439] = i[48];
  assign o[12440] = i[48];
  assign o[12441] = i[48];
  assign o[12442] = i[48];
  assign o[12443] = i[48];
  assign o[12444] = i[48];
  assign o[12445] = i[48];
  assign o[12446] = i[48];
  assign o[12447] = i[48];
  assign o[12448] = i[48];
  assign o[12449] = i[48];
  assign o[12450] = i[48];
  assign o[12451] = i[48];
  assign o[12452] = i[48];
  assign o[12453] = i[48];
  assign o[12454] = i[48];
  assign o[12455] = i[48];
  assign o[12456] = i[48];
  assign o[12457] = i[48];
  assign o[12458] = i[48];
  assign o[12459] = i[48];
  assign o[12460] = i[48];
  assign o[12461] = i[48];
  assign o[12462] = i[48];
  assign o[12463] = i[48];
  assign o[12464] = i[48];
  assign o[12465] = i[48];
  assign o[12466] = i[48];
  assign o[12467] = i[48];
  assign o[12468] = i[48];
  assign o[12469] = i[48];
  assign o[12470] = i[48];
  assign o[12471] = i[48];
  assign o[12472] = i[48];
  assign o[12473] = i[48];
  assign o[12474] = i[48];
  assign o[12475] = i[48];
  assign o[12476] = i[48];
  assign o[12477] = i[48];
  assign o[12478] = i[48];
  assign o[12479] = i[48];
  assign o[12480] = i[48];
  assign o[12481] = i[48];
  assign o[12482] = i[48];
  assign o[12483] = i[48];
  assign o[12484] = i[48];
  assign o[12485] = i[48];
  assign o[12486] = i[48];
  assign o[12487] = i[48];
  assign o[12488] = i[48];
  assign o[12489] = i[48];
  assign o[12490] = i[48];
  assign o[12491] = i[48];
  assign o[12492] = i[48];
  assign o[12493] = i[48];
  assign o[12494] = i[48];
  assign o[12495] = i[48];
  assign o[12496] = i[48];
  assign o[12497] = i[48];
  assign o[12498] = i[48];
  assign o[12499] = i[48];
  assign o[12500] = i[48];
  assign o[12501] = i[48];
  assign o[12502] = i[48];
  assign o[12503] = i[48];
  assign o[12504] = i[48];
  assign o[12505] = i[48];
  assign o[12506] = i[48];
  assign o[12507] = i[48];
  assign o[12508] = i[48];
  assign o[12509] = i[48];
  assign o[12510] = i[48];
  assign o[12511] = i[48];
  assign o[12512] = i[48];
  assign o[12513] = i[48];
  assign o[12514] = i[48];
  assign o[12515] = i[48];
  assign o[12516] = i[48];
  assign o[12517] = i[48];
  assign o[12518] = i[48];
  assign o[12519] = i[48];
  assign o[12520] = i[48];
  assign o[12521] = i[48];
  assign o[12522] = i[48];
  assign o[12523] = i[48];
  assign o[12524] = i[48];
  assign o[12525] = i[48];
  assign o[12526] = i[48];
  assign o[12527] = i[48];
  assign o[12528] = i[48];
  assign o[12529] = i[48];
  assign o[12530] = i[48];
  assign o[12531] = i[48];
  assign o[12532] = i[48];
  assign o[12533] = i[48];
  assign o[12534] = i[48];
  assign o[12535] = i[48];
  assign o[12536] = i[48];
  assign o[12537] = i[48];
  assign o[12538] = i[48];
  assign o[12539] = i[48];
  assign o[12540] = i[48];
  assign o[12541] = i[48];
  assign o[12542] = i[48];
  assign o[12543] = i[48];
  assign o[12032] = i[47];
  assign o[12033] = i[47];
  assign o[12034] = i[47];
  assign o[12035] = i[47];
  assign o[12036] = i[47];
  assign o[12037] = i[47];
  assign o[12038] = i[47];
  assign o[12039] = i[47];
  assign o[12040] = i[47];
  assign o[12041] = i[47];
  assign o[12042] = i[47];
  assign o[12043] = i[47];
  assign o[12044] = i[47];
  assign o[12045] = i[47];
  assign o[12046] = i[47];
  assign o[12047] = i[47];
  assign o[12048] = i[47];
  assign o[12049] = i[47];
  assign o[12050] = i[47];
  assign o[12051] = i[47];
  assign o[12052] = i[47];
  assign o[12053] = i[47];
  assign o[12054] = i[47];
  assign o[12055] = i[47];
  assign o[12056] = i[47];
  assign o[12057] = i[47];
  assign o[12058] = i[47];
  assign o[12059] = i[47];
  assign o[12060] = i[47];
  assign o[12061] = i[47];
  assign o[12062] = i[47];
  assign o[12063] = i[47];
  assign o[12064] = i[47];
  assign o[12065] = i[47];
  assign o[12066] = i[47];
  assign o[12067] = i[47];
  assign o[12068] = i[47];
  assign o[12069] = i[47];
  assign o[12070] = i[47];
  assign o[12071] = i[47];
  assign o[12072] = i[47];
  assign o[12073] = i[47];
  assign o[12074] = i[47];
  assign o[12075] = i[47];
  assign o[12076] = i[47];
  assign o[12077] = i[47];
  assign o[12078] = i[47];
  assign o[12079] = i[47];
  assign o[12080] = i[47];
  assign o[12081] = i[47];
  assign o[12082] = i[47];
  assign o[12083] = i[47];
  assign o[12084] = i[47];
  assign o[12085] = i[47];
  assign o[12086] = i[47];
  assign o[12087] = i[47];
  assign o[12088] = i[47];
  assign o[12089] = i[47];
  assign o[12090] = i[47];
  assign o[12091] = i[47];
  assign o[12092] = i[47];
  assign o[12093] = i[47];
  assign o[12094] = i[47];
  assign o[12095] = i[47];
  assign o[12096] = i[47];
  assign o[12097] = i[47];
  assign o[12098] = i[47];
  assign o[12099] = i[47];
  assign o[12100] = i[47];
  assign o[12101] = i[47];
  assign o[12102] = i[47];
  assign o[12103] = i[47];
  assign o[12104] = i[47];
  assign o[12105] = i[47];
  assign o[12106] = i[47];
  assign o[12107] = i[47];
  assign o[12108] = i[47];
  assign o[12109] = i[47];
  assign o[12110] = i[47];
  assign o[12111] = i[47];
  assign o[12112] = i[47];
  assign o[12113] = i[47];
  assign o[12114] = i[47];
  assign o[12115] = i[47];
  assign o[12116] = i[47];
  assign o[12117] = i[47];
  assign o[12118] = i[47];
  assign o[12119] = i[47];
  assign o[12120] = i[47];
  assign o[12121] = i[47];
  assign o[12122] = i[47];
  assign o[12123] = i[47];
  assign o[12124] = i[47];
  assign o[12125] = i[47];
  assign o[12126] = i[47];
  assign o[12127] = i[47];
  assign o[12128] = i[47];
  assign o[12129] = i[47];
  assign o[12130] = i[47];
  assign o[12131] = i[47];
  assign o[12132] = i[47];
  assign o[12133] = i[47];
  assign o[12134] = i[47];
  assign o[12135] = i[47];
  assign o[12136] = i[47];
  assign o[12137] = i[47];
  assign o[12138] = i[47];
  assign o[12139] = i[47];
  assign o[12140] = i[47];
  assign o[12141] = i[47];
  assign o[12142] = i[47];
  assign o[12143] = i[47];
  assign o[12144] = i[47];
  assign o[12145] = i[47];
  assign o[12146] = i[47];
  assign o[12147] = i[47];
  assign o[12148] = i[47];
  assign o[12149] = i[47];
  assign o[12150] = i[47];
  assign o[12151] = i[47];
  assign o[12152] = i[47];
  assign o[12153] = i[47];
  assign o[12154] = i[47];
  assign o[12155] = i[47];
  assign o[12156] = i[47];
  assign o[12157] = i[47];
  assign o[12158] = i[47];
  assign o[12159] = i[47];
  assign o[12160] = i[47];
  assign o[12161] = i[47];
  assign o[12162] = i[47];
  assign o[12163] = i[47];
  assign o[12164] = i[47];
  assign o[12165] = i[47];
  assign o[12166] = i[47];
  assign o[12167] = i[47];
  assign o[12168] = i[47];
  assign o[12169] = i[47];
  assign o[12170] = i[47];
  assign o[12171] = i[47];
  assign o[12172] = i[47];
  assign o[12173] = i[47];
  assign o[12174] = i[47];
  assign o[12175] = i[47];
  assign o[12176] = i[47];
  assign o[12177] = i[47];
  assign o[12178] = i[47];
  assign o[12179] = i[47];
  assign o[12180] = i[47];
  assign o[12181] = i[47];
  assign o[12182] = i[47];
  assign o[12183] = i[47];
  assign o[12184] = i[47];
  assign o[12185] = i[47];
  assign o[12186] = i[47];
  assign o[12187] = i[47];
  assign o[12188] = i[47];
  assign o[12189] = i[47];
  assign o[12190] = i[47];
  assign o[12191] = i[47];
  assign o[12192] = i[47];
  assign o[12193] = i[47];
  assign o[12194] = i[47];
  assign o[12195] = i[47];
  assign o[12196] = i[47];
  assign o[12197] = i[47];
  assign o[12198] = i[47];
  assign o[12199] = i[47];
  assign o[12200] = i[47];
  assign o[12201] = i[47];
  assign o[12202] = i[47];
  assign o[12203] = i[47];
  assign o[12204] = i[47];
  assign o[12205] = i[47];
  assign o[12206] = i[47];
  assign o[12207] = i[47];
  assign o[12208] = i[47];
  assign o[12209] = i[47];
  assign o[12210] = i[47];
  assign o[12211] = i[47];
  assign o[12212] = i[47];
  assign o[12213] = i[47];
  assign o[12214] = i[47];
  assign o[12215] = i[47];
  assign o[12216] = i[47];
  assign o[12217] = i[47];
  assign o[12218] = i[47];
  assign o[12219] = i[47];
  assign o[12220] = i[47];
  assign o[12221] = i[47];
  assign o[12222] = i[47];
  assign o[12223] = i[47];
  assign o[12224] = i[47];
  assign o[12225] = i[47];
  assign o[12226] = i[47];
  assign o[12227] = i[47];
  assign o[12228] = i[47];
  assign o[12229] = i[47];
  assign o[12230] = i[47];
  assign o[12231] = i[47];
  assign o[12232] = i[47];
  assign o[12233] = i[47];
  assign o[12234] = i[47];
  assign o[12235] = i[47];
  assign o[12236] = i[47];
  assign o[12237] = i[47];
  assign o[12238] = i[47];
  assign o[12239] = i[47];
  assign o[12240] = i[47];
  assign o[12241] = i[47];
  assign o[12242] = i[47];
  assign o[12243] = i[47];
  assign o[12244] = i[47];
  assign o[12245] = i[47];
  assign o[12246] = i[47];
  assign o[12247] = i[47];
  assign o[12248] = i[47];
  assign o[12249] = i[47];
  assign o[12250] = i[47];
  assign o[12251] = i[47];
  assign o[12252] = i[47];
  assign o[12253] = i[47];
  assign o[12254] = i[47];
  assign o[12255] = i[47];
  assign o[12256] = i[47];
  assign o[12257] = i[47];
  assign o[12258] = i[47];
  assign o[12259] = i[47];
  assign o[12260] = i[47];
  assign o[12261] = i[47];
  assign o[12262] = i[47];
  assign o[12263] = i[47];
  assign o[12264] = i[47];
  assign o[12265] = i[47];
  assign o[12266] = i[47];
  assign o[12267] = i[47];
  assign o[12268] = i[47];
  assign o[12269] = i[47];
  assign o[12270] = i[47];
  assign o[12271] = i[47];
  assign o[12272] = i[47];
  assign o[12273] = i[47];
  assign o[12274] = i[47];
  assign o[12275] = i[47];
  assign o[12276] = i[47];
  assign o[12277] = i[47];
  assign o[12278] = i[47];
  assign o[12279] = i[47];
  assign o[12280] = i[47];
  assign o[12281] = i[47];
  assign o[12282] = i[47];
  assign o[12283] = i[47];
  assign o[12284] = i[47];
  assign o[12285] = i[47];
  assign o[12286] = i[47];
  assign o[12287] = i[47];
  assign o[11776] = i[46];
  assign o[11777] = i[46];
  assign o[11778] = i[46];
  assign o[11779] = i[46];
  assign o[11780] = i[46];
  assign o[11781] = i[46];
  assign o[11782] = i[46];
  assign o[11783] = i[46];
  assign o[11784] = i[46];
  assign o[11785] = i[46];
  assign o[11786] = i[46];
  assign o[11787] = i[46];
  assign o[11788] = i[46];
  assign o[11789] = i[46];
  assign o[11790] = i[46];
  assign o[11791] = i[46];
  assign o[11792] = i[46];
  assign o[11793] = i[46];
  assign o[11794] = i[46];
  assign o[11795] = i[46];
  assign o[11796] = i[46];
  assign o[11797] = i[46];
  assign o[11798] = i[46];
  assign o[11799] = i[46];
  assign o[11800] = i[46];
  assign o[11801] = i[46];
  assign o[11802] = i[46];
  assign o[11803] = i[46];
  assign o[11804] = i[46];
  assign o[11805] = i[46];
  assign o[11806] = i[46];
  assign o[11807] = i[46];
  assign o[11808] = i[46];
  assign o[11809] = i[46];
  assign o[11810] = i[46];
  assign o[11811] = i[46];
  assign o[11812] = i[46];
  assign o[11813] = i[46];
  assign o[11814] = i[46];
  assign o[11815] = i[46];
  assign o[11816] = i[46];
  assign o[11817] = i[46];
  assign o[11818] = i[46];
  assign o[11819] = i[46];
  assign o[11820] = i[46];
  assign o[11821] = i[46];
  assign o[11822] = i[46];
  assign o[11823] = i[46];
  assign o[11824] = i[46];
  assign o[11825] = i[46];
  assign o[11826] = i[46];
  assign o[11827] = i[46];
  assign o[11828] = i[46];
  assign o[11829] = i[46];
  assign o[11830] = i[46];
  assign o[11831] = i[46];
  assign o[11832] = i[46];
  assign o[11833] = i[46];
  assign o[11834] = i[46];
  assign o[11835] = i[46];
  assign o[11836] = i[46];
  assign o[11837] = i[46];
  assign o[11838] = i[46];
  assign o[11839] = i[46];
  assign o[11840] = i[46];
  assign o[11841] = i[46];
  assign o[11842] = i[46];
  assign o[11843] = i[46];
  assign o[11844] = i[46];
  assign o[11845] = i[46];
  assign o[11846] = i[46];
  assign o[11847] = i[46];
  assign o[11848] = i[46];
  assign o[11849] = i[46];
  assign o[11850] = i[46];
  assign o[11851] = i[46];
  assign o[11852] = i[46];
  assign o[11853] = i[46];
  assign o[11854] = i[46];
  assign o[11855] = i[46];
  assign o[11856] = i[46];
  assign o[11857] = i[46];
  assign o[11858] = i[46];
  assign o[11859] = i[46];
  assign o[11860] = i[46];
  assign o[11861] = i[46];
  assign o[11862] = i[46];
  assign o[11863] = i[46];
  assign o[11864] = i[46];
  assign o[11865] = i[46];
  assign o[11866] = i[46];
  assign o[11867] = i[46];
  assign o[11868] = i[46];
  assign o[11869] = i[46];
  assign o[11870] = i[46];
  assign o[11871] = i[46];
  assign o[11872] = i[46];
  assign o[11873] = i[46];
  assign o[11874] = i[46];
  assign o[11875] = i[46];
  assign o[11876] = i[46];
  assign o[11877] = i[46];
  assign o[11878] = i[46];
  assign o[11879] = i[46];
  assign o[11880] = i[46];
  assign o[11881] = i[46];
  assign o[11882] = i[46];
  assign o[11883] = i[46];
  assign o[11884] = i[46];
  assign o[11885] = i[46];
  assign o[11886] = i[46];
  assign o[11887] = i[46];
  assign o[11888] = i[46];
  assign o[11889] = i[46];
  assign o[11890] = i[46];
  assign o[11891] = i[46];
  assign o[11892] = i[46];
  assign o[11893] = i[46];
  assign o[11894] = i[46];
  assign o[11895] = i[46];
  assign o[11896] = i[46];
  assign o[11897] = i[46];
  assign o[11898] = i[46];
  assign o[11899] = i[46];
  assign o[11900] = i[46];
  assign o[11901] = i[46];
  assign o[11902] = i[46];
  assign o[11903] = i[46];
  assign o[11904] = i[46];
  assign o[11905] = i[46];
  assign o[11906] = i[46];
  assign o[11907] = i[46];
  assign o[11908] = i[46];
  assign o[11909] = i[46];
  assign o[11910] = i[46];
  assign o[11911] = i[46];
  assign o[11912] = i[46];
  assign o[11913] = i[46];
  assign o[11914] = i[46];
  assign o[11915] = i[46];
  assign o[11916] = i[46];
  assign o[11917] = i[46];
  assign o[11918] = i[46];
  assign o[11919] = i[46];
  assign o[11920] = i[46];
  assign o[11921] = i[46];
  assign o[11922] = i[46];
  assign o[11923] = i[46];
  assign o[11924] = i[46];
  assign o[11925] = i[46];
  assign o[11926] = i[46];
  assign o[11927] = i[46];
  assign o[11928] = i[46];
  assign o[11929] = i[46];
  assign o[11930] = i[46];
  assign o[11931] = i[46];
  assign o[11932] = i[46];
  assign o[11933] = i[46];
  assign o[11934] = i[46];
  assign o[11935] = i[46];
  assign o[11936] = i[46];
  assign o[11937] = i[46];
  assign o[11938] = i[46];
  assign o[11939] = i[46];
  assign o[11940] = i[46];
  assign o[11941] = i[46];
  assign o[11942] = i[46];
  assign o[11943] = i[46];
  assign o[11944] = i[46];
  assign o[11945] = i[46];
  assign o[11946] = i[46];
  assign o[11947] = i[46];
  assign o[11948] = i[46];
  assign o[11949] = i[46];
  assign o[11950] = i[46];
  assign o[11951] = i[46];
  assign o[11952] = i[46];
  assign o[11953] = i[46];
  assign o[11954] = i[46];
  assign o[11955] = i[46];
  assign o[11956] = i[46];
  assign o[11957] = i[46];
  assign o[11958] = i[46];
  assign o[11959] = i[46];
  assign o[11960] = i[46];
  assign o[11961] = i[46];
  assign o[11962] = i[46];
  assign o[11963] = i[46];
  assign o[11964] = i[46];
  assign o[11965] = i[46];
  assign o[11966] = i[46];
  assign o[11967] = i[46];
  assign o[11968] = i[46];
  assign o[11969] = i[46];
  assign o[11970] = i[46];
  assign o[11971] = i[46];
  assign o[11972] = i[46];
  assign o[11973] = i[46];
  assign o[11974] = i[46];
  assign o[11975] = i[46];
  assign o[11976] = i[46];
  assign o[11977] = i[46];
  assign o[11978] = i[46];
  assign o[11979] = i[46];
  assign o[11980] = i[46];
  assign o[11981] = i[46];
  assign o[11982] = i[46];
  assign o[11983] = i[46];
  assign o[11984] = i[46];
  assign o[11985] = i[46];
  assign o[11986] = i[46];
  assign o[11987] = i[46];
  assign o[11988] = i[46];
  assign o[11989] = i[46];
  assign o[11990] = i[46];
  assign o[11991] = i[46];
  assign o[11992] = i[46];
  assign o[11993] = i[46];
  assign o[11994] = i[46];
  assign o[11995] = i[46];
  assign o[11996] = i[46];
  assign o[11997] = i[46];
  assign o[11998] = i[46];
  assign o[11999] = i[46];
  assign o[12000] = i[46];
  assign o[12001] = i[46];
  assign o[12002] = i[46];
  assign o[12003] = i[46];
  assign o[12004] = i[46];
  assign o[12005] = i[46];
  assign o[12006] = i[46];
  assign o[12007] = i[46];
  assign o[12008] = i[46];
  assign o[12009] = i[46];
  assign o[12010] = i[46];
  assign o[12011] = i[46];
  assign o[12012] = i[46];
  assign o[12013] = i[46];
  assign o[12014] = i[46];
  assign o[12015] = i[46];
  assign o[12016] = i[46];
  assign o[12017] = i[46];
  assign o[12018] = i[46];
  assign o[12019] = i[46];
  assign o[12020] = i[46];
  assign o[12021] = i[46];
  assign o[12022] = i[46];
  assign o[12023] = i[46];
  assign o[12024] = i[46];
  assign o[12025] = i[46];
  assign o[12026] = i[46];
  assign o[12027] = i[46];
  assign o[12028] = i[46];
  assign o[12029] = i[46];
  assign o[12030] = i[46];
  assign o[12031] = i[46];
  assign o[11520] = i[45];
  assign o[11521] = i[45];
  assign o[11522] = i[45];
  assign o[11523] = i[45];
  assign o[11524] = i[45];
  assign o[11525] = i[45];
  assign o[11526] = i[45];
  assign o[11527] = i[45];
  assign o[11528] = i[45];
  assign o[11529] = i[45];
  assign o[11530] = i[45];
  assign o[11531] = i[45];
  assign o[11532] = i[45];
  assign o[11533] = i[45];
  assign o[11534] = i[45];
  assign o[11535] = i[45];
  assign o[11536] = i[45];
  assign o[11537] = i[45];
  assign o[11538] = i[45];
  assign o[11539] = i[45];
  assign o[11540] = i[45];
  assign o[11541] = i[45];
  assign o[11542] = i[45];
  assign o[11543] = i[45];
  assign o[11544] = i[45];
  assign o[11545] = i[45];
  assign o[11546] = i[45];
  assign o[11547] = i[45];
  assign o[11548] = i[45];
  assign o[11549] = i[45];
  assign o[11550] = i[45];
  assign o[11551] = i[45];
  assign o[11552] = i[45];
  assign o[11553] = i[45];
  assign o[11554] = i[45];
  assign o[11555] = i[45];
  assign o[11556] = i[45];
  assign o[11557] = i[45];
  assign o[11558] = i[45];
  assign o[11559] = i[45];
  assign o[11560] = i[45];
  assign o[11561] = i[45];
  assign o[11562] = i[45];
  assign o[11563] = i[45];
  assign o[11564] = i[45];
  assign o[11565] = i[45];
  assign o[11566] = i[45];
  assign o[11567] = i[45];
  assign o[11568] = i[45];
  assign o[11569] = i[45];
  assign o[11570] = i[45];
  assign o[11571] = i[45];
  assign o[11572] = i[45];
  assign o[11573] = i[45];
  assign o[11574] = i[45];
  assign o[11575] = i[45];
  assign o[11576] = i[45];
  assign o[11577] = i[45];
  assign o[11578] = i[45];
  assign o[11579] = i[45];
  assign o[11580] = i[45];
  assign o[11581] = i[45];
  assign o[11582] = i[45];
  assign o[11583] = i[45];
  assign o[11584] = i[45];
  assign o[11585] = i[45];
  assign o[11586] = i[45];
  assign o[11587] = i[45];
  assign o[11588] = i[45];
  assign o[11589] = i[45];
  assign o[11590] = i[45];
  assign o[11591] = i[45];
  assign o[11592] = i[45];
  assign o[11593] = i[45];
  assign o[11594] = i[45];
  assign o[11595] = i[45];
  assign o[11596] = i[45];
  assign o[11597] = i[45];
  assign o[11598] = i[45];
  assign o[11599] = i[45];
  assign o[11600] = i[45];
  assign o[11601] = i[45];
  assign o[11602] = i[45];
  assign o[11603] = i[45];
  assign o[11604] = i[45];
  assign o[11605] = i[45];
  assign o[11606] = i[45];
  assign o[11607] = i[45];
  assign o[11608] = i[45];
  assign o[11609] = i[45];
  assign o[11610] = i[45];
  assign o[11611] = i[45];
  assign o[11612] = i[45];
  assign o[11613] = i[45];
  assign o[11614] = i[45];
  assign o[11615] = i[45];
  assign o[11616] = i[45];
  assign o[11617] = i[45];
  assign o[11618] = i[45];
  assign o[11619] = i[45];
  assign o[11620] = i[45];
  assign o[11621] = i[45];
  assign o[11622] = i[45];
  assign o[11623] = i[45];
  assign o[11624] = i[45];
  assign o[11625] = i[45];
  assign o[11626] = i[45];
  assign o[11627] = i[45];
  assign o[11628] = i[45];
  assign o[11629] = i[45];
  assign o[11630] = i[45];
  assign o[11631] = i[45];
  assign o[11632] = i[45];
  assign o[11633] = i[45];
  assign o[11634] = i[45];
  assign o[11635] = i[45];
  assign o[11636] = i[45];
  assign o[11637] = i[45];
  assign o[11638] = i[45];
  assign o[11639] = i[45];
  assign o[11640] = i[45];
  assign o[11641] = i[45];
  assign o[11642] = i[45];
  assign o[11643] = i[45];
  assign o[11644] = i[45];
  assign o[11645] = i[45];
  assign o[11646] = i[45];
  assign o[11647] = i[45];
  assign o[11648] = i[45];
  assign o[11649] = i[45];
  assign o[11650] = i[45];
  assign o[11651] = i[45];
  assign o[11652] = i[45];
  assign o[11653] = i[45];
  assign o[11654] = i[45];
  assign o[11655] = i[45];
  assign o[11656] = i[45];
  assign o[11657] = i[45];
  assign o[11658] = i[45];
  assign o[11659] = i[45];
  assign o[11660] = i[45];
  assign o[11661] = i[45];
  assign o[11662] = i[45];
  assign o[11663] = i[45];
  assign o[11664] = i[45];
  assign o[11665] = i[45];
  assign o[11666] = i[45];
  assign o[11667] = i[45];
  assign o[11668] = i[45];
  assign o[11669] = i[45];
  assign o[11670] = i[45];
  assign o[11671] = i[45];
  assign o[11672] = i[45];
  assign o[11673] = i[45];
  assign o[11674] = i[45];
  assign o[11675] = i[45];
  assign o[11676] = i[45];
  assign o[11677] = i[45];
  assign o[11678] = i[45];
  assign o[11679] = i[45];
  assign o[11680] = i[45];
  assign o[11681] = i[45];
  assign o[11682] = i[45];
  assign o[11683] = i[45];
  assign o[11684] = i[45];
  assign o[11685] = i[45];
  assign o[11686] = i[45];
  assign o[11687] = i[45];
  assign o[11688] = i[45];
  assign o[11689] = i[45];
  assign o[11690] = i[45];
  assign o[11691] = i[45];
  assign o[11692] = i[45];
  assign o[11693] = i[45];
  assign o[11694] = i[45];
  assign o[11695] = i[45];
  assign o[11696] = i[45];
  assign o[11697] = i[45];
  assign o[11698] = i[45];
  assign o[11699] = i[45];
  assign o[11700] = i[45];
  assign o[11701] = i[45];
  assign o[11702] = i[45];
  assign o[11703] = i[45];
  assign o[11704] = i[45];
  assign o[11705] = i[45];
  assign o[11706] = i[45];
  assign o[11707] = i[45];
  assign o[11708] = i[45];
  assign o[11709] = i[45];
  assign o[11710] = i[45];
  assign o[11711] = i[45];
  assign o[11712] = i[45];
  assign o[11713] = i[45];
  assign o[11714] = i[45];
  assign o[11715] = i[45];
  assign o[11716] = i[45];
  assign o[11717] = i[45];
  assign o[11718] = i[45];
  assign o[11719] = i[45];
  assign o[11720] = i[45];
  assign o[11721] = i[45];
  assign o[11722] = i[45];
  assign o[11723] = i[45];
  assign o[11724] = i[45];
  assign o[11725] = i[45];
  assign o[11726] = i[45];
  assign o[11727] = i[45];
  assign o[11728] = i[45];
  assign o[11729] = i[45];
  assign o[11730] = i[45];
  assign o[11731] = i[45];
  assign o[11732] = i[45];
  assign o[11733] = i[45];
  assign o[11734] = i[45];
  assign o[11735] = i[45];
  assign o[11736] = i[45];
  assign o[11737] = i[45];
  assign o[11738] = i[45];
  assign o[11739] = i[45];
  assign o[11740] = i[45];
  assign o[11741] = i[45];
  assign o[11742] = i[45];
  assign o[11743] = i[45];
  assign o[11744] = i[45];
  assign o[11745] = i[45];
  assign o[11746] = i[45];
  assign o[11747] = i[45];
  assign o[11748] = i[45];
  assign o[11749] = i[45];
  assign o[11750] = i[45];
  assign o[11751] = i[45];
  assign o[11752] = i[45];
  assign o[11753] = i[45];
  assign o[11754] = i[45];
  assign o[11755] = i[45];
  assign o[11756] = i[45];
  assign o[11757] = i[45];
  assign o[11758] = i[45];
  assign o[11759] = i[45];
  assign o[11760] = i[45];
  assign o[11761] = i[45];
  assign o[11762] = i[45];
  assign o[11763] = i[45];
  assign o[11764] = i[45];
  assign o[11765] = i[45];
  assign o[11766] = i[45];
  assign o[11767] = i[45];
  assign o[11768] = i[45];
  assign o[11769] = i[45];
  assign o[11770] = i[45];
  assign o[11771] = i[45];
  assign o[11772] = i[45];
  assign o[11773] = i[45];
  assign o[11774] = i[45];
  assign o[11775] = i[45];
  assign o[11264] = i[44];
  assign o[11265] = i[44];
  assign o[11266] = i[44];
  assign o[11267] = i[44];
  assign o[11268] = i[44];
  assign o[11269] = i[44];
  assign o[11270] = i[44];
  assign o[11271] = i[44];
  assign o[11272] = i[44];
  assign o[11273] = i[44];
  assign o[11274] = i[44];
  assign o[11275] = i[44];
  assign o[11276] = i[44];
  assign o[11277] = i[44];
  assign o[11278] = i[44];
  assign o[11279] = i[44];
  assign o[11280] = i[44];
  assign o[11281] = i[44];
  assign o[11282] = i[44];
  assign o[11283] = i[44];
  assign o[11284] = i[44];
  assign o[11285] = i[44];
  assign o[11286] = i[44];
  assign o[11287] = i[44];
  assign o[11288] = i[44];
  assign o[11289] = i[44];
  assign o[11290] = i[44];
  assign o[11291] = i[44];
  assign o[11292] = i[44];
  assign o[11293] = i[44];
  assign o[11294] = i[44];
  assign o[11295] = i[44];
  assign o[11296] = i[44];
  assign o[11297] = i[44];
  assign o[11298] = i[44];
  assign o[11299] = i[44];
  assign o[11300] = i[44];
  assign o[11301] = i[44];
  assign o[11302] = i[44];
  assign o[11303] = i[44];
  assign o[11304] = i[44];
  assign o[11305] = i[44];
  assign o[11306] = i[44];
  assign o[11307] = i[44];
  assign o[11308] = i[44];
  assign o[11309] = i[44];
  assign o[11310] = i[44];
  assign o[11311] = i[44];
  assign o[11312] = i[44];
  assign o[11313] = i[44];
  assign o[11314] = i[44];
  assign o[11315] = i[44];
  assign o[11316] = i[44];
  assign o[11317] = i[44];
  assign o[11318] = i[44];
  assign o[11319] = i[44];
  assign o[11320] = i[44];
  assign o[11321] = i[44];
  assign o[11322] = i[44];
  assign o[11323] = i[44];
  assign o[11324] = i[44];
  assign o[11325] = i[44];
  assign o[11326] = i[44];
  assign o[11327] = i[44];
  assign o[11328] = i[44];
  assign o[11329] = i[44];
  assign o[11330] = i[44];
  assign o[11331] = i[44];
  assign o[11332] = i[44];
  assign o[11333] = i[44];
  assign o[11334] = i[44];
  assign o[11335] = i[44];
  assign o[11336] = i[44];
  assign o[11337] = i[44];
  assign o[11338] = i[44];
  assign o[11339] = i[44];
  assign o[11340] = i[44];
  assign o[11341] = i[44];
  assign o[11342] = i[44];
  assign o[11343] = i[44];
  assign o[11344] = i[44];
  assign o[11345] = i[44];
  assign o[11346] = i[44];
  assign o[11347] = i[44];
  assign o[11348] = i[44];
  assign o[11349] = i[44];
  assign o[11350] = i[44];
  assign o[11351] = i[44];
  assign o[11352] = i[44];
  assign o[11353] = i[44];
  assign o[11354] = i[44];
  assign o[11355] = i[44];
  assign o[11356] = i[44];
  assign o[11357] = i[44];
  assign o[11358] = i[44];
  assign o[11359] = i[44];
  assign o[11360] = i[44];
  assign o[11361] = i[44];
  assign o[11362] = i[44];
  assign o[11363] = i[44];
  assign o[11364] = i[44];
  assign o[11365] = i[44];
  assign o[11366] = i[44];
  assign o[11367] = i[44];
  assign o[11368] = i[44];
  assign o[11369] = i[44];
  assign o[11370] = i[44];
  assign o[11371] = i[44];
  assign o[11372] = i[44];
  assign o[11373] = i[44];
  assign o[11374] = i[44];
  assign o[11375] = i[44];
  assign o[11376] = i[44];
  assign o[11377] = i[44];
  assign o[11378] = i[44];
  assign o[11379] = i[44];
  assign o[11380] = i[44];
  assign o[11381] = i[44];
  assign o[11382] = i[44];
  assign o[11383] = i[44];
  assign o[11384] = i[44];
  assign o[11385] = i[44];
  assign o[11386] = i[44];
  assign o[11387] = i[44];
  assign o[11388] = i[44];
  assign o[11389] = i[44];
  assign o[11390] = i[44];
  assign o[11391] = i[44];
  assign o[11392] = i[44];
  assign o[11393] = i[44];
  assign o[11394] = i[44];
  assign o[11395] = i[44];
  assign o[11396] = i[44];
  assign o[11397] = i[44];
  assign o[11398] = i[44];
  assign o[11399] = i[44];
  assign o[11400] = i[44];
  assign o[11401] = i[44];
  assign o[11402] = i[44];
  assign o[11403] = i[44];
  assign o[11404] = i[44];
  assign o[11405] = i[44];
  assign o[11406] = i[44];
  assign o[11407] = i[44];
  assign o[11408] = i[44];
  assign o[11409] = i[44];
  assign o[11410] = i[44];
  assign o[11411] = i[44];
  assign o[11412] = i[44];
  assign o[11413] = i[44];
  assign o[11414] = i[44];
  assign o[11415] = i[44];
  assign o[11416] = i[44];
  assign o[11417] = i[44];
  assign o[11418] = i[44];
  assign o[11419] = i[44];
  assign o[11420] = i[44];
  assign o[11421] = i[44];
  assign o[11422] = i[44];
  assign o[11423] = i[44];
  assign o[11424] = i[44];
  assign o[11425] = i[44];
  assign o[11426] = i[44];
  assign o[11427] = i[44];
  assign o[11428] = i[44];
  assign o[11429] = i[44];
  assign o[11430] = i[44];
  assign o[11431] = i[44];
  assign o[11432] = i[44];
  assign o[11433] = i[44];
  assign o[11434] = i[44];
  assign o[11435] = i[44];
  assign o[11436] = i[44];
  assign o[11437] = i[44];
  assign o[11438] = i[44];
  assign o[11439] = i[44];
  assign o[11440] = i[44];
  assign o[11441] = i[44];
  assign o[11442] = i[44];
  assign o[11443] = i[44];
  assign o[11444] = i[44];
  assign o[11445] = i[44];
  assign o[11446] = i[44];
  assign o[11447] = i[44];
  assign o[11448] = i[44];
  assign o[11449] = i[44];
  assign o[11450] = i[44];
  assign o[11451] = i[44];
  assign o[11452] = i[44];
  assign o[11453] = i[44];
  assign o[11454] = i[44];
  assign o[11455] = i[44];
  assign o[11456] = i[44];
  assign o[11457] = i[44];
  assign o[11458] = i[44];
  assign o[11459] = i[44];
  assign o[11460] = i[44];
  assign o[11461] = i[44];
  assign o[11462] = i[44];
  assign o[11463] = i[44];
  assign o[11464] = i[44];
  assign o[11465] = i[44];
  assign o[11466] = i[44];
  assign o[11467] = i[44];
  assign o[11468] = i[44];
  assign o[11469] = i[44];
  assign o[11470] = i[44];
  assign o[11471] = i[44];
  assign o[11472] = i[44];
  assign o[11473] = i[44];
  assign o[11474] = i[44];
  assign o[11475] = i[44];
  assign o[11476] = i[44];
  assign o[11477] = i[44];
  assign o[11478] = i[44];
  assign o[11479] = i[44];
  assign o[11480] = i[44];
  assign o[11481] = i[44];
  assign o[11482] = i[44];
  assign o[11483] = i[44];
  assign o[11484] = i[44];
  assign o[11485] = i[44];
  assign o[11486] = i[44];
  assign o[11487] = i[44];
  assign o[11488] = i[44];
  assign o[11489] = i[44];
  assign o[11490] = i[44];
  assign o[11491] = i[44];
  assign o[11492] = i[44];
  assign o[11493] = i[44];
  assign o[11494] = i[44];
  assign o[11495] = i[44];
  assign o[11496] = i[44];
  assign o[11497] = i[44];
  assign o[11498] = i[44];
  assign o[11499] = i[44];
  assign o[11500] = i[44];
  assign o[11501] = i[44];
  assign o[11502] = i[44];
  assign o[11503] = i[44];
  assign o[11504] = i[44];
  assign o[11505] = i[44];
  assign o[11506] = i[44];
  assign o[11507] = i[44];
  assign o[11508] = i[44];
  assign o[11509] = i[44];
  assign o[11510] = i[44];
  assign o[11511] = i[44];
  assign o[11512] = i[44];
  assign o[11513] = i[44];
  assign o[11514] = i[44];
  assign o[11515] = i[44];
  assign o[11516] = i[44];
  assign o[11517] = i[44];
  assign o[11518] = i[44];
  assign o[11519] = i[44];
  assign o[11008] = i[43];
  assign o[11009] = i[43];
  assign o[11010] = i[43];
  assign o[11011] = i[43];
  assign o[11012] = i[43];
  assign o[11013] = i[43];
  assign o[11014] = i[43];
  assign o[11015] = i[43];
  assign o[11016] = i[43];
  assign o[11017] = i[43];
  assign o[11018] = i[43];
  assign o[11019] = i[43];
  assign o[11020] = i[43];
  assign o[11021] = i[43];
  assign o[11022] = i[43];
  assign o[11023] = i[43];
  assign o[11024] = i[43];
  assign o[11025] = i[43];
  assign o[11026] = i[43];
  assign o[11027] = i[43];
  assign o[11028] = i[43];
  assign o[11029] = i[43];
  assign o[11030] = i[43];
  assign o[11031] = i[43];
  assign o[11032] = i[43];
  assign o[11033] = i[43];
  assign o[11034] = i[43];
  assign o[11035] = i[43];
  assign o[11036] = i[43];
  assign o[11037] = i[43];
  assign o[11038] = i[43];
  assign o[11039] = i[43];
  assign o[11040] = i[43];
  assign o[11041] = i[43];
  assign o[11042] = i[43];
  assign o[11043] = i[43];
  assign o[11044] = i[43];
  assign o[11045] = i[43];
  assign o[11046] = i[43];
  assign o[11047] = i[43];
  assign o[11048] = i[43];
  assign o[11049] = i[43];
  assign o[11050] = i[43];
  assign o[11051] = i[43];
  assign o[11052] = i[43];
  assign o[11053] = i[43];
  assign o[11054] = i[43];
  assign o[11055] = i[43];
  assign o[11056] = i[43];
  assign o[11057] = i[43];
  assign o[11058] = i[43];
  assign o[11059] = i[43];
  assign o[11060] = i[43];
  assign o[11061] = i[43];
  assign o[11062] = i[43];
  assign o[11063] = i[43];
  assign o[11064] = i[43];
  assign o[11065] = i[43];
  assign o[11066] = i[43];
  assign o[11067] = i[43];
  assign o[11068] = i[43];
  assign o[11069] = i[43];
  assign o[11070] = i[43];
  assign o[11071] = i[43];
  assign o[11072] = i[43];
  assign o[11073] = i[43];
  assign o[11074] = i[43];
  assign o[11075] = i[43];
  assign o[11076] = i[43];
  assign o[11077] = i[43];
  assign o[11078] = i[43];
  assign o[11079] = i[43];
  assign o[11080] = i[43];
  assign o[11081] = i[43];
  assign o[11082] = i[43];
  assign o[11083] = i[43];
  assign o[11084] = i[43];
  assign o[11085] = i[43];
  assign o[11086] = i[43];
  assign o[11087] = i[43];
  assign o[11088] = i[43];
  assign o[11089] = i[43];
  assign o[11090] = i[43];
  assign o[11091] = i[43];
  assign o[11092] = i[43];
  assign o[11093] = i[43];
  assign o[11094] = i[43];
  assign o[11095] = i[43];
  assign o[11096] = i[43];
  assign o[11097] = i[43];
  assign o[11098] = i[43];
  assign o[11099] = i[43];
  assign o[11100] = i[43];
  assign o[11101] = i[43];
  assign o[11102] = i[43];
  assign o[11103] = i[43];
  assign o[11104] = i[43];
  assign o[11105] = i[43];
  assign o[11106] = i[43];
  assign o[11107] = i[43];
  assign o[11108] = i[43];
  assign o[11109] = i[43];
  assign o[11110] = i[43];
  assign o[11111] = i[43];
  assign o[11112] = i[43];
  assign o[11113] = i[43];
  assign o[11114] = i[43];
  assign o[11115] = i[43];
  assign o[11116] = i[43];
  assign o[11117] = i[43];
  assign o[11118] = i[43];
  assign o[11119] = i[43];
  assign o[11120] = i[43];
  assign o[11121] = i[43];
  assign o[11122] = i[43];
  assign o[11123] = i[43];
  assign o[11124] = i[43];
  assign o[11125] = i[43];
  assign o[11126] = i[43];
  assign o[11127] = i[43];
  assign o[11128] = i[43];
  assign o[11129] = i[43];
  assign o[11130] = i[43];
  assign o[11131] = i[43];
  assign o[11132] = i[43];
  assign o[11133] = i[43];
  assign o[11134] = i[43];
  assign o[11135] = i[43];
  assign o[11136] = i[43];
  assign o[11137] = i[43];
  assign o[11138] = i[43];
  assign o[11139] = i[43];
  assign o[11140] = i[43];
  assign o[11141] = i[43];
  assign o[11142] = i[43];
  assign o[11143] = i[43];
  assign o[11144] = i[43];
  assign o[11145] = i[43];
  assign o[11146] = i[43];
  assign o[11147] = i[43];
  assign o[11148] = i[43];
  assign o[11149] = i[43];
  assign o[11150] = i[43];
  assign o[11151] = i[43];
  assign o[11152] = i[43];
  assign o[11153] = i[43];
  assign o[11154] = i[43];
  assign o[11155] = i[43];
  assign o[11156] = i[43];
  assign o[11157] = i[43];
  assign o[11158] = i[43];
  assign o[11159] = i[43];
  assign o[11160] = i[43];
  assign o[11161] = i[43];
  assign o[11162] = i[43];
  assign o[11163] = i[43];
  assign o[11164] = i[43];
  assign o[11165] = i[43];
  assign o[11166] = i[43];
  assign o[11167] = i[43];
  assign o[11168] = i[43];
  assign o[11169] = i[43];
  assign o[11170] = i[43];
  assign o[11171] = i[43];
  assign o[11172] = i[43];
  assign o[11173] = i[43];
  assign o[11174] = i[43];
  assign o[11175] = i[43];
  assign o[11176] = i[43];
  assign o[11177] = i[43];
  assign o[11178] = i[43];
  assign o[11179] = i[43];
  assign o[11180] = i[43];
  assign o[11181] = i[43];
  assign o[11182] = i[43];
  assign o[11183] = i[43];
  assign o[11184] = i[43];
  assign o[11185] = i[43];
  assign o[11186] = i[43];
  assign o[11187] = i[43];
  assign o[11188] = i[43];
  assign o[11189] = i[43];
  assign o[11190] = i[43];
  assign o[11191] = i[43];
  assign o[11192] = i[43];
  assign o[11193] = i[43];
  assign o[11194] = i[43];
  assign o[11195] = i[43];
  assign o[11196] = i[43];
  assign o[11197] = i[43];
  assign o[11198] = i[43];
  assign o[11199] = i[43];
  assign o[11200] = i[43];
  assign o[11201] = i[43];
  assign o[11202] = i[43];
  assign o[11203] = i[43];
  assign o[11204] = i[43];
  assign o[11205] = i[43];
  assign o[11206] = i[43];
  assign o[11207] = i[43];
  assign o[11208] = i[43];
  assign o[11209] = i[43];
  assign o[11210] = i[43];
  assign o[11211] = i[43];
  assign o[11212] = i[43];
  assign o[11213] = i[43];
  assign o[11214] = i[43];
  assign o[11215] = i[43];
  assign o[11216] = i[43];
  assign o[11217] = i[43];
  assign o[11218] = i[43];
  assign o[11219] = i[43];
  assign o[11220] = i[43];
  assign o[11221] = i[43];
  assign o[11222] = i[43];
  assign o[11223] = i[43];
  assign o[11224] = i[43];
  assign o[11225] = i[43];
  assign o[11226] = i[43];
  assign o[11227] = i[43];
  assign o[11228] = i[43];
  assign o[11229] = i[43];
  assign o[11230] = i[43];
  assign o[11231] = i[43];
  assign o[11232] = i[43];
  assign o[11233] = i[43];
  assign o[11234] = i[43];
  assign o[11235] = i[43];
  assign o[11236] = i[43];
  assign o[11237] = i[43];
  assign o[11238] = i[43];
  assign o[11239] = i[43];
  assign o[11240] = i[43];
  assign o[11241] = i[43];
  assign o[11242] = i[43];
  assign o[11243] = i[43];
  assign o[11244] = i[43];
  assign o[11245] = i[43];
  assign o[11246] = i[43];
  assign o[11247] = i[43];
  assign o[11248] = i[43];
  assign o[11249] = i[43];
  assign o[11250] = i[43];
  assign o[11251] = i[43];
  assign o[11252] = i[43];
  assign o[11253] = i[43];
  assign o[11254] = i[43];
  assign o[11255] = i[43];
  assign o[11256] = i[43];
  assign o[11257] = i[43];
  assign o[11258] = i[43];
  assign o[11259] = i[43];
  assign o[11260] = i[43];
  assign o[11261] = i[43];
  assign o[11262] = i[43];
  assign o[11263] = i[43];
  assign o[10752] = i[42];
  assign o[10753] = i[42];
  assign o[10754] = i[42];
  assign o[10755] = i[42];
  assign o[10756] = i[42];
  assign o[10757] = i[42];
  assign o[10758] = i[42];
  assign o[10759] = i[42];
  assign o[10760] = i[42];
  assign o[10761] = i[42];
  assign o[10762] = i[42];
  assign o[10763] = i[42];
  assign o[10764] = i[42];
  assign o[10765] = i[42];
  assign o[10766] = i[42];
  assign o[10767] = i[42];
  assign o[10768] = i[42];
  assign o[10769] = i[42];
  assign o[10770] = i[42];
  assign o[10771] = i[42];
  assign o[10772] = i[42];
  assign o[10773] = i[42];
  assign o[10774] = i[42];
  assign o[10775] = i[42];
  assign o[10776] = i[42];
  assign o[10777] = i[42];
  assign o[10778] = i[42];
  assign o[10779] = i[42];
  assign o[10780] = i[42];
  assign o[10781] = i[42];
  assign o[10782] = i[42];
  assign o[10783] = i[42];
  assign o[10784] = i[42];
  assign o[10785] = i[42];
  assign o[10786] = i[42];
  assign o[10787] = i[42];
  assign o[10788] = i[42];
  assign o[10789] = i[42];
  assign o[10790] = i[42];
  assign o[10791] = i[42];
  assign o[10792] = i[42];
  assign o[10793] = i[42];
  assign o[10794] = i[42];
  assign o[10795] = i[42];
  assign o[10796] = i[42];
  assign o[10797] = i[42];
  assign o[10798] = i[42];
  assign o[10799] = i[42];
  assign o[10800] = i[42];
  assign o[10801] = i[42];
  assign o[10802] = i[42];
  assign o[10803] = i[42];
  assign o[10804] = i[42];
  assign o[10805] = i[42];
  assign o[10806] = i[42];
  assign o[10807] = i[42];
  assign o[10808] = i[42];
  assign o[10809] = i[42];
  assign o[10810] = i[42];
  assign o[10811] = i[42];
  assign o[10812] = i[42];
  assign o[10813] = i[42];
  assign o[10814] = i[42];
  assign o[10815] = i[42];
  assign o[10816] = i[42];
  assign o[10817] = i[42];
  assign o[10818] = i[42];
  assign o[10819] = i[42];
  assign o[10820] = i[42];
  assign o[10821] = i[42];
  assign o[10822] = i[42];
  assign o[10823] = i[42];
  assign o[10824] = i[42];
  assign o[10825] = i[42];
  assign o[10826] = i[42];
  assign o[10827] = i[42];
  assign o[10828] = i[42];
  assign o[10829] = i[42];
  assign o[10830] = i[42];
  assign o[10831] = i[42];
  assign o[10832] = i[42];
  assign o[10833] = i[42];
  assign o[10834] = i[42];
  assign o[10835] = i[42];
  assign o[10836] = i[42];
  assign o[10837] = i[42];
  assign o[10838] = i[42];
  assign o[10839] = i[42];
  assign o[10840] = i[42];
  assign o[10841] = i[42];
  assign o[10842] = i[42];
  assign o[10843] = i[42];
  assign o[10844] = i[42];
  assign o[10845] = i[42];
  assign o[10846] = i[42];
  assign o[10847] = i[42];
  assign o[10848] = i[42];
  assign o[10849] = i[42];
  assign o[10850] = i[42];
  assign o[10851] = i[42];
  assign o[10852] = i[42];
  assign o[10853] = i[42];
  assign o[10854] = i[42];
  assign o[10855] = i[42];
  assign o[10856] = i[42];
  assign o[10857] = i[42];
  assign o[10858] = i[42];
  assign o[10859] = i[42];
  assign o[10860] = i[42];
  assign o[10861] = i[42];
  assign o[10862] = i[42];
  assign o[10863] = i[42];
  assign o[10864] = i[42];
  assign o[10865] = i[42];
  assign o[10866] = i[42];
  assign o[10867] = i[42];
  assign o[10868] = i[42];
  assign o[10869] = i[42];
  assign o[10870] = i[42];
  assign o[10871] = i[42];
  assign o[10872] = i[42];
  assign o[10873] = i[42];
  assign o[10874] = i[42];
  assign o[10875] = i[42];
  assign o[10876] = i[42];
  assign o[10877] = i[42];
  assign o[10878] = i[42];
  assign o[10879] = i[42];
  assign o[10880] = i[42];
  assign o[10881] = i[42];
  assign o[10882] = i[42];
  assign o[10883] = i[42];
  assign o[10884] = i[42];
  assign o[10885] = i[42];
  assign o[10886] = i[42];
  assign o[10887] = i[42];
  assign o[10888] = i[42];
  assign o[10889] = i[42];
  assign o[10890] = i[42];
  assign o[10891] = i[42];
  assign o[10892] = i[42];
  assign o[10893] = i[42];
  assign o[10894] = i[42];
  assign o[10895] = i[42];
  assign o[10896] = i[42];
  assign o[10897] = i[42];
  assign o[10898] = i[42];
  assign o[10899] = i[42];
  assign o[10900] = i[42];
  assign o[10901] = i[42];
  assign o[10902] = i[42];
  assign o[10903] = i[42];
  assign o[10904] = i[42];
  assign o[10905] = i[42];
  assign o[10906] = i[42];
  assign o[10907] = i[42];
  assign o[10908] = i[42];
  assign o[10909] = i[42];
  assign o[10910] = i[42];
  assign o[10911] = i[42];
  assign o[10912] = i[42];
  assign o[10913] = i[42];
  assign o[10914] = i[42];
  assign o[10915] = i[42];
  assign o[10916] = i[42];
  assign o[10917] = i[42];
  assign o[10918] = i[42];
  assign o[10919] = i[42];
  assign o[10920] = i[42];
  assign o[10921] = i[42];
  assign o[10922] = i[42];
  assign o[10923] = i[42];
  assign o[10924] = i[42];
  assign o[10925] = i[42];
  assign o[10926] = i[42];
  assign o[10927] = i[42];
  assign o[10928] = i[42];
  assign o[10929] = i[42];
  assign o[10930] = i[42];
  assign o[10931] = i[42];
  assign o[10932] = i[42];
  assign o[10933] = i[42];
  assign o[10934] = i[42];
  assign o[10935] = i[42];
  assign o[10936] = i[42];
  assign o[10937] = i[42];
  assign o[10938] = i[42];
  assign o[10939] = i[42];
  assign o[10940] = i[42];
  assign o[10941] = i[42];
  assign o[10942] = i[42];
  assign o[10943] = i[42];
  assign o[10944] = i[42];
  assign o[10945] = i[42];
  assign o[10946] = i[42];
  assign o[10947] = i[42];
  assign o[10948] = i[42];
  assign o[10949] = i[42];
  assign o[10950] = i[42];
  assign o[10951] = i[42];
  assign o[10952] = i[42];
  assign o[10953] = i[42];
  assign o[10954] = i[42];
  assign o[10955] = i[42];
  assign o[10956] = i[42];
  assign o[10957] = i[42];
  assign o[10958] = i[42];
  assign o[10959] = i[42];
  assign o[10960] = i[42];
  assign o[10961] = i[42];
  assign o[10962] = i[42];
  assign o[10963] = i[42];
  assign o[10964] = i[42];
  assign o[10965] = i[42];
  assign o[10966] = i[42];
  assign o[10967] = i[42];
  assign o[10968] = i[42];
  assign o[10969] = i[42];
  assign o[10970] = i[42];
  assign o[10971] = i[42];
  assign o[10972] = i[42];
  assign o[10973] = i[42];
  assign o[10974] = i[42];
  assign o[10975] = i[42];
  assign o[10976] = i[42];
  assign o[10977] = i[42];
  assign o[10978] = i[42];
  assign o[10979] = i[42];
  assign o[10980] = i[42];
  assign o[10981] = i[42];
  assign o[10982] = i[42];
  assign o[10983] = i[42];
  assign o[10984] = i[42];
  assign o[10985] = i[42];
  assign o[10986] = i[42];
  assign o[10987] = i[42];
  assign o[10988] = i[42];
  assign o[10989] = i[42];
  assign o[10990] = i[42];
  assign o[10991] = i[42];
  assign o[10992] = i[42];
  assign o[10993] = i[42];
  assign o[10994] = i[42];
  assign o[10995] = i[42];
  assign o[10996] = i[42];
  assign o[10997] = i[42];
  assign o[10998] = i[42];
  assign o[10999] = i[42];
  assign o[11000] = i[42];
  assign o[11001] = i[42];
  assign o[11002] = i[42];
  assign o[11003] = i[42];
  assign o[11004] = i[42];
  assign o[11005] = i[42];
  assign o[11006] = i[42];
  assign o[11007] = i[42];
  assign o[10496] = i[41];
  assign o[10497] = i[41];
  assign o[10498] = i[41];
  assign o[10499] = i[41];
  assign o[10500] = i[41];
  assign o[10501] = i[41];
  assign o[10502] = i[41];
  assign o[10503] = i[41];
  assign o[10504] = i[41];
  assign o[10505] = i[41];
  assign o[10506] = i[41];
  assign o[10507] = i[41];
  assign o[10508] = i[41];
  assign o[10509] = i[41];
  assign o[10510] = i[41];
  assign o[10511] = i[41];
  assign o[10512] = i[41];
  assign o[10513] = i[41];
  assign o[10514] = i[41];
  assign o[10515] = i[41];
  assign o[10516] = i[41];
  assign o[10517] = i[41];
  assign o[10518] = i[41];
  assign o[10519] = i[41];
  assign o[10520] = i[41];
  assign o[10521] = i[41];
  assign o[10522] = i[41];
  assign o[10523] = i[41];
  assign o[10524] = i[41];
  assign o[10525] = i[41];
  assign o[10526] = i[41];
  assign o[10527] = i[41];
  assign o[10528] = i[41];
  assign o[10529] = i[41];
  assign o[10530] = i[41];
  assign o[10531] = i[41];
  assign o[10532] = i[41];
  assign o[10533] = i[41];
  assign o[10534] = i[41];
  assign o[10535] = i[41];
  assign o[10536] = i[41];
  assign o[10537] = i[41];
  assign o[10538] = i[41];
  assign o[10539] = i[41];
  assign o[10540] = i[41];
  assign o[10541] = i[41];
  assign o[10542] = i[41];
  assign o[10543] = i[41];
  assign o[10544] = i[41];
  assign o[10545] = i[41];
  assign o[10546] = i[41];
  assign o[10547] = i[41];
  assign o[10548] = i[41];
  assign o[10549] = i[41];
  assign o[10550] = i[41];
  assign o[10551] = i[41];
  assign o[10552] = i[41];
  assign o[10553] = i[41];
  assign o[10554] = i[41];
  assign o[10555] = i[41];
  assign o[10556] = i[41];
  assign o[10557] = i[41];
  assign o[10558] = i[41];
  assign o[10559] = i[41];
  assign o[10560] = i[41];
  assign o[10561] = i[41];
  assign o[10562] = i[41];
  assign o[10563] = i[41];
  assign o[10564] = i[41];
  assign o[10565] = i[41];
  assign o[10566] = i[41];
  assign o[10567] = i[41];
  assign o[10568] = i[41];
  assign o[10569] = i[41];
  assign o[10570] = i[41];
  assign o[10571] = i[41];
  assign o[10572] = i[41];
  assign o[10573] = i[41];
  assign o[10574] = i[41];
  assign o[10575] = i[41];
  assign o[10576] = i[41];
  assign o[10577] = i[41];
  assign o[10578] = i[41];
  assign o[10579] = i[41];
  assign o[10580] = i[41];
  assign o[10581] = i[41];
  assign o[10582] = i[41];
  assign o[10583] = i[41];
  assign o[10584] = i[41];
  assign o[10585] = i[41];
  assign o[10586] = i[41];
  assign o[10587] = i[41];
  assign o[10588] = i[41];
  assign o[10589] = i[41];
  assign o[10590] = i[41];
  assign o[10591] = i[41];
  assign o[10592] = i[41];
  assign o[10593] = i[41];
  assign o[10594] = i[41];
  assign o[10595] = i[41];
  assign o[10596] = i[41];
  assign o[10597] = i[41];
  assign o[10598] = i[41];
  assign o[10599] = i[41];
  assign o[10600] = i[41];
  assign o[10601] = i[41];
  assign o[10602] = i[41];
  assign o[10603] = i[41];
  assign o[10604] = i[41];
  assign o[10605] = i[41];
  assign o[10606] = i[41];
  assign o[10607] = i[41];
  assign o[10608] = i[41];
  assign o[10609] = i[41];
  assign o[10610] = i[41];
  assign o[10611] = i[41];
  assign o[10612] = i[41];
  assign o[10613] = i[41];
  assign o[10614] = i[41];
  assign o[10615] = i[41];
  assign o[10616] = i[41];
  assign o[10617] = i[41];
  assign o[10618] = i[41];
  assign o[10619] = i[41];
  assign o[10620] = i[41];
  assign o[10621] = i[41];
  assign o[10622] = i[41];
  assign o[10623] = i[41];
  assign o[10624] = i[41];
  assign o[10625] = i[41];
  assign o[10626] = i[41];
  assign o[10627] = i[41];
  assign o[10628] = i[41];
  assign o[10629] = i[41];
  assign o[10630] = i[41];
  assign o[10631] = i[41];
  assign o[10632] = i[41];
  assign o[10633] = i[41];
  assign o[10634] = i[41];
  assign o[10635] = i[41];
  assign o[10636] = i[41];
  assign o[10637] = i[41];
  assign o[10638] = i[41];
  assign o[10639] = i[41];
  assign o[10640] = i[41];
  assign o[10641] = i[41];
  assign o[10642] = i[41];
  assign o[10643] = i[41];
  assign o[10644] = i[41];
  assign o[10645] = i[41];
  assign o[10646] = i[41];
  assign o[10647] = i[41];
  assign o[10648] = i[41];
  assign o[10649] = i[41];
  assign o[10650] = i[41];
  assign o[10651] = i[41];
  assign o[10652] = i[41];
  assign o[10653] = i[41];
  assign o[10654] = i[41];
  assign o[10655] = i[41];
  assign o[10656] = i[41];
  assign o[10657] = i[41];
  assign o[10658] = i[41];
  assign o[10659] = i[41];
  assign o[10660] = i[41];
  assign o[10661] = i[41];
  assign o[10662] = i[41];
  assign o[10663] = i[41];
  assign o[10664] = i[41];
  assign o[10665] = i[41];
  assign o[10666] = i[41];
  assign o[10667] = i[41];
  assign o[10668] = i[41];
  assign o[10669] = i[41];
  assign o[10670] = i[41];
  assign o[10671] = i[41];
  assign o[10672] = i[41];
  assign o[10673] = i[41];
  assign o[10674] = i[41];
  assign o[10675] = i[41];
  assign o[10676] = i[41];
  assign o[10677] = i[41];
  assign o[10678] = i[41];
  assign o[10679] = i[41];
  assign o[10680] = i[41];
  assign o[10681] = i[41];
  assign o[10682] = i[41];
  assign o[10683] = i[41];
  assign o[10684] = i[41];
  assign o[10685] = i[41];
  assign o[10686] = i[41];
  assign o[10687] = i[41];
  assign o[10688] = i[41];
  assign o[10689] = i[41];
  assign o[10690] = i[41];
  assign o[10691] = i[41];
  assign o[10692] = i[41];
  assign o[10693] = i[41];
  assign o[10694] = i[41];
  assign o[10695] = i[41];
  assign o[10696] = i[41];
  assign o[10697] = i[41];
  assign o[10698] = i[41];
  assign o[10699] = i[41];
  assign o[10700] = i[41];
  assign o[10701] = i[41];
  assign o[10702] = i[41];
  assign o[10703] = i[41];
  assign o[10704] = i[41];
  assign o[10705] = i[41];
  assign o[10706] = i[41];
  assign o[10707] = i[41];
  assign o[10708] = i[41];
  assign o[10709] = i[41];
  assign o[10710] = i[41];
  assign o[10711] = i[41];
  assign o[10712] = i[41];
  assign o[10713] = i[41];
  assign o[10714] = i[41];
  assign o[10715] = i[41];
  assign o[10716] = i[41];
  assign o[10717] = i[41];
  assign o[10718] = i[41];
  assign o[10719] = i[41];
  assign o[10720] = i[41];
  assign o[10721] = i[41];
  assign o[10722] = i[41];
  assign o[10723] = i[41];
  assign o[10724] = i[41];
  assign o[10725] = i[41];
  assign o[10726] = i[41];
  assign o[10727] = i[41];
  assign o[10728] = i[41];
  assign o[10729] = i[41];
  assign o[10730] = i[41];
  assign o[10731] = i[41];
  assign o[10732] = i[41];
  assign o[10733] = i[41];
  assign o[10734] = i[41];
  assign o[10735] = i[41];
  assign o[10736] = i[41];
  assign o[10737] = i[41];
  assign o[10738] = i[41];
  assign o[10739] = i[41];
  assign o[10740] = i[41];
  assign o[10741] = i[41];
  assign o[10742] = i[41];
  assign o[10743] = i[41];
  assign o[10744] = i[41];
  assign o[10745] = i[41];
  assign o[10746] = i[41];
  assign o[10747] = i[41];
  assign o[10748] = i[41];
  assign o[10749] = i[41];
  assign o[10750] = i[41];
  assign o[10751] = i[41];
  assign o[10240] = i[40];
  assign o[10241] = i[40];
  assign o[10242] = i[40];
  assign o[10243] = i[40];
  assign o[10244] = i[40];
  assign o[10245] = i[40];
  assign o[10246] = i[40];
  assign o[10247] = i[40];
  assign o[10248] = i[40];
  assign o[10249] = i[40];
  assign o[10250] = i[40];
  assign o[10251] = i[40];
  assign o[10252] = i[40];
  assign o[10253] = i[40];
  assign o[10254] = i[40];
  assign o[10255] = i[40];
  assign o[10256] = i[40];
  assign o[10257] = i[40];
  assign o[10258] = i[40];
  assign o[10259] = i[40];
  assign o[10260] = i[40];
  assign o[10261] = i[40];
  assign o[10262] = i[40];
  assign o[10263] = i[40];
  assign o[10264] = i[40];
  assign o[10265] = i[40];
  assign o[10266] = i[40];
  assign o[10267] = i[40];
  assign o[10268] = i[40];
  assign o[10269] = i[40];
  assign o[10270] = i[40];
  assign o[10271] = i[40];
  assign o[10272] = i[40];
  assign o[10273] = i[40];
  assign o[10274] = i[40];
  assign o[10275] = i[40];
  assign o[10276] = i[40];
  assign o[10277] = i[40];
  assign o[10278] = i[40];
  assign o[10279] = i[40];
  assign o[10280] = i[40];
  assign o[10281] = i[40];
  assign o[10282] = i[40];
  assign o[10283] = i[40];
  assign o[10284] = i[40];
  assign o[10285] = i[40];
  assign o[10286] = i[40];
  assign o[10287] = i[40];
  assign o[10288] = i[40];
  assign o[10289] = i[40];
  assign o[10290] = i[40];
  assign o[10291] = i[40];
  assign o[10292] = i[40];
  assign o[10293] = i[40];
  assign o[10294] = i[40];
  assign o[10295] = i[40];
  assign o[10296] = i[40];
  assign o[10297] = i[40];
  assign o[10298] = i[40];
  assign o[10299] = i[40];
  assign o[10300] = i[40];
  assign o[10301] = i[40];
  assign o[10302] = i[40];
  assign o[10303] = i[40];
  assign o[10304] = i[40];
  assign o[10305] = i[40];
  assign o[10306] = i[40];
  assign o[10307] = i[40];
  assign o[10308] = i[40];
  assign o[10309] = i[40];
  assign o[10310] = i[40];
  assign o[10311] = i[40];
  assign o[10312] = i[40];
  assign o[10313] = i[40];
  assign o[10314] = i[40];
  assign o[10315] = i[40];
  assign o[10316] = i[40];
  assign o[10317] = i[40];
  assign o[10318] = i[40];
  assign o[10319] = i[40];
  assign o[10320] = i[40];
  assign o[10321] = i[40];
  assign o[10322] = i[40];
  assign o[10323] = i[40];
  assign o[10324] = i[40];
  assign o[10325] = i[40];
  assign o[10326] = i[40];
  assign o[10327] = i[40];
  assign o[10328] = i[40];
  assign o[10329] = i[40];
  assign o[10330] = i[40];
  assign o[10331] = i[40];
  assign o[10332] = i[40];
  assign o[10333] = i[40];
  assign o[10334] = i[40];
  assign o[10335] = i[40];
  assign o[10336] = i[40];
  assign o[10337] = i[40];
  assign o[10338] = i[40];
  assign o[10339] = i[40];
  assign o[10340] = i[40];
  assign o[10341] = i[40];
  assign o[10342] = i[40];
  assign o[10343] = i[40];
  assign o[10344] = i[40];
  assign o[10345] = i[40];
  assign o[10346] = i[40];
  assign o[10347] = i[40];
  assign o[10348] = i[40];
  assign o[10349] = i[40];
  assign o[10350] = i[40];
  assign o[10351] = i[40];
  assign o[10352] = i[40];
  assign o[10353] = i[40];
  assign o[10354] = i[40];
  assign o[10355] = i[40];
  assign o[10356] = i[40];
  assign o[10357] = i[40];
  assign o[10358] = i[40];
  assign o[10359] = i[40];
  assign o[10360] = i[40];
  assign o[10361] = i[40];
  assign o[10362] = i[40];
  assign o[10363] = i[40];
  assign o[10364] = i[40];
  assign o[10365] = i[40];
  assign o[10366] = i[40];
  assign o[10367] = i[40];
  assign o[10368] = i[40];
  assign o[10369] = i[40];
  assign o[10370] = i[40];
  assign o[10371] = i[40];
  assign o[10372] = i[40];
  assign o[10373] = i[40];
  assign o[10374] = i[40];
  assign o[10375] = i[40];
  assign o[10376] = i[40];
  assign o[10377] = i[40];
  assign o[10378] = i[40];
  assign o[10379] = i[40];
  assign o[10380] = i[40];
  assign o[10381] = i[40];
  assign o[10382] = i[40];
  assign o[10383] = i[40];
  assign o[10384] = i[40];
  assign o[10385] = i[40];
  assign o[10386] = i[40];
  assign o[10387] = i[40];
  assign o[10388] = i[40];
  assign o[10389] = i[40];
  assign o[10390] = i[40];
  assign o[10391] = i[40];
  assign o[10392] = i[40];
  assign o[10393] = i[40];
  assign o[10394] = i[40];
  assign o[10395] = i[40];
  assign o[10396] = i[40];
  assign o[10397] = i[40];
  assign o[10398] = i[40];
  assign o[10399] = i[40];
  assign o[10400] = i[40];
  assign o[10401] = i[40];
  assign o[10402] = i[40];
  assign o[10403] = i[40];
  assign o[10404] = i[40];
  assign o[10405] = i[40];
  assign o[10406] = i[40];
  assign o[10407] = i[40];
  assign o[10408] = i[40];
  assign o[10409] = i[40];
  assign o[10410] = i[40];
  assign o[10411] = i[40];
  assign o[10412] = i[40];
  assign o[10413] = i[40];
  assign o[10414] = i[40];
  assign o[10415] = i[40];
  assign o[10416] = i[40];
  assign o[10417] = i[40];
  assign o[10418] = i[40];
  assign o[10419] = i[40];
  assign o[10420] = i[40];
  assign o[10421] = i[40];
  assign o[10422] = i[40];
  assign o[10423] = i[40];
  assign o[10424] = i[40];
  assign o[10425] = i[40];
  assign o[10426] = i[40];
  assign o[10427] = i[40];
  assign o[10428] = i[40];
  assign o[10429] = i[40];
  assign o[10430] = i[40];
  assign o[10431] = i[40];
  assign o[10432] = i[40];
  assign o[10433] = i[40];
  assign o[10434] = i[40];
  assign o[10435] = i[40];
  assign o[10436] = i[40];
  assign o[10437] = i[40];
  assign o[10438] = i[40];
  assign o[10439] = i[40];
  assign o[10440] = i[40];
  assign o[10441] = i[40];
  assign o[10442] = i[40];
  assign o[10443] = i[40];
  assign o[10444] = i[40];
  assign o[10445] = i[40];
  assign o[10446] = i[40];
  assign o[10447] = i[40];
  assign o[10448] = i[40];
  assign o[10449] = i[40];
  assign o[10450] = i[40];
  assign o[10451] = i[40];
  assign o[10452] = i[40];
  assign o[10453] = i[40];
  assign o[10454] = i[40];
  assign o[10455] = i[40];
  assign o[10456] = i[40];
  assign o[10457] = i[40];
  assign o[10458] = i[40];
  assign o[10459] = i[40];
  assign o[10460] = i[40];
  assign o[10461] = i[40];
  assign o[10462] = i[40];
  assign o[10463] = i[40];
  assign o[10464] = i[40];
  assign o[10465] = i[40];
  assign o[10466] = i[40];
  assign o[10467] = i[40];
  assign o[10468] = i[40];
  assign o[10469] = i[40];
  assign o[10470] = i[40];
  assign o[10471] = i[40];
  assign o[10472] = i[40];
  assign o[10473] = i[40];
  assign o[10474] = i[40];
  assign o[10475] = i[40];
  assign o[10476] = i[40];
  assign o[10477] = i[40];
  assign o[10478] = i[40];
  assign o[10479] = i[40];
  assign o[10480] = i[40];
  assign o[10481] = i[40];
  assign o[10482] = i[40];
  assign o[10483] = i[40];
  assign o[10484] = i[40];
  assign o[10485] = i[40];
  assign o[10486] = i[40];
  assign o[10487] = i[40];
  assign o[10488] = i[40];
  assign o[10489] = i[40];
  assign o[10490] = i[40];
  assign o[10491] = i[40];
  assign o[10492] = i[40];
  assign o[10493] = i[40];
  assign o[10494] = i[40];
  assign o[10495] = i[40];
  assign o[9984] = i[39];
  assign o[9985] = i[39];
  assign o[9986] = i[39];
  assign o[9987] = i[39];
  assign o[9988] = i[39];
  assign o[9989] = i[39];
  assign o[9990] = i[39];
  assign o[9991] = i[39];
  assign o[9992] = i[39];
  assign o[9993] = i[39];
  assign o[9994] = i[39];
  assign o[9995] = i[39];
  assign o[9996] = i[39];
  assign o[9997] = i[39];
  assign o[9998] = i[39];
  assign o[9999] = i[39];
  assign o[10000] = i[39];
  assign o[10001] = i[39];
  assign o[10002] = i[39];
  assign o[10003] = i[39];
  assign o[10004] = i[39];
  assign o[10005] = i[39];
  assign o[10006] = i[39];
  assign o[10007] = i[39];
  assign o[10008] = i[39];
  assign o[10009] = i[39];
  assign o[10010] = i[39];
  assign o[10011] = i[39];
  assign o[10012] = i[39];
  assign o[10013] = i[39];
  assign o[10014] = i[39];
  assign o[10015] = i[39];
  assign o[10016] = i[39];
  assign o[10017] = i[39];
  assign o[10018] = i[39];
  assign o[10019] = i[39];
  assign o[10020] = i[39];
  assign o[10021] = i[39];
  assign o[10022] = i[39];
  assign o[10023] = i[39];
  assign o[10024] = i[39];
  assign o[10025] = i[39];
  assign o[10026] = i[39];
  assign o[10027] = i[39];
  assign o[10028] = i[39];
  assign o[10029] = i[39];
  assign o[10030] = i[39];
  assign o[10031] = i[39];
  assign o[10032] = i[39];
  assign o[10033] = i[39];
  assign o[10034] = i[39];
  assign o[10035] = i[39];
  assign o[10036] = i[39];
  assign o[10037] = i[39];
  assign o[10038] = i[39];
  assign o[10039] = i[39];
  assign o[10040] = i[39];
  assign o[10041] = i[39];
  assign o[10042] = i[39];
  assign o[10043] = i[39];
  assign o[10044] = i[39];
  assign o[10045] = i[39];
  assign o[10046] = i[39];
  assign o[10047] = i[39];
  assign o[10048] = i[39];
  assign o[10049] = i[39];
  assign o[10050] = i[39];
  assign o[10051] = i[39];
  assign o[10052] = i[39];
  assign o[10053] = i[39];
  assign o[10054] = i[39];
  assign o[10055] = i[39];
  assign o[10056] = i[39];
  assign o[10057] = i[39];
  assign o[10058] = i[39];
  assign o[10059] = i[39];
  assign o[10060] = i[39];
  assign o[10061] = i[39];
  assign o[10062] = i[39];
  assign o[10063] = i[39];
  assign o[10064] = i[39];
  assign o[10065] = i[39];
  assign o[10066] = i[39];
  assign o[10067] = i[39];
  assign o[10068] = i[39];
  assign o[10069] = i[39];
  assign o[10070] = i[39];
  assign o[10071] = i[39];
  assign o[10072] = i[39];
  assign o[10073] = i[39];
  assign o[10074] = i[39];
  assign o[10075] = i[39];
  assign o[10076] = i[39];
  assign o[10077] = i[39];
  assign o[10078] = i[39];
  assign o[10079] = i[39];
  assign o[10080] = i[39];
  assign o[10081] = i[39];
  assign o[10082] = i[39];
  assign o[10083] = i[39];
  assign o[10084] = i[39];
  assign o[10085] = i[39];
  assign o[10086] = i[39];
  assign o[10087] = i[39];
  assign o[10088] = i[39];
  assign o[10089] = i[39];
  assign o[10090] = i[39];
  assign o[10091] = i[39];
  assign o[10092] = i[39];
  assign o[10093] = i[39];
  assign o[10094] = i[39];
  assign o[10095] = i[39];
  assign o[10096] = i[39];
  assign o[10097] = i[39];
  assign o[10098] = i[39];
  assign o[10099] = i[39];
  assign o[10100] = i[39];
  assign o[10101] = i[39];
  assign o[10102] = i[39];
  assign o[10103] = i[39];
  assign o[10104] = i[39];
  assign o[10105] = i[39];
  assign o[10106] = i[39];
  assign o[10107] = i[39];
  assign o[10108] = i[39];
  assign o[10109] = i[39];
  assign o[10110] = i[39];
  assign o[10111] = i[39];
  assign o[10112] = i[39];
  assign o[10113] = i[39];
  assign o[10114] = i[39];
  assign o[10115] = i[39];
  assign o[10116] = i[39];
  assign o[10117] = i[39];
  assign o[10118] = i[39];
  assign o[10119] = i[39];
  assign o[10120] = i[39];
  assign o[10121] = i[39];
  assign o[10122] = i[39];
  assign o[10123] = i[39];
  assign o[10124] = i[39];
  assign o[10125] = i[39];
  assign o[10126] = i[39];
  assign o[10127] = i[39];
  assign o[10128] = i[39];
  assign o[10129] = i[39];
  assign o[10130] = i[39];
  assign o[10131] = i[39];
  assign o[10132] = i[39];
  assign o[10133] = i[39];
  assign o[10134] = i[39];
  assign o[10135] = i[39];
  assign o[10136] = i[39];
  assign o[10137] = i[39];
  assign o[10138] = i[39];
  assign o[10139] = i[39];
  assign o[10140] = i[39];
  assign o[10141] = i[39];
  assign o[10142] = i[39];
  assign o[10143] = i[39];
  assign o[10144] = i[39];
  assign o[10145] = i[39];
  assign o[10146] = i[39];
  assign o[10147] = i[39];
  assign o[10148] = i[39];
  assign o[10149] = i[39];
  assign o[10150] = i[39];
  assign o[10151] = i[39];
  assign o[10152] = i[39];
  assign o[10153] = i[39];
  assign o[10154] = i[39];
  assign o[10155] = i[39];
  assign o[10156] = i[39];
  assign o[10157] = i[39];
  assign o[10158] = i[39];
  assign o[10159] = i[39];
  assign o[10160] = i[39];
  assign o[10161] = i[39];
  assign o[10162] = i[39];
  assign o[10163] = i[39];
  assign o[10164] = i[39];
  assign o[10165] = i[39];
  assign o[10166] = i[39];
  assign o[10167] = i[39];
  assign o[10168] = i[39];
  assign o[10169] = i[39];
  assign o[10170] = i[39];
  assign o[10171] = i[39];
  assign o[10172] = i[39];
  assign o[10173] = i[39];
  assign o[10174] = i[39];
  assign o[10175] = i[39];
  assign o[10176] = i[39];
  assign o[10177] = i[39];
  assign o[10178] = i[39];
  assign o[10179] = i[39];
  assign o[10180] = i[39];
  assign o[10181] = i[39];
  assign o[10182] = i[39];
  assign o[10183] = i[39];
  assign o[10184] = i[39];
  assign o[10185] = i[39];
  assign o[10186] = i[39];
  assign o[10187] = i[39];
  assign o[10188] = i[39];
  assign o[10189] = i[39];
  assign o[10190] = i[39];
  assign o[10191] = i[39];
  assign o[10192] = i[39];
  assign o[10193] = i[39];
  assign o[10194] = i[39];
  assign o[10195] = i[39];
  assign o[10196] = i[39];
  assign o[10197] = i[39];
  assign o[10198] = i[39];
  assign o[10199] = i[39];
  assign o[10200] = i[39];
  assign o[10201] = i[39];
  assign o[10202] = i[39];
  assign o[10203] = i[39];
  assign o[10204] = i[39];
  assign o[10205] = i[39];
  assign o[10206] = i[39];
  assign o[10207] = i[39];
  assign o[10208] = i[39];
  assign o[10209] = i[39];
  assign o[10210] = i[39];
  assign o[10211] = i[39];
  assign o[10212] = i[39];
  assign o[10213] = i[39];
  assign o[10214] = i[39];
  assign o[10215] = i[39];
  assign o[10216] = i[39];
  assign o[10217] = i[39];
  assign o[10218] = i[39];
  assign o[10219] = i[39];
  assign o[10220] = i[39];
  assign o[10221] = i[39];
  assign o[10222] = i[39];
  assign o[10223] = i[39];
  assign o[10224] = i[39];
  assign o[10225] = i[39];
  assign o[10226] = i[39];
  assign o[10227] = i[39];
  assign o[10228] = i[39];
  assign o[10229] = i[39];
  assign o[10230] = i[39];
  assign o[10231] = i[39];
  assign o[10232] = i[39];
  assign o[10233] = i[39];
  assign o[10234] = i[39];
  assign o[10235] = i[39];
  assign o[10236] = i[39];
  assign o[10237] = i[39];
  assign o[10238] = i[39];
  assign o[10239] = i[39];
  assign o[9728] = i[38];
  assign o[9729] = i[38];
  assign o[9730] = i[38];
  assign o[9731] = i[38];
  assign o[9732] = i[38];
  assign o[9733] = i[38];
  assign o[9734] = i[38];
  assign o[9735] = i[38];
  assign o[9736] = i[38];
  assign o[9737] = i[38];
  assign o[9738] = i[38];
  assign o[9739] = i[38];
  assign o[9740] = i[38];
  assign o[9741] = i[38];
  assign o[9742] = i[38];
  assign o[9743] = i[38];
  assign o[9744] = i[38];
  assign o[9745] = i[38];
  assign o[9746] = i[38];
  assign o[9747] = i[38];
  assign o[9748] = i[38];
  assign o[9749] = i[38];
  assign o[9750] = i[38];
  assign o[9751] = i[38];
  assign o[9752] = i[38];
  assign o[9753] = i[38];
  assign o[9754] = i[38];
  assign o[9755] = i[38];
  assign o[9756] = i[38];
  assign o[9757] = i[38];
  assign o[9758] = i[38];
  assign o[9759] = i[38];
  assign o[9760] = i[38];
  assign o[9761] = i[38];
  assign o[9762] = i[38];
  assign o[9763] = i[38];
  assign o[9764] = i[38];
  assign o[9765] = i[38];
  assign o[9766] = i[38];
  assign o[9767] = i[38];
  assign o[9768] = i[38];
  assign o[9769] = i[38];
  assign o[9770] = i[38];
  assign o[9771] = i[38];
  assign o[9772] = i[38];
  assign o[9773] = i[38];
  assign o[9774] = i[38];
  assign o[9775] = i[38];
  assign o[9776] = i[38];
  assign o[9777] = i[38];
  assign o[9778] = i[38];
  assign o[9779] = i[38];
  assign o[9780] = i[38];
  assign o[9781] = i[38];
  assign o[9782] = i[38];
  assign o[9783] = i[38];
  assign o[9784] = i[38];
  assign o[9785] = i[38];
  assign o[9786] = i[38];
  assign o[9787] = i[38];
  assign o[9788] = i[38];
  assign o[9789] = i[38];
  assign o[9790] = i[38];
  assign o[9791] = i[38];
  assign o[9792] = i[38];
  assign o[9793] = i[38];
  assign o[9794] = i[38];
  assign o[9795] = i[38];
  assign o[9796] = i[38];
  assign o[9797] = i[38];
  assign o[9798] = i[38];
  assign o[9799] = i[38];
  assign o[9800] = i[38];
  assign o[9801] = i[38];
  assign o[9802] = i[38];
  assign o[9803] = i[38];
  assign o[9804] = i[38];
  assign o[9805] = i[38];
  assign o[9806] = i[38];
  assign o[9807] = i[38];
  assign o[9808] = i[38];
  assign o[9809] = i[38];
  assign o[9810] = i[38];
  assign o[9811] = i[38];
  assign o[9812] = i[38];
  assign o[9813] = i[38];
  assign o[9814] = i[38];
  assign o[9815] = i[38];
  assign o[9816] = i[38];
  assign o[9817] = i[38];
  assign o[9818] = i[38];
  assign o[9819] = i[38];
  assign o[9820] = i[38];
  assign o[9821] = i[38];
  assign o[9822] = i[38];
  assign o[9823] = i[38];
  assign o[9824] = i[38];
  assign o[9825] = i[38];
  assign o[9826] = i[38];
  assign o[9827] = i[38];
  assign o[9828] = i[38];
  assign o[9829] = i[38];
  assign o[9830] = i[38];
  assign o[9831] = i[38];
  assign o[9832] = i[38];
  assign o[9833] = i[38];
  assign o[9834] = i[38];
  assign o[9835] = i[38];
  assign o[9836] = i[38];
  assign o[9837] = i[38];
  assign o[9838] = i[38];
  assign o[9839] = i[38];
  assign o[9840] = i[38];
  assign o[9841] = i[38];
  assign o[9842] = i[38];
  assign o[9843] = i[38];
  assign o[9844] = i[38];
  assign o[9845] = i[38];
  assign o[9846] = i[38];
  assign o[9847] = i[38];
  assign o[9848] = i[38];
  assign o[9849] = i[38];
  assign o[9850] = i[38];
  assign o[9851] = i[38];
  assign o[9852] = i[38];
  assign o[9853] = i[38];
  assign o[9854] = i[38];
  assign o[9855] = i[38];
  assign o[9856] = i[38];
  assign o[9857] = i[38];
  assign o[9858] = i[38];
  assign o[9859] = i[38];
  assign o[9860] = i[38];
  assign o[9861] = i[38];
  assign o[9862] = i[38];
  assign o[9863] = i[38];
  assign o[9864] = i[38];
  assign o[9865] = i[38];
  assign o[9866] = i[38];
  assign o[9867] = i[38];
  assign o[9868] = i[38];
  assign o[9869] = i[38];
  assign o[9870] = i[38];
  assign o[9871] = i[38];
  assign o[9872] = i[38];
  assign o[9873] = i[38];
  assign o[9874] = i[38];
  assign o[9875] = i[38];
  assign o[9876] = i[38];
  assign o[9877] = i[38];
  assign o[9878] = i[38];
  assign o[9879] = i[38];
  assign o[9880] = i[38];
  assign o[9881] = i[38];
  assign o[9882] = i[38];
  assign o[9883] = i[38];
  assign o[9884] = i[38];
  assign o[9885] = i[38];
  assign o[9886] = i[38];
  assign o[9887] = i[38];
  assign o[9888] = i[38];
  assign o[9889] = i[38];
  assign o[9890] = i[38];
  assign o[9891] = i[38];
  assign o[9892] = i[38];
  assign o[9893] = i[38];
  assign o[9894] = i[38];
  assign o[9895] = i[38];
  assign o[9896] = i[38];
  assign o[9897] = i[38];
  assign o[9898] = i[38];
  assign o[9899] = i[38];
  assign o[9900] = i[38];
  assign o[9901] = i[38];
  assign o[9902] = i[38];
  assign o[9903] = i[38];
  assign o[9904] = i[38];
  assign o[9905] = i[38];
  assign o[9906] = i[38];
  assign o[9907] = i[38];
  assign o[9908] = i[38];
  assign o[9909] = i[38];
  assign o[9910] = i[38];
  assign o[9911] = i[38];
  assign o[9912] = i[38];
  assign o[9913] = i[38];
  assign o[9914] = i[38];
  assign o[9915] = i[38];
  assign o[9916] = i[38];
  assign o[9917] = i[38];
  assign o[9918] = i[38];
  assign o[9919] = i[38];
  assign o[9920] = i[38];
  assign o[9921] = i[38];
  assign o[9922] = i[38];
  assign o[9923] = i[38];
  assign o[9924] = i[38];
  assign o[9925] = i[38];
  assign o[9926] = i[38];
  assign o[9927] = i[38];
  assign o[9928] = i[38];
  assign o[9929] = i[38];
  assign o[9930] = i[38];
  assign o[9931] = i[38];
  assign o[9932] = i[38];
  assign o[9933] = i[38];
  assign o[9934] = i[38];
  assign o[9935] = i[38];
  assign o[9936] = i[38];
  assign o[9937] = i[38];
  assign o[9938] = i[38];
  assign o[9939] = i[38];
  assign o[9940] = i[38];
  assign o[9941] = i[38];
  assign o[9942] = i[38];
  assign o[9943] = i[38];
  assign o[9944] = i[38];
  assign o[9945] = i[38];
  assign o[9946] = i[38];
  assign o[9947] = i[38];
  assign o[9948] = i[38];
  assign o[9949] = i[38];
  assign o[9950] = i[38];
  assign o[9951] = i[38];
  assign o[9952] = i[38];
  assign o[9953] = i[38];
  assign o[9954] = i[38];
  assign o[9955] = i[38];
  assign o[9956] = i[38];
  assign o[9957] = i[38];
  assign o[9958] = i[38];
  assign o[9959] = i[38];
  assign o[9960] = i[38];
  assign o[9961] = i[38];
  assign o[9962] = i[38];
  assign o[9963] = i[38];
  assign o[9964] = i[38];
  assign o[9965] = i[38];
  assign o[9966] = i[38];
  assign o[9967] = i[38];
  assign o[9968] = i[38];
  assign o[9969] = i[38];
  assign o[9970] = i[38];
  assign o[9971] = i[38];
  assign o[9972] = i[38];
  assign o[9973] = i[38];
  assign o[9974] = i[38];
  assign o[9975] = i[38];
  assign o[9976] = i[38];
  assign o[9977] = i[38];
  assign o[9978] = i[38];
  assign o[9979] = i[38];
  assign o[9980] = i[38];
  assign o[9981] = i[38];
  assign o[9982] = i[38];
  assign o[9983] = i[38];
  assign o[9472] = i[37];
  assign o[9473] = i[37];
  assign o[9474] = i[37];
  assign o[9475] = i[37];
  assign o[9476] = i[37];
  assign o[9477] = i[37];
  assign o[9478] = i[37];
  assign o[9479] = i[37];
  assign o[9480] = i[37];
  assign o[9481] = i[37];
  assign o[9482] = i[37];
  assign o[9483] = i[37];
  assign o[9484] = i[37];
  assign o[9485] = i[37];
  assign o[9486] = i[37];
  assign o[9487] = i[37];
  assign o[9488] = i[37];
  assign o[9489] = i[37];
  assign o[9490] = i[37];
  assign o[9491] = i[37];
  assign o[9492] = i[37];
  assign o[9493] = i[37];
  assign o[9494] = i[37];
  assign o[9495] = i[37];
  assign o[9496] = i[37];
  assign o[9497] = i[37];
  assign o[9498] = i[37];
  assign o[9499] = i[37];
  assign o[9500] = i[37];
  assign o[9501] = i[37];
  assign o[9502] = i[37];
  assign o[9503] = i[37];
  assign o[9504] = i[37];
  assign o[9505] = i[37];
  assign o[9506] = i[37];
  assign o[9507] = i[37];
  assign o[9508] = i[37];
  assign o[9509] = i[37];
  assign o[9510] = i[37];
  assign o[9511] = i[37];
  assign o[9512] = i[37];
  assign o[9513] = i[37];
  assign o[9514] = i[37];
  assign o[9515] = i[37];
  assign o[9516] = i[37];
  assign o[9517] = i[37];
  assign o[9518] = i[37];
  assign o[9519] = i[37];
  assign o[9520] = i[37];
  assign o[9521] = i[37];
  assign o[9522] = i[37];
  assign o[9523] = i[37];
  assign o[9524] = i[37];
  assign o[9525] = i[37];
  assign o[9526] = i[37];
  assign o[9527] = i[37];
  assign o[9528] = i[37];
  assign o[9529] = i[37];
  assign o[9530] = i[37];
  assign o[9531] = i[37];
  assign o[9532] = i[37];
  assign o[9533] = i[37];
  assign o[9534] = i[37];
  assign o[9535] = i[37];
  assign o[9536] = i[37];
  assign o[9537] = i[37];
  assign o[9538] = i[37];
  assign o[9539] = i[37];
  assign o[9540] = i[37];
  assign o[9541] = i[37];
  assign o[9542] = i[37];
  assign o[9543] = i[37];
  assign o[9544] = i[37];
  assign o[9545] = i[37];
  assign o[9546] = i[37];
  assign o[9547] = i[37];
  assign o[9548] = i[37];
  assign o[9549] = i[37];
  assign o[9550] = i[37];
  assign o[9551] = i[37];
  assign o[9552] = i[37];
  assign o[9553] = i[37];
  assign o[9554] = i[37];
  assign o[9555] = i[37];
  assign o[9556] = i[37];
  assign o[9557] = i[37];
  assign o[9558] = i[37];
  assign o[9559] = i[37];
  assign o[9560] = i[37];
  assign o[9561] = i[37];
  assign o[9562] = i[37];
  assign o[9563] = i[37];
  assign o[9564] = i[37];
  assign o[9565] = i[37];
  assign o[9566] = i[37];
  assign o[9567] = i[37];
  assign o[9568] = i[37];
  assign o[9569] = i[37];
  assign o[9570] = i[37];
  assign o[9571] = i[37];
  assign o[9572] = i[37];
  assign o[9573] = i[37];
  assign o[9574] = i[37];
  assign o[9575] = i[37];
  assign o[9576] = i[37];
  assign o[9577] = i[37];
  assign o[9578] = i[37];
  assign o[9579] = i[37];
  assign o[9580] = i[37];
  assign o[9581] = i[37];
  assign o[9582] = i[37];
  assign o[9583] = i[37];
  assign o[9584] = i[37];
  assign o[9585] = i[37];
  assign o[9586] = i[37];
  assign o[9587] = i[37];
  assign o[9588] = i[37];
  assign o[9589] = i[37];
  assign o[9590] = i[37];
  assign o[9591] = i[37];
  assign o[9592] = i[37];
  assign o[9593] = i[37];
  assign o[9594] = i[37];
  assign o[9595] = i[37];
  assign o[9596] = i[37];
  assign o[9597] = i[37];
  assign o[9598] = i[37];
  assign o[9599] = i[37];
  assign o[9600] = i[37];
  assign o[9601] = i[37];
  assign o[9602] = i[37];
  assign o[9603] = i[37];
  assign o[9604] = i[37];
  assign o[9605] = i[37];
  assign o[9606] = i[37];
  assign o[9607] = i[37];
  assign o[9608] = i[37];
  assign o[9609] = i[37];
  assign o[9610] = i[37];
  assign o[9611] = i[37];
  assign o[9612] = i[37];
  assign o[9613] = i[37];
  assign o[9614] = i[37];
  assign o[9615] = i[37];
  assign o[9616] = i[37];
  assign o[9617] = i[37];
  assign o[9618] = i[37];
  assign o[9619] = i[37];
  assign o[9620] = i[37];
  assign o[9621] = i[37];
  assign o[9622] = i[37];
  assign o[9623] = i[37];
  assign o[9624] = i[37];
  assign o[9625] = i[37];
  assign o[9626] = i[37];
  assign o[9627] = i[37];
  assign o[9628] = i[37];
  assign o[9629] = i[37];
  assign o[9630] = i[37];
  assign o[9631] = i[37];
  assign o[9632] = i[37];
  assign o[9633] = i[37];
  assign o[9634] = i[37];
  assign o[9635] = i[37];
  assign o[9636] = i[37];
  assign o[9637] = i[37];
  assign o[9638] = i[37];
  assign o[9639] = i[37];
  assign o[9640] = i[37];
  assign o[9641] = i[37];
  assign o[9642] = i[37];
  assign o[9643] = i[37];
  assign o[9644] = i[37];
  assign o[9645] = i[37];
  assign o[9646] = i[37];
  assign o[9647] = i[37];
  assign o[9648] = i[37];
  assign o[9649] = i[37];
  assign o[9650] = i[37];
  assign o[9651] = i[37];
  assign o[9652] = i[37];
  assign o[9653] = i[37];
  assign o[9654] = i[37];
  assign o[9655] = i[37];
  assign o[9656] = i[37];
  assign o[9657] = i[37];
  assign o[9658] = i[37];
  assign o[9659] = i[37];
  assign o[9660] = i[37];
  assign o[9661] = i[37];
  assign o[9662] = i[37];
  assign o[9663] = i[37];
  assign o[9664] = i[37];
  assign o[9665] = i[37];
  assign o[9666] = i[37];
  assign o[9667] = i[37];
  assign o[9668] = i[37];
  assign o[9669] = i[37];
  assign o[9670] = i[37];
  assign o[9671] = i[37];
  assign o[9672] = i[37];
  assign o[9673] = i[37];
  assign o[9674] = i[37];
  assign o[9675] = i[37];
  assign o[9676] = i[37];
  assign o[9677] = i[37];
  assign o[9678] = i[37];
  assign o[9679] = i[37];
  assign o[9680] = i[37];
  assign o[9681] = i[37];
  assign o[9682] = i[37];
  assign o[9683] = i[37];
  assign o[9684] = i[37];
  assign o[9685] = i[37];
  assign o[9686] = i[37];
  assign o[9687] = i[37];
  assign o[9688] = i[37];
  assign o[9689] = i[37];
  assign o[9690] = i[37];
  assign o[9691] = i[37];
  assign o[9692] = i[37];
  assign o[9693] = i[37];
  assign o[9694] = i[37];
  assign o[9695] = i[37];
  assign o[9696] = i[37];
  assign o[9697] = i[37];
  assign o[9698] = i[37];
  assign o[9699] = i[37];
  assign o[9700] = i[37];
  assign o[9701] = i[37];
  assign o[9702] = i[37];
  assign o[9703] = i[37];
  assign o[9704] = i[37];
  assign o[9705] = i[37];
  assign o[9706] = i[37];
  assign o[9707] = i[37];
  assign o[9708] = i[37];
  assign o[9709] = i[37];
  assign o[9710] = i[37];
  assign o[9711] = i[37];
  assign o[9712] = i[37];
  assign o[9713] = i[37];
  assign o[9714] = i[37];
  assign o[9715] = i[37];
  assign o[9716] = i[37];
  assign o[9717] = i[37];
  assign o[9718] = i[37];
  assign o[9719] = i[37];
  assign o[9720] = i[37];
  assign o[9721] = i[37];
  assign o[9722] = i[37];
  assign o[9723] = i[37];
  assign o[9724] = i[37];
  assign o[9725] = i[37];
  assign o[9726] = i[37];
  assign o[9727] = i[37];
  assign o[9216] = i[36];
  assign o[9217] = i[36];
  assign o[9218] = i[36];
  assign o[9219] = i[36];
  assign o[9220] = i[36];
  assign o[9221] = i[36];
  assign o[9222] = i[36];
  assign o[9223] = i[36];
  assign o[9224] = i[36];
  assign o[9225] = i[36];
  assign o[9226] = i[36];
  assign o[9227] = i[36];
  assign o[9228] = i[36];
  assign o[9229] = i[36];
  assign o[9230] = i[36];
  assign o[9231] = i[36];
  assign o[9232] = i[36];
  assign o[9233] = i[36];
  assign o[9234] = i[36];
  assign o[9235] = i[36];
  assign o[9236] = i[36];
  assign o[9237] = i[36];
  assign o[9238] = i[36];
  assign o[9239] = i[36];
  assign o[9240] = i[36];
  assign o[9241] = i[36];
  assign o[9242] = i[36];
  assign o[9243] = i[36];
  assign o[9244] = i[36];
  assign o[9245] = i[36];
  assign o[9246] = i[36];
  assign o[9247] = i[36];
  assign o[9248] = i[36];
  assign o[9249] = i[36];
  assign o[9250] = i[36];
  assign o[9251] = i[36];
  assign o[9252] = i[36];
  assign o[9253] = i[36];
  assign o[9254] = i[36];
  assign o[9255] = i[36];
  assign o[9256] = i[36];
  assign o[9257] = i[36];
  assign o[9258] = i[36];
  assign o[9259] = i[36];
  assign o[9260] = i[36];
  assign o[9261] = i[36];
  assign o[9262] = i[36];
  assign o[9263] = i[36];
  assign o[9264] = i[36];
  assign o[9265] = i[36];
  assign o[9266] = i[36];
  assign o[9267] = i[36];
  assign o[9268] = i[36];
  assign o[9269] = i[36];
  assign o[9270] = i[36];
  assign o[9271] = i[36];
  assign o[9272] = i[36];
  assign o[9273] = i[36];
  assign o[9274] = i[36];
  assign o[9275] = i[36];
  assign o[9276] = i[36];
  assign o[9277] = i[36];
  assign o[9278] = i[36];
  assign o[9279] = i[36];
  assign o[9280] = i[36];
  assign o[9281] = i[36];
  assign o[9282] = i[36];
  assign o[9283] = i[36];
  assign o[9284] = i[36];
  assign o[9285] = i[36];
  assign o[9286] = i[36];
  assign o[9287] = i[36];
  assign o[9288] = i[36];
  assign o[9289] = i[36];
  assign o[9290] = i[36];
  assign o[9291] = i[36];
  assign o[9292] = i[36];
  assign o[9293] = i[36];
  assign o[9294] = i[36];
  assign o[9295] = i[36];
  assign o[9296] = i[36];
  assign o[9297] = i[36];
  assign o[9298] = i[36];
  assign o[9299] = i[36];
  assign o[9300] = i[36];
  assign o[9301] = i[36];
  assign o[9302] = i[36];
  assign o[9303] = i[36];
  assign o[9304] = i[36];
  assign o[9305] = i[36];
  assign o[9306] = i[36];
  assign o[9307] = i[36];
  assign o[9308] = i[36];
  assign o[9309] = i[36];
  assign o[9310] = i[36];
  assign o[9311] = i[36];
  assign o[9312] = i[36];
  assign o[9313] = i[36];
  assign o[9314] = i[36];
  assign o[9315] = i[36];
  assign o[9316] = i[36];
  assign o[9317] = i[36];
  assign o[9318] = i[36];
  assign o[9319] = i[36];
  assign o[9320] = i[36];
  assign o[9321] = i[36];
  assign o[9322] = i[36];
  assign o[9323] = i[36];
  assign o[9324] = i[36];
  assign o[9325] = i[36];
  assign o[9326] = i[36];
  assign o[9327] = i[36];
  assign o[9328] = i[36];
  assign o[9329] = i[36];
  assign o[9330] = i[36];
  assign o[9331] = i[36];
  assign o[9332] = i[36];
  assign o[9333] = i[36];
  assign o[9334] = i[36];
  assign o[9335] = i[36];
  assign o[9336] = i[36];
  assign o[9337] = i[36];
  assign o[9338] = i[36];
  assign o[9339] = i[36];
  assign o[9340] = i[36];
  assign o[9341] = i[36];
  assign o[9342] = i[36];
  assign o[9343] = i[36];
  assign o[9344] = i[36];
  assign o[9345] = i[36];
  assign o[9346] = i[36];
  assign o[9347] = i[36];
  assign o[9348] = i[36];
  assign o[9349] = i[36];
  assign o[9350] = i[36];
  assign o[9351] = i[36];
  assign o[9352] = i[36];
  assign o[9353] = i[36];
  assign o[9354] = i[36];
  assign o[9355] = i[36];
  assign o[9356] = i[36];
  assign o[9357] = i[36];
  assign o[9358] = i[36];
  assign o[9359] = i[36];
  assign o[9360] = i[36];
  assign o[9361] = i[36];
  assign o[9362] = i[36];
  assign o[9363] = i[36];
  assign o[9364] = i[36];
  assign o[9365] = i[36];
  assign o[9366] = i[36];
  assign o[9367] = i[36];
  assign o[9368] = i[36];
  assign o[9369] = i[36];
  assign o[9370] = i[36];
  assign o[9371] = i[36];
  assign o[9372] = i[36];
  assign o[9373] = i[36];
  assign o[9374] = i[36];
  assign o[9375] = i[36];
  assign o[9376] = i[36];
  assign o[9377] = i[36];
  assign o[9378] = i[36];
  assign o[9379] = i[36];
  assign o[9380] = i[36];
  assign o[9381] = i[36];
  assign o[9382] = i[36];
  assign o[9383] = i[36];
  assign o[9384] = i[36];
  assign o[9385] = i[36];
  assign o[9386] = i[36];
  assign o[9387] = i[36];
  assign o[9388] = i[36];
  assign o[9389] = i[36];
  assign o[9390] = i[36];
  assign o[9391] = i[36];
  assign o[9392] = i[36];
  assign o[9393] = i[36];
  assign o[9394] = i[36];
  assign o[9395] = i[36];
  assign o[9396] = i[36];
  assign o[9397] = i[36];
  assign o[9398] = i[36];
  assign o[9399] = i[36];
  assign o[9400] = i[36];
  assign o[9401] = i[36];
  assign o[9402] = i[36];
  assign o[9403] = i[36];
  assign o[9404] = i[36];
  assign o[9405] = i[36];
  assign o[9406] = i[36];
  assign o[9407] = i[36];
  assign o[9408] = i[36];
  assign o[9409] = i[36];
  assign o[9410] = i[36];
  assign o[9411] = i[36];
  assign o[9412] = i[36];
  assign o[9413] = i[36];
  assign o[9414] = i[36];
  assign o[9415] = i[36];
  assign o[9416] = i[36];
  assign o[9417] = i[36];
  assign o[9418] = i[36];
  assign o[9419] = i[36];
  assign o[9420] = i[36];
  assign o[9421] = i[36];
  assign o[9422] = i[36];
  assign o[9423] = i[36];
  assign o[9424] = i[36];
  assign o[9425] = i[36];
  assign o[9426] = i[36];
  assign o[9427] = i[36];
  assign o[9428] = i[36];
  assign o[9429] = i[36];
  assign o[9430] = i[36];
  assign o[9431] = i[36];
  assign o[9432] = i[36];
  assign o[9433] = i[36];
  assign o[9434] = i[36];
  assign o[9435] = i[36];
  assign o[9436] = i[36];
  assign o[9437] = i[36];
  assign o[9438] = i[36];
  assign o[9439] = i[36];
  assign o[9440] = i[36];
  assign o[9441] = i[36];
  assign o[9442] = i[36];
  assign o[9443] = i[36];
  assign o[9444] = i[36];
  assign o[9445] = i[36];
  assign o[9446] = i[36];
  assign o[9447] = i[36];
  assign o[9448] = i[36];
  assign o[9449] = i[36];
  assign o[9450] = i[36];
  assign o[9451] = i[36];
  assign o[9452] = i[36];
  assign o[9453] = i[36];
  assign o[9454] = i[36];
  assign o[9455] = i[36];
  assign o[9456] = i[36];
  assign o[9457] = i[36];
  assign o[9458] = i[36];
  assign o[9459] = i[36];
  assign o[9460] = i[36];
  assign o[9461] = i[36];
  assign o[9462] = i[36];
  assign o[9463] = i[36];
  assign o[9464] = i[36];
  assign o[9465] = i[36];
  assign o[9466] = i[36];
  assign o[9467] = i[36];
  assign o[9468] = i[36];
  assign o[9469] = i[36];
  assign o[9470] = i[36];
  assign o[9471] = i[36];
  assign o[8960] = i[35];
  assign o[8961] = i[35];
  assign o[8962] = i[35];
  assign o[8963] = i[35];
  assign o[8964] = i[35];
  assign o[8965] = i[35];
  assign o[8966] = i[35];
  assign o[8967] = i[35];
  assign o[8968] = i[35];
  assign o[8969] = i[35];
  assign o[8970] = i[35];
  assign o[8971] = i[35];
  assign o[8972] = i[35];
  assign o[8973] = i[35];
  assign o[8974] = i[35];
  assign o[8975] = i[35];
  assign o[8976] = i[35];
  assign o[8977] = i[35];
  assign o[8978] = i[35];
  assign o[8979] = i[35];
  assign o[8980] = i[35];
  assign o[8981] = i[35];
  assign o[8982] = i[35];
  assign o[8983] = i[35];
  assign o[8984] = i[35];
  assign o[8985] = i[35];
  assign o[8986] = i[35];
  assign o[8987] = i[35];
  assign o[8988] = i[35];
  assign o[8989] = i[35];
  assign o[8990] = i[35];
  assign o[8991] = i[35];
  assign o[8992] = i[35];
  assign o[8993] = i[35];
  assign o[8994] = i[35];
  assign o[8995] = i[35];
  assign o[8996] = i[35];
  assign o[8997] = i[35];
  assign o[8998] = i[35];
  assign o[8999] = i[35];
  assign o[9000] = i[35];
  assign o[9001] = i[35];
  assign o[9002] = i[35];
  assign o[9003] = i[35];
  assign o[9004] = i[35];
  assign o[9005] = i[35];
  assign o[9006] = i[35];
  assign o[9007] = i[35];
  assign o[9008] = i[35];
  assign o[9009] = i[35];
  assign o[9010] = i[35];
  assign o[9011] = i[35];
  assign o[9012] = i[35];
  assign o[9013] = i[35];
  assign o[9014] = i[35];
  assign o[9015] = i[35];
  assign o[9016] = i[35];
  assign o[9017] = i[35];
  assign o[9018] = i[35];
  assign o[9019] = i[35];
  assign o[9020] = i[35];
  assign o[9021] = i[35];
  assign o[9022] = i[35];
  assign o[9023] = i[35];
  assign o[9024] = i[35];
  assign o[9025] = i[35];
  assign o[9026] = i[35];
  assign o[9027] = i[35];
  assign o[9028] = i[35];
  assign o[9029] = i[35];
  assign o[9030] = i[35];
  assign o[9031] = i[35];
  assign o[9032] = i[35];
  assign o[9033] = i[35];
  assign o[9034] = i[35];
  assign o[9035] = i[35];
  assign o[9036] = i[35];
  assign o[9037] = i[35];
  assign o[9038] = i[35];
  assign o[9039] = i[35];
  assign o[9040] = i[35];
  assign o[9041] = i[35];
  assign o[9042] = i[35];
  assign o[9043] = i[35];
  assign o[9044] = i[35];
  assign o[9045] = i[35];
  assign o[9046] = i[35];
  assign o[9047] = i[35];
  assign o[9048] = i[35];
  assign o[9049] = i[35];
  assign o[9050] = i[35];
  assign o[9051] = i[35];
  assign o[9052] = i[35];
  assign o[9053] = i[35];
  assign o[9054] = i[35];
  assign o[9055] = i[35];
  assign o[9056] = i[35];
  assign o[9057] = i[35];
  assign o[9058] = i[35];
  assign o[9059] = i[35];
  assign o[9060] = i[35];
  assign o[9061] = i[35];
  assign o[9062] = i[35];
  assign o[9063] = i[35];
  assign o[9064] = i[35];
  assign o[9065] = i[35];
  assign o[9066] = i[35];
  assign o[9067] = i[35];
  assign o[9068] = i[35];
  assign o[9069] = i[35];
  assign o[9070] = i[35];
  assign o[9071] = i[35];
  assign o[9072] = i[35];
  assign o[9073] = i[35];
  assign o[9074] = i[35];
  assign o[9075] = i[35];
  assign o[9076] = i[35];
  assign o[9077] = i[35];
  assign o[9078] = i[35];
  assign o[9079] = i[35];
  assign o[9080] = i[35];
  assign o[9081] = i[35];
  assign o[9082] = i[35];
  assign o[9083] = i[35];
  assign o[9084] = i[35];
  assign o[9085] = i[35];
  assign o[9086] = i[35];
  assign o[9087] = i[35];
  assign o[9088] = i[35];
  assign o[9089] = i[35];
  assign o[9090] = i[35];
  assign o[9091] = i[35];
  assign o[9092] = i[35];
  assign o[9093] = i[35];
  assign o[9094] = i[35];
  assign o[9095] = i[35];
  assign o[9096] = i[35];
  assign o[9097] = i[35];
  assign o[9098] = i[35];
  assign o[9099] = i[35];
  assign o[9100] = i[35];
  assign o[9101] = i[35];
  assign o[9102] = i[35];
  assign o[9103] = i[35];
  assign o[9104] = i[35];
  assign o[9105] = i[35];
  assign o[9106] = i[35];
  assign o[9107] = i[35];
  assign o[9108] = i[35];
  assign o[9109] = i[35];
  assign o[9110] = i[35];
  assign o[9111] = i[35];
  assign o[9112] = i[35];
  assign o[9113] = i[35];
  assign o[9114] = i[35];
  assign o[9115] = i[35];
  assign o[9116] = i[35];
  assign o[9117] = i[35];
  assign o[9118] = i[35];
  assign o[9119] = i[35];
  assign o[9120] = i[35];
  assign o[9121] = i[35];
  assign o[9122] = i[35];
  assign o[9123] = i[35];
  assign o[9124] = i[35];
  assign o[9125] = i[35];
  assign o[9126] = i[35];
  assign o[9127] = i[35];
  assign o[9128] = i[35];
  assign o[9129] = i[35];
  assign o[9130] = i[35];
  assign o[9131] = i[35];
  assign o[9132] = i[35];
  assign o[9133] = i[35];
  assign o[9134] = i[35];
  assign o[9135] = i[35];
  assign o[9136] = i[35];
  assign o[9137] = i[35];
  assign o[9138] = i[35];
  assign o[9139] = i[35];
  assign o[9140] = i[35];
  assign o[9141] = i[35];
  assign o[9142] = i[35];
  assign o[9143] = i[35];
  assign o[9144] = i[35];
  assign o[9145] = i[35];
  assign o[9146] = i[35];
  assign o[9147] = i[35];
  assign o[9148] = i[35];
  assign o[9149] = i[35];
  assign o[9150] = i[35];
  assign o[9151] = i[35];
  assign o[9152] = i[35];
  assign o[9153] = i[35];
  assign o[9154] = i[35];
  assign o[9155] = i[35];
  assign o[9156] = i[35];
  assign o[9157] = i[35];
  assign o[9158] = i[35];
  assign o[9159] = i[35];
  assign o[9160] = i[35];
  assign o[9161] = i[35];
  assign o[9162] = i[35];
  assign o[9163] = i[35];
  assign o[9164] = i[35];
  assign o[9165] = i[35];
  assign o[9166] = i[35];
  assign o[9167] = i[35];
  assign o[9168] = i[35];
  assign o[9169] = i[35];
  assign o[9170] = i[35];
  assign o[9171] = i[35];
  assign o[9172] = i[35];
  assign o[9173] = i[35];
  assign o[9174] = i[35];
  assign o[9175] = i[35];
  assign o[9176] = i[35];
  assign o[9177] = i[35];
  assign o[9178] = i[35];
  assign o[9179] = i[35];
  assign o[9180] = i[35];
  assign o[9181] = i[35];
  assign o[9182] = i[35];
  assign o[9183] = i[35];
  assign o[9184] = i[35];
  assign o[9185] = i[35];
  assign o[9186] = i[35];
  assign o[9187] = i[35];
  assign o[9188] = i[35];
  assign o[9189] = i[35];
  assign o[9190] = i[35];
  assign o[9191] = i[35];
  assign o[9192] = i[35];
  assign o[9193] = i[35];
  assign o[9194] = i[35];
  assign o[9195] = i[35];
  assign o[9196] = i[35];
  assign o[9197] = i[35];
  assign o[9198] = i[35];
  assign o[9199] = i[35];
  assign o[9200] = i[35];
  assign o[9201] = i[35];
  assign o[9202] = i[35];
  assign o[9203] = i[35];
  assign o[9204] = i[35];
  assign o[9205] = i[35];
  assign o[9206] = i[35];
  assign o[9207] = i[35];
  assign o[9208] = i[35];
  assign o[9209] = i[35];
  assign o[9210] = i[35];
  assign o[9211] = i[35];
  assign o[9212] = i[35];
  assign o[9213] = i[35];
  assign o[9214] = i[35];
  assign o[9215] = i[35];
  assign o[8704] = i[34];
  assign o[8705] = i[34];
  assign o[8706] = i[34];
  assign o[8707] = i[34];
  assign o[8708] = i[34];
  assign o[8709] = i[34];
  assign o[8710] = i[34];
  assign o[8711] = i[34];
  assign o[8712] = i[34];
  assign o[8713] = i[34];
  assign o[8714] = i[34];
  assign o[8715] = i[34];
  assign o[8716] = i[34];
  assign o[8717] = i[34];
  assign o[8718] = i[34];
  assign o[8719] = i[34];
  assign o[8720] = i[34];
  assign o[8721] = i[34];
  assign o[8722] = i[34];
  assign o[8723] = i[34];
  assign o[8724] = i[34];
  assign o[8725] = i[34];
  assign o[8726] = i[34];
  assign o[8727] = i[34];
  assign o[8728] = i[34];
  assign o[8729] = i[34];
  assign o[8730] = i[34];
  assign o[8731] = i[34];
  assign o[8732] = i[34];
  assign o[8733] = i[34];
  assign o[8734] = i[34];
  assign o[8735] = i[34];
  assign o[8736] = i[34];
  assign o[8737] = i[34];
  assign o[8738] = i[34];
  assign o[8739] = i[34];
  assign o[8740] = i[34];
  assign o[8741] = i[34];
  assign o[8742] = i[34];
  assign o[8743] = i[34];
  assign o[8744] = i[34];
  assign o[8745] = i[34];
  assign o[8746] = i[34];
  assign o[8747] = i[34];
  assign o[8748] = i[34];
  assign o[8749] = i[34];
  assign o[8750] = i[34];
  assign o[8751] = i[34];
  assign o[8752] = i[34];
  assign o[8753] = i[34];
  assign o[8754] = i[34];
  assign o[8755] = i[34];
  assign o[8756] = i[34];
  assign o[8757] = i[34];
  assign o[8758] = i[34];
  assign o[8759] = i[34];
  assign o[8760] = i[34];
  assign o[8761] = i[34];
  assign o[8762] = i[34];
  assign o[8763] = i[34];
  assign o[8764] = i[34];
  assign o[8765] = i[34];
  assign o[8766] = i[34];
  assign o[8767] = i[34];
  assign o[8768] = i[34];
  assign o[8769] = i[34];
  assign o[8770] = i[34];
  assign o[8771] = i[34];
  assign o[8772] = i[34];
  assign o[8773] = i[34];
  assign o[8774] = i[34];
  assign o[8775] = i[34];
  assign o[8776] = i[34];
  assign o[8777] = i[34];
  assign o[8778] = i[34];
  assign o[8779] = i[34];
  assign o[8780] = i[34];
  assign o[8781] = i[34];
  assign o[8782] = i[34];
  assign o[8783] = i[34];
  assign o[8784] = i[34];
  assign o[8785] = i[34];
  assign o[8786] = i[34];
  assign o[8787] = i[34];
  assign o[8788] = i[34];
  assign o[8789] = i[34];
  assign o[8790] = i[34];
  assign o[8791] = i[34];
  assign o[8792] = i[34];
  assign o[8793] = i[34];
  assign o[8794] = i[34];
  assign o[8795] = i[34];
  assign o[8796] = i[34];
  assign o[8797] = i[34];
  assign o[8798] = i[34];
  assign o[8799] = i[34];
  assign o[8800] = i[34];
  assign o[8801] = i[34];
  assign o[8802] = i[34];
  assign o[8803] = i[34];
  assign o[8804] = i[34];
  assign o[8805] = i[34];
  assign o[8806] = i[34];
  assign o[8807] = i[34];
  assign o[8808] = i[34];
  assign o[8809] = i[34];
  assign o[8810] = i[34];
  assign o[8811] = i[34];
  assign o[8812] = i[34];
  assign o[8813] = i[34];
  assign o[8814] = i[34];
  assign o[8815] = i[34];
  assign o[8816] = i[34];
  assign o[8817] = i[34];
  assign o[8818] = i[34];
  assign o[8819] = i[34];
  assign o[8820] = i[34];
  assign o[8821] = i[34];
  assign o[8822] = i[34];
  assign o[8823] = i[34];
  assign o[8824] = i[34];
  assign o[8825] = i[34];
  assign o[8826] = i[34];
  assign o[8827] = i[34];
  assign o[8828] = i[34];
  assign o[8829] = i[34];
  assign o[8830] = i[34];
  assign o[8831] = i[34];
  assign o[8832] = i[34];
  assign o[8833] = i[34];
  assign o[8834] = i[34];
  assign o[8835] = i[34];
  assign o[8836] = i[34];
  assign o[8837] = i[34];
  assign o[8838] = i[34];
  assign o[8839] = i[34];
  assign o[8840] = i[34];
  assign o[8841] = i[34];
  assign o[8842] = i[34];
  assign o[8843] = i[34];
  assign o[8844] = i[34];
  assign o[8845] = i[34];
  assign o[8846] = i[34];
  assign o[8847] = i[34];
  assign o[8848] = i[34];
  assign o[8849] = i[34];
  assign o[8850] = i[34];
  assign o[8851] = i[34];
  assign o[8852] = i[34];
  assign o[8853] = i[34];
  assign o[8854] = i[34];
  assign o[8855] = i[34];
  assign o[8856] = i[34];
  assign o[8857] = i[34];
  assign o[8858] = i[34];
  assign o[8859] = i[34];
  assign o[8860] = i[34];
  assign o[8861] = i[34];
  assign o[8862] = i[34];
  assign o[8863] = i[34];
  assign o[8864] = i[34];
  assign o[8865] = i[34];
  assign o[8866] = i[34];
  assign o[8867] = i[34];
  assign o[8868] = i[34];
  assign o[8869] = i[34];
  assign o[8870] = i[34];
  assign o[8871] = i[34];
  assign o[8872] = i[34];
  assign o[8873] = i[34];
  assign o[8874] = i[34];
  assign o[8875] = i[34];
  assign o[8876] = i[34];
  assign o[8877] = i[34];
  assign o[8878] = i[34];
  assign o[8879] = i[34];
  assign o[8880] = i[34];
  assign o[8881] = i[34];
  assign o[8882] = i[34];
  assign o[8883] = i[34];
  assign o[8884] = i[34];
  assign o[8885] = i[34];
  assign o[8886] = i[34];
  assign o[8887] = i[34];
  assign o[8888] = i[34];
  assign o[8889] = i[34];
  assign o[8890] = i[34];
  assign o[8891] = i[34];
  assign o[8892] = i[34];
  assign o[8893] = i[34];
  assign o[8894] = i[34];
  assign o[8895] = i[34];
  assign o[8896] = i[34];
  assign o[8897] = i[34];
  assign o[8898] = i[34];
  assign o[8899] = i[34];
  assign o[8900] = i[34];
  assign o[8901] = i[34];
  assign o[8902] = i[34];
  assign o[8903] = i[34];
  assign o[8904] = i[34];
  assign o[8905] = i[34];
  assign o[8906] = i[34];
  assign o[8907] = i[34];
  assign o[8908] = i[34];
  assign o[8909] = i[34];
  assign o[8910] = i[34];
  assign o[8911] = i[34];
  assign o[8912] = i[34];
  assign o[8913] = i[34];
  assign o[8914] = i[34];
  assign o[8915] = i[34];
  assign o[8916] = i[34];
  assign o[8917] = i[34];
  assign o[8918] = i[34];
  assign o[8919] = i[34];
  assign o[8920] = i[34];
  assign o[8921] = i[34];
  assign o[8922] = i[34];
  assign o[8923] = i[34];
  assign o[8924] = i[34];
  assign o[8925] = i[34];
  assign o[8926] = i[34];
  assign o[8927] = i[34];
  assign o[8928] = i[34];
  assign o[8929] = i[34];
  assign o[8930] = i[34];
  assign o[8931] = i[34];
  assign o[8932] = i[34];
  assign o[8933] = i[34];
  assign o[8934] = i[34];
  assign o[8935] = i[34];
  assign o[8936] = i[34];
  assign o[8937] = i[34];
  assign o[8938] = i[34];
  assign o[8939] = i[34];
  assign o[8940] = i[34];
  assign o[8941] = i[34];
  assign o[8942] = i[34];
  assign o[8943] = i[34];
  assign o[8944] = i[34];
  assign o[8945] = i[34];
  assign o[8946] = i[34];
  assign o[8947] = i[34];
  assign o[8948] = i[34];
  assign o[8949] = i[34];
  assign o[8950] = i[34];
  assign o[8951] = i[34];
  assign o[8952] = i[34];
  assign o[8953] = i[34];
  assign o[8954] = i[34];
  assign o[8955] = i[34];
  assign o[8956] = i[34];
  assign o[8957] = i[34];
  assign o[8958] = i[34];
  assign o[8959] = i[34];
  assign o[8448] = i[33];
  assign o[8449] = i[33];
  assign o[8450] = i[33];
  assign o[8451] = i[33];
  assign o[8452] = i[33];
  assign o[8453] = i[33];
  assign o[8454] = i[33];
  assign o[8455] = i[33];
  assign o[8456] = i[33];
  assign o[8457] = i[33];
  assign o[8458] = i[33];
  assign o[8459] = i[33];
  assign o[8460] = i[33];
  assign o[8461] = i[33];
  assign o[8462] = i[33];
  assign o[8463] = i[33];
  assign o[8464] = i[33];
  assign o[8465] = i[33];
  assign o[8466] = i[33];
  assign o[8467] = i[33];
  assign o[8468] = i[33];
  assign o[8469] = i[33];
  assign o[8470] = i[33];
  assign o[8471] = i[33];
  assign o[8472] = i[33];
  assign o[8473] = i[33];
  assign o[8474] = i[33];
  assign o[8475] = i[33];
  assign o[8476] = i[33];
  assign o[8477] = i[33];
  assign o[8478] = i[33];
  assign o[8479] = i[33];
  assign o[8480] = i[33];
  assign o[8481] = i[33];
  assign o[8482] = i[33];
  assign o[8483] = i[33];
  assign o[8484] = i[33];
  assign o[8485] = i[33];
  assign o[8486] = i[33];
  assign o[8487] = i[33];
  assign o[8488] = i[33];
  assign o[8489] = i[33];
  assign o[8490] = i[33];
  assign o[8491] = i[33];
  assign o[8492] = i[33];
  assign o[8493] = i[33];
  assign o[8494] = i[33];
  assign o[8495] = i[33];
  assign o[8496] = i[33];
  assign o[8497] = i[33];
  assign o[8498] = i[33];
  assign o[8499] = i[33];
  assign o[8500] = i[33];
  assign o[8501] = i[33];
  assign o[8502] = i[33];
  assign o[8503] = i[33];
  assign o[8504] = i[33];
  assign o[8505] = i[33];
  assign o[8506] = i[33];
  assign o[8507] = i[33];
  assign o[8508] = i[33];
  assign o[8509] = i[33];
  assign o[8510] = i[33];
  assign o[8511] = i[33];
  assign o[8512] = i[33];
  assign o[8513] = i[33];
  assign o[8514] = i[33];
  assign o[8515] = i[33];
  assign o[8516] = i[33];
  assign o[8517] = i[33];
  assign o[8518] = i[33];
  assign o[8519] = i[33];
  assign o[8520] = i[33];
  assign o[8521] = i[33];
  assign o[8522] = i[33];
  assign o[8523] = i[33];
  assign o[8524] = i[33];
  assign o[8525] = i[33];
  assign o[8526] = i[33];
  assign o[8527] = i[33];
  assign o[8528] = i[33];
  assign o[8529] = i[33];
  assign o[8530] = i[33];
  assign o[8531] = i[33];
  assign o[8532] = i[33];
  assign o[8533] = i[33];
  assign o[8534] = i[33];
  assign o[8535] = i[33];
  assign o[8536] = i[33];
  assign o[8537] = i[33];
  assign o[8538] = i[33];
  assign o[8539] = i[33];
  assign o[8540] = i[33];
  assign o[8541] = i[33];
  assign o[8542] = i[33];
  assign o[8543] = i[33];
  assign o[8544] = i[33];
  assign o[8545] = i[33];
  assign o[8546] = i[33];
  assign o[8547] = i[33];
  assign o[8548] = i[33];
  assign o[8549] = i[33];
  assign o[8550] = i[33];
  assign o[8551] = i[33];
  assign o[8552] = i[33];
  assign o[8553] = i[33];
  assign o[8554] = i[33];
  assign o[8555] = i[33];
  assign o[8556] = i[33];
  assign o[8557] = i[33];
  assign o[8558] = i[33];
  assign o[8559] = i[33];
  assign o[8560] = i[33];
  assign o[8561] = i[33];
  assign o[8562] = i[33];
  assign o[8563] = i[33];
  assign o[8564] = i[33];
  assign o[8565] = i[33];
  assign o[8566] = i[33];
  assign o[8567] = i[33];
  assign o[8568] = i[33];
  assign o[8569] = i[33];
  assign o[8570] = i[33];
  assign o[8571] = i[33];
  assign o[8572] = i[33];
  assign o[8573] = i[33];
  assign o[8574] = i[33];
  assign o[8575] = i[33];
  assign o[8576] = i[33];
  assign o[8577] = i[33];
  assign o[8578] = i[33];
  assign o[8579] = i[33];
  assign o[8580] = i[33];
  assign o[8581] = i[33];
  assign o[8582] = i[33];
  assign o[8583] = i[33];
  assign o[8584] = i[33];
  assign o[8585] = i[33];
  assign o[8586] = i[33];
  assign o[8587] = i[33];
  assign o[8588] = i[33];
  assign o[8589] = i[33];
  assign o[8590] = i[33];
  assign o[8591] = i[33];
  assign o[8592] = i[33];
  assign o[8593] = i[33];
  assign o[8594] = i[33];
  assign o[8595] = i[33];
  assign o[8596] = i[33];
  assign o[8597] = i[33];
  assign o[8598] = i[33];
  assign o[8599] = i[33];
  assign o[8600] = i[33];
  assign o[8601] = i[33];
  assign o[8602] = i[33];
  assign o[8603] = i[33];
  assign o[8604] = i[33];
  assign o[8605] = i[33];
  assign o[8606] = i[33];
  assign o[8607] = i[33];
  assign o[8608] = i[33];
  assign o[8609] = i[33];
  assign o[8610] = i[33];
  assign o[8611] = i[33];
  assign o[8612] = i[33];
  assign o[8613] = i[33];
  assign o[8614] = i[33];
  assign o[8615] = i[33];
  assign o[8616] = i[33];
  assign o[8617] = i[33];
  assign o[8618] = i[33];
  assign o[8619] = i[33];
  assign o[8620] = i[33];
  assign o[8621] = i[33];
  assign o[8622] = i[33];
  assign o[8623] = i[33];
  assign o[8624] = i[33];
  assign o[8625] = i[33];
  assign o[8626] = i[33];
  assign o[8627] = i[33];
  assign o[8628] = i[33];
  assign o[8629] = i[33];
  assign o[8630] = i[33];
  assign o[8631] = i[33];
  assign o[8632] = i[33];
  assign o[8633] = i[33];
  assign o[8634] = i[33];
  assign o[8635] = i[33];
  assign o[8636] = i[33];
  assign o[8637] = i[33];
  assign o[8638] = i[33];
  assign o[8639] = i[33];
  assign o[8640] = i[33];
  assign o[8641] = i[33];
  assign o[8642] = i[33];
  assign o[8643] = i[33];
  assign o[8644] = i[33];
  assign o[8645] = i[33];
  assign o[8646] = i[33];
  assign o[8647] = i[33];
  assign o[8648] = i[33];
  assign o[8649] = i[33];
  assign o[8650] = i[33];
  assign o[8651] = i[33];
  assign o[8652] = i[33];
  assign o[8653] = i[33];
  assign o[8654] = i[33];
  assign o[8655] = i[33];
  assign o[8656] = i[33];
  assign o[8657] = i[33];
  assign o[8658] = i[33];
  assign o[8659] = i[33];
  assign o[8660] = i[33];
  assign o[8661] = i[33];
  assign o[8662] = i[33];
  assign o[8663] = i[33];
  assign o[8664] = i[33];
  assign o[8665] = i[33];
  assign o[8666] = i[33];
  assign o[8667] = i[33];
  assign o[8668] = i[33];
  assign o[8669] = i[33];
  assign o[8670] = i[33];
  assign o[8671] = i[33];
  assign o[8672] = i[33];
  assign o[8673] = i[33];
  assign o[8674] = i[33];
  assign o[8675] = i[33];
  assign o[8676] = i[33];
  assign o[8677] = i[33];
  assign o[8678] = i[33];
  assign o[8679] = i[33];
  assign o[8680] = i[33];
  assign o[8681] = i[33];
  assign o[8682] = i[33];
  assign o[8683] = i[33];
  assign o[8684] = i[33];
  assign o[8685] = i[33];
  assign o[8686] = i[33];
  assign o[8687] = i[33];
  assign o[8688] = i[33];
  assign o[8689] = i[33];
  assign o[8690] = i[33];
  assign o[8691] = i[33];
  assign o[8692] = i[33];
  assign o[8693] = i[33];
  assign o[8694] = i[33];
  assign o[8695] = i[33];
  assign o[8696] = i[33];
  assign o[8697] = i[33];
  assign o[8698] = i[33];
  assign o[8699] = i[33];
  assign o[8700] = i[33];
  assign o[8701] = i[33];
  assign o[8702] = i[33];
  assign o[8703] = i[33];
  assign o[8192] = i[32];
  assign o[8193] = i[32];
  assign o[8194] = i[32];
  assign o[8195] = i[32];
  assign o[8196] = i[32];
  assign o[8197] = i[32];
  assign o[8198] = i[32];
  assign o[8199] = i[32];
  assign o[8200] = i[32];
  assign o[8201] = i[32];
  assign o[8202] = i[32];
  assign o[8203] = i[32];
  assign o[8204] = i[32];
  assign o[8205] = i[32];
  assign o[8206] = i[32];
  assign o[8207] = i[32];
  assign o[8208] = i[32];
  assign o[8209] = i[32];
  assign o[8210] = i[32];
  assign o[8211] = i[32];
  assign o[8212] = i[32];
  assign o[8213] = i[32];
  assign o[8214] = i[32];
  assign o[8215] = i[32];
  assign o[8216] = i[32];
  assign o[8217] = i[32];
  assign o[8218] = i[32];
  assign o[8219] = i[32];
  assign o[8220] = i[32];
  assign o[8221] = i[32];
  assign o[8222] = i[32];
  assign o[8223] = i[32];
  assign o[8224] = i[32];
  assign o[8225] = i[32];
  assign o[8226] = i[32];
  assign o[8227] = i[32];
  assign o[8228] = i[32];
  assign o[8229] = i[32];
  assign o[8230] = i[32];
  assign o[8231] = i[32];
  assign o[8232] = i[32];
  assign o[8233] = i[32];
  assign o[8234] = i[32];
  assign o[8235] = i[32];
  assign o[8236] = i[32];
  assign o[8237] = i[32];
  assign o[8238] = i[32];
  assign o[8239] = i[32];
  assign o[8240] = i[32];
  assign o[8241] = i[32];
  assign o[8242] = i[32];
  assign o[8243] = i[32];
  assign o[8244] = i[32];
  assign o[8245] = i[32];
  assign o[8246] = i[32];
  assign o[8247] = i[32];
  assign o[8248] = i[32];
  assign o[8249] = i[32];
  assign o[8250] = i[32];
  assign o[8251] = i[32];
  assign o[8252] = i[32];
  assign o[8253] = i[32];
  assign o[8254] = i[32];
  assign o[8255] = i[32];
  assign o[8256] = i[32];
  assign o[8257] = i[32];
  assign o[8258] = i[32];
  assign o[8259] = i[32];
  assign o[8260] = i[32];
  assign o[8261] = i[32];
  assign o[8262] = i[32];
  assign o[8263] = i[32];
  assign o[8264] = i[32];
  assign o[8265] = i[32];
  assign o[8266] = i[32];
  assign o[8267] = i[32];
  assign o[8268] = i[32];
  assign o[8269] = i[32];
  assign o[8270] = i[32];
  assign o[8271] = i[32];
  assign o[8272] = i[32];
  assign o[8273] = i[32];
  assign o[8274] = i[32];
  assign o[8275] = i[32];
  assign o[8276] = i[32];
  assign o[8277] = i[32];
  assign o[8278] = i[32];
  assign o[8279] = i[32];
  assign o[8280] = i[32];
  assign o[8281] = i[32];
  assign o[8282] = i[32];
  assign o[8283] = i[32];
  assign o[8284] = i[32];
  assign o[8285] = i[32];
  assign o[8286] = i[32];
  assign o[8287] = i[32];
  assign o[8288] = i[32];
  assign o[8289] = i[32];
  assign o[8290] = i[32];
  assign o[8291] = i[32];
  assign o[8292] = i[32];
  assign o[8293] = i[32];
  assign o[8294] = i[32];
  assign o[8295] = i[32];
  assign o[8296] = i[32];
  assign o[8297] = i[32];
  assign o[8298] = i[32];
  assign o[8299] = i[32];
  assign o[8300] = i[32];
  assign o[8301] = i[32];
  assign o[8302] = i[32];
  assign o[8303] = i[32];
  assign o[8304] = i[32];
  assign o[8305] = i[32];
  assign o[8306] = i[32];
  assign o[8307] = i[32];
  assign o[8308] = i[32];
  assign o[8309] = i[32];
  assign o[8310] = i[32];
  assign o[8311] = i[32];
  assign o[8312] = i[32];
  assign o[8313] = i[32];
  assign o[8314] = i[32];
  assign o[8315] = i[32];
  assign o[8316] = i[32];
  assign o[8317] = i[32];
  assign o[8318] = i[32];
  assign o[8319] = i[32];
  assign o[8320] = i[32];
  assign o[8321] = i[32];
  assign o[8322] = i[32];
  assign o[8323] = i[32];
  assign o[8324] = i[32];
  assign o[8325] = i[32];
  assign o[8326] = i[32];
  assign o[8327] = i[32];
  assign o[8328] = i[32];
  assign o[8329] = i[32];
  assign o[8330] = i[32];
  assign o[8331] = i[32];
  assign o[8332] = i[32];
  assign o[8333] = i[32];
  assign o[8334] = i[32];
  assign o[8335] = i[32];
  assign o[8336] = i[32];
  assign o[8337] = i[32];
  assign o[8338] = i[32];
  assign o[8339] = i[32];
  assign o[8340] = i[32];
  assign o[8341] = i[32];
  assign o[8342] = i[32];
  assign o[8343] = i[32];
  assign o[8344] = i[32];
  assign o[8345] = i[32];
  assign o[8346] = i[32];
  assign o[8347] = i[32];
  assign o[8348] = i[32];
  assign o[8349] = i[32];
  assign o[8350] = i[32];
  assign o[8351] = i[32];
  assign o[8352] = i[32];
  assign o[8353] = i[32];
  assign o[8354] = i[32];
  assign o[8355] = i[32];
  assign o[8356] = i[32];
  assign o[8357] = i[32];
  assign o[8358] = i[32];
  assign o[8359] = i[32];
  assign o[8360] = i[32];
  assign o[8361] = i[32];
  assign o[8362] = i[32];
  assign o[8363] = i[32];
  assign o[8364] = i[32];
  assign o[8365] = i[32];
  assign o[8366] = i[32];
  assign o[8367] = i[32];
  assign o[8368] = i[32];
  assign o[8369] = i[32];
  assign o[8370] = i[32];
  assign o[8371] = i[32];
  assign o[8372] = i[32];
  assign o[8373] = i[32];
  assign o[8374] = i[32];
  assign o[8375] = i[32];
  assign o[8376] = i[32];
  assign o[8377] = i[32];
  assign o[8378] = i[32];
  assign o[8379] = i[32];
  assign o[8380] = i[32];
  assign o[8381] = i[32];
  assign o[8382] = i[32];
  assign o[8383] = i[32];
  assign o[8384] = i[32];
  assign o[8385] = i[32];
  assign o[8386] = i[32];
  assign o[8387] = i[32];
  assign o[8388] = i[32];
  assign o[8389] = i[32];
  assign o[8390] = i[32];
  assign o[8391] = i[32];
  assign o[8392] = i[32];
  assign o[8393] = i[32];
  assign o[8394] = i[32];
  assign o[8395] = i[32];
  assign o[8396] = i[32];
  assign o[8397] = i[32];
  assign o[8398] = i[32];
  assign o[8399] = i[32];
  assign o[8400] = i[32];
  assign o[8401] = i[32];
  assign o[8402] = i[32];
  assign o[8403] = i[32];
  assign o[8404] = i[32];
  assign o[8405] = i[32];
  assign o[8406] = i[32];
  assign o[8407] = i[32];
  assign o[8408] = i[32];
  assign o[8409] = i[32];
  assign o[8410] = i[32];
  assign o[8411] = i[32];
  assign o[8412] = i[32];
  assign o[8413] = i[32];
  assign o[8414] = i[32];
  assign o[8415] = i[32];
  assign o[8416] = i[32];
  assign o[8417] = i[32];
  assign o[8418] = i[32];
  assign o[8419] = i[32];
  assign o[8420] = i[32];
  assign o[8421] = i[32];
  assign o[8422] = i[32];
  assign o[8423] = i[32];
  assign o[8424] = i[32];
  assign o[8425] = i[32];
  assign o[8426] = i[32];
  assign o[8427] = i[32];
  assign o[8428] = i[32];
  assign o[8429] = i[32];
  assign o[8430] = i[32];
  assign o[8431] = i[32];
  assign o[8432] = i[32];
  assign o[8433] = i[32];
  assign o[8434] = i[32];
  assign o[8435] = i[32];
  assign o[8436] = i[32];
  assign o[8437] = i[32];
  assign o[8438] = i[32];
  assign o[8439] = i[32];
  assign o[8440] = i[32];
  assign o[8441] = i[32];
  assign o[8442] = i[32];
  assign o[8443] = i[32];
  assign o[8444] = i[32];
  assign o[8445] = i[32];
  assign o[8446] = i[32];
  assign o[8447] = i[32];
  assign o[7936] = i[31];
  assign o[7937] = i[31];
  assign o[7938] = i[31];
  assign o[7939] = i[31];
  assign o[7940] = i[31];
  assign o[7941] = i[31];
  assign o[7942] = i[31];
  assign o[7943] = i[31];
  assign o[7944] = i[31];
  assign o[7945] = i[31];
  assign o[7946] = i[31];
  assign o[7947] = i[31];
  assign o[7948] = i[31];
  assign o[7949] = i[31];
  assign o[7950] = i[31];
  assign o[7951] = i[31];
  assign o[7952] = i[31];
  assign o[7953] = i[31];
  assign o[7954] = i[31];
  assign o[7955] = i[31];
  assign o[7956] = i[31];
  assign o[7957] = i[31];
  assign o[7958] = i[31];
  assign o[7959] = i[31];
  assign o[7960] = i[31];
  assign o[7961] = i[31];
  assign o[7962] = i[31];
  assign o[7963] = i[31];
  assign o[7964] = i[31];
  assign o[7965] = i[31];
  assign o[7966] = i[31];
  assign o[7967] = i[31];
  assign o[7968] = i[31];
  assign o[7969] = i[31];
  assign o[7970] = i[31];
  assign o[7971] = i[31];
  assign o[7972] = i[31];
  assign o[7973] = i[31];
  assign o[7974] = i[31];
  assign o[7975] = i[31];
  assign o[7976] = i[31];
  assign o[7977] = i[31];
  assign o[7978] = i[31];
  assign o[7979] = i[31];
  assign o[7980] = i[31];
  assign o[7981] = i[31];
  assign o[7982] = i[31];
  assign o[7983] = i[31];
  assign o[7984] = i[31];
  assign o[7985] = i[31];
  assign o[7986] = i[31];
  assign o[7987] = i[31];
  assign o[7988] = i[31];
  assign o[7989] = i[31];
  assign o[7990] = i[31];
  assign o[7991] = i[31];
  assign o[7992] = i[31];
  assign o[7993] = i[31];
  assign o[7994] = i[31];
  assign o[7995] = i[31];
  assign o[7996] = i[31];
  assign o[7997] = i[31];
  assign o[7998] = i[31];
  assign o[7999] = i[31];
  assign o[8000] = i[31];
  assign o[8001] = i[31];
  assign o[8002] = i[31];
  assign o[8003] = i[31];
  assign o[8004] = i[31];
  assign o[8005] = i[31];
  assign o[8006] = i[31];
  assign o[8007] = i[31];
  assign o[8008] = i[31];
  assign o[8009] = i[31];
  assign o[8010] = i[31];
  assign o[8011] = i[31];
  assign o[8012] = i[31];
  assign o[8013] = i[31];
  assign o[8014] = i[31];
  assign o[8015] = i[31];
  assign o[8016] = i[31];
  assign o[8017] = i[31];
  assign o[8018] = i[31];
  assign o[8019] = i[31];
  assign o[8020] = i[31];
  assign o[8021] = i[31];
  assign o[8022] = i[31];
  assign o[8023] = i[31];
  assign o[8024] = i[31];
  assign o[8025] = i[31];
  assign o[8026] = i[31];
  assign o[8027] = i[31];
  assign o[8028] = i[31];
  assign o[8029] = i[31];
  assign o[8030] = i[31];
  assign o[8031] = i[31];
  assign o[8032] = i[31];
  assign o[8033] = i[31];
  assign o[8034] = i[31];
  assign o[8035] = i[31];
  assign o[8036] = i[31];
  assign o[8037] = i[31];
  assign o[8038] = i[31];
  assign o[8039] = i[31];
  assign o[8040] = i[31];
  assign o[8041] = i[31];
  assign o[8042] = i[31];
  assign o[8043] = i[31];
  assign o[8044] = i[31];
  assign o[8045] = i[31];
  assign o[8046] = i[31];
  assign o[8047] = i[31];
  assign o[8048] = i[31];
  assign o[8049] = i[31];
  assign o[8050] = i[31];
  assign o[8051] = i[31];
  assign o[8052] = i[31];
  assign o[8053] = i[31];
  assign o[8054] = i[31];
  assign o[8055] = i[31];
  assign o[8056] = i[31];
  assign o[8057] = i[31];
  assign o[8058] = i[31];
  assign o[8059] = i[31];
  assign o[8060] = i[31];
  assign o[8061] = i[31];
  assign o[8062] = i[31];
  assign o[8063] = i[31];
  assign o[8064] = i[31];
  assign o[8065] = i[31];
  assign o[8066] = i[31];
  assign o[8067] = i[31];
  assign o[8068] = i[31];
  assign o[8069] = i[31];
  assign o[8070] = i[31];
  assign o[8071] = i[31];
  assign o[8072] = i[31];
  assign o[8073] = i[31];
  assign o[8074] = i[31];
  assign o[8075] = i[31];
  assign o[8076] = i[31];
  assign o[8077] = i[31];
  assign o[8078] = i[31];
  assign o[8079] = i[31];
  assign o[8080] = i[31];
  assign o[8081] = i[31];
  assign o[8082] = i[31];
  assign o[8083] = i[31];
  assign o[8084] = i[31];
  assign o[8085] = i[31];
  assign o[8086] = i[31];
  assign o[8087] = i[31];
  assign o[8088] = i[31];
  assign o[8089] = i[31];
  assign o[8090] = i[31];
  assign o[8091] = i[31];
  assign o[8092] = i[31];
  assign o[8093] = i[31];
  assign o[8094] = i[31];
  assign o[8095] = i[31];
  assign o[8096] = i[31];
  assign o[8097] = i[31];
  assign o[8098] = i[31];
  assign o[8099] = i[31];
  assign o[8100] = i[31];
  assign o[8101] = i[31];
  assign o[8102] = i[31];
  assign o[8103] = i[31];
  assign o[8104] = i[31];
  assign o[8105] = i[31];
  assign o[8106] = i[31];
  assign o[8107] = i[31];
  assign o[8108] = i[31];
  assign o[8109] = i[31];
  assign o[8110] = i[31];
  assign o[8111] = i[31];
  assign o[8112] = i[31];
  assign o[8113] = i[31];
  assign o[8114] = i[31];
  assign o[8115] = i[31];
  assign o[8116] = i[31];
  assign o[8117] = i[31];
  assign o[8118] = i[31];
  assign o[8119] = i[31];
  assign o[8120] = i[31];
  assign o[8121] = i[31];
  assign o[8122] = i[31];
  assign o[8123] = i[31];
  assign o[8124] = i[31];
  assign o[8125] = i[31];
  assign o[8126] = i[31];
  assign o[8127] = i[31];
  assign o[8128] = i[31];
  assign o[8129] = i[31];
  assign o[8130] = i[31];
  assign o[8131] = i[31];
  assign o[8132] = i[31];
  assign o[8133] = i[31];
  assign o[8134] = i[31];
  assign o[8135] = i[31];
  assign o[8136] = i[31];
  assign o[8137] = i[31];
  assign o[8138] = i[31];
  assign o[8139] = i[31];
  assign o[8140] = i[31];
  assign o[8141] = i[31];
  assign o[8142] = i[31];
  assign o[8143] = i[31];
  assign o[8144] = i[31];
  assign o[8145] = i[31];
  assign o[8146] = i[31];
  assign o[8147] = i[31];
  assign o[8148] = i[31];
  assign o[8149] = i[31];
  assign o[8150] = i[31];
  assign o[8151] = i[31];
  assign o[8152] = i[31];
  assign o[8153] = i[31];
  assign o[8154] = i[31];
  assign o[8155] = i[31];
  assign o[8156] = i[31];
  assign o[8157] = i[31];
  assign o[8158] = i[31];
  assign o[8159] = i[31];
  assign o[8160] = i[31];
  assign o[8161] = i[31];
  assign o[8162] = i[31];
  assign o[8163] = i[31];
  assign o[8164] = i[31];
  assign o[8165] = i[31];
  assign o[8166] = i[31];
  assign o[8167] = i[31];
  assign o[8168] = i[31];
  assign o[8169] = i[31];
  assign o[8170] = i[31];
  assign o[8171] = i[31];
  assign o[8172] = i[31];
  assign o[8173] = i[31];
  assign o[8174] = i[31];
  assign o[8175] = i[31];
  assign o[8176] = i[31];
  assign o[8177] = i[31];
  assign o[8178] = i[31];
  assign o[8179] = i[31];
  assign o[8180] = i[31];
  assign o[8181] = i[31];
  assign o[8182] = i[31];
  assign o[8183] = i[31];
  assign o[8184] = i[31];
  assign o[8185] = i[31];
  assign o[8186] = i[31];
  assign o[8187] = i[31];
  assign o[8188] = i[31];
  assign o[8189] = i[31];
  assign o[8190] = i[31];
  assign o[8191] = i[31];
  assign o[7680] = i[30];
  assign o[7681] = i[30];
  assign o[7682] = i[30];
  assign o[7683] = i[30];
  assign o[7684] = i[30];
  assign o[7685] = i[30];
  assign o[7686] = i[30];
  assign o[7687] = i[30];
  assign o[7688] = i[30];
  assign o[7689] = i[30];
  assign o[7690] = i[30];
  assign o[7691] = i[30];
  assign o[7692] = i[30];
  assign o[7693] = i[30];
  assign o[7694] = i[30];
  assign o[7695] = i[30];
  assign o[7696] = i[30];
  assign o[7697] = i[30];
  assign o[7698] = i[30];
  assign o[7699] = i[30];
  assign o[7700] = i[30];
  assign o[7701] = i[30];
  assign o[7702] = i[30];
  assign o[7703] = i[30];
  assign o[7704] = i[30];
  assign o[7705] = i[30];
  assign o[7706] = i[30];
  assign o[7707] = i[30];
  assign o[7708] = i[30];
  assign o[7709] = i[30];
  assign o[7710] = i[30];
  assign o[7711] = i[30];
  assign o[7712] = i[30];
  assign o[7713] = i[30];
  assign o[7714] = i[30];
  assign o[7715] = i[30];
  assign o[7716] = i[30];
  assign o[7717] = i[30];
  assign o[7718] = i[30];
  assign o[7719] = i[30];
  assign o[7720] = i[30];
  assign o[7721] = i[30];
  assign o[7722] = i[30];
  assign o[7723] = i[30];
  assign o[7724] = i[30];
  assign o[7725] = i[30];
  assign o[7726] = i[30];
  assign o[7727] = i[30];
  assign o[7728] = i[30];
  assign o[7729] = i[30];
  assign o[7730] = i[30];
  assign o[7731] = i[30];
  assign o[7732] = i[30];
  assign o[7733] = i[30];
  assign o[7734] = i[30];
  assign o[7735] = i[30];
  assign o[7736] = i[30];
  assign o[7737] = i[30];
  assign o[7738] = i[30];
  assign o[7739] = i[30];
  assign o[7740] = i[30];
  assign o[7741] = i[30];
  assign o[7742] = i[30];
  assign o[7743] = i[30];
  assign o[7744] = i[30];
  assign o[7745] = i[30];
  assign o[7746] = i[30];
  assign o[7747] = i[30];
  assign o[7748] = i[30];
  assign o[7749] = i[30];
  assign o[7750] = i[30];
  assign o[7751] = i[30];
  assign o[7752] = i[30];
  assign o[7753] = i[30];
  assign o[7754] = i[30];
  assign o[7755] = i[30];
  assign o[7756] = i[30];
  assign o[7757] = i[30];
  assign o[7758] = i[30];
  assign o[7759] = i[30];
  assign o[7760] = i[30];
  assign o[7761] = i[30];
  assign o[7762] = i[30];
  assign o[7763] = i[30];
  assign o[7764] = i[30];
  assign o[7765] = i[30];
  assign o[7766] = i[30];
  assign o[7767] = i[30];
  assign o[7768] = i[30];
  assign o[7769] = i[30];
  assign o[7770] = i[30];
  assign o[7771] = i[30];
  assign o[7772] = i[30];
  assign o[7773] = i[30];
  assign o[7774] = i[30];
  assign o[7775] = i[30];
  assign o[7776] = i[30];
  assign o[7777] = i[30];
  assign o[7778] = i[30];
  assign o[7779] = i[30];
  assign o[7780] = i[30];
  assign o[7781] = i[30];
  assign o[7782] = i[30];
  assign o[7783] = i[30];
  assign o[7784] = i[30];
  assign o[7785] = i[30];
  assign o[7786] = i[30];
  assign o[7787] = i[30];
  assign o[7788] = i[30];
  assign o[7789] = i[30];
  assign o[7790] = i[30];
  assign o[7791] = i[30];
  assign o[7792] = i[30];
  assign o[7793] = i[30];
  assign o[7794] = i[30];
  assign o[7795] = i[30];
  assign o[7796] = i[30];
  assign o[7797] = i[30];
  assign o[7798] = i[30];
  assign o[7799] = i[30];
  assign o[7800] = i[30];
  assign o[7801] = i[30];
  assign o[7802] = i[30];
  assign o[7803] = i[30];
  assign o[7804] = i[30];
  assign o[7805] = i[30];
  assign o[7806] = i[30];
  assign o[7807] = i[30];
  assign o[7808] = i[30];
  assign o[7809] = i[30];
  assign o[7810] = i[30];
  assign o[7811] = i[30];
  assign o[7812] = i[30];
  assign o[7813] = i[30];
  assign o[7814] = i[30];
  assign o[7815] = i[30];
  assign o[7816] = i[30];
  assign o[7817] = i[30];
  assign o[7818] = i[30];
  assign o[7819] = i[30];
  assign o[7820] = i[30];
  assign o[7821] = i[30];
  assign o[7822] = i[30];
  assign o[7823] = i[30];
  assign o[7824] = i[30];
  assign o[7825] = i[30];
  assign o[7826] = i[30];
  assign o[7827] = i[30];
  assign o[7828] = i[30];
  assign o[7829] = i[30];
  assign o[7830] = i[30];
  assign o[7831] = i[30];
  assign o[7832] = i[30];
  assign o[7833] = i[30];
  assign o[7834] = i[30];
  assign o[7835] = i[30];
  assign o[7836] = i[30];
  assign o[7837] = i[30];
  assign o[7838] = i[30];
  assign o[7839] = i[30];
  assign o[7840] = i[30];
  assign o[7841] = i[30];
  assign o[7842] = i[30];
  assign o[7843] = i[30];
  assign o[7844] = i[30];
  assign o[7845] = i[30];
  assign o[7846] = i[30];
  assign o[7847] = i[30];
  assign o[7848] = i[30];
  assign o[7849] = i[30];
  assign o[7850] = i[30];
  assign o[7851] = i[30];
  assign o[7852] = i[30];
  assign o[7853] = i[30];
  assign o[7854] = i[30];
  assign o[7855] = i[30];
  assign o[7856] = i[30];
  assign o[7857] = i[30];
  assign o[7858] = i[30];
  assign o[7859] = i[30];
  assign o[7860] = i[30];
  assign o[7861] = i[30];
  assign o[7862] = i[30];
  assign o[7863] = i[30];
  assign o[7864] = i[30];
  assign o[7865] = i[30];
  assign o[7866] = i[30];
  assign o[7867] = i[30];
  assign o[7868] = i[30];
  assign o[7869] = i[30];
  assign o[7870] = i[30];
  assign o[7871] = i[30];
  assign o[7872] = i[30];
  assign o[7873] = i[30];
  assign o[7874] = i[30];
  assign o[7875] = i[30];
  assign o[7876] = i[30];
  assign o[7877] = i[30];
  assign o[7878] = i[30];
  assign o[7879] = i[30];
  assign o[7880] = i[30];
  assign o[7881] = i[30];
  assign o[7882] = i[30];
  assign o[7883] = i[30];
  assign o[7884] = i[30];
  assign o[7885] = i[30];
  assign o[7886] = i[30];
  assign o[7887] = i[30];
  assign o[7888] = i[30];
  assign o[7889] = i[30];
  assign o[7890] = i[30];
  assign o[7891] = i[30];
  assign o[7892] = i[30];
  assign o[7893] = i[30];
  assign o[7894] = i[30];
  assign o[7895] = i[30];
  assign o[7896] = i[30];
  assign o[7897] = i[30];
  assign o[7898] = i[30];
  assign o[7899] = i[30];
  assign o[7900] = i[30];
  assign o[7901] = i[30];
  assign o[7902] = i[30];
  assign o[7903] = i[30];
  assign o[7904] = i[30];
  assign o[7905] = i[30];
  assign o[7906] = i[30];
  assign o[7907] = i[30];
  assign o[7908] = i[30];
  assign o[7909] = i[30];
  assign o[7910] = i[30];
  assign o[7911] = i[30];
  assign o[7912] = i[30];
  assign o[7913] = i[30];
  assign o[7914] = i[30];
  assign o[7915] = i[30];
  assign o[7916] = i[30];
  assign o[7917] = i[30];
  assign o[7918] = i[30];
  assign o[7919] = i[30];
  assign o[7920] = i[30];
  assign o[7921] = i[30];
  assign o[7922] = i[30];
  assign o[7923] = i[30];
  assign o[7924] = i[30];
  assign o[7925] = i[30];
  assign o[7926] = i[30];
  assign o[7927] = i[30];
  assign o[7928] = i[30];
  assign o[7929] = i[30];
  assign o[7930] = i[30];
  assign o[7931] = i[30];
  assign o[7932] = i[30];
  assign o[7933] = i[30];
  assign o[7934] = i[30];
  assign o[7935] = i[30];
  assign o[7424] = i[29];
  assign o[7425] = i[29];
  assign o[7426] = i[29];
  assign o[7427] = i[29];
  assign o[7428] = i[29];
  assign o[7429] = i[29];
  assign o[7430] = i[29];
  assign o[7431] = i[29];
  assign o[7432] = i[29];
  assign o[7433] = i[29];
  assign o[7434] = i[29];
  assign o[7435] = i[29];
  assign o[7436] = i[29];
  assign o[7437] = i[29];
  assign o[7438] = i[29];
  assign o[7439] = i[29];
  assign o[7440] = i[29];
  assign o[7441] = i[29];
  assign o[7442] = i[29];
  assign o[7443] = i[29];
  assign o[7444] = i[29];
  assign o[7445] = i[29];
  assign o[7446] = i[29];
  assign o[7447] = i[29];
  assign o[7448] = i[29];
  assign o[7449] = i[29];
  assign o[7450] = i[29];
  assign o[7451] = i[29];
  assign o[7452] = i[29];
  assign o[7453] = i[29];
  assign o[7454] = i[29];
  assign o[7455] = i[29];
  assign o[7456] = i[29];
  assign o[7457] = i[29];
  assign o[7458] = i[29];
  assign o[7459] = i[29];
  assign o[7460] = i[29];
  assign o[7461] = i[29];
  assign o[7462] = i[29];
  assign o[7463] = i[29];
  assign o[7464] = i[29];
  assign o[7465] = i[29];
  assign o[7466] = i[29];
  assign o[7467] = i[29];
  assign o[7468] = i[29];
  assign o[7469] = i[29];
  assign o[7470] = i[29];
  assign o[7471] = i[29];
  assign o[7472] = i[29];
  assign o[7473] = i[29];
  assign o[7474] = i[29];
  assign o[7475] = i[29];
  assign o[7476] = i[29];
  assign o[7477] = i[29];
  assign o[7478] = i[29];
  assign o[7479] = i[29];
  assign o[7480] = i[29];
  assign o[7481] = i[29];
  assign o[7482] = i[29];
  assign o[7483] = i[29];
  assign o[7484] = i[29];
  assign o[7485] = i[29];
  assign o[7486] = i[29];
  assign o[7487] = i[29];
  assign o[7488] = i[29];
  assign o[7489] = i[29];
  assign o[7490] = i[29];
  assign o[7491] = i[29];
  assign o[7492] = i[29];
  assign o[7493] = i[29];
  assign o[7494] = i[29];
  assign o[7495] = i[29];
  assign o[7496] = i[29];
  assign o[7497] = i[29];
  assign o[7498] = i[29];
  assign o[7499] = i[29];
  assign o[7500] = i[29];
  assign o[7501] = i[29];
  assign o[7502] = i[29];
  assign o[7503] = i[29];
  assign o[7504] = i[29];
  assign o[7505] = i[29];
  assign o[7506] = i[29];
  assign o[7507] = i[29];
  assign o[7508] = i[29];
  assign o[7509] = i[29];
  assign o[7510] = i[29];
  assign o[7511] = i[29];
  assign o[7512] = i[29];
  assign o[7513] = i[29];
  assign o[7514] = i[29];
  assign o[7515] = i[29];
  assign o[7516] = i[29];
  assign o[7517] = i[29];
  assign o[7518] = i[29];
  assign o[7519] = i[29];
  assign o[7520] = i[29];
  assign o[7521] = i[29];
  assign o[7522] = i[29];
  assign o[7523] = i[29];
  assign o[7524] = i[29];
  assign o[7525] = i[29];
  assign o[7526] = i[29];
  assign o[7527] = i[29];
  assign o[7528] = i[29];
  assign o[7529] = i[29];
  assign o[7530] = i[29];
  assign o[7531] = i[29];
  assign o[7532] = i[29];
  assign o[7533] = i[29];
  assign o[7534] = i[29];
  assign o[7535] = i[29];
  assign o[7536] = i[29];
  assign o[7537] = i[29];
  assign o[7538] = i[29];
  assign o[7539] = i[29];
  assign o[7540] = i[29];
  assign o[7541] = i[29];
  assign o[7542] = i[29];
  assign o[7543] = i[29];
  assign o[7544] = i[29];
  assign o[7545] = i[29];
  assign o[7546] = i[29];
  assign o[7547] = i[29];
  assign o[7548] = i[29];
  assign o[7549] = i[29];
  assign o[7550] = i[29];
  assign o[7551] = i[29];
  assign o[7552] = i[29];
  assign o[7553] = i[29];
  assign o[7554] = i[29];
  assign o[7555] = i[29];
  assign o[7556] = i[29];
  assign o[7557] = i[29];
  assign o[7558] = i[29];
  assign o[7559] = i[29];
  assign o[7560] = i[29];
  assign o[7561] = i[29];
  assign o[7562] = i[29];
  assign o[7563] = i[29];
  assign o[7564] = i[29];
  assign o[7565] = i[29];
  assign o[7566] = i[29];
  assign o[7567] = i[29];
  assign o[7568] = i[29];
  assign o[7569] = i[29];
  assign o[7570] = i[29];
  assign o[7571] = i[29];
  assign o[7572] = i[29];
  assign o[7573] = i[29];
  assign o[7574] = i[29];
  assign o[7575] = i[29];
  assign o[7576] = i[29];
  assign o[7577] = i[29];
  assign o[7578] = i[29];
  assign o[7579] = i[29];
  assign o[7580] = i[29];
  assign o[7581] = i[29];
  assign o[7582] = i[29];
  assign o[7583] = i[29];
  assign o[7584] = i[29];
  assign o[7585] = i[29];
  assign o[7586] = i[29];
  assign o[7587] = i[29];
  assign o[7588] = i[29];
  assign o[7589] = i[29];
  assign o[7590] = i[29];
  assign o[7591] = i[29];
  assign o[7592] = i[29];
  assign o[7593] = i[29];
  assign o[7594] = i[29];
  assign o[7595] = i[29];
  assign o[7596] = i[29];
  assign o[7597] = i[29];
  assign o[7598] = i[29];
  assign o[7599] = i[29];
  assign o[7600] = i[29];
  assign o[7601] = i[29];
  assign o[7602] = i[29];
  assign o[7603] = i[29];
  assign o[7604] = i[29];
  assign o[7605] = i[29];
  assign o[7606] = i[29];
  assign o[7607] = i[29];
  assign o[7608] = i[29];
  assign o[7609] = i[29];
  assign o[7610] = i[29];
  assign o[7611] = i[29];
  assign o[7612] = i[29];
  assign o[7613] = i[29];
  assign o[7614] = i[29];
  assign o[7615] = i[29];
  assign o[7616] = i[29];
  assign o[7617] = i[29];
  assign o[7618] = i[29];
  assign o[7619] = i[29];
  assign o[7620] = i[29];
  assign o[7621] = i[29];
  assign o[7622] = i[29];
  assign o[7623] = i[29];
  assign o[7624] = i[29];
  assign o[7625] = i[29];
  assign o[7626] = i[29];
  assign o[7627] = i[29];
  assign o[7628] = i[29];
  assign o[7629] = i[29];
  assign o[7630] = i[29];
  assign o[7631] = i[29];
  assign o[7632] = i[29];
  assign o[7633] = i[29];
  assign o[7634] = i[29];
  assign o[7635] = i[29];
  assign o[7636] = i[29];
  assign o[7637] = i[29];
  assign o[7638] = i[29];
  assign o[7639] = i[29];
  assign o[7640] = i[29];
  assign o[7641] = i[29];
  assign o[7642] = i[29];
  assign o[7643] = i[29];
  assign o[7644] = i[29];
  assign o[7645] = i[29];
  assign o[7646] = i[29];
  assign o[7647] = i[29];
  assign o[7648] = i[29];
  assign o[7649] = i[29];
  assign o[7650] = i[29];
  assign o[7651] = i[29];
  assign o[7652] = i[29];
  assign o[7653] = i[29];
  assign o[7654] = i[29];
  assign o[7655] = i[29];
  assign o[7656] = i[29];
  assign o[7657] = i[29];
  assign o[7658] = i[29];
  assign o[7659] = i[29];
  assign o[7660] = i[29];
  assign o[7661] = i[29];
  assign o[7662] = i[29];
  assign o[7663] = i[29];
  assign o[7664] = i[29];
  assign o[7665] = i[29];
  assign o[7666] = i[29];
  assign o[7667] = i[29];
  assign o[7668] = i[29];
  assign o[7669] = i[29];
  assign o[7670] = i[29];
  assign o[7671] = i[29];
  assign o[7672] = i[29];
  assign o[7673] = i[29];
  assign o[7674] = i[29];
  assign o[7675] = i[29];
  assign o[7676] = i[29];
  assign o[7677] = i[29];
  assign o[7678] = i[29];
  assign o[7679] = i[29];
  assign o[7168] = i[28];
  assign o[7169] = i[28];
  assign o[7170] = i[28];
  assign o[7171] = i[28];
  assign o[7172] = i[28];
  assign o[7173] = i[28];
  assign o[7174] = i[28];
  assign o[7175] = i[28];
  assign o[7176] = i[28];
  assign o[7177] = i[28];
  assign o[7178] = i[28];
  assign o[7179] = i[28];
  assign o[7180] = i[28];
  assign o[7181] = i[28];
  assign o[7182] = i[28];
  assign o[7183] = i[28];
  assign o[7184] = i[28];
  assign o[7185] = i[28];
  assign o[7186] = i[28];
  assign o[7187] = i[28];
  assign o[7188] = i[28];
  assign o[7189] = i[28];
  assign o[7190] = i[28];
  assign o[7191] = i[28];
  assign o[7192] = i[28];
  assign o[7193] = i[28];
  assign o[7194] = i[28];
  assign o[7195] = i[28];
  assign o[7196] = i[28];
  assign o[7197] = i[28];
  assign o[7198] = i[28];
  assign o[7199] = i[28];
  assign o[7200] = i[28];
  assign o[7201] = i[28];
  assign o[7202] = i[28];
  assign o[7203] = i[28];
  assign o[7204] = i[28];
  assign o[7205] = i[28];
  assign o[7206] = i[28];
  assign o[7207] = i[28];
  assign o[7208] = i[28];
  assign o[7209] = i[28];
  assign o[7210] = i[28];
  assign o[7211] = i[28];
  assign o[7212] = i[28];
  assign o[7213] = i[28];
  assign o[7214] = i[28];
  assign o[7215] = i[28];
  assign o[7216] = i[28];
  assign o[7217] = i[28];
  assign o[7218] = i[28];
  assign o[7219] = i[28];
  assign o[7220] = i[28];
  assign o[7221] = i[28];
  assign o[7222] = i[28];
  assign o[7223] = i[28];
  assign o[7224] = i[28];
  assign o[7225] = i[28];
  assign o[7226] = i[28];
  assign o[7227] = i[28];
  assign o[7228] = i[28];
  assign o[7229] = i[28];
  assign o[7230] = i[28];
  assign o[7231] = i[28];
  assign o[7232] = i[28];
  assign o[7233] = i[28];
  assign o[7234] = i[28];
  assign o[7235] = i[28];
  assign o[7236] = i[28];
  assign o[7237] = i[28];
  assign o[7238] = i[28];
  assign o[7239] = i[28];
  assign o[7240] = i[28];
  assign o[7241] = i[28];
  assign o[7242] = i[28];
  assign o[7243] = i[28];
  assign o[7244] = i[28];
  assign o[7245] = i[28];
  assign o[7246] = i[28];
  assign o[7247] = i[28];
  assign o[7248] = i[28];
  assign o[7249] = i[28];
  assign o[7250] = i[28];
  assign o[7251] = i[28];
  assign o[7252] = i[28];
  assign o[7253] = i[28];
  assign o[7254] = i[28];
  assign o[7255] = i[28];
  assign o[7256] = i[28];
  assign o[7257] = i[28];
  assign o[7258] = i[28];
  assign o[7259] = i[28];
  assign o[7260] = i[28];
  assign o[7261] = i[28];
  assign o[7262] = i[28];
  assign o[7263] = i[28];
  assign o[7264] = i[28];
  assign o[7265] = i[28];
  assign o[7266] = i[28];
  assign o[7267] = i[28];
  assign o[7268] = i[28];
  assign o[7269] = i[28];
  assign o[7270] = i[28];
  assign o[7271] = i[28];
  assign o[7272] = i[28];
  assign o[7273] = i[28];
  assign o[7274] = i[28];
  assign o[7275] = i[28];
  assign o[7276] = i[28];
  assign o[7277] = i[28];
  assign o[7278] = i[28];
  assign o[7279] = i[28];
  assign o[7280] = i[28];
  assign o[7281] = i[28];
  assign o[7282] = i[28];
  assign o[7283] = i[28];
  assign o[7284] = i[28];
  assign o[7285] = i[28];
  assign o[7286] = i[28];
  assign o[7287] = i[28];
  assign o[7288] = i[28];
  assign o[7289] = i[28];
  assign o[7290] = i[28];
  assign o[7291] = i[28];
  assign o[7292] = i[28];
  assign o[7293] = i[28];
  assign o[7294] = i[28];
  assign o[7295] = i[28];
  assign o[7296] = i[28];
  assign o[7297] = i[28];
  assign o[7298] = i[28];
  assign o[7299] = i[28];
  assign o[7300] = i[28];
  assign o[7301] = i[28];
  assign o[7302] = i[28];
  assign o[7303] = i[28];
  assign o[7304] = i[28];
  assign o[7305] = i[28];
  assign o[7306] = i[28];
  assign o[7307] = i[28];
  assign o[7308] = i[28];
  assign o[7309] = i[28];
  assign o[7310] = i[28];
  assign o[7311] = i[28];
  assign o[7312] = i[28];
  assign o[7313] = i[28];
  assign o[7314] = i[28];
  assign o[7315] = i[28];
  assign o[7316] = i[28];
  assign o[7317] = i[28];
  assign o[7318] = i[28];
  assign o[7319] = i[28];
  assign o[7320] = i[28];
  assign o[7321] = i[28];
  assign o[7322] = i[28];
  assign o[7323] = i[28];
  assign o[7324] = i[28];
  assign o[7325] = i[28];
  assign o[7326] = i[28];
  assign o[7327] = i[28];
  assign o[7328] = i[28];
  assign o[7329] = i[28];
  assign o[7330] = i[28];
  assign o[7331] = i[28];
  assign o[7332] = i[28];
  assign o[7333] = i[28];
  assign o[7334] = i[28];
  assign o[7335] = i[28];
  assign o[7336] = i[28];
  assign o[7337] = i[28];
  assign o[7338] = i[28];
  assign o[7339] = i[28];
  assign o[7340] = i[28];
  assign o[7341] = i[28];
  assign o[7342] = i[28];
  assign o[7343] = i[28];
  assign o[7344] = i[28];
  assign o[7345] = i[28];
  assign o[7346] = i[28];
  assign o[7347] = i[28];
  assign o[7348] = i[28];
  assign o[7349] = i[28];
  assign o[7350] = i[28];
  assign o[7351] = i[28];
  assign o[7352] = i[28];
  assign o[7353] = i[28];
  assign o[7354] = i[28];
  assign o[7355] = i[28];
  assign o[7356] = i[28];
  assign o[7357] = i[28];
  assign o[7358] = i[28];
  assign o[7359] = i[28];
  assign o[7360] = i[28];
  assign o[7361] = i[28];
  assign o[7362] = i[28];
  assign o[7363] = i[28];
  assign o[7364] = i[28];
  assign o[7365] = i[28];
  assign o[7366] = i[28];
  assign o[7367] = i[28];
  assign o[7368] = i[28];
  assign o[7369] = i[28];
  assign o[7370] = i[28];
  assign o[7371] = i[28];
  assign o[7372] = i[28];
  assign o[7373] = i[28];
  assign o[7374] = i[28];
  assign o[7375] = i[28];
  assign o[7376] = i[28];
  assign o[7377] = i[28];
  assign o[7378] = i[28];
  assign o[7379] = i[28];
  assign o[7380] = i[28];
  assign o[7381] = i[28];
  assign o[7382] = i[28];
  assign o[7383] = i[28];
  assign o[7384] = i[28];
  assign o[7385] = i[28];
  assign o[7386] = i[28];
  assign o[7387] = i[28];
  assign o[7388] = i[28];
  assign o[7389] = i[28];
  assign o[7390] = i[28];
  assign o[7391] = i[28];
  assign o[7392] = i[28];
  assign o[7393] = i[28];
  assign o[7394] = i[28];
  assign o[7395] = i[28];
  assign o[7396] = i[28];
  assign o[7397] = i[28];
  assign o[7398] = i[28];
  assign o[7399] = i[28];
  assign o[7400] = i[28];
  assign o[7401] = i[28];
  assign o[7402] = i[28];
  assign o[7403] = i[28];
  assign o[7404] = i[28];
  assign o[7405] = i[28];
  assign o[7406] = i[28];
  assign o[7407] = i[28];
  assign o[7408] = i[28];
  assign o[7409] = i[28];
  assign o[7410] = i[28];
  assign o[7411] = i[28];
  assign o[7412] = i[28];
  assign o[7413] = i[28];
  assign o[7414] = i[28];
  assign o[7415] = i[28];
  assign o[7416] = i[28];
  assign o[7417] = i[28];
  assign o[7418] = i[28];
  assign o[7419] = i[28];
  assign o[7420] = i[28];
  assign o[7421] = i[28];
  assign o[7422] = i[28];
  assign o[7423] = i[28];
  assign o[6912] = i[27];
  assign o[6913] = i[27];
  assign o[6914] = i[27];
  assign o[6915] = i[27];
  assign o[6916] = i[27];
  assign o[6917] = i[27];
  assign o[6918] = i[27];
  assign o[6919] = i[27];
  assign o[6920] = i[27];
  assign o[6921] = i[27];
  assign o[6922] = i[27];
  assign o[6923] = i[27];
  assign o[6924] = i[27];
  assign o[6925] = i[27];
  assign o[6926] = i[27];
  assign o[6927] = i[27];
  assign o[6928] = i[27];
  assign o[6929] = i[27];
  assign o[6930] = i[27];
  assign o[6931] = i[27];
  assign o[6932] = i[27];
  assign o[6933] = i[27];
  assign o[6934] = i[27];
  assign o[6935] = i[27];
  assign o[6936] = i[27];
  assign o[6937] = i[27];
  assign o[6938] = i[27];
  assign o[6939] = i[27];
  assign o[6940] = i[27];
  assign o[6941] = i[27];
  assign o[6942] = i[27];
  assign o[6943] = i[27];
  assign o[6944] = i[27];
  assign o[6945] = i[27];
  assign o[6946] = i[27];
  assign o[6947] = i[27];
  assign o[6948] = i[27];
  assign o[6949] = i[27];
  assign o[6950] = i[27];
  assign o[6951] = i[27];
  assign o[6952] = i[27];
  assign o[6953] = i[27];
  assign o[6954] = i[27];
  assign o[6955] = i[27];
  assign o[6956] = i[27];
  assign o[6957] = i[27];
  assign o[6958] = i[27];
  assign o[6959] = i[27];
  assign o[6960] = i[27];
  assign o[6961] = i[27];
  assign o[6962] = i[27];
  assign o[6963] = i[27];
  assign o[6964] = i[27];
  assign o[6965] = i[27];
  assign o[6966] = i[27];
  assign o[6967] = i[27];
  assign o[6968] = i[27];
  assign o[6969] = i[27];
  assign o[6970] = i[27];
  assign o[6971] = i[27];
  assign o[6972] = i[27];
  assign o[6973] = i[27];
  assign o[6974] = i[27];
  assign o[6975] = i[27];
  assign o[6976] = i[27];
  assign o[6977] = i[27];
  assign o[6978] = i[27];
  assign o[6979] = i[27];
  assign o[6980] = i[27];
  assign o[6981] = i[27];
  assign o[6982] = i[27];
  assign o[6983] = i[27];
  assign o[6984] = i[27];
  assign o[6985] = i[27];
  assign o[6986] = i[27];
  assign o[6987] = i[27];
  assign o[6988] = i[27];
  assign o[6989] = i[27];
  assign o[6990] = i[27];
  assign o[6991] = i[27];
  assign o[6992] = i[27];
  assign o[6993] = i[27];
  assign o[6994] = i[27];
  assign o[6995] = i[27];
  assign o[6996] = i[27];
  assign o[6997] = i[27];
  assign o[6998] = i[27];
  assign o[6999] = i[27];
  assign o[7000] = i[27];
  assign o[7001] = i[27];
  assign o[7002] = i[27];
  assign o[7003] = i[27];
  assign o[7004] = i[27];
  assign o[7005] = i[27];
  assign o[7006] = i[27];
  assign o[7007] = i[27];
  assign o[7008] = i[27];
  assign o[7009] = i[27];
  assign o[7010] = i[27];
  assign o[7011] = i[27];
  assign o[7012] = i[27];
  assign o[7013] = i[27];
  assign o[7014] = i[27];
  assign o[7015] = i[27];
  assign o[7016] = i[27];
  assign o[7017] = i[27];
  assign o[7018] = i[27];
  assign o[7019] = i[27];
  assign o[7020] = i[27];
  assign o[7021] = i[27];
  assign o[7022] = i[27];
  assign o[7023] = i[27];
  assign o[7024] = i[27];
  assign o[7025] = i[27];
  assign o[7026] = i[27];
  assign o[7027] = i[27];
  assign o[7028] = i[27];
  assign o[7029] = i[27];
  assign o[7030] = i[27];
  assign o[7031] = i[27];
  assign o[7032] = i[27];
  assign o[7033] = i[27];
  assign o[7034] = i[27];
  assign o[7035] = i[27];
  assign o[7036] = i[27];
  assign o[7037] = i[27];
  assign o[7038] = i[27];
  assign o[7039] = i[27];
  assign o[7040] = i[27];
  assign o[7041] = i[27];
  assign o[7042] = i[27];
  assign o[7043] = i[27];
  assign o[7044] = i[27];
  assign o[7045] = i[27];
  assign o[7046] = i[27];
  assign o[7047] = i[27];
  assign o[7048] = i[27];
  assign o[7049] = i[27];
  assign o[7050] = i[27];
  assign o[7051] = i[27];
  assign o[7052] = i[27];
  assign o[7053] = i[27];
  assign o[7054] = i[27];
  assign o[7055] = i[27];
  assign o[7056] = i[27];
  assign o[7057] = i[27];
  assign o[7058] = i[27];
  assign o[7059] = i[27];
  assign o[7060] = i[27];
  assign o[7061] = i[27];
  assign o[7062] = i[27];
  assign o[7063] = i[27];
  assign o[7064] = i[27];
  assign o[7065] = i[27];
  assign o[7066] = i[27];
  assign o[7067] = i[27];
  assign o[7068] = i[27];
  assign o[7069] = i[27];
  assign o[7070] = i[27];
  assign o[7071] = i[27];
  assign o[7072] = i[27];
  assign o[7073] = i[27];
  assign o[7074] = i[27];
  assign o[7075] = i[27];
  assign o[7076] = i[27];
  assign o[7077] = i[27];
  assign o[7078] = i[27];
  assign o[7079] = i[27];
  assign o[7080] = i[27];
  assign o[7081] = i[27];
  assign o[7082] = i[27];
  assign o[7083] = i[27];
  assign o[7084] = i[27];
  assign o[7085] = i[27];
  assign o[7086] = i[27];
  assign o[7087] = i[27];
  assign o[7088] = i[27];
  assign o[7089] = i[27];
  assign o[7090] = i[27];
  assign o[7091] = i[27];
  assign o[7092] = i[27];
  assign o[7093] = i[27];
  assign o[7094] = i[27];
  assign o[7095] = i[27];
  assign o[7096] = i[27];
  assign o[7097] = i[27];
  assign o[7098] = i[27];
  assign o[7099] = i[27];
  assign o[7100] = i[27];
  assign o[7101] = i[27];
  assign o[7102] = i[27];
  assign o[7103] = i[27];
  assign o[7104] = i[27];
  assign o[7105] = i[27];
  assign o[7106] = i[27];
  assign o[7107] = i[27];
  assign o[7108] = i[27];
  assign o[7109] = i[27];
  assign o[7110] = i[27];
  assign o[7111] = i[27];
  assign o[7112] = i[27];
  assign o[7113] = i[27];
  assign o[7114] = i[27];
  assign o[7115] = i[27];
  assign o[7116] = i[27];
  assign o[7117] = i[27];
  assign o[7118] = i[27];
  assign o[7119] = i[27];
  assign o[7120] = i[27];
  assign o[7121] = i[27];
  assign o[7122] = i[27];
  assign o[7123] = i[27];
  assign o[7124] = i[27];
  assign o[7125] = i[27];
  assign o[7126] = i[27];
  assign o[7127] = i[27];
  assign o[7128] = i[27];
  assign o[7129] = i[27];
  assign o[7130] = i[27];
  assign o[7131] = i[27];
  assign o[7132] = i[27];
  assign o[7133] = i[27];
  assign o[7134] = i[27];
  assign o[7135] = i[27];
  assign o[7136] = i[27];
  assign o[7137] = i[27];
  assign o[7138] = i[27];
  assign o[7139] = i[27];
  assign o[7140] = i[27];
  assign o[7141] = i[27];
  assign o[7142] = i[27];
  assign o[7143] = i[27];
  assign o[7144] = i[27];
  assign o[7145] = i[27];
  assign o[7146] = i[27];
  assign o[7147] = i[27];
  assign o[7148] = i[27];
  assign o[7149] = i[27];
  assign o[7150] = i[27];
  assign o[7151] = i[27];
  assign o[7152] = i[27];
  assign o[7153] = i[27];
  assign o[7154] = i[27];
  assign o[7155] = i[27];
  assign o[7156] = i[27];
  assign o[7157] = i[27];
  assign o[7158] = i[27];
  assign o[7159] = i[27];
  assign o[7160] = i[27];
  assign o[7161] = i[27];
  assign o[7162] = i[27];
  assign o[7163] = i[27];
  assign o[7164] = i[27];
  assign o[7165] = i[27];
  assign o[7166] = i[27];
  assign o[7167] = i[27];
  assign o[6656] = i[26];
  assign o[6657] = i[26];
  assign o[6658] = i[26];
  assign o[6659] = i[26];
  assign o[6660] = i[26];
  assign o[6661] = i[26];
  assign o[6662] = i[26];
  assign o[6663] = i[26];
  assign o[6664] = i[26];
  assign o[6665] = i[26];
  assign o[6666] = i[26];
  assign o[6667] = i[26];
  assign o[6668] = i[26];
  assign o[6669] = i[26];
  assign o[6670] = i[26];
  assign o[6671] = i[26];
  assign o[6672] = i[26];
  assign o[6673] = i[26];
  assign o[6674] = i[26];
  assign o[6675] = i[26];
  assign o[6676] = i[26];
  assign o[6677] = i[26];
  assign o[6678] = i[26];
  assign o[6679] = i[26];
  assign o[6680] = i[26];
  assign o[6681] = i[26];
  assign o[6682] = i[26];
  assign o[6683] = i[26];
  assign o[6684] = i[26];
  assign o[6685] = i[26];
  assign o[6686] = i[26];
  assign o[6687] = i[26];
  assign o[6688] = i[26];
  assign o[6689] = i[26];
  assign o[6690] = i[26];
  assign o[6691] = i[26];
  assign o[6692] = i[26];
  assign o[6693] = i[26];
  assign o[6694] = i[26];
  assign o[6695] = i[26];
  assign o[6696] = i[26];
  assign o[6697] = i[26];
  assign o[6698] = i[26];
  assign o[6699] = i[26];
  assign o[6700] = i[26];
  assign o[6701] = i[26];
  assign o[6702] = i[26];
  assign o[6703] = i[26];
  assign o[6704] = i[26];
  assign o[6705] = i[26];
  assign o[6706] = i[26];
  assign o[6707] = i[26];
  assign o[6708] = i[26];
  assign o[6709] = i[26];
  assign o[6710] = i[26];
  assign o[6711] = i[26];
  assign o[6712] = i[26];
  assign o[6713] = i[26];
  assign o[6714] = i[26];
  assign o[6715] = i[26];
  assign o[6716] = i[26];
  assign o[6717] = i[26];
  assign o[6718] = i[26];
  assign o[6719] = i[26];
  assign o[6720] = i[26];
  assign o[6721] = i[26];
  assign o[6722] = i[26];
  assign o[6723] = i[26];
  assign o[6724] = i[26];
  assign o[6725] = i[26];
  assign o[6726] = i[26];
  assign o[6727] = i[26];
  assign o[6728] = i[26];
  assign o[6729] = i[26];
  assign o[6730] = i[26];
  assign o[6731] = i[26];
  assign o[6732] = i[26];
  assign o[6733] = i[26];
  assign o[6734] = i[26];
  assign o[6735] = i[26];
  assign o[6736] = i[26];
  assign o[6737] = i[26];
  assign o[6738] = i[26];
  assign o[6739] = i[26];
  assign o[6740] = i[26];
  assign o[6741] = i[26];
  assign o[6742] = i[26];
  assign o[6743] = i[26];
  assign o[6744] = i[26];
  assign o[6745] = i[26];
  assign o[6746] = i[26];
  assign o[6747] = i[26];
  assign o[6748] = i[26];
  assign o[6749] = i[26];
  assign o[6750] = i[26];
  assign o[6751] = i[26];
  assign o[6752] = i[26];
  assign o[6753] = i[26];
  assign o[6754] = i[26];
  assign o[6755] = i[26];
  assign o[6756] = i[26];
  assign o[6757] = i[26];
  assign o[6758] = i[26];
  assign o[6759] = i[26];
  assign o[6760] = i[26];
  assign o[6761] = i[26];
  assign o[6762] = i[26];
  assign o[6763] = i[26];
  assign o[6764] = i[26];
  assign o[6765] = i[26];
  assign o[6766] = i[26];
  assign o[6767] = i[26];
  assign o[6768] = i[26];
  assign o[6769] = i[26];
  assign o[6770] = i[26];
  assign o[6771] = i[26];
  assign o[6772] = i[26];
  assign o[6773] = i[26];
  assign o[6774] = i[26];
  assign o[6775] = i[26];
  assign o[6776] = i[26];
  assign o[6777] = i[26];
  assign o[6778] = i[26];
  assign o[6779] = i[26];
  assign o[6780] = i[26];
  assign o[6781] = i[26];
  assign o[6782] = i[26];
  assign o[6783] = i[26];
  assign o[6784] = i[26];
  assign o[6785] = i[26];
  assign o[6786] = i[26];
  assign o[6787] = i[26];
  assign o[6788] = i[26];
  assign o[6789] = i[26];
  assign o[6790] = i[26];
  assign o[6791] = i[26];
  assign o[6792] = i[26];
  assign o[6793] = i[26];
  assign o[6794] = i[26];
  assign o[6795] = i[26];
  assign o[6796] = i[26];
  assign o[6797] = i[26];
  assign o[6798] = i[26];
  assign o[6799] = i[26];
  assign o[6800] = i[26];
  assign o[6801] = i[26];
  assign o[6802] = i[26];
  assign o[6803] = i[26];
  assign o[6804] = i[26];
  assign o[6805] = i[26];
  assign o[6806] = i[26];
  assign o[6807] = i[26];
  assign o[6808] = i[26];
  assign o[6809] = i[26];
  assign o[6810] = i[26];
  assign o[6811] = i[26];
  assign o[6812] = i[26];
  assign o[6813] = i[26];
  assign o[6814] = i[26];
  assign o[6815] = i[26];
  assign o[6816] = i[26];
  assign o[6817] = i[26];
  assign o[6818] = i[26];
  assign o[6819] = i[26];
  assign o[6820] = i[26];
  assign o[6821] = i[26];
  assign o[6822] = i[26];
  assign o[6823] = i[26];
  assign o[6824] = i[26];
  assign o[6825] = i[26];
  assign o[6826] = i[26];
  assign o[6827] = i[26];
  assign o[6828] = i[26];
  assign o[6829] = i[26];
  assign o[6830] = i[26];
  assign o[6831] = i[26];
  assign o[6832] = i[26];
  assign o[6833] = i[26];
  assign o[6834] = i[26];
  assign o[6835] = i[26];
  assign o[6836] = i[26];
  assign o[6837] = i[26];
  assign o[6838] = i[26];
  assign o[6839] = i[26];
  assign o[6840] = i[26];
  assign o[6841] = i[26];
  assign o[6842] = i[26];
  assign o[6843] = i[26];
  assign o[6844] = i[26];
  assign o[6845] = i[26];
  assign o[6846] = i[26];
  assign o[6847] = i[26];
  assign o[6848] = i[26];
  assign o[6849] = i[26];
  assign o[6850] = i[26];
  assign o[6851] = i[26];
  assign o[6852] = i[26];
  assign o[6853] = i[26];
  assign o[6854] = i[26];
  assign o[6855] = i[26];
  assign o[6856] = i[26];
  assign o[6857] = i[26];
  assign o[6858] = i[26];
  assign o[6859] = i[26];
  assign o[6860] = i[26];
  assign o[6861] = i[26];
  assign o[6862] = i[26];
  assign o[6863] = i[26];
  assign o[6864] = i[26];
  assign o[6865] = i[26];
  assign o[6866] = i[26];
  assign o[6867] = i[26];
  assign o[6868] = i[26];
  assign o[6869] = i[26];
  assign o[6870] = i[26];
  assign o[6871] = i[26];
  assign o[6872] = i[26];
  assign o[6873] = i[26];
  assign o[6874] = i[26];
  assign o[6875] = i[26];
  assign o[6876] = i[26];
  assign o[6877] = i[26];
  assign o[6878] = i[26];
  assign o[6879] = i[26];
  assign o[6880] = i[26];
  assign o[6881] = i[26];
  assign o[6882] = i[26];
  assign o[6883] = i[26];
  assign o[6884] = i[26];
  assign o[6885] = i[26];
  assign o[6886] = i[26];
  assign o[6887] = i[26];
  assign o[6888] = i[26];
  assign o[6889] = i[26];
  assign o[6890] = i[26];
  assign o[6891] = i[26];
  assign o[6892] = i[26];
  assign o[6893] = i[26];
  assign o[6894] = i[26];
  assign o[6895] = i[26];
  assign o[6896] = i[26];
  assign o[6897] = i[26];
  assign o[6898] = i[26];
  assign o[6899] = i[26];
  assign o[6900] = i[26];
  assign o[6901] = i[26];
  assign o[6902] = i[26];
  assign o[6903] = i[26];
  assign o[6904] = i[26];
  assign o[6905] = i[26];
  assign o[6906] = i[26];
  assign o[6907] = i[26];
  assign o[6908] = i[26];
  assign o[6909] = i[26];
  assign o[6910] = i[26];
  assign o[6911] = i[26];
  assign o[6400] = i[25];
  assign o[6401] = i[25];
  assign o[6402] = i[25];
  assign o[6403] = i[25];
  assign o[6404] = i[25];
  assign o[6405] = i[25];
  assign o[6406] = i[25];
  assign o[6407] = i[25];
  assign o[6408] = i[25];
  assign o[6409] = i[25];
  assign o[6410] = i[25];
  assign o[6411] = i[25];
  assign o[6412] = i[25];
  assign o[6413] = i[25];
  assign o[6414] = i[25];
  assign o[6415] = i[25];
  assign o[6416] = i[25];
  assign o[6417] = i[25];
  assign o[6418] = i[25];
  assign o[6419] = i[25];
  assign o[6420] = i[25];
  assign o[6421] = i[25];
  assign o[6422] = i[25];
  assign o[6423] = i[25];
  assign o[6424] = i[25];
  assign o[6425] = i[25];
  assign o[6426] = i[25];
  assign o[6427] = i[25];
  assign o[6428] = i[25];
  assign o[6429] = i[25];
  assign o[6430] = i[25];
  assign o[6431] = i[25];
  assign o[6432] = i[25];
  assign o[6433] = i[25];
  assign o[6434] = i[25];
  assign o[6435] = i[25];
  assign o[6436] = i[25];
  assign o[6437] = i[25];
  assign o[6438] = i[25];
  assign o[6439] = i[25];
  assign o[6440] = i[25];
  assign o[6441] = i[25];
  assign o[6442] = i[25];
  assign o[6443] = i[25];
  assign o[6444] = i[25];
  assign o[6445] = i[25];
  assign o[6446] = i[25];
  assign o[6447] = i[25];
  assign o[6448] = i[25];
  assign o[6449] = i[25];
  assign o[6450] = i[25];
  assign o[6451] = i[25];
  assign o[6452] = i[25];
  assign o[6453] = i[25];
  assign o[6454] = i[25];
  assign o[6455] = i[25];
  assign o[6456] = i[25];
  assign o[6457] = i[25];
  assign o[6458] = i[25];
  assign o[6459] = i[25];
  assign o[6460] = i[25];
  assign o[6461] = i[25];
  assign o[6462] = i[25];
  assign o[6463] = i[25];
  assign o[6464] = i[25];
  assign o[6465] = i[25];
  assign o[6466] = i[25];
  assign o[6467] = i[25];
  assign o[6468] = i[25];
  assign o[6469] = i[25];
  assign o[6470] = i[25];
  assign o[6471] = i[25];
  assign o[6472] = i[25];
  assign o[6473] = i[25];
  assign o[6474] = i[25];
  assign o[6475] = i[25];
  assign o[6476] = i[25];
  assign o[6477] = i[25];
  assign o[6478] = i[25];
  assign o[6479] = i[25];
  assign o[6480] = i[25];
  assign o[6481] = i[25];
  assign o[6482] = i[25];
  assign o[6483] = i[25];
  assign o[6484] = i[25];
  assign o[6485] = i[25];
  assign o[6486] = i[25];
  assign o[6487] = i[25];
  assign o[6488] = i[25];
  assign o[6489] = i[25];
  assign o[6490] = i[25];
  assign o[6491] = i[25];
  assign o[6492] = i[25];
  assign o[6493] = i[25];
  assign o[6494] = i[25];
  assign o[6495] = i[25];
  assign o[6496] = i[25];
  assign o[6497] = i[25];
  assign o[6498] = i[25];
  assign o[6499] = i[25];
  assign o[6500] = i[25];
  assign o[6501] = i[25];
  assign o[6502] = i[25];
  assign o[6503] = i[25];
  assign o[6504] = i[25];
  assign o[6505] = i[25];
  assign o[6506] = i[25];
  assign o[6507] = i[25];
  assign o[6508] = i[25];
  assign o[6509] = i[25];
  assign o[6510] = i[25];
  assign o[6511] = i[25];
  assign o[6512] = i[25];
  assign o[6513] = i[25];
  assign o[6514] = i[25];
  assign o[6515] = i[25];
  assign o[6516] = i[25];
  assign o[6517] = i[25];
  assign o[6518] = i[25];
  assign o[6519] = i[25];
  assign o[6520] = i[25];
  assign o[6521] = i[25];
  assign o[6522] = i[25];
  assign o[6523] = i[25];
  assign o[6524] = i[25];
  assign o[6525] = i[25];
  assign o[6526] = i[25];
  assign o[6527] = i[25];
  assign o[6528] = i[25];
  assign o[6529] = i[25];
  assign o[6530] = i[25];
  assign o[6531] = i[25];
  assign o[6532] = i[25];
  assign o[6533] = i[25];
  assign o[6534] = i[25];
  assign o[6535] = i[25];
  assign o[6536] = i[25];
  assign o[6537] = i[25];
  assign o[6538] = i[25];
  assign o[6539] = i[25];
  assign o[6540] = i[25];
  assign o[6541] = i[25];
  assign o[6542] = i[25];
  assign o[6543] = i[25];
  assign o[6544] = i[25];
  assign o[6545] = i[25];
  assign o[6546] = i[25];
  assign o[6547] = i[25];
  assign o[6548] = i[25];
  assign o[6549] = i[25];
  assign o[6550] = i[25];
  assign o[6551] = i[25];
  assign o[6552] = i[25];
  assign o[6553] = i[25];
  assign o[6554] = i[25];
  assign o[6555] = i[25];
  assign o[6556] = i[25];
  assign o[6557] = i[25];
  assign o[6558] = i[25];
  assign o[6559] = i[25];
  assign o[6560] = i[25];
  assign o[6561] = i[25];
  assign o[6562] = i[25];
  assign o[6563] = i[25];
  assign o[6564] = i[25];
  assign o[6565] = i[25];
  assign o[6566] = i[25];
  assign o[6567] = i[25];
  assign o[6568] = i[25];
  assign o[6569] = i[25];
  assign o[6570] = i[25];
  assign o[6571] = i[25];
  assign o[6572] = i[25];
  assign o[6573] = i[25];
  assign o[6574] = i[25];
  assign o[6575] = i[25];
  assign o[6576] = i[25];
  assign o[6577] = i[25];
  assign o[6578] = i[25];
  assign o[6579] = i[25];
  assign o[6580] = i[25];
  assign o[6581] = i[25];
  assign o[6582] = i[25];
  assign o[6583] = i[25];
  assign o[6584] = i[25];
  assign o[6585] = i[25];
  assign o[6586] = i[25];
  assign o[6587] = i[25];
  assign o[6588] = i[25];
  assign o[6589] = i[25];
  assign o[6590] = i[25];
  assign o[6591] = i[25];
  assign o[6592] = i[25];
  assign o[6593] = i[25];
  assign o[6594] = i[25];
  assign o[6595] = i[25];
  assign o[6596] = i[25];
  assign o[6597] = i[25];
  assign o[6598] = i[25];
  assign o[6599] = i[25];
  assign o[6600] = i[25];
  assign o[6601] = i[25];
  assign o[6602] = i[25];
  assign o[6603] = i[25];
  assign o[6604] = i[25];
  assign o[6605] = i[25];
  assign o[6606] = i[25];
  assign o[6607] = i[25];
  assign o[6608] = i[25];
  assign o[6609] = i[25];
  assign o[6610] = i[25];
  assign o[6611] = i[25];
  assign o[6612] = i[25];
  assign o[6613] = i[25];
  assign o[6614] = i[25];
  assign o[6615] = i[25];
  assign o[6616] = i[25];
  assign o[6617] = i[25];
  assign o[6618] = i[25];
  assign o[6619] = i[25];
  assign o[6620] = i[25];
  assign o[6621] = i[25];
  assign o[6622] = i[25];
  assign o[6623] = i[25];
  assign o[6624] = i[25];
  assign o[6625] = i[25];
  assign o[6626] = i[25];
  assign o[6627] = i[25];
  assign o[6628] = i[25];
  assign o[6629] = i[25];
  assign o[6630] = i[25];
  assign o[6631] = i[25];
  assign o[6632] = i[25];
  assign o[6633] = i[25];
  assign o[6634] = i[25];
  assign o[6635] = i[25];
  assign o[6636] = i[25];
  assign o[6637] = i[25];
  assign o[6638] = i[25];
  assign o[6639] = i[25];
  assign o[6640] = i[25];
  assign o[6641] = i[25];
  assign o[6642] = i[25];
  assign o[6643] = i[25];
  assign o[6644] = i[25];
  assign o[6645] = i[25];
  assign o[6646] = i[25];
  assign o[6647] = i[25];
  assign o[6648] = i[25];
  assign o[6649] = i[25];
  assign o[6650] = i[25];
  assign o[6651] = i[25];
  assign o[6652] = i[25];
  assign o[6653] = i[25];
  assign o[6654] = i[25];
  assign o[6655] = i[25];
  assign o[6144] = i[24];
  assign o[6145] = i[24];
  assign o[6146] = i[24];
  assign o[6147] = i[24];
  assign o[6148] = i[24];
  assign o[6149] = i[24];
  assign o[6150] = i[24];
  assign o[6151] = i[24];
  assign o[6152] = i[24];
  assign o[6153] = i[24];
  assign o[6154] = i[24];
  assign o[6155] = i[24];
  assign o[6156] = i[24];
  assign o[6157] = i[24];
  assign o[6158] = i[24];
  assign o[6159] = i[24];
  assign o[6160] = i[24];
  assign o[6161] = i[24];
  assign o[6162] = i[24];
  assign o[6163] = i[24];
  assign o[6164] = i[24];
  assign o[6165] = i[24];
  assign o[6166] = i[24];
  assign o[6167] = i[24];
  assign o[6168] = i[24];
  assign o[6169] = i[24];
  assign o[6170] = i[24];
  assign o[6171] = i[24];
  assign o[6172] = i[24];
  assign o[6173] = i[24];
  assign o[6174] = i[24];
  assign o[6175] = i[24];
  assign o[6176] = i[24];
  assign o[6177] = i[24];
  assign o[6178] = i[24];
  assign o[6179] = i[24];
  assign o[6180] = i[24];
  assign o[6181] = i[24];
  assign o[6182] = i[24];
  assign o[6183] = i[24];
  assign o[6184] = i[24];
  assign o[6185] = i[24];
  assign o[6186] = i[24];
  assign o[6187] = i[24];
  assign o[6188] = i[24];
  assign o[6189] = i[24];
  assign o[6190] = i[24];
  assign o[6191] = i[24];
  assign o[6192] = i[24];
  assign o[6193] = i[24];
  assign o[6194] = i[24];
  assign o[6195] = i[24];
  assign o[6196] = i[24];
  assign o[6197] = i[24];
  assign o[6198] = i[24];
  assign o[6199] = i[24];
  assign o[6200] = i[24];
  assign o[6201] = i[24];
  assign o[6202] = i[24];
  assign o[6203] = i[24];
  assign o[6204] = i[24];
  assign o[6205] = i[24];
  assign o[6206] = i[24];
  assign o[6207] = i[24];
  assign o[6208] = i[24];
  assign o[6209] = i[24];
  assign o[6210] = i[24];
  assign o[6211] = i[24];
  assign o[6212] = i[24];
  assign o[6213] = i[24];
  assign o[6214] = i[24];
  assign o[6215] = i[24];
  assign o[6216] = i[24];
  assign o[6217] = i[24];
  assign o[6218] = i[24];
  assign o[6219] = i[24];
  assign o[6220] = i[24];
  assign o[6221] = i[24];
  assign o[6222] = i[24];
  assign o[6223] = i[24];
  assign o[6224] = i[24];
  assign o[6225] = i[24];
  assign o[6226] = i[24];
  assign o[6227] = i[24];
  assign o[6228] = i[24];
  assign o[6229] = i[24];
  assign o[6230] = i[24];
  assign o[6231] = i[24];
  assign o[6232] = i[24];
  assign o[6233] = i[24];
  assign o[6234] = i[24];
  assign o[6235] = i[24];
  assign o[6236] = i[24];
  assign o[6237] = i[24];
  assign o[6238] = i[24];
  assign o[6239] = i[24];
  assign o[6240] = i[24];
  assign o[6241] = i[24];
  assign o[6242] = i[24];
  assign o[6243] = i[24];
  assign o[6244] = i[24];
  assign o[6245] = i[24];
  assign o[6246] = i[24];
  assign o[6247] = i[24];
  assign o[6248] = i[24];
  assign o[6249] = i[24];
  assign o[6250] = i[24];
  assign o[6251] = i[24];
  assign o[6252] = i[24];
  assign o[6253] = i[24];
  assign o[6254] = i[24];
  assign o[6255] = i[24];
  assign o[6256] = i[24];
  assign o[6257] = i[24];
  assign o[6258] = i[24];
  assign o[6259] = i[24];
  assign o[6260] = i[24];
  assign o[6261] = i[24];
  assign o[6262] = i[24];
  assign o[6263] = i[24];
  assign o[6264] = i[24];
  assign o[6265] = i[24];
  assign o[6266] = i[24];
  assign o[6267] = i[24];
  assign o[6268] = i[24];
  assign o[6269] = i[24];
  assign o[6270] = i[24];
  assign o[6271] = i[24];
  assign o[6272] = i[24];
  assign o[6273] = i[24];
  assign o[6274] = i[24];
  assign o[6275] = i[24];
  assign o[6276] = i[24];
  assign o[6277] = i[24];
  assign o[6278] = i[24];
  assign o[6279] = i[24];
  assign o[6280] = i[24];
  assign o[6281] = i[24];
  assign o[6282] = i[24];
  assign o[6283] = i[24];
  assign o[6284] = i[24];
  assign o[6285] = i[24];
  assign o[6286] = i[24];
  assign o[6287] = i[24];
  assign o[6288] = i[24];
  assign o[6289] = i[24];
  assign o[6290] = i[24];
  assign o[6291] = i[24];
  assign o[6292] = i[24];
  assign o[6293] = i[24];
  assign o[6294] = i[24];
  assign o[6295] = i[24];
  assign o[6296] = i[24];
  assign o[6297] = i[24];
  assign o[6298] = i[24];
  assign o[6299] = i[24];
  assign o[6300] = i[24];
  assign o[6301] = i[24];
  assign o[6302] = i[24];
  assign o[6303] = i[24];
  assign o[6304] = i[24];
  assign o[6305] = i[24];
  assign o[6306] = i[24];
  assign o[6307] = i[24];
  assign o[6308] = i[24];
  assign o[6309] = i[24];
  assign o[6310] = i[24];
  assign o[6311] = i[24];
  assign o[6312] = i[24];
  assign o[6313] = i[24];
  assign o[6314] = i[24];
  assign o[6315] = i[24];
  assign o[6316] = i[24];
  assign o[6317] = i[24];
  assign o[6318] = i[24];
  assign o[6319] = i[24];
  assign o[6320] = i[24];
  assign o[6321] = i[24];
  assign o[6322] = i[24];
  assign o[6323] = i[24];
  assign o[6324] = i[24];
  assign o[6325] = i[24];
  assign o[6326] = i[24];
  assign o[6327] = i[24];
  assign o[6328] = i[24];
  assign o[6329] = i[24];
  assign o[6330] = i[24];
  assign o[6331] = i[24];
  assign o[6332] = i[24];
  assign o[6333] = i[24];
  assign o[6334] = i[24];
  assign o[6335] = i[24];
  assign o[6336] = i[24];
  assign o[6337] = i[24];
  assign o[6338] = i[24];
  assign o[6339] = i[24];
  assign o[6340] = i[24];
  assign o[6341] = i[24];
  assign o[6342] = i[24];
  assign o[6343] = i[24];
  assign o[6344] = i[24];
  assign o[6345] = i[24];
  assign o[6346] = i[24];
  assign o[6347] = i[24];
  assign o[6348] = i[24];
  assign o[6349] = i[24];
  assign o[6350] = i[24];
  assign o[6351] = i[24];
  assign o[6352] = i[24];
  assign o[6353] = i[24];
  assign o[6354] = i[24];
  assign o[6355] = i[24];
  assign o[6356] = i[24];
  assign o[6357] = i[24];
  assign o[6358] = i[24];
  assign o[6359] = i[24];
  assign o[6360] = i[24];
  assign o[6361] = i[24];
  assign o[6362] = i[24];
  assign o[6363] = i[24];
  assign o[6364] = i[24];
  assign o[6365] = i[24];
  assign o[6366] = i[24];
  assign o[6367] = i[24];
  assign o[6368] = i[24];
  assign o[6369] = i[24];
  assign o[6370] = i[24];
  assign o[6371] = i[24];
  assign o[6372] = i[24];
  assign o[6373] = i[24];
  assign o[6374] = i[24];
  assign o[6375] = i[24];
  assign o[6376] = i[24];
  assign o[6377] = i[24];
  assign o[6378] = i[24];
  assign o[6379] = i[24];
  assign o[6380] = i[24];
  assign o[6381] = i[24];
  assign o[6382] = i[24];
  assign o[6383] = i[24];
  assign o[6384] = i[24];
  assign o[6385] = i[24];
  assign o[6386] = i[24];
  assign o[6387] = i[24];
  assign o[6388] = i[24];
  assign o[6389] = i[24];
  assign o[6390] = i[24];
  assign o[6391] = i[24];
  assign o[6392] = i[24];
  assign o[6393] = i[24];
  assign o[6394] = i[24];
  assign o[6395] = i[24];
  assign o[6396] = i[24];
  assign o[6397] = i[24];
  assign o[6398] = i[24];
  assign o[6399] = i[24];
  assign o[5888] = i[23];
  assign o[5889] = i[23];
  assign o[5890] = i[23];
  assign o[5891] = i[23];
  assign o[5892] = i[23];
  assign o[5893] = i[23];
  assign o[5894] = i[23];
  assign o[5895] = i[23];
  assign o[5896] = i[23];
  assign o[5897] = i[23];
  assign o[5898] = i[23];
  assign o[5899] = i[23];
  assign o[5900] = i[23];
  assign o[5901] = i[23];
  assign o[5902] = i[23];
  assign o[5903] = i[23];
  assign o[5904] = i[23];
  assign o[5905] = i[23];
  assign o[5906] = i[23];
  assign o[5907] = i[23];
  assign o[5908] = i[23];
  assign o[5909] = i[23];
  assign o[5910] = i[23];
  assign o[5911] = i[23];
  assign o[5912] = i[23];
  assign o[5913] = i[23];
  assign o[5914] = i[23];
  assign o[5915] = i[23];
  assign o[5916] = i[23];
  assign o[5917] = i[23];
  assign o[5918] = i[23];
  assign o[5919] = i[23];
  assign o[5920] = i[23];
  assign o[5921] = i[23];
  assign o[5922] = i[23];
  assign o[5923] = i[23];
  assign o[5924] = i[23];
  assign o[5925] = i[23];
  assign o[5926] = i[23];
  assign o[5927] = i[23];
  assign o[5928] = i[23];
  assign o[5929] = i[23];
  assign o[5930] = i[23];
  assign o[5931] = i[23];
  assign o[5932] = i[23];
  assign o[5933] = i[23];
  assign o[5934] = i[23];
  assign o[5935] = i[23];
  assign o[5936] = i[23];
  assign o[5937] = i[23];
  assign o[5938] = i[23];
  assign o[5939] = i[23];
  assign o[5940] = i[23];
  assign o[5941] = i[23];
  assign o[5942] = i[23];
  assign o[5943] = i[23];
  assign o[5944] = i[23];
  assign o[5945] = i[23];
  assign o[5946] = i[23];
  assign o[5947] = i[23];
  assign o[5948] = i[23];
  assign o[5949] = i[23];
  assign o[5950] = i[23];
  assign o[5951] = i[23];
  assign o[5952] = i[23];
  assign o[5953] = i[23];
  assign o[5954] = i[23];
  assign o[5955] = i[23];
  assign o[5956] = i[23];
  assign o[5957] = i[23];
  assign o[5958] = i[23];
  assign o[5959] = i[23];
  assign o[5960] = i[23];
  assign o[5961] = i[23];
  assign o[5962] = i[23];
  assign o[5963] = i[23];
  assign o[5964] = i[23];
  assign o[5965] = i[23];
  assign o[5966] = i[23];
  assign o[5967] = i[23];
  assign o[5968] = i[23];
  assign o[5969] = i[23];
  assign o[5970] = i[23];
  assign o[5971] = i[23];
  assign o[5972] = i[23];
  assign o[5973] = i[23];
  assign o[5974] = i[23];
  assign o[5975] = i[23];
  assign o[5976] = i[23];
  assign o[5977] = i[23];
  assign o[5978] = i[23];
  assign o[5979] = i[23];
  assign o[5980] = i[23];
  assign o[5981] = i[23];
  assign o[5982] = i[23];
  assign o[5983] = i[23];
  assign o[5984] = i[23];
  assign o[5985] = i[23];
  assign o[5986] = i[23];
  assign o[5987] = i[23];
  assign o[5988] = i[23];
  assign o[5989] = i[23];
  assign o[5990] = i[23];
  assign o[5991] = i[23];
  assign o[5992] = i[23];
  assign o[5993] = i[23];
  assign o[5994] = i[23];
  assign o[5995] = i[23];
  assign o[5996] = i[23];
  assign o[5997] = i[23];
  assign o[5998] = i[23];
  assign o[5999] = i[23];
  assign o[6000] = i[23];
  assign o[6001] = i[23];
  assign o[6002] = i[23];
  assign o[6003] = i[23];
  assign o[6004] = i[23];
  assign o[6005] = i[23];
  assign o[6006] = i[23];
  assign o[6007] = i[23];
  assign o[6008] = i[23];
  assign o[6009] = i[23];
  assign o[6010] = i[23];
  assign o[6011] = i[23];
  assign o[6012] = i[23];
  assign o[6013] = i[23];
  assign o[6014] = i[23];
  assign o[6015] = i[23];
  assign o[6016] = i[23];
  assign o[6017] = i[23];
  assign o[6018] = i[23];
  assign o[6019] = i[23];
  assign o[6020] = i[23];
  assign o[6021] = i[23];
  assign o[6022] = i[23];
  assign o[6023] = i[23];
  assign o[6024] = i[23];
  assign o[6025] = i[23];
  assign o[6026] = i[23];
  assign o[6027] = i[23];
  assign o[6028] = i[23];
  assign o[6029] = i[23];
  assign o[6030] = i[23];
  assign o[6031] = i[23];
  assign o[6032] = i[23];
  assign o[6033] = i[23];
  assign o[6034] = i[23];
  assign o[6035] = i[23];
  assign o[6036] = i[23];
  assign o[6037] = i[23];
  assign o[6038] = i[23];
  assign o[6039] = i[23];
  assign o[6040] = i[23];
  assign o[6041] = i[23];
  assign o[6042] = i[23];
  assign o[6043] = i[23];
  assign o[6044] = i[23];
  assign o[6045] = i[23];
  assign o[6046] = i[23];
  assign o[6047] = i[23];
  assign o[6048] = i[23];
  assign o[6049] = i[23];
  assign o[6050] = i[23];
  assign o[6051] = i[23];
  assign o[6052] = i[23];
  assign o[6053] = i[23];
  assign o[6054] = i[23];
  assign o[6055] = i[23];
  assign o[6056] = i[23];
  assign o[6057] = i[23];
  assign o[6058] = i[23];
  assign o[6059] = i[23];
  assign o[6060] = i[23];
  assign o[6061] = i[23];
  assign o[6062] = i[23];
  assign o[6063] = i[23];
  assign o[6064] = i[23];
  assign o[6065] = i[23];
  assign o[6066] = i[23];
  assign o[6067] = i[23];
  assign o[6068] = i[23];
  assign o[6069] = i[23];
  assign o[6070] = i[23];
  assign o[6071] = i[23];
  assign o[6072] = i[23];
  assign o[6073] = i[23];
  assign o[6074] = i[23];
  assign o[6075] = i[23];
  assign o[6076] = i[23];
  assign o[6077] = i[23];
  assign o[6078] = i[23];
  assign o[6079] = i[23];
  assign o[6080] = i[23];
  assign o[6081] = i[23];
  assign o[6082] = i[23];
  assign o[6083] = i[23];
  assign o[6084] = i[23];
  assign o[6085] = i[23];
  assign o[6086] = i[23];
  assign o[6087] = i[23];
  assign o[6088] = i[23];
  assign o[6089] = i[23];
  assign o[6090] = i[23];
  assign o[6091] = i[23];
  assign o[6092] = i[23];
  assign o[6093] = i[23];
  assign o[6094] = i[23];
  assign o[6095] = i[23];
  assign o[6096] = i[23];
  assign o[6097] = i[23];
  assign o[6098] = i[23];
  assign o[6099] = i[23];
  assign o[6100] = i[23];
  assign o[6101] = i[23];
  assign o[6102] = i[23];
  assign o[6103] = i[23];
  assign o[6104] = i[23];
  assign o[6105] = i[23];
  assign o[6106] = i[23];
  assign o[6107] = i[23];
  assign o[6108] = i[23];
  assign o[6109] = i[23];
  assign o[6110] = i[23];
  assign o[6111] = i[23];
  assign o[6112] = i[23];
  assign o[6113] = i[23];
  assign o[6114] = i[23];
  assign o[6115] = i[23];
  assign o[6116] = i[23];
  assign o[6117] = i[23];
  assign o[6118] = i[23];
  assign o[6119] = i[23];
  assign o[6120] = i[23];
  assign o[6121] = i[23];
  assign o[6122] = i[23];
  assign o[6123] = i[23];
  assign o[6124] = i[23];
  assign o[6125] = i[23];
  assign o[6126] = i[23];
  assign o[6127] = i[23];
  assign o[6128] = i[23];
  assign o[6129] = i[23];
  assign o[6130] = i[23];
  assign o[6131] = i[23];
  assign o[6132] = i[23];
  assign o[6133] = i[23];
  assign o[6134] = i[23];
  assign o[6135] = i[23];
  assign o[6136] = i[23];
  assign o[6137] = i[23];
  assign o[6138] = i[23];
  assign o[6139] = i[23];
  assign o[6140] = i[23];
  assign o[6141] = i[23];
  assign o[6142] = i[23];
  assign o[6143] = i[23];
  assign o[5632] = i[22];
  assign o[5633] = i[22];
  assign o[5634] = i[22];
  assign o[5635] = i[22];
  assign o[5636] = i[22];
  assign o[5637] = i[22];
  assign o[5638] = i[22];
  assign o[5639] = i[22];
  assign o[5640] = i[22];
  assign o[5641] = i[22];
  assign o[5642] = i[22];
  assign o[5643] = i[22];
  assign o[5644] = i[22];
  assign o[5645] = i[22];
  assign o[5646] = i[22];
  assign o[5647] = i[22];
  assign o[5648] = i[22];
  assign o[5649] = i[22];
  assign o[5650] = i[22];
  assign o[5651] = i[22];
  assign o[5652] = i[22];
  assign o[5653] = i[22];
  assign o[5654] = i[22];
  assign o[5655] = i[22];
  assign o[5656] = i[22];
  assign o[5657] = i[22];
  assign o[5658] = i[22];
  assign o[5659] = i[22];
  assign o[5660] = i[22];
  assign o[5661] = i[22];
  assign o[5662] = i[22];
  assign o[5663] = i[22];
  assign o[5664] = i[22];
  assign o[5665] = i[22];
  assign o[5666] = i[22];
  assign o[5667] = i[22];
  assign o[5668] = i[22];
  assign o[5669] = i[22];
  assign o[5670] = i[22];
  assign o[5671] = i[22];
  assign o[5672] = i[22];
  assign o[5673] = i[22];
  assign o[5674] = i[22];
  assign o[5675] = i[22];
  assign o[5676] = i[22];
  assign o[5677] = i[22];
  assign o[5678] = i[22];
  assign o[5679] = i[22];
  assign o[5680] = i[22];
  assign o[5681] = i[22];
  assign o[5682] = i[22];
  assign o[5683] = i[22];
  assign o[5684] = i[22];
  assign o[5685] = i[22];
  assign o[5686] = i[22];
  assign o[5687] = i[22];
  assign o[5688] = i[22];
  assign o[5689] = i[22];
  assign o[5690] = i[22];
  assign o[5691] = i[22];
  assign o[5692] = i[22];
  assign o[5693] = i[22];
  assign o[5694] = i[22];
  assign o[5695] = i[22];
  assign o[5696] = i[22];
  assign o[5697] = i[22];
  assign o[5698] = i[22];
  assign o[5699] = i[22];
  assign o[5700] = i[22];
  assign o[5701] = i[22];
  assign o[5702] = i[22];
  assign o[5703] = i[22];
  assign o[5704] = i[22];
  assign o[5705] = i[22];
  assign o[5706] = i[22];
  assign o[5707] = i[22];
  assign o[5708] = i[22];
  assign o[5709] = i[22];
  assign o[5710] = i[22];
  assign o[5711] = i[22];
  assign o[5712] = i[22];
  assign o[5713] = i[22];
  assign o[5714] = i[22];
  assign o[5715] = i[22];
  assign o[5716] = i[22];
  assign o[5717] = i[22];
  assign o[5718] = i[22];
  assign o[5719] = i[22];
  assign o[5720] = i[22];
  assign o[5721] = i[22];
  assign o[5722] = i[22];
  assign o[5723] = i[22];
  assign o[5724] = i[22];
  assign o[5725] = i[22];
  assign o[5726] = i[22];
  assign o[5727] = i[22];
  assign o[5728] = i[22];
  assign o[5729] = i[22];
  assign o[5730] = i[22];
  assign o[5731] = i[22];
  assign o[5732] = i[22];
  assign o[5733] = i[22];
  assign o[5734] = i[22];
  assign o[5735] = i[22];
  assign o[5736] = i[22];
  assign o[5737] = i[22];
  assign o[5738] = i[22];
  assign o[5739] = i[22];
  assign o[5740] = i[22];
  assign o[5741] = i[22];
  assign o[5742] = i[22];
  assign o[5743] = i[22];
  assign o[5744] = i[22];
  assign o[5745] = i[22];
  assign o[5746] = i[22];
  assign o[5747] = i[22];
  assign o[5748] = i[22];
  assign o[5749] = i[22];
  assign o[5750] = i[22];
  assign o[5751] = i[22];
  assign o[5752] = i[22];
  assign o[5753] = i[22];
  assign o[5754] = i[22];
  assign o[5755] = i[22];
  assign o[5756] = i[22];
  assign o[5757] = i[22];
  assign o[5758] = i[22];
  assign o[5759] = i[22];
  assign o[5760] = i[22];
  assign o[5761] = i[22];
  assign o[5762] = i[22];
  assign o[5763] = i[22];
  assign o[5764] = i[22];
  assign o[5765] = i[22];
  assign o[5766] = i[22];
  assign o[5767] = i[22];
  assign o[5768] = i[22];
  assign o[5769] = i[22];
  assign o[5770] = i[22];
  assign o[5771] = i[22];
  assign o[5772] = i[22];
  assign o[5773] = i[22];
  assign o[5774] = i[22];
  assign o[5775] = i[22];
  assign o[5776] = i[22];
  assign o[5777] = i[22];
  assign o[5778] = i[22];
  assign o[5779] = i[22];
  assign o[5780] = i[22];
  assign o[5781] = i[22];
  assign o[5782] = i[22];
  assign o[5783] = i[22];
  assign o[5784] = i[22];
  assign o[5785] = i[22];
  assign o[5786] = i[22];
  assign o[5787] = i[22];
  assign o[5788] = i[22];
  assign o[5789] = i[22];
  assign o[5790] = i[22];
  assign o[5791] = i[22];
  assign o[5792] = i[22];
  assign o[5793] = i[22];
  assign o[5794] = i[22];
  assign o[5795] = i[22];
  assign o[5796] = i[22];
  assign o[5797] = i[22];
  assign o[5798] = i[22];
  assign o[5799] = i[22];
  assign o[5800] = i[22];
  assign o[5801] = i[22];
  assign o[5802] = i[22];
  assign o[5803] = i[22];
  assign o[5804] = i[22];
  assign o[5805] = i[22];
  assign o[5806] = i[22];
  assign o[5807] = i[22];
  assign o[5808] = i[22];
  assign o[5809] = i[22];
  assign o[5810] = i[22];
  assign o[5811] = i[22];
  assign o[5812] = i[22];
  assign o[5813] = i[22];
  assign o[5814] = i[22];
  assign o[5815] = i[22];
  assign o[5816] = i[22];
  assign o[5817] = i[22];
  assign o[5818] = i[22];
  assign o[5819] = i[22];
  assign o[5820] = i[22];
  assign o[5821] = i[22];
  assign o[5822] = i[22];
  assign o[5823] = i[22];
  assign o[5824] = i[22];
  assign o[5825] = i[22];
  assign o[5826] = i[22];
  assign o[5827] = i[22];
  assign o[5828] = i[22];
  assign o[5829] = i[22];
  assign o[5830] = i[22];
  assign o[5831] = i[22];
  assign o[5832] = i[22];
  assign o[5833] = i[22];
  assign o[5834] = i[22];
  assign o[5835] = i[22];
  assign o[5836] = i[22];
  assign o[5837] = i[22];
  assign o[5838] = i[22];
  assign o[5839] = i[22];
  assign o[5840] = i[22];
  assign o[5841] = i[22];
  assign o[5842] = i[22];
  assign o[5843] = i[22];
  assign o[5844] = i[22];
  assign o[5845] = i[22];
  assign o[5846] = i[22];
  assign o[5847] = i[22];
  assign o[5848] = i[22];
  assign o[5849] = i[22];
  assign o[5850] = i[22];
  assign o[5851] = i[22];
  assign o[5852] = i[22];
  assign o[5853] = i[22];
  assign o[5854] = i[22];
  assign o[5855] = i[22];
  assign o[5856] = i[22];
  assign o[5857] = i[22];
  assign o[5858] = i[22];
  assign o[5859] = i[22];
  assign o[5860] = i[22];
  assign o[5861] = i[22];
  assign o[5862] = i[22];
  assign o[5863] = i[22];
  assign o[5864] = i[22];
  assign o[5865] = i[22];
  assign o[5866] = i[22];
  assign o[5867] = i[22];
  assign o[5868] = i[22];
  assign o[5869] = i[22];
  assign o[5870] = i[22];
  assign o[5871] = i[22];
  assign o[5872] = i[22];
  assign o[5873] = i[22];
  assign o[5874] = i[22];
  assign o[5875] = i[22];
  assign o[5876] = i[22];
  assign o[5877] = i[22];
  assign o[5878] = i[22];
  assign o[5879] = i[22];
  assign o[5880] = i[22];
  assign o[5881] = i[22];
  assign o[5882] = i[22];
  assign o[5883] = i[22];
  assign o[5884] = i[22];
  assign o[5885] = i[22];
  assign o[5886] = i[22];
  assign o[5887] = i[22];
  assign o[5376] = i[21];
  assign o[5377] = i[21];
  assign o[5378] = i[21];
  assign o[5379] = i[21];
  assign o[5380] = i[21];
  assign o[5381] = i[21];
  assign o[5382] = i[21];
  assign o[5383] = i[21];
  assign o[5384] = i[21];
  assign o[5385] = i[21];
  assign o[5386] = i[21];
  assign o[5387] = i[21];
  assign o[5388] = i[21];
  assign o[5389] = i[21];
  assign o[5390] = i[21];
  assign o[5391] = i[21];
  assign o[5392] = i[21];
  assign o[5393] = i[21];
  assign o[5394] = i[21];
  assign o[5395] = i[21];
  assign o[5396] = i[21];
  assign o[5397] = i[21];
  assign o[5398] = i[21];
  assign o[5399] = i[21];
  assign o[5400] = i[21];
  assign o[5401] = i[21];
  assign o[5402] = i[21];
  assign o[5403] = i[21];
  assign o[5404] = i[21];
  assign o[5405] = i[21];
  assign o[5406] = i[21];
  assign o[5407] = i[21];
  assign o[5408] = i[21];
  assign o[5409] = i[21];
  assign o[5410] = i[21];
  assign o[5411] = i[21];
  assign o[5412] = i[21];
  assign o[5413] = i[21];
  assign o[5414] = i[21];
  assign o[5415] = i[21];
  assign o[5416] = i[21];
  assign o[5417] = i[21];
  assign o[5418] = i[21];
  assign o[5419] = i[21];
  assign o[5420] = i[21];
  assign o[5421] = i[21];
  assign o[5422] = i[21];
  assign o[5423] = i[21];
  assign o[5424] = i[21];
  assign o[5425] = i[21];
  assign o[5426] = i[21];
  assign o[5427] = i[21];
  assign o[5428] = i[21];
  assign o[5429] = i[21];
  assign o[5430] = i[21];
  assign o[5431] = i[21];
  assign o[5432] = i[21];
  assign o[5433] = i[21];
  assign o[5434] = i[21];
  assign o[5435] = i[21];
  assign o[5436] = i[21];
  assign o[5437] = i[21];
  assign o[5438] = i[21];
  assign o[5439] = i[21];
  assign o[5440] = i[21];
  assign o[5441] = i[21];
  assign o[5442] = i[21];
  assign o[5443] = i[21];
  assign o[5444] = i[21];
  assign o[5445] = i[21];
  assign o[5446] = i[21];
  assign o[5447] = i[21];
  assign o[5448] = i[21];
  assign o[5449] = i[21];
  assign o[5450] = i[21];
  assign o[5451] = i[21];
  assign o[5452] = i[21];
  assign o[5453] = i[21];
  assign o[5454] = i[21];
  assign o[5455] = i[21];
  assign o[5456] = i[21];
  assign o[5457] = i[21];
  assign o[5458] = i[21];
  assign o[5459] = i[21];
  assign o[5460] = i[21];
  assign o[5461] = i[21];
  assign o[5462] = i[21];
  assign o[5463] = i[21];
  assign o[5464] = i[21];
  assign o[5465] = i[21];
  assign o[5466] = i[21];
  assign o[5467] = i[21];
  assign o[5468] = i[21];
  assign o[5469] = i[21];
  assign o[5470] = i[21];
  assign o[5471] = i[21];
  assign o[5472] = i[21];
  assign o[5473] = i[21];
  assign o[5474] = i[21];
  assign o[5475] = i[21];
  assign o[5476] = i[21];
  assign o[5477] = i[21];
  assign o[5478] = i[21];
  assign o[5479] = i[21];
  assign o[5480] = i[21];
  assign o[5481] = i[21];
  assign o[5482] = i[21];
  assign o[5483] = i[21];
  assign o[5484] = i[21];
  assign o[5485] = i[21];
  assign o[5486] = i[21];
  assign o[5487] = i[21];
  assign o[5488] = i[21];
  assign o[5489] = i[21];
  assign o[5490] = i[21];
  assign o[5491] = i[21];
  assign o[5492] = i[21];
  assign o[5493] = i[21];
  assign o[5494] = i[21];
  assign o[5495] = i[21];
  assign o[5496] = i[21];
  assign o[5497] = i[21];
  assign o[5498] = i[21];
  assign o[5499] = i[21];
  assign o[5500] = i[21];
  assign o[5501] = i[21];
  assign o[5502] = i[21];
  assign o[5503] = i[21];
  assign o[5504] = i[21];
  assign o[5505] = i[21];
  assign o[5506] = i[21];
  assign o[5507] = i[21];
  assign o[5508] = i[21];
  assign o[5509] = i[21];
  assign o[5510] = i[21];
  assign o[5511] = i[21];
  assign o[5512] = i[21];
  assign o[5513] = i[21];
  assign o[5514] = i[21];
  assign o[5515] = i[21];
  assign o[5516] = i[21];
  assign o[5517] = i[21];
  assign o[5518] = i[21];
  assign o[5519] = i[21];
  assign o[5520] = i[21];
  assign o[5521] = i[21];
  assign o[5522] = i[21];
  assign o[5523] = i[21];
  assign o[5524] = i[21];
  assign o[5525] = i[21];
  assign o[5526] = i[21];
  assign o[5527] = i[21];
  assign o[5528] = i[21];
  assign o[5529] = i[21];
  assign o[5530] = i[21];
  assign o[5531] = i[21];
  assign o[5532] = i[21];
  assign o[5533] = i[21];
  assign o[5534] = i[21];
  assign o[5535] = i[21];
  assign o[5536] = i[21];
  assign o[5537] = i[21];
  assign o[5538] = i[21];
  assign o[5539] = i[21];
  assign o[5540] = i[21];
  assign o[5541] = i[21];
  assign o[5542] = i[21];
  assign o[5543] = i[21];
  assign o[5544] = i[21];
  assign o[5545] = i[21];
  assign o[5546] = i[21];
  assign o[5547] = i[21];
  assign o[5548] = i[21];
  assign o[5549] = i[21];
  assign o[5550] = i[21];
  assign o[5551] = i[21];
  assign o[5552] = i[21];
  assign o[5553] = i[21];
  assign o[5554] = i[21];
  assign o[5555] = i[21];
  assign o[5556] = i[21];
  assign o[5557] = i[21];
  assign o[5558] = i[21];
  assign o[5559] = i[21];
  assign o[5560] = i[21];
  assign o[5561] = i[21];
  assign o[5562] = i[21];
  assign o[5563] = i[21];
  assign o[5564] = i[21];
  assign o[5565] = i[21];
  assign o[5566] = i[21];
  assign o[5567] = i[21];
  assign o[5568] = i[21];
  assign o[5569] = i[21];
  assign o[5570] = i[21];
  assign o[5571] = i[21];
  assign o[5572] = i[21];
  assign o[5573] = i[21];
  assign o[5574] = i[21];
  assign o[5575] = i[21];
  assign o[5576] = i[21];
  assign o[5577] = i[21];
  assign o[5578] = i[21];
  assign o[5579] = i[21];
  assign o[5580] = i[21];
  assign o[5581] = i[21];
  assign o[5582] = i[21];
  assign o[5583] = i[21];
  assign o[5584] = i[21];
  assign o[5585] = i[21];
  assign o[5586] = i[21];
  assign o[5587] = i[21];
  assign o[5588] = i[21];
  assign o[5589] = i[21];
  assign o[5590] = i[21];
  assign o[5591] = i[21];
  assign o[5592] = i[21];
  assign o[5593] = i[21];
  assign o[5594] = i[21];
  assign o[5595] = i[21];
  assign o[5596] = i[21];
  assign o[5597] = i[21];
  assign o[5598] = i[21];
  assign o[5599] = i[21];
  assign o[5600] = i[21];
  assign o[5601] = i[21];
  assign o[5602] = i[21];
  assign o[5603] = i[21];
  assign o[5604] = i[21];
  assign o[5605] = i[21];
  assign o[5606] = i[21];
  assign o[5607] = i[21];
  assign o[5608] = i[21];
  assign o[5609] = i[21];
  assign o[5610] = i[21];
  assign o[5611] = i[21];
  assign o[5612] = i[21];
  assign o[5613] = i[21];
  assign o[5614] = i[21];
  assign o[5615] = i[21];
  assign o[5616] = i[21];
  assign o[5617] = i[21];
  assign o[5618] = i[21];
  assign o[5619] = i[21];
  assign o[5620] = i[21];
  assign o[5621] = i[21];
  assign o[5622] = i[21];
  assign o[5623] = i[21];
  assign o[5624] = i[21];
  assign o[5625] = i[21];
  assign o[5626] = i[21];
  assign o[5627] = i[21];
  assign o[5628] = i[21];
  assign o[5629] = i[21];
  assign o[5630] = i[21];
  assign o[5631] = i[21];
  assign o[5120] = i[20];
  assign o[5121] = i[20];
  assign o[5122] = i[20];
  assign o[5123] = i[20];
  assign o[5124] = i[20];
  assign o[5125] = i[20];
  assign o[5126] = i[20];
  assign o[5127] = i[20];
  assign o[5128] = i[20];
  assign o[5129] = i[20];
  assign o[5130] = i[20];
  assign o[5131] = i[20];
  assign o[5132] = i[20];
  assign o[5133] = i[20];
  assign o[5134] = i[20];
  assign o[5135] = i[20];
  assign o[5136] = i[20];
  assign o[5137] = i[20];
  assign o[5138] = i[20];
  assign o[5139] = i[20];
  assign o[5140] = i[20];
  assign o[5141] = i[20];
  assign o[5142] = i[20];
  assign o[5143] = i[20];
  assign o[5144] = i[20];
  assign o[5145] = i[20];
  assign o[5146] = i[20];
  assign o[5147] = i[20];
  assign o[5148] = i[20];
  assign o[5149] = i[20];
  assign o[5150] = i[20];
  assign o[5151] = i[20];
  assign o[5152] = i[20];
  assign o[5153] = i[20];
  assign o[5154] = i[20];
  assign o[5155] = i[20];
  assign o[5156] = i[20];
  assign o[5157] = i[20];
  assign o[5158] = i[20];
  assign o[5159] = i[20];
  assign o[5160] = i[20];
  assign o[5161] = i[20];
  assign o[5162] = i[20];
  assign o[5163] = i[20];
  assign o[5164] = i[20];
  assign o[5165] = i[20];
  assign o[5166] = i[20];
  assign o[5167] = i[20];
  assign o[5168] = i[20];
  assign o[5169] = i[20];
  assign o[5170] = i[20];
  assign o[5171] = i[20];
  assign o[5172] = i[20];
  assign o[5173] = i[20];
  assign o[5174] = i[20];
  assign o[5175] = i[20];
  assign o[5176] = i[20];
  assign o[5177] = i[20];
  assign o[5178] = i[20];
  assign o[5179] = i[20];
  assign o[5180] = i[20];
  assign o[5181] = i[20];
  assign o[5182] = i[20];
  assign o[5183] = i[20];
  assign o[5184] = i[20];
  assign o[5185] = i[20];
  assign o[5186] = i[20];
  assign o[5187] = i[20];
  assign o[5188] = i[20];
  assign o[5189] = i[20];
  assign o[5190] = i[20];
  assign o[5191] = i[20];
  assign o[5192] = i[20];
  assign o[5193] = i[20];
  assign o[5194] = i[20];
  assign o[5195] = i[20];
  assign o[5196] = i[20];
  assign o[5197] = i[20];
  assign o[5198] = i[20];
  assign o[5199] = i[20];
  assign o[5200] = i[20];
  assign o[5201] = i[20];
  assign o[5202] = i[20];
  assign o[5203] = i[20];
  assign o[5204] = i[20];
  assign o[5205] = i[20];
  assign o[5206] = i[20];
  assign o[5207] = i[20];
  assign o[5208] = i[20];
  assign o[5209] = i[20];
  assign o[5210] = i[20];
  assign o[5211] = i[20];
  assign o[5212] = i[20];
  assign o[5213] = i[20];
  assign o[5214] = i[20];
  assign o[5215] = i[20];
  assign o[5216] = i[20];
  assign o[5217] = i[20];
  assign o[5218] = i[20];
  assign o[5219] = i[20];
  assign o[5220] = i[20];
  assign o[5221] = i[20];
  assign o[5222] = i[20];
  assign o[5223] = i[20];
  assign o[5224] = i[20];
  assign o[5225] = i[20];
  assign o[5226] = i[20];
  assign o[5227] = i[20];
  assign o[5228] = i[20];
  assign o[5229] = i[20];
  assign o[5230] = i[20];
  assign o[5231] = i[20];
  assign o[5232] = i[20];
  assign o[5233] = i[20];
  assign o[5234] = i[20];
  assign o[5235] = i[20];
  assign o[5236] = i[20];
  assign o[5237] = i[20];
  assign o[5238] = i[20];
  assign o[5239] = i[20];
  assign o[5240] = i[20];
  assign o[5241] = i[20];
  assign o[5242] = i[20];
  assign o[5243] = i[20];
  assign o[5244] = i[20];
  assign o[5245] = i[20];
  assign o[5246] = i[20];
  assign o[5247] = i[20];
  assign o[5248] = i[20];
  assign o[5249] = i[20];
  assign o[5250] = i[20];
  assign o[5251] = i[20];
  assign o[5252] = i[20];
  assign o[5253] = i[20];
  assign o[5254] = i[20];
  assign o[5255] = i[20];
  assign o[5256] = i[20];
  assign o[5257] = i[20];
  assign o[5258] = i[20];
  assign o[5259] = i[20];
  assign o[5260] = i[20];
  assign o[5261] = i[20];
  assign o[5262] = i[20];
  assign o[5263] = i[20];
  assign o[5264] = i[20];
  assign o[5265] = i[20];
  assign o[5266] = i[20];
  assign o[5267] = i[20];
  assign o[5268] = i[20];
  assign o[5269] = i[20];
  assign o[5270] = i[20];
  assign o[5271] = i[20];
  assign o[5272] = i[20];
  assign o[5273] = i[20];
  assign o[5274] = i[20];
  assign o[5275] = i[20];
  assign o[5276] = i[20];
  assign o[5277] = i[20];
  assign o[5278] = i[20];
  assign o[5279] = i[20];
  assign o[5280] = i[20];
  assign o[5281] = i[20];
  assign o[5282] = i[20];
  assign o[5283] = i[20];
  assign o[5284] = i[20];
  assign o[5285] = i[20];
  assign o[5286] = i[20];
  assign o[5287] = i[20];
  assign o[5288] = i[20];
  assign o[5289] = i[20];
  assign o[5290] = i[20];
  assign o[5291] = i[20];
  assign o[5292] = i[20];
  assign o[5293] = i[20];
  assign o[5294] = i[20];
  assign o[5295] = i[20];
  assign o[5296] = i[20];
  assign o[5297] = i[20];
  assign o[5298] = i[20];
  assign o[5299] = i[20];
  assign o[5300] = i[20];
  assign o[5301] = i[20];
  assign o[5302] = i[20];
  assign o[5303] = i[20];
  assign o[5304] = i[20];
  assign o[5305] = i[20];
  assign o[5306] = i[20];
  assign o[5307] = i[20];
  assign o[5308] = i[20];
  assign o[5309] = i[20];
  assign o[5310] = i[20];
  assign o[5311] = i[20];
  assign o[5312] = i[20];
  assign o[5313] = i[20];
  assign o[5314] = i[20];
  assign o[5315] = i[20];
  assign o[5316] = i[20];
  assign o[5317] = i[20];
  assign o[5318] = i[20];
  assign o[5319] = i[20];
  assign o[5320] = i[20];
  assign o[5321] = i[20];
  assign o[5322] = i[20];
  assign o[5323] = i[20];
  assign o[5324] = i[20];
  assign o[5325] = i[20];
  assign o[5326] = i[20];
  assign o[5327] = i[20];
  assign o[5328] = i[20];
  assign o[5329] = i[20];
  assign o[5330] = i[20];
  assign o[5331] = i[20];
  assign o[5332] = i[20];
  assign o[5333] = i[20];
  assign o[5334] = i[20];
  assign o[5335] = i[20];
  assign o[5336] = i[20];
  assign o[5337] = i[20];
  assign o[5338] = i[20];
  assign o[5339] = i[20];
  assign o[5340] = i[20];
  assign o[5341] = i[20];
  assign o[5342] = i[20];
  assign o[5343] = i[20];
  assign o[5344] = i[20];
  assign o[5345] = i[20];
  assign o[5346] = i[20];
  assign o[5347] = i[20];
  assign o[5348] = i[20];
  assign o[5349] = i[20];
  assign o[5350] = i[20];
  assign o[5351] = i[20];
  assign o[5352] = i[20];
  assign o[5353] = i[20];
  assign o[5354] = i[20];
  assign o[5355] = i[20];
  assign o[5356] = i[20];
  assign o[5357] = i[20];
  assign o[5358] = i[20];
  assign o[5359] = i[20];
  assign o[5360] = i[20];
  assign o[5361] = i[20];
  assign o[5362] = i[20];
  assign o[5363] = i[20];
  assign o[5364] = i[20];
  assign o[5365] = i[20];
  assign o[5366] = i[20];
  assign o[5367] = i[20];
  assign o[5368] = i[20];
  assign o[5369] = i[20];
  assign o[5370] = i[20];
  assign o[5371] = i[20];
  assign o[5372] = i[20];
  assign o[5373] = i[20];
  assign o[5374] = i[20];
  assign o[5375] = i[20];
  assign o[4864] = i[19];
  assign o[4865] = i[19];
  assign o[4866] = i[19];
  assign o[4867] = i[19];
  assign o[4868] = i[19];
  assign o[4869] = i[19];
  assign o[4870] = i[19];
  assign o[4871] = i[19];
  assign o[4872] = i[19];
  assign o[4873] = i[19];
  assign o[4874] = i[19];
  assign o[4875] = i[19];
  assign o[4876] = i[19];
  assign o[4877] = i[19];
  assign o[4878] = i[19];
  assign o[4879] = i[19];
  assign o[4880] = i[19];
  assign o[4881] = i[19];
  assign o[4882] = i[19];
  assign o[4883] = i[19];
  assign o[4884] = i[19];
  assign o[4885] = i[19];
  assign o[4886] = i[19];
  assign o[4887] = i[19];
  assign o[4888] = i[19];
  assign o[4889] = i[19];
  assign o[4890] = i[19];
  assign o[4891] = i[19];
  assign o[4892] = i[19];
  assign o[4893] = i[19];
  assign o[4894] = i[19];
  assign o[4895] = i[19];
  assign o[4896] = i[19];
  assign o[4897] = i[19];
  assign o[4898] = i[19];
  assign o[4899] = i[19];
  assign o[4900] = i[19];
  assign o[4901] = i[19];
  assign o[4902] = i[19];
  assign o[4903] = i[19];
  assign o[4904] = i[19];
  assign o[4905] = i[19];
  assign o[4906] = i[19];
  assign o[4907] = i[19];
  assign o[4908] = i[19];
  assign o[4909] = i[19];
  assign o[4910] = i[19];
  assign o[4911] = i[19];
  assign o[4912] = i[19];
  assign o[4913] = i[19];
  assign o[4914] = i[19];
  assign o[4915] = i[19];
  assign o[4916] = i[19];
  assign o[4917] = i[19];
  assign o[4918] = i[19];
  assign o[4919] = i[19];
  assign o[4920] = i[19];
  assign o[4921] = i[19];
  assign o[4922] = i[19];
  assign o[4923] = i[19];
  assign o[4924] = i[19];
  assign o[4925] = i[19];
  assign o[4926] = i[19];
  assign o[4927] = i[19];
  assign o[4928] = i[19];
  assign o[4929] = i[19];
  assign o[4930] = i[19];
  assign o[4931] = i[19];
  assign o[4932] = i[19];
  assign o[4933] = i[19];
  assign o[4934] = i[19];
  assign o[4935] = i[19];
  assign o[4936] = i[19];
  assign o[4937] = i[19];
  assign o[4938] = i[19];
  assign o[4939] = i[19];
  assign o[4940] = i[19];
  assign o[4941] = i[19];
  assign o[4942] = i[19];
  assign o[4943] = i[19];
  assign o[4944] = i[19];
  assign o[4945] = i[19];
  assign o[4946] = i[19];
  assign o[4947] = i[19];
  assign o[4948] = i[19];
  assign o[4949] = i[19];
  assign o[4950] = i[19];
  assign o[4951] = i[19];
  assign o[4952] = i[19];
  assign o[4953] = i[19];
  assign o[4954] = i[19];
  assign o[4955] = i[19];
  assign o[4956] = i[19];
  assign o[4957] = i[19];
  assign o[4958] = i[19];
  assign o[4959] = i[19];
  assign o[4960] = i[19];
  assign o[4961] = i[19];
  assign o[4962] = i[19];
  assign o[4963] = i[19];
  assign o[4964] = i[19];
  assign o[4965] = i[19];
  assign o[4966] = i[19];
  assign o[4967] = i[19];
  assign o[4968] = i[19];
  assign o[4969] = i[19];
  assign o[4970] = i[19];
  assign o[4971] = i[19];
  assign o[4972] = i[19];
  assign o[4973] = i[19];
  assign o[4974] = i[19];
  assign o[4975] = i[19];
  assign o[4976] = i[19];
  assign o[4977] = i[19];
  assign o[4978] = i[19];
  assign o[4979] = i[19];
  assign o[4980] = i[19];
  assign o[4981] = i[19];
  assign o[4982] = i[19];
  assign o[4983] = i[19];
  assign o[4984] = i[19];
  assign o[4985] = i[19];
  assign o[4986] = i[19];
  assign o[4987] = i[19];
  assign o[4988] = i[19];
  assign o[4989] = i[19];
  assign o[4990] = i[19];
  assign o[4991] = i[19];
  assign o[4992] = i[19];
  assign o[4993] = i[19];
  assign o[4994] = i[19];
  assign o[4995] = i[19];
  assign o[4996] = i[19];
  assign o[4997] = i[19];
  assign o[4998] = i[19];
  assign o[4999] = i[19];
  assign o[5000] = i[19];
  assign o[5001] = i[19];
  assign o[5002] = i[19];
  assign o[5003] = i[19];
  assign o[5004] = i[19];
  assign o[5005] = i[19];
  assign o[5006] = i[19];
  assign o[5007] = i[19];
  assign o[5008] = i[19];
  assign o[5009] = i[19];
  assign o[5010] = i[19];
  assign o[5011] = i[19];
  assign o[5012] = i[19];
  assign o[5013] = i[19];
  assign o[5014] = i[19];
  assign o[5015] = i[19];
  assign o[5016] = i[19];
  assign o[5017] = i[19];
  assign o[5018] = i[19];
  assign o[5019] = i[19];
  assign o[5020] = i[19];
  assign o[5021] = i[19];
  assign o[5022] = i[19];
  assign o[5023] = i[19];
  assign o[5024] = i[19];
  assign o[5025] = i[19];
  assign o[5026] = i[19];
  assign o[5027] = i[19];
  assign o[5028] = i[19];
  assign o[5029] = i[19];
  assign o[5030] = i[19];
  assign o[5031] = i[19];
  assign o[5032] = i[19];
  assign o[5033] = i[19];
  assign o[5034] = i[19];
  assign o[5035] = i[19];
  assign o[5036] = i[19];
  assign o[5037] = i[19];
  assign o[5038] = i[19];
  assign o[5039] = i[19];
  assign o[5040] = i[19];
  assign o[5041] = i[19];
  assign o[5042] = i[19];
  assign o[5043] = i[19];
  assign o[5044] = i[19];
  assign o[5045] = i[19];
  assign o[5046] = i[19];
  assign o[5047] = i[19];
  assign o[5048] = i[19];
  assign o[5049] = i[19];
  assign o[5050] = i[19];
  assign o[5051] = i[19];
  assign o[5052] = i[19];
  assign o[5053] = i[19];
  assign o[5054] = i[19];
  assign o[5055] = i[19];
  assign o[5056] = i[19];
  assign o[5057] = i[19];
  assign o[5058] = i[19];
  assign o[5059] = i[19];
  assign o[5060] = i[19];
  assign o[5061] = i[19];
  assign o[5062] = i[19];
  assign o[5063] = i[19];
  assign o[5064] = i[19];
  assign o[5065] = i[19];
  assign o[5066] = i[19];
  assign o[5067] = i[19];
  assign o[5068] = i[19];
  assign o[5069] = i[19];
  assign o[5070] = i[19];
  assign o[5071] = i[19];
  assign o[5072] = i[19];
  assign o[5073] = i[19];
  assign o[5074] = i[19];
  assign o[5075] = i[19];
  assign o[5076] = i[19];
  assign o[5077] = i[19];
  assign o[5078] = i[19];
  assign o[5079] = i[19];
  assign o[5080] = i[19];
  assign o[5081] = i[19];
  assign o[5082] = i[19];
  assign o[5083] = i[19];
  assign o[5084] = i[19];
  assign o[5085] = i[19];
  assign o[5086] = i[19];
  assign o[5087] = i[19];
  assign o[5088] = i[19];
  assign o[5089] = i[19];
  assign o[5090] = i[19];
  assign o[5091] = i[19];
  assign o[5092] = i[19];
  assign o[5093] = i[19];
  assign o[5094] = i[19];
  assign o[5095] = i[19];
  assign o[5096] = i[19];
  assign o[5097] = i[19];
  assign o[5098] = i[19];
  assign o[5099] = i[19];
  assign o[5100] = i[19];
  assign o[5101] = i[19];
  assign o[5102] = i[19];
  assign o[5103] = i[19];
  assign o[5104] = i[19];
  assign o[5105] = i[19];
  assign o[5106] = i[19];
  assign o[5107] = i[19];
  assign o[5108] = i[19];
  assign o[5109] = i[19];
  assign o[5110] = i[19];
  assign o[5111] = i[19];
  assign o[5112] = i[19];
  assign o[5113] = i[19];
  assign o[5114] = i[19];
  assign o[5115] = i[19];
  assign o[5116] = i[19];
  assign o[5117] = i[19];
  assign o[5118] = i[19];
  assign o[5119] = i[19];
  assign o[4608] = i[18];
  assign o[4609] = i[18];
  assign o[4610] = i[18];
  assign o[4611] = i[18];
  assign o[4612] = i[18];
  assign o[4613] = i[18];
  assign o[4614] = i[18];
  assign o[4615] = i[18];
  assign o[4616] = i[18];
  assign o[4617] = i[18];
  assign o[4618] = i[18];
  assign o[4619] = i[18];
  assign o[4620] = i[18];
  assign o[4621] = i[18];
  assign o[4622] = i[18];
  assign o[4623] = i[18];
  assign o[4624] = i[18];
  assign o[4625] = i[18];
  assign o[4626] = i[18];
  assign o[4627] = i[18];
  assign o[4628] = i[18];
  assign o[4629] = i[18];
  assign o[4630] = i[18];
  assign o[4631] = i[18];
  assign o[4632] = i[18];
  assign o[4633] = i[18];
  assign o[4634] = i[18];
  assign o[4635] = i[18];
  assign o[4636] = i[18];
  assign o[4637] = i[18];
  assign o[4638] = i[18];
  assign o[4639] = i[18];
  assign o[4640] = i[18];
  assign o[4641] = i[18];
  assign o[4642] = i[18];
  assign o[4643] = i[18];
  assign o[4644] = i[18];
  assign o[4645] = i[18];
  assign o[4646] = i[18];
  assign o[4647] = i[18];
  assign o[4648] = i[18];
  assign o[4649] = i[18];
  assign o[4650] = i[18];
  assign o[4651] = i[18];
  assign o[4652] = i[18];
  assign o[4653] = i[18];
  assign o[4654] = i[18];
  assign o[4655] = i[18];
  assign o[4656] = i[18];
  assign o[4657] = i[18];
  assign o[4658] = i[18];
  assign o[4659] = i[18];
  assign o[4660] = i[18];
  assign o[4661] = i[18];
  assign o[4662] = i[18];
  assign o[4663] = i[18];
  assign o[4664] = i[18];
  assign o[4665] = i[18];
  assign o[4666] = i[18];
  assign o[4667] = i[18];
  assign o[4668] = i[18];
  assign o[4669] = i[18];
  assign o[4670] = i[18];
  assign o[4671] = i[18];
  assign o[4672] = i[18];
  assign o[4673] = i[18];
  assign o[4674] = i[18];
  assign o[4675] = i[18];
  assign o[4676] = i[18];
  assign o[4677] = i[18];
  assign o[4678] = i[18];
  assign o[4679] = i[18];
  assign o[4680] = i[18];
  assign o[4681] = i[18];
  assign o[4682] = i[18];
  assign o[4683] = i[18];
  assign o[4684] = i[18];
  assign o[4685] = i[18];
  assign o[4686] = i[18];
  assign o[4687] = i[18];
  assign o[4688] = i[18];
  assign o[4689] = i[18];
  assign o[4690] = i[18];
  assign o[4691] = i[18];
  assign o[4692] = i[18];
  assign o[4693] = i[18];
  assign o[4694] = i[18];
  assign o[4695] = i[18];
  assign o[4696] = i[18];
  assign o[4697] = i[18];
  assign o[4698] = i[18];
  assign o[4699] = i[18];
  assign o[4700] = i[18];
  assign o[4701] = i[18];
  assign o[4702] = i[18];
  assign o[4703] = i[18];
  assign o[4704] = i[18];
  assign o[4705] = i[18];
  assign o[4706] = i[18];
  assign o[4707] = i[18];
  assign o[4708] = i[18];
  assign o[4709] = i[18];
  assign o[4710] = i[18];
  assign o[4711] = i[18];
  assign o[4712] = i[18];
  assign o[4713] = i[18];
  assign o[4714] = i[18];
  assign o[4715] = i[18];
  assign o[4716] = i[18];
  assign o[4717] = i[18];
  assign o[4718] = i[18];
  assign o[4719] = i[18];
  assign o[4720] = i[18];
  assign o[4721] = i[18];
  assign o[4722] = i[18];
  assign o[4723] = i[18];
  assign o[4724] = i[18];
  assign o[4725] = i[18];
  assign o[4726] = i[18];
  assign o[4727] = i[18];
  assign o[4728] = i[18];
  assign o[4729] = i[18];
  assign o[4730] = i[18];
  assign o[4731] = i[18];
  assign o[4732] = i[18];
  assign o[4733] = i[18];
  assign o[4734] = i[18];
  assign o[4735] = i[18];
  assign o[4736] = i[18];
  assign o[4737] = i[18];
  assign o[4738] = i[18];
  assign o[4739] = i[18];
  assign o[4740] = i[18];
  assign o[4741] = i[18];
  assign o[4742] = i[18];
  assign o[4743] = i[18];
  assign o[4744] = i[18];
  assign o[4745] = i[18];
  assign o[4746] = i[18];
  assign o[4747] = i[18];
  assign o[4748] = i[18];
  assign o[4749] = i[18];
  assign o[4750] = i[18];
  assign o[4751] = i[18];
  assign o[4752] = i[18];
  assign o[4753] = i[18];
  assign o[4754] = i[18];
  assign o[4755] = i[18];
  assign o[4756] = i[18];
  assign o[4757] = i[18];
  assign o[4758] = i[18];
  assign o[4759] = i[18];
  assign o[4760] = i[18];
  assign o[4761] = i[18];
  assign o[4762] = i[18];
  assign o[4763] = i[18];
  assign o[4764] = i[18];
  assign o[4765] = i[18];
  assign o[4766] = i[18];
  assign o[4767] = i[18];
  assign o[4768] = i[18];
  assign o[4769] = i[18];
  assign o[4770] = i[18];
  assign o[4771] = i[18];
  assign o[4772] = i[18];
  assign o[4773] = i[18];
  assign o[4774] = i[18];
  assign o[4775] = i[18];
  assign o[4776] = i[18];
  assign o[4777] = i[18];
  assign o[4778] = i[18];
  assign o[4779] = i[18];
  assign o[4780] = i[18];
  assign o[4781] = i[18];
  assign o[4782] = i[18];
  assign o[4783] = i[18];
  assign o[4784] = i[18];
  assign o[4785] = i[18];
  assign o[4786] = i[18];
  assign o[4787] = i[18];
  assign o[4788] = i[18];
  assign o[4789] = i[18];
  assign o[4790] = i[18];
  assign o[4791] = i[18];
  assign o[4792] = i[18];
  assign o[4793] = i[18];
  assign o[4794] = i[18];
  assign o[4795] = i[18];
  assign o[4796] = i[18];
  assign o[4797] = i[18];
  assign o[4798] = i[18];
  assign o[4799] = i[18];
  assign o[4800] = i[18];
  assign o[4801] = i[18];
  assign o[4802] = i[18];
  assign o[4803] = i[18];
  assign o[4804] = i[18];
  assign o[4805] = i[18];
  assign o[4806] = i[18];
  assign o[4807] = i[18];
  assign o[4808] = i[18];
  assign o[4809] = i[18];
  assign o[4810] = i[18];
  assign o[4811] = i[18];
  assign o[4812] = i[18];
  assign o[4813] = i[18];
  assign o[4814] = i[18];
  assign o[4815] = i[18];
  assign o[4816] = i[18];
  assign o[4817] = i[18];
  assign o[4818] = i[18];
  assign o[4819] = i[18];
  assign o[4820] = i[18];
  assign o[4821] = i[18];
  assign o[4822] = i[18];
  assign o[4823] = i[18];
  assign o[4824] = i[18];
  assign o[4825] = i[18];
  assign o[4826] = i[18];
  assign o[4827] = i[18];
  assign o[4828] = i[18];
  assign o[4829] = i[18];
  assign o[4830] = i[18];
  assign o[4831] = i[18];
  assign o[4832] = i[18];
  assign o[4833] = i[18];
  assign o[4834] = i[18];
  assign o[4835] = i[18];
  assign o[4836] = i[18];
  assign o[4837] = i[18];
  assign o[4838] = i[18];
  assign o[4839] = i[18];
  assign o[4840] = i[18];
  assign o[4841] = i[18];
  assign o[4842] = i[18];
  assign o[4843] = i[18];
  assign o[4844] = i[18];
  assign o[4845] = i[18];
  assign o[4846] = i[18];
  assign o[4847] = i[18];
  assign o[4848] = i[18];
  assign o[4849] = i[18];
  assign o[4850] = i[18];
  assign o[4851] = i[18];
  assign o[4852] = i[18];
  assign o[4853] = i[18];
  assign o[4854] = i[18];
  assign o[4855] = i[18];
  assign o[4856] = i[18];
  assign o[4857] = i[18];
  assign o[4858] = i[18];
  assign o[4859] = i[18];
  assign o[4860] = i[18];
  assign o[4861] = i[18];
  assign o[4862] = i[18];
  assign o[4863] = i[18];
  assign o[4352] = i[17];
  assign o[4353] = i[17];
  assign o[4354] = i[17];
  assign o[4355] = i[17];
  assign o[4356] = i[17];
  assign o[4357] = i[17];
  assign o[4358] = i[17];
  assign o[4359] = i[17];
  assign o[4360] = i[17];
  assign o[4361] = i[17];
  assign o[4362] = i[17];
  assign o[4363] = i[17];
  assign o[4364] = i[17];
  assign o[4365] = i[17];
  assign o[4366] = i[17];
  assign o[4367] = i[17];
  assign o[4368] = i[17];
  assign o[4369] = i[17];
  assign o[4370] = i[17];
  assign o[4371] = i[17];
  assign o[4372] = i[17];
  assign o[4373] = i[17];
  assign o[4374] = i[17];
  assign o[4375] = i[17];
  assign o[4376] = i[17];
  assign o[4377] = i[17];
  assign o[4378] = i[17];
  assign o[4379] = i[17];
  assign o[4380] = i[17];
  assign o[4381] = i[17];
  assign o[4382] = i[17];
  assign o[4383] = i[17];
  assign o[4384] = i[17];
  assign o[4385] = i[17];
  assign o[4386] = i[17];
  assign o[4387] = i[17];
  assign o[4388] = i[17];
  assign o[4389] = i[17];
  assign o[4390] = i[17];
  assign o[4391] = i[17];
  assign o[4392] = i[17];
  assign o[4393] = i[17];
  assign o[4394] = i[17];
  assign o[4395] = i[17];
  assign o[4396] = i[17];
  assign o[4397] = i[17];
  assign o[4398] = i[17];
  assign o[4399] = i[17];
  assign o[4400] = i[17];
  assign o[4401] = i[17];
  assign o[4402] = i[17];
  assign o[4403] = i[17];
  assign o[4404] = i[17];
  assign o[4405] = i[17];
  assign o[4406] = i[17];
  assign o[4407] = i[17];
  assign o[4408] = i[17];
  assign o[4409] = i[17];
  assign o[4410] = i[17];
  assign o[4411] = i[17];
  assign o[4412] = i[17];
  assign o[4413] = i[17];
  assign o[4414] = i[17];
  assign o[4415] = i[17];
  assign o[4416] = i[17];
  assign o[4417] = i[17];
  assign o[4418] = i[17];
  assign o[4419] = i[17];
  assign o[4420] = i[17];
  assign o[4421] = i[17];
  assign o[4422] = i[17];
  assign o[4423] = i[17];
  assign o[4424] = i[17];
  assign o[4425] = i[17];
  assign o[4426] = i[17];
  assign o[4427] = i[17];
  assign o[4428] = i[17];
  assign o[4429] = i[17];
  assign o[4430] = i[17];
  assign o[4431] = i[17];
  assign o[4432] = i[17];
  assign o[4433] = i[17];
  assign o[4434] = i[17];
  assign o[4435] = i[17];
  assign o[4436] = i[17];
  assign o[4437] = i[17];
  assign o[4438] = i[17];
  assign o[4439] = i[17];
  assign o[4440] = i[17];
  assign o[4441] = i[17];
  assign o[4442] = i[17];
  assign o[4443] = i[17];
  assign o[4444] = i[17];
  assign o[4445] = i[17];
  assign o[4446] = i[17];
  assign o[4447] = i[17];
  assign o[4448] = i[17];
  assign o[4449] = i[17];
  assign o[4450] = i[17];
  assign o[4451] = i[17];
  assign o[4452] = i[17];
  assign o[4453] = i[17];
  assign o[4454] = i[17];
  assign o[4455] = i[17];
  assign o[4456] = i[17];
  assign o[4457] = i[17];
  assign o[4458] = i[17];
  assign o[4459] = i[17];
  assign o[4460] = i[17];
  assign o[4461] = i[17];
  assign o[4462] = i[17];
  assign o[4463] = i[17];
  assign o[4464] = i[17];
  assign o[4465] = i[17];
  assign o[4466] = i[17];
  assign o[4467] = i[17];
  assign o[4468] = i[17];
  assign o[4469] = i[17];
  assign o[4470] = i[17];
  assign o[4471] = i[17];
  assign o[4472] = i[17];
  assign o[4473] = i[17];
  assign o[4474] = i[17];
  assign o[4475] = i[17];
  assign o[4476] = i[17];
  assign o[4477] = i[17];
  assign o[4478] = i[17];
  assign o[4479] = i[17];
  assign o[4480] = i[17];
  assign o[4481] = i[17];
  assign o[4482] = i[17];
  assign o[4483] = i[17];
  assign o[4484] = i[17];
  assign o[4485] = i[17];
  assign o[4486] = i[17];
  assign o[4487] = i[17];
  assign o[4488] = i[17];
  assign o[4489] = i[17];
  assign o[4490] = i[17];
  assign o[4491] = i[17];
  assign o[4492] = i[17];
  assign o[4493] = i[17];
  assign o[4494] = i[17];
  assign o[4495] = i[17];
  assign o[4496] = i[17];
  assign o[4497] = i[17];
  assign o[4498] = i[17];
  assign o[4499] = i[17];
  assign o[4500] = i[17];
  assign o[4501] = i[17];
  assign o[4502] = i[17];
  assign o[4503] = i[17];
  assign o[4504] = i[17];
  assign o[4505] = i[17];
  assign o[4506] = i[17];
  assign o[4507] = i[17];
  assign o[4508] = i[17];
  assign o[4509] = i[17];
  assign o[4510] = i[17];
  assign o[4511] = i[17];
  assign o[4512] = i[17];
  assign o[4513] = i[17];
  assign o[4514] = i[17];
  assign o[4515] = i[17];
  assign o[4516] = i[17];
  assign o[4517] = i[17];
  assign o[4518] = i[17];
  assign o[4519] = i[17];
  assign o[4520] = i[17];
  assign o[4521] = i[17];
  assign o[4522] = i[17];
  assign o[4523] = i[17];
  assign o[4524] = i[17];
  assign o[4525] = i[17];
  assign o[4526] = i[17];
  assign o[4527] = i[17];
  assign o[4528] = i[17];
  assign o[4529] = i[17];
  assign o[4530] = i[17];
  assign o[4531] = i[17];
  assign o[4532] = i[17];
  assign o[4533] = i[17];
  assign o[4534] = i[17];
  assign o[4535] = i[17];
  assign o[4536] = i[17];
  assign o[4537] = i[17];
  assign o[4538] = i[17];
  assign o[4539] = i[17];
  assign o[4540] = i[17];
  assign o[4541] = i[17];
  assign o[4542] = i[17];
  assign o[4543] = i[17];
  assign o[4544] = i[17];
  assign o[4545] = i[17];
  assign o[4546] = i[17];
  assign o[4547] = i[17];
  assign o[4548] = i[17];
  assign o[4549] = i[17];
  assign o[4550] = i[17];
  assign o[4551] = i[17];
  assign o[4552] = i[17];
  assign o[4553] = i[17];
  assign o[4554] = i[17];
  assign o[4555] = i[17];
  assign o[4556] = i[17];
  assign o[4557] = i[17];
  assign o[4558] = i[17];
  assign o[4559] = i[17];
  assign o[4560] = i[17];
  assign o[4561] = i[17];
  assign o[4562] = i[17];
  assign o[4563] = i[17];
  assign o[4564] = i[17];
  assign o[4565] = i[17];
  assign o[4566] = i[17];
  assign o[4567] = i[17];
  assign o[4568] = i[17];
  assign o[4569] = i[17];
  assign o[4570] = i[17];
  assign o[4571] = i[17];
  assign o[4572] = i[17];
  assign o[4573] = i[17];
  assign o[4574] = i[17];
  assign o[4575] = i[17];
  assign o[4576] = i[17];
  assign o[4577] = i[17];
  assign o[4578] = i[17];
  assign o[4579] = i[17];
  assign o[4580] = i[17];
  assign o[4581] = i[17];
  assign o[4582] = i[17];
  assign o[4583] = i[17];
  assign o[4584] = i[17];
  assign o[4585] = i[17];
  assign o[4586] = i[17];
  assign o[4587] = i[17];
  assign o[4588] = i[17];
  assign o[4589] = i[17];
  assign o[4590] = i[17];
  assign o[4591] = i[17];
  assign o[4592] = i[17];
  assign o[4593] = i[17];
  assign o[4594] = i[17];
  assign o[4595] = i[17];
  assign o[4596] = i[17];
  assign o[4597] = i[17];
  assign o[4598] = i[17];
  assign o[4599] = i[17];
  assign o[4600] = i[17];
  assign o[4601] = i[17];
  assign o[4602] = i[17];
  assign o[4603] = i[17];
  assign o[4604] = i[17];
  assign o[4605] = i[17];
  assign o[4606] = i[17];
  assign o[4607] = i[17];
  assign o[4096] = i[16];
  assign o[4097] = i[16];
  assign o[4098] = i[16];
  assign o[4099] = i[16];
  assign o[4100] = i[16];
  assign o[4101] = i[16];
  assign o[4102] = i[16];
  assign o[4103] = i[16];
  assign o[4104] = i[16];
  assign o[4105] = i[16];
  assign o[4106] = i[16];
  assign o[4107] = i[16];
  assign o[4108] = i[16];
  assign o[4109] = i[16];
  assign o[4110] = i[16];
  assign o[4111] = i[16];
  assign o[4112] = i[16];
  assign o[4113] = i[16];
  assign o[4114] = i[16];
  assign o[4115] = i[16];
  assign o[4116] = i[16];
  assign o[4117] = i[16];
  assign o[4118] = i[16];
  assign o[4119] = i[16];
  assign o[4120] = i[16];
  assign o[4121] = i[16];
  assign o[4122] = i[16];
  assign o[4123] = i[16];
  assign o[4124] = i[16];
  assign o[4125] = i[16];
  assign o[4126] = i[16];
  assign o[4127] = i[16];
  assign o[4128] = i[16];
  assign o[4129] = i[16];
  assign o[4130] = i[16];
  assign o[4131] = i[16];
  assign o[4132] = i[16];
  assign o[4133] = i[16];
  assign o[4134] = i[16];
  assign o[4135] = i[16];
  assign o[4136] = i[16];
  assign o[4137] = i[16];
  assign o[4138] = i[16];
  assign o[4139] = i[16];
  assign o[4140] = i[16];
  assign o[4141] = i[16];
  assign o[4142] = i[16];
  assign o[4143] = i[16];
  assign o[4144] = i[16];
  assign o[4145] = i[16];
  assign o[4146] = i[16];
  assign o[4147] = i[16];
  assign o[4148] = i[16];
  assign o[4149] = i[16];
  assign o[4150] = i[16];
  assign o[4151] = i[16];
  assign o[4152] = i[16];
  assign o[4153] = i[16];
  assign o[4154] = i[16];
  assign o[4155] = i[16];
  assign o[4156] = i[16];
  assign o[4157] = i[16];
  assign o[4158] = i[16];
  assign o[4159] = i[16];
  assign o[4160] = i[16];
  assign o[4161] = i[16];
  assign o[4162] = i[16];
  assign o[4163] = i[16];
  assign o[4164] = i[16];
  assign o[4165] = i[16];
  assign o[4166] = i[16];
  assign o[4167] = i[16];
  assign o[4168] = i[16];
  assign o[4169] = i[16];
  assign o[4170] = i[16];
  assign o[4171] = i[16];
  assign o[4172] = i[16];
  assign o[4173] = i[16];
  assign o[4174] = i[16];
  assign o[4175] = i[16];
  assign o[4176] = i[16];
  assign o[4177] = i[16];
  assign o[4178] = i[16];
  assign o[4179] = i[16];
  assign o[4180] = i[16];
  assign o[4181] = i[16];
  assign o[4182] = i[16];
  assign o[4183] = i[16];
  assign o[4184] = i[16];
  assign o[4185] = i[16];
  assign o[4186] = i[16];
  assign o[4187] = i[16];
  assign o[4188] = i[16];
  assign o[4189] = i[16];
  assign o[4190] = i[16];
  assign o[4191] = i[16];
  assign o[4192] = i[16];
  assign o[4193] = i[16];
  assign o[4194] = i[16];
  assign o[4195] = i[16];
  assign o[4196] = i[16];
  assign o[4197] = i[16];
  assign o[4198] = i[16];
  assign o[4199] = i[16];
  assign o[4200] = i[16];
  assign o[4201] = i[16];
  assign o[4202] = i[16];
  assign o[4203] = i[16];
  assign o[4204] = i[16];
  assign o[4205] = i[16];
  assign o[4206] = i[16];
  assign o[4207] = i[16];
  assign o[4208] = i[16];
  assign o[4209] = i[16];
  assign o[4210] = i[16];
  assign o[4211] = i[16];
  assign o[4212] = i[16];
  assign o[4213] = i[16];
  assign o[4214] = i[16];
  assign o[4215] = i[16];
  assign o[4216] = i[16];
  assign o[4217] = i[16];
  assign o[4218] = i[16];
  assign o[4219] = i[16];
  assign o[4220] = i[16];
  assign o[4221] = i[16];
  assign o[4222] = i[16];
  assign o[4223] = i[16];
  assign o[4224] = i[16];
  assign o[4225] = i[16];
  assign o[4226] = i[16];
  assign o[4227] = i[16];
  assign o[4228] = i[16];
  assign o[4229] = i[16];
  assign o[4230] = i[16];
  assign o[4231] = i[16];
  assign o[4232] = i[16];
  assign o[4233] = i[16];
  assign o[4234] = i[16];
  assign o[4235] = i[16];
  assign o[4236] = i[16];
  assign o[4237] = i[16];
  assign o[4238] = i[16];
  assign o[4239] = i[16];
  assign o[4240] = i[16];
  assign o[4241] = i[16];
  assign o[4242] = i[16];
  assign o[4243] = i[16];
  assign o[4244] = i[16];
  assign o[4245] = i[16];
  assign o[4246] = i[16];
  assign o[4247] = i[16];
  assign o[4248] = i[16];
  assign o[4249] = i[16];
  assign o[4250] = i[16];
  assign o[4251] = i[16];
  assign o[4252] = i[16];
  assign o[4253] = i[16];
  assign o[4254] = i[16];
  assign o[4255] = i[16];
  assign o[4256] = i[16];
  assign o[4257] = i[16];
  assign o[4258] = i[16];
  assign o[4259] = i[16];
  assign o[4260] = i[16];
  assign o[4261] = i[16];
  assign o[4262] = i[16];
  assign o[4263] = i[16];
  assign o[4264] = i[16];
  assign o[4265] = i[16];
  assign o[4266] = i[16];
  assign o[4267] = i[16];
  assign o[4268] = i[16];
  assign o[4269] = i[16];
  assign o[4270] = i[16];
  assign o[4271] = i[16];
  assign o[4272] = i[16];
  assign o[4273] = i[16];
  assign o[4274] = i[16];
  assign o[4275] = i[16];
  assign o[4276] = i[16];
  assign o[4277] = i[16];
  assign o[4278] = i[16];
  assign o[4279] = i[16];
  assign o[4280] = i[16];
  assign o[4281] = i[16];
  assign o[4282] = i[16];
  assign o[4283] = i[16];
  assign o[4284] = i[16];
  assign o[4285] = i[16];
  assign o[4286] = i[16];
  assign o[4287] = i[16];
  assign o[4288] = i[16];
  assign o[4289] = i[16];
  assign o[4290] = i[16];
  assign o[4291] = i[16];
  assign o[4292] = i[16];
  assign o[4293] = i[16];
  assign o[4294] = i[16];
  assign o[4295] = i[16];
  assign o[4296] = i[16];
  assign o[4297] = i[16];
  assign o[4298] = i[16];
  assign o[4299] = i[16];
  assign o[4300] = i[16];
  assign o[4301] = i[16];
  assign o[4302] = i[16];
  assign o[4303] = i[16];
  assign o[4304] = i[16];
  assign o[4305] = i[16];
  assign o[4306] = i[16];
  assign o[4307] = i[16];
  assign o[4308] = i[16];
  assign o[4309] = i[16];
  assign o[4310] = i[16];
  assign o[4311] = i[16];
  assign o[4312] = i[16];
  assign o[4313] = i[16];
  assign o[4314] = i[16];
  assign o[4315] = i[16];
  assign o[4316] = i[16];
  assign o[4317] = i[16];
  assign o[4318] = i[16];
  assign o[4319] = i[16];
  assign o[4320] = i[16];
  assign o[4321] = i[16];
  assign o[4322] = i[16];
  assign o[4323] = i[16];
  assign o[4324] = i[16];
  assign o[4325] = i[16];
  assign o[4326] = i[16];
  assign o[4327] = i[16];
  assign o[4328] = i[16];
  assign o[4329] = i[16];
  assign o[4330] = i[16];
  assign o[4331] = i[16];
  assign o[4332] = i[16];
  assign o[4333] = i[16];
  assign o[4334] = i[16];
  assign o[4335] = i[16];
  assign o[4336] = i[16];
  assign o[4337] = i[16];
  assign o[4338] = i[16];
  assign o[4339] = i[16];
  assign o[4340] = i[16];
  assign o[4341] = i[16];
  assign o[4342] = i[16];
  assign o[4343] = i[16];
  assign o[4344] = i[16];
  assign o[4345] = i[16];
  assign o[4346] = i[16];
  assign o[4347] = i[16];
  assign o[4348] = i[16];
  assign o[4349] = i[16];
  assign o[4350] = i[16];
  assign o[4351] = i[16];
  assign o[3840] = i[15];
  assign o[3841] = i[15];
  assign o[3842] = i[15];
  assign o[3843] = i[15];
  assign o[3844] = i[15];
  assign o[3845] = i[15];
  assign o[3846] = i[15];
  assign o[3847] = i[15];
  assign o[3848] = i[15];
  assign o[3849] = i[15];
  assign o[3850] = i[15];
  assign o[3851] = i[15];
  assign o[3852] = i[15];
  assign o[3853] = i[15];
  assign o[3854] = i[15];
  assign o[3855] = i[15];
  assign o[3856] = i[15];
  assign o[3857] = i[15];
  assign o[3858] = i[15];
  assign o[3859] = i[15];
  assign o[3860] = i[15];
  assign o[3861] = i[15];
  assign o[3862] = i[15];
  assign o[3863] = i[15];
  assign o[3864] = i[15];
  assign o[3865] = i[15];
  assign o[3866] = i[15];
  assign o[3867] = i[15];
  assign o[3868] = i[15];
  assign o[3869] = i[15];
  assign o[3870] = i[15];
  assign o[3871] = i[15];
  assign o[3872] = i[15];
  assign o[3873] = i[15];
  assign o[3874] = i[15];
  assign o[3875] = i[15];
  assign o[3876] = i[15];
  assign o[3877] = i[15];
  assign o[3878] = i[15];
  assign o[3879] = i[15];
  assign o[3880] = i[15];
  assign o[3881] = i[15];
  assign o[3882] = i[15];
  assign o[3883] = i[15];
  assign o[3884] = i[15];
  assign o[3885] = i[15];
  assign o[3886] = i[15];
  assign o[3887] = i[15];
  assign o[3888] = i[15];
  assign o[3889] = i[15];
  assign o[3890] = i[15];
  assign o[3891] = i[15];
  assign o[3892] = i[15];
  assign o[3893] = i[15];
  assign o[3894] = i[15];
  assign o[3895] = i[15];
  assign o[3896] = i[15];
  assign o[3897] = i[15];
  assign o[3898] = i[15];
  assign o[3899] = i[15];
  assign o[3900] = i[15];
  assign o[3901] = i[15];
  assign o[3902] = i[15];
  assign o[3903] = i[15];
  assign o[3904] = i[15];
  assign o[3905] = i[15];
  assign o[3906] = i[15];
  assign o[3907] = i[15];
  assign o[3908] = i[15];
  assign o[3909] = i[15];
  assign o[3910] = i[15];
  assign o[3911] = i[15];
  assign o[3912] = i[15];
  assign o[3913] = i[15];
  assign o[3914] = i[15];
  assign o[3915] = i[15];
  assign o[3916] = i[15];
  assign o[3917] = i[15];
  assign o[3918] = i[15];
  assign o[3919] = i[15];
  assign o[3920] = i[15];
  assign o[3921] = i[15];
  assign o[3922] = i[15];
  assign o[3923] = i[15];
  assign o[3924] = i[15];
  assign o[3925] = i[15];
  assign o[3926] = i[15];
  assign o[3927] = i[15];
  assign o[3928] = i[15];
  assign o[3929] = i[15];
  assign o[3930] = i[15];
  assign o[3931] = i[15];
  assign o[3932] = i[15];
  assign o[3933] = i[15];
  assign o[3934] = i[15];
  assign o[3935] = i[15];
  assign o[3936] = i[15];
  assign o[3937] = i[15];
  assign o[3938] = i[15];
  assign o[3939] = i[15];
  assign o[3940] = i[15];
  assign o[3941] = i[15];
  assign o[3942] = i[15];
  assign o[3943] = i[15];
  assign o[3944] = i[15];
  assign o[3945] = i[15];
  assign o[3946] = i[15];
  assign o[3947] = i[15];
  assign o[3948] = i[15];
  assign o[3949] = i[15];
  assign o[3950] = i[15];
  assign o[3951] = i[15];
  assign o[3952] = i[15];
  assign o[3953] = i[15];
  assign o[3954] = i[15];
  assign o[3955] = i[15];
  assign o[3956] = i[15];
  assign o[3957] = i[15];
  assign o[3958] = i[15];
  assign o[3959] = i[15];
  assign o[3960] = i[15];
  assign o[3961] = i[15];
  assign o[3962] = i[15];
  assign o[3963] = i[15];
  assign o[3964] = i[15];
  assign o[3965] = i[15];
  assign o[3966] = i[15];
  assign o[3967] = i[15];
  assign o[3968] = i[15];
  assign o[3969] = i[15];
  assign o[3970] = i[15];
  assign o[3971] = i[15];
  assign o[3972] = i[15];
  assign o[3973] = i[15];
  assign o[3974] = i[15];
  assign o[3975] = i[15];
  assign o[3976] = i[15];
  assign o[3977] = i[15];
  assign o[3978] = i[15];
  assign o[3979] = i[15];
  assign o[3980] = i[15];
  assign o[3981] = i[15];
  assign o[3982] = i[15];
  assign o[3983] = i[15];
  assign o[3984] = i[15];
  assign o[3985] = i[15];
  assign o[3986] = i[15];
  assign o[3987] = i[15];
  assign o[3988] = i[15];
  assign o[3989] = i[15];
  assign o[3990] = i[15];
  assign o[3991] = i[15];
  assign o[3992] = i[15];
  assign o[3993] = i[15];
  assign o[3994] = i[15];
  assign o[3995] = i[15];
  assign o[3996] = i[15];
  assign o[3997] = i[15];
  assign o[3998] = i[15];
  assign o[3999] = i[15];
  assign o[4000] = i[15];
  assign o[4001] = i[15];
  assign o[4002] = i[15];
  assign o[4003] = i[15];
  assign o[4004] = i[15];
  assign o[4005] = i[15];
  assign o[4006] = i[15];
  assign o[4007] = i[15];
  assign o[4008] = i[15];
  assign o[4009] = i[15];
  assign o[4010] = i[15];
  assign o[4011] = i[15];
  assign o[4012] = i[15];
  assign o[4013] = i[15];
  assign o[4014] = i[15];
  assign o[4015] = i[15];
  assign o[4016] = i[15];
  assign o[4017] = i[15];
  assign o[4018] = i[15];
  assign o[4019] = i[15];
  assign o[4020] = i[15];
  assign o[4021] = i[15];
  assign o[4022] = i[15];
  assign o[4023] = i[15];
  assign o[4024] = i[15];
  assign o[4025] = i[15];
  assign o[4026] = i[15];
  assign o[4027] = i[15];
  assign o[4028] = i[15];
  assign o[4029] = i[15];
  assign o[4030] = i[15];
  assign o[4031] = i[15];
  assign o[4032] = i[15];
  assign o[4033] = i[15];
  assign o[4034] = i[15];
  assign o[4035] = i[15];
  assign o[4036] = i[15];
  assign o[4037] = i[15];
  assign o[4038] = i[15];
  assign o[4039] = i[15];
  assign o[4040] = i[15];
  assign o[4041] = i[15];
  assign o[4042] = i[15];
  assign o[4043] = i[15];
  assign o[4044] = i[15];
  assign o[4045] = i[15];
  assign o[4046] = i[15];
  assign o[4047] = i[15];
  assign o[4048] = i[15];
  assign o[4049] = i[15];
  assign o[4050] = i[15];
  assign o[4051] = i[15];
  assign o[4052] = i[15];
  assign o[4053] = i[15];
  assign o[4054] = i[15];
  assign o[4055] = i[15];
  assign o[4056] = i[15];
  assign o[4057] = i[15];
  assign o[4058] = i[15];
  assign o[4059] = i[15];
  assign o[4060] = i[15];
  assign o[4061] = i[15];
  assign o[4062] = i[15];
  assign o[4063] = i[15];
  assign o[4064] = i[15];
  assign o[4065] = i[15];
  assign o[4066] = i[15];
  assign o[4067] = i[15];
  assign o[4068] = i[15];
  assign o[4069] = i[15];
  assign o[4070] = i[15];
  assign o[4071] = i[15];
  assign o[4072] = i[15];
  assign o[4073] = i[15];
  assign o[4074] = i[15];
  assign o[4075] = i[15];
  assign o[4076] = i[15];
  assign o[4077] = i[15];
  assign o[4078] = i[15];
  assign o[4079] = i[15];
  assign o[4080] = i[15];
  assign o[4081] = i[15];
  assign o[4082] = i[15];
  assign o[4083] = i[15];
  assign o[4084] = i[15];
  assign o[4085] = i[15];
  assign o[4086] = i[15];
  assign o[4087] = i[15];
  assign o[4088] = i[15];
  assign o[4089] = i[15];
  assign o[4090] = i[15];
  assign o[4091] = i[15];
  assign o[4092] = i[15];
  assign o[4093] = i[15];
  assign o[4094] = i[15];
  assign o[4095] = i[15];
  assign o[3584] = i[14];
  assign o[3585] = i[14];
  assign o[3586] = i[14];
  assign o[3587] = i[14];
  assign o[3588] = i[14];
  assign o[3589] = i[14];
  assign o[3590] = i[14];
  assign o[3591] = i[14];
  assign o[3592] = i[14];
  assign o[3593] = i[14];
  assign o[3594] = i[14];
  assign o[3595] = i[14];
  assign o[3596] = i[14];
  assign o[3597] = i[14];
  assign o[3598] = i[14];
  assign o[3599] = i[14];
  assign o[3600] = i[14];
  assign o[3601] = i[14];
  assign o[3602] = i[14];
  assign o[3603] = i[14];
  assign o[3604] = i[14];
  assign o[3605] = i[14];
  assign o[3606] = i[14];
  assign o[3607] = i[14];
  assign o[3608] = i[14];
  assign o[3609] = i[14];
  assign o[3610] = i[14];
  assign o[3611] = i[14];
  assign o[3612] = i[14];
  assign o[3613] = i[14];
  assign o[3614] = i[14];
  assign o[3615] = i[14];
  assign o[3616] = i[14];
  assign o[3617] = i[14];
  assign o[3618] = i[14];
  assign o[3619] = i[14];
  assign o[3620] = i[14];
  assign o[3621] = i[14];
  assign o[3622] = i[14];
  assign o[3623] = i[14];
  assign o[3624] = i[14];
  assign o[3625] = i[14];
  assign o[3626] = i[14];
  assign o[3627] = i[14];
  assign o[3628] = i[14];
  assign o[3629] = i[14];
  assign o[3630] = i[14];
  assign o[3631] = i[14];
  assign o[3632] = i[14];
  assign o[3633] = i[14];
  assign o[3634] = i[14];
  assign o[3635] = i[14];
  assign o[3636] = i[14];
  assign o[3637] = i[14];
  assign o[3638] = i[14];
  assign o[3639] = i[14];
  assign o[3640] = i[14];
  assign o[3641] = i[14];
  assign o[3642] = i[14];
  assign o[3643] = i[14];
  assign o[3644] = i[14];
  assign o[3645] = i[14];
  assign o[3646] = i[14];
  assign o[3647] = i[14];
  assign o[3648] = i[14];
  assign o[3649] = i[14];
  assign o[3650] = i[14];
  assign o[3651] = i[14];
  assign o[3652] = i[14];
  assign o[3653] = i[14];
  assign o[3654] = i[14];
  assign o[3655] = i[14];
  assign o[3656] = i[14];
  assign o[3657] = i[14];
  assign o[3658] = i[14];
  assign o[3659] = i[14];
  assign o[3660] = i[14];
  assign o[3661] = i[14];
  assign o[3662] = i[14];
  assign o[3663] = i[14];
  assign o[3664] = i[14];
  assign o[3665] = i[14];
  assign o[3666] = i[14];
  assign o[3667] = i[14];
  assign o[3668] = i[14];
  assign o[3669] = i[14];
  assign o[3670] = i[14];
  assign o[3671] = i[14];
  assign o[3672] = i[14];
  assign o[3673] = i[14];
  assign o[3674] = i[14];
  assign o[3675] = i[14];
  assign o[3676] = i[14];
  assign o[3677] = i[14];
  assign o[3678] = i[14];
  assign o[3679] = i[14];
  assign o[3680] = i[14];
  assign o[3681] = i[14];
  assign o[3682] = i[14];
  assign o[3683] = i[14];
  assign o[3684] = i[14];
  assign o[3685] = i[14];
  assign o[3686] = i[14];
  assign o[3687] = i[14];
  assign o[3688] = i[14];
  assign o[3689] = i[14];
  assign o[3690] = i[14];
  assign o[3691] = i[14];
  assign o[3692] = i[14];
  assign o[3693] = i[14];
  assign o[3694] = i[14];
  assign o[3695] = i[14];
  assign o[3696] = i[14];
  assign o[3697] = i[14];
  assign o[3698] = i[14];
  assign o[3699] = i[14];
  assign o[3700] = i[14];
  assign o[3701] = i[14];
  assign o[3702] = i[14];
  assign o[3703] = i[14];
  assign o[3704] = i[14];
  assign o[3705] = i[14];
  assign o[3706] = i[14];
  assign o[3707] = i[14];
  assign o[3708] = i[14];
  assign o[3709] = i[14];
  assign o[3710] = i[14];
  assign o[3711] = i[14];
  assign o[3712] = i[14];
  assign o[3713] = i[14];
  assign o[3714] = i[14];
  assign o[3715] = i[14];
  assign o[3716] = i[14];
  assign o[3717] = i[14];
  assign o[3718] = i[14];
  assign o[3719] = i[14];
  assign o[3720] = i[14];
  assign o[3721] = i[14];
  assign o[3722] = i[14];
  assign o[3723] = i[14];
  assign o[3724] = i[14];
  assign o[3725] = i[14];
  assign o[3726] = i[14];
  assign o[3727] = i[14];
  assign o[3728] = i[14];
  assign o[3729] = i[14];
  assign o[3730] = i[14];
  assign o[3731] = i[14];
  assign o[3732] = i[14];
  assign o[3733] = i[14];
  assign o[3734] = i[14];
  assign o[3735] = i[14];
  assign o[3736] = i[14];
  assign o[3737] = i[14];
  assign o[3738] = i[14];
  assign o[3739] = i[14];
  assign o[3740] = i[14];
  assign o[3741] = i[14];
  assign o[3742] = i[14];
  assign o[3743] = i[14];
  assign o[3744] = i[14];
  assign o[3745] = i[14];
  assign o[3746] = i[14];
  assign o[3747] = i[14];
  assign o[3748] = i[14];
  assign o[3749] = i[14];
  assign o[3750] = i[14];
  assign o[3751] = i[14];
  assign o[3752] = i[14];
  assign o[3753] = i[14];
  assign o[3754] = i[14];
  assign o[3755] = i[14];
  assign o[3756] = i[14];
  assign o[3757] = i[14];
  assign o[3758] = i[14];
  assign o[3759] = i[14];
  assign o[3760] = i[14];
  assign o[3761] = i[14];
  assign o[3762] = i[14];
  assign o[3763] = i[14];
  assign o[3764] = i[14];
  assign o[3765] = i[14];
  assign o[3766] = i[14];
  assign o[3767] = i[14];
  assign o[3768] = i[14];
  assign o[3769] = i[14];
  assign o[3770] = i[14];
  assign o[3771] = i[14];
  assign o[3772] = i[14];
  assign o[3773] = i[14];
  assign o[3774] = i[14];
  assign o[3775] = i[14];
  assign o[3776] = i[14];
  assign o[3777] = i[14];
  assign o[3778] = i[14];
  assign o[3779] = i[14];
  assign o[3780] = i[14];
  assign o[3781] = i[14];
  assign o[3782] = i[14];
  assign o[3783] = i[14];
  assign o[3784] = i[14];
  assign o[3785] = i[14];
  assign o[3786] = i[14];
  assign o[3787] = i[14];
  assign o[3788] = i[14];
  assign o[3789] = i[14];
  assign o[3790] = i[14];
  assign o[3791] = i[14];
  assign o[3792] = i[14];
  assign o[3793] = i[14];
  assign o[3794] = i[14];
  assign o[3795] = i[14];
  assign o[3796] = i[14];
  assign o[3797] = i[14];
  assign o[3798] = i[14];
  assign o[3799] = i[14];
  assign o[3800] = i[14];
  assign o[3801] = i[14];
  assign o[3802] = i[14];
  assign o[3803] = i[14];
  assign o[3804] = i[14];
  assign o[3805] = i[14];
  assign o[3806] = i[14];
  assign o[3807] = i[14];
  assign o[3808] = i[14];
  assign o[3809] = i[14];
  assign o[3810] = i[14];
  assign o[3811] = i[14];
  assign o[3812] = i[14];
  assign o[3813] = i[14];
  assign o[3814] = i[14];
  assign o[3815] = i[14];
  assign o[3816] = i[14];
  assign o[3817] = i[14];
  assign o[3818] = i[14];
  assign o[3819] = i[14];
  assign o[3820] = i[14];
  assign o[3821] = i[14];
  assign o[3822] = i[14];
  assign o[3823] = i[14];
  assign o[3824] = i[14];
  assign o[3825] = i[14];
  assign o[3826] = i[14];
  assign o[3827] = i[14];
  assign o[3828] = i[14];
  assign o[3829] = i[14];
  assign o[3830] = i[14];
  assign o[3831] = i[14];
  assign o[3832] = i[14];
  assign o[3833] = i[14];
  assign o[3834] = i[14];
  assign o[3835] = i[14];
  assign o[3836] = i[14];
  assign o[3837] = i[14];
  assign o[3838] = i[14];
  assign o[3839] = i[14];
  assign o[3328] = i[13];
  assign o[3329] = i[13];
  assign o[3330] = i[13];
  assign o[3331] = i[13];
  assign o[3332] = i[13];
  assign o[3333] = i[13];
  assign o[3334] = i[13];
  assign o[3335] = i[13];
  assign o[3336] = i[13];
  assign o[3337] = i[13];
  assign o[3338] = i[13];
  assign o[3339] = i[13];
  assign o[3340] = i[13];
  assign o[3341] = i[13];
  assign o[3342] = i[13];
  assign o[3343] = i[13];
  assign o[3344] = i[13];
  assign o[3345] = i[13];
  assign o[3346] = i[13];
  assign o[3347] = i[13];
  assign o[3348] = i[13];
  assign o[3349] = i[13];
  assign o[3350] = i[13];
  assign o[3351] = i[13];
  assign o[3352] = i[13];
  assign o[3353] = i[13];
  assign o[3354] = i[13];
  assign o[3355] = i[13];
  assign o[3356] = i[13];
  assign o[3357] = i[13];
  assign o[3358] = i[13];
  assign o[3359] = i[13];
  assign o[3360] = i[13];
  assign o[3361] = i[13];
  assign o[3362] = i[13];
  assign o[3363] = i[13];
  assign o[3364] = i[13];
  assign o[3365] = i[13];
  assign o[3366] = i[13];
  assign o[3367] = i[13];
  assign o[3368] = i[13];
  assign o[3369] = i[13];
  assign o[3370] = i[13];
  assign o[3371] = i[13];
  assign o[3372] = i[13];
  assign o[3373] = i[13];
  assign o[3374] = i[13];
  assign o[3375] = i[13];
  assign o[3376] = i[13];
  assign o[3377] = i[13];
  assign o[3378] = i[13];
  assign o[3379] = i[13];
  assign o[3380] = i[13];
  assign o[3381] = i[13];
  assign o[3382] = i[13];
  assign o[3383] = i[13];
  assign o[3384] = i[13];
  assign o[3385] = i[13];
  assign o[3386] = i[13];
  assign o[3387] = i[13];
  assign o[3388] = i[13];
  assign o[3389] = i[13];
  assign o[3390] = i[13];
  assign o[3391] = i[13];
  assign o[3392] = i[13];
  assign o[3393] = i[13];
  assign o[3394] = i[13];
  assign o[3395] = i[13];
  assign o[3396] = i[13];
  assign o[3397] = i[13];
  assign o[3398] = i[13];
  assign o[3399] = i[13];
  assign o[3400] = i[13];
  assign o[3401] = i[13];
  assign o[3402] = i[13];
  assign o[3403] = i[13];
  assign o[3404] = i[13];
  assign o[3405] = i[13];
  assign o[3406] = i[13];
  assign o[3407] = i[13];
  assign o[3408] = i[13];
  assign o[3409] = i[13];
  assign o[3410] = i[13];
  assign o[3411] = i[13];
  assign o[3412] = i[13];
  assign o[3413] = i[13];
  assign o[3414] = i[13];
  assign o[3415] = i[13];
  assign o[3416] = i[13];
  assign o[3417] = i[13];
  assign o[3418] = i[13];
  assign o[3419] = i[13];
  assign o[3420] = i[13];
  assign o[3421] = i[13];
  assign o[3422] = i[13];
  assign o[3423] = i[13];
  assign o[3424] = i[13];
  assign o[3425] = i[13];
  assign o[3426] = i[13];
  assign o[3427] = i[13];
  assign o[3428] = i[13];
  assign o[3429] = i[13];
  assign o[3430] = i[13];
  assign o[3431] = i[13];
  assign o[3432] = i[13];
  assign o[3433] = i[13];
  assign o[3434] = i[13];
  assign o[3435] = i[13];
  assign o[3436] = i[13];
  assign o[3437] = i[13];
  assign o[3438] = i[13];
  assign o[3439] = i[13];
  assign o[3440] = i[13];
  assign o[3441] = i[13];
  assign o[3442] = i[13];
  assign o[3443] = i[13];
  assign o[3444] = i[13];
  assign o[3445] = i[13];
  assign o[3446] = i[13];
  assign o[3447] = i[13];
  assign o[3448] = i[13];
  assign o[3449] = i[13];
  assign o[3450] = i[13];
  assign o[3451] = i[13];
  assign o[3452] = i[13];
  assign o[3453] = i[13];
  assign o[3454] = i[13];
  assign o[3455] = i[13];
  assign o[3456] = i[13];
  assign o[3457] = i[13];
  assign o[3458] = i[13];
  assign o[3459] = i[13];
  assign o[3460] = i[13];
  assign o[3461] = i[13];
  assign o[3462] = i[13];
  assign o[3463] = i[13];
  assign o[3464] = i[13];
  assign o[3465] = i[13];
  assign o[3466] = i[13];
  assign o[3467] = i[13];
  assign o[3468] = i[13];
  assign o[3469] = i[13];
  assign o[3470] = i[13];
  assign o[3471] = i[13];
  assign o[3472] = i[13];
  assign o[3473] = i[13];
  assign o[3474] = i[13];
  assign o[3475] = i[13];
  assign o[3476] = i[13];
  assign o[3477] = i[13];
  assign o[3478] = i[13];
  assign o[3479] = i[13];
  assign o[3480] = i[13];
  assign o[3481] = i[13];
  assign o[3482] = i[13];
  assign o[3483] = i[13];
  assign o[3484] = i[13];
  assign o[3485] = i[13];
  assign o[3486] = i[13];
  assign o[3487] = i[13];
  assign o[3488] = i[13];
  assign o[3489] = i[13];
  assign o[3490] = i[13];
  assign o[3491] = i[13];
  assign o[3492] = i[13];
  assign o[3493] = i[13];
  assign o[3494] = i[13];
  assign o[3495] = i[13];
  assign o[3496] = i[13];
  assign o[3497] = i[13];
  assign o[3498] = i[13];
  assign o[3499] = i[13];
  assign o[3500] = i[13];
  assign o[3501] = i[13];
  assign o[3502] = i[13];
  assign o[3503] = i[13];
  assign o[3504] = i[13];
  assign o[3505] = i[13];
  assign o[3506] = i[13];
  assign o[3507] = i[13];
  assign o[3508] = i[13];
  assign o[3509] = i[13];
  assign o[3510] = i[13];
  assign o[3511] = i[13];
  assign o[3512] = i[13];
  assign o[3513] = i[13];
  assign o[3514] = i[13];
  assign o[3515] = i[13];
  assign o[3516] = i[13];
  assign o[3517] = i[13];
  assign o[3518] = i[13];
  assign o[3519] = i[13];
  assign o[3520] = i[13];
  assign o[3521] = i[13];
  assign o[3522] = i[13];
  assign o[3523] = i[13];
  assign o[3524] = i[13];
  assign o[3525] = i[13];
  assign o[3526] = i[13];
  assign o[3527] = i[13];
  assign o[3528] = i[13];
  assign o[3529] = i[13];
  assign o[3530] = i[13];
  assign o[3531] = i[13];
  assign o[3532] = i[13];
  assign o[3533] = i[13];
  assign o[3534] = i[13];
  assign o[3535] = i[13];
  assign o[3536] = i[13];
  assign o[3537] = i[13];
  assign o[3538] = i[13];
  assign o[3539] = i[13];
  assign o[3540] = i[13];
  assign o[3541] = i[13];
  assign o[3542] = i[13];
  assign o[3543] = i[13];
  assign o[3544] = i[13];
  assign o[3545] = i[13];
  assign o[3546] = i[13];
  assign o[3547] = i[13];
  assign o[3548] = i[13];
  assign o[3549] = i[13];
  assign o[3550] = i[13];
  assign o[3551] = i[13];
  assign o[3552] = i[13];
  assign o[3553] = i[13];
  assign o[3554] = i[13];
  assign o[3555] = i[13];
  assign o[3556] = i[13];
  assign o[3557] = i[13];
  assign o[3558] = i[13];
  assign o[3559] = i[13];
  assign o[3560] = i[13];
  assign o[3561] = i[13];
  assign o[3562] = i[13];
  assign o[3563] = i[13];
  assign o[3564] = i[13];
  assign o[3565] = i[13];
  assign o[3566] = i[13];
  assign o[3567] = i[13];
  assign o[3568] = i[13];
  assign o[3569] = i[13];
  assign o[3570] = i[13];
  assign o[3571] = i[13];
  assign o[3572] = i[13];
  assign o[3573] = i[13];
  assign o[3574] = i[13];
  assign o[3575] = i[13];
  assign o[3576] = i[13];
  assign o[3577] = i[13];
  assign o[3578] = i[13];
  assign o[3579] = i[13];
  assign o[3580] = i[13];
  assign o[3581] = i[13];
  assign o[3582] = i[13];
  assign o[3583] = i[13];
  assign o[3072] = i[12];
  assign o[3073] = i[12];
  assign o[3074] = i[12];
  assign o[3075] = i[12];
  assign o[3076] = i[12];
  assign o[3077] = i[12];
  assign o[3078] = i[12];
  assign o[3079] = i[12];
  assign o[3080] = i[12];
  assign o[3081] = i[12];
  assign o[3082] = i[12];
  assign o[3083] = i[12];
  assign o[3084] = i[12];
  assign o[3085] = i[12];
  assign o[3086] = i[12];
  assign o[3087] = i[12];
  assign o[3088] = i[12];
  assign o[3089] = i[12];
  assign o[3090] = i[12];
  assign o[3091] = i[12];
  assign o[3092] = i[12];
  assign o[3093] = i[12];
  assign o[3094] = i[12];
  assign o[3095] = i[12];
  assign o[3096] = i[12];
  assign o[3097] = i[12];
  assign o[3098] = i[12];
  assign o[3099] = i[12];
  assign o[3100] = i[12];
  assign o[3101] = i[12];
  assign o[3102] = i[12];
  assign o[3103] = i[12];
  assign o[3104] = i[12];
  assign o[3105] = i[12];
  assign o[3106] = i[12];
  assign o[3107] = i[12];
  assign o[3108] = i[12];
  assign o[3109] = i[12];
  assign o[3110] = i[12];
  assign o[3111] = i[12];
  assign o[3112] = i[12];
  assign o[3113] = i[12];
  assign o[3114] = i[12];
  assign o[3115] = i[12];
  assign o[3116] = i[12];
  assign o[3117] = i[12];
  assign o[3118] = i[12];
  assign o[3119] = i[12];
  assign o[3120] = i[12];
  assign o[3121] = i[12];
  assign o[3122] = i[12];
  assign o[3123] = i[12];
  assign o[3124] = i[12];
  assign o[3125] = i[12];
  assign o[3126] = i[12];
  assign o[3127] = i[12];
  assign o[3128] = i[12];
  assign o[3129] = i[12];
  assign o[3130] = i[12];
  assign o[3131] = i[12];
  assign o[3132] = i[12];
  assign o[3133] = i[12];
  assign o[3134] = i[12];
  assign o[3135] = i[12];
  assign o[3136] = i[12];
  assign o[3137] = i[12];
  assign o[3138] = i[12];
  assign o[3139] = i[12];
  assign o[3140] = i[12];
  assign o[3141] = i[12];
  assign o[3142] = i[12];
  assign o[3143] = i[12];
  assign o[3144] = i[12];
  assign o[3145] = i[12];
  assign o[3146] = i[12];
  assign o[3147] = i[12];
  assign o[3148] = i[12];
  assign o[3149] = i[12];
  assign o[3150] = i[12];
  assign o[3151] = i[12];
  assign o[3152] = i[12];
  assign o[3153] = i[12];
  assign o[3154] = i[12];
  assign o[3155] = i[12];
  assign o[3156] = i[12];
  assign o[3157] = i[12];
  assign o[3158] = i[12];
  assign o[3159] = i[12];
  assign o[3160] = i[12];
  assign o[3161] = i[12];
  assign o[3162] = i[12];
  assign o[3163] = i[12];
  assign o[3164] = i[12];
  assign o[3165] = i[12];
  assign o[3166] = i[12];
  assign o[3167] = i[12];
  assign o[3168] = i[12];
  assign o[3169] = i[12];
  assign o[3170] = i[12];
  assign o[3171] = i[12];
  assign o[3172] = i[12];
  assign o[3173] = i[12];
  assign o[3174] = i[12];
  assign o[3175] = i[12];
  assign o[3176] = i[12];
  assign o[3177] = i[12];
  assign o[3178] = i[12];
  assign o[3179] = i[12];
  assign o[3180] = i[12];
  assign o[3181] = i[12];
  assign o[3182] = i[12];
  assign o[3183] = i[12];
  assign o[3184] = i[12];
  assign o[3185] = i[12];
  assign o[3186] = i[12];
  assign o[3187] = i[12];
  assign o[3188] = i[12];
  assign o[3189] = i[12];
  assign o[3190] = i[12];
  assign o[3191] = i[12];
  assign o[3192] = i[12];
  assign o[3193] = i[12];
  assign o[3194] = i[12];
  assign o[3195] = i[12];
  assign o[3196] = i[12];
  assign o[3197] = i[12];
  assign o[3198] = i[12];
  assign o[3199] = i[12];
  assign o[3200] = i[12];
  assign o[3201] = i[12];
  assign o[3202] = i[12];
  assign o[3203] = i[12];
  assign o[3204] = i[12];
  assign o[3205] = i[12];
  assign o[3206] = i[12];
  assign o[3207] = i[12];
  assign o[3208] = i[12];
  assign o[3209] = i[12];
  assign o[3210] = i[12];
  assign o[3211] = i[12];
  assign o[3212] = i[12];
  assign o[3213] = i[12];
  assign o[3214] = i[12];
  assign o[3215] = i[12];
  assign o[3216] = i[12];
  assign o[3217] = i[12];
  assign o[3218] = i[12];
  assign o[3219] = i[12];
  assign o[3220] = i[12];
  assign o[3221] = i[12];
  assign o[3222] = i[12];
  assign o[3223] = i[12];
  assign o[3224] = i[12];
  assign o[3225] = i[12];
  assign o[3226] = i[12];
  assign o[3227] = i[12];
  assign o[3228] = i[12];
  assign o[3229] = i[12];
  assign o[3230] = i[12];
  assign o[3231] = i[12];
  assign o[3232] = i[12];
  assign o[3233] = i[12];
  assign o[3234] = i[12];
  assign o[3235] = i[12];
  assign o[3236] = i[12];
  assign o[3237] = i[12];
  assign o[3238] = i[12];
  assign o[3239] = i[12];
  assign o[3240] = i[12];
  assign o[3241] = i[12];
  assign o[3242] = i[12];
  assign o[3243] = i[12];
  assign o[3244] = i[12];
  assign o[3245] = i[12];
  assign o[3246] = i[12];
  assign o[3247] = i[12];
  assign o[3248] = i[12];
  assign o[3249] = i[12];
  assign o[3250] = i[12];
  assign o[3251] = i[12];
  assign o[3252] = i[12];
  assign o[3253] = i[12];
  assign o[3254] = i[12];
  assign o[3255] = i[12];
  assign o[3256] = i[12];
  assign o[3257] = i[12];
  assign o[3258] = i[12];
  assign o[3259] = i[12];
  assign o[3260] = i[12];
  assign o[3261] = i[12];
  assign o[3262] = i[12];
  assign o[3263] = i[12];
  assign o[3264] = i[12];
  assign o[3265] = i[12];
  assign o[3266] = i[12];
  assign o[3267] = i[12];
  assign o[3268] = i[12];
  assign o[3269] = i[12];
  assign o[3270] = i[12];
  assign o[3271] = i[12];
  assign o[3272] = i[12];
  assign o[3273] = i[12];
  assign o[3274] = i[12];
  assign o[3275] = i[12];
  assign o[3276] = i[12];
  assign o[3277] = i[12];
  assign o[3278] = i[12];
  assign o[3279] = i[12];
  assign o[3280] = i[12];
  assign o[3281] = i[12];
  assign o[3282] = i[12];
  assign o[3283] = i[12];
  assign o[3284] = i[12];
  assign o[3285] = i[12];
  assign o[3286] = i[12];
  assign o[3287] = i[12];
  assign o[3288] = i[12];
  assign o[3289] = i[12];
  assign o[3290] = i[12];
  assign o[3291] = i[12];
  assign o[3292] = i[12];
  assign o[3293] = i[12];
  assign o[3294] = i[12];
  assign o[3295] = i[12];
  assign o[3296] = i[12];
  assign o[3297] = i[12];
  assign o[3298] = i[12];
  assign o[3299] = i[12];
  assign o[3300] = i[12];
  assign o[3301] = i[12];
  assign o[3302] = i[12];
  assign o[3303] = i[12];
  assign o[3304] = i[12];
  assign o[3305] = i[12];
  assign o[3306] = i[12];
  assign o[3307] = i[12];
  assign o[3308] = i[12];
  assign o[3309] = i[12];
  assign o[3310] = i[12];
  assign o[3311] = i[12];
  assign o[3312] = i[12];
  assign o[3313] = i[12];
  assign o[3314] = i[12];
  assign o[3315] = i[12];
  assign o[3316] = i[12];
  assign o[3317] = i[12];
  assign o[3318] = i[12];
  assign o[3319] = i[12];
  assign o[3320] = i[12];
  assign o[3321] = i[12];
  assign o[3322] = i[12];
  assign o[3323] = i[12];
  assign o[3324] = i[12];
  assign o[3325] = i[12];
  assign o[3326] = i[12];
  assign o[3327] = i[12];
  assign o[2816] = i[11];
  assign o[2817] = i[11];
  assign o[2818] = i[11];
  assign o[2819] = i[11];
  assign o[2820] = i[11];
  assign o[2821] = i[11];
  assign o[2822] = i[11];
  assign o[2823] = i[11];
  assign o[2824] = i[11];
  assign o[2825] = i[11];
  assign o[2826] = i[11];
  assign o[2827] = i[11];
  assign o[2828] = i[11];
  assign o[2829] = i[11];
  assign o[2830] = i[11];
  assign o[2831] = i[11];
  assign o[2832] = i[11];
  assign o[2833] = i[11];
  assign o[2834] = i[11];
  assign o[2835] = i[11];
  assign o[2836] = i[11];
  assign o[2837] = i[11];
  assign o[2838] = i[11];
  assign o[2839] = i[11];
  assign o[2840] = i[11];
  assign o[2841] = i[11];
  assign o[2842] = i[11];
  assign o[2843] = i[11];
  assign o[2844] = i[11];
  assign o[2845] = i[11];
  assign o[2846] = i[11];
  assign o[2847] = i[11];
  assign o[2848] = i[11];
  assign o[2849] = i[11];
  assign o[2850] = i[11];
  assign o[2851] = i[11];
  assign o[2852] = i[11];
  assign o[2853] = i[11];
  assign o[2854] = i[11];
  assign o[2855] = i[11];
  assign o[2856] = i[11];
  assign o[2857] = i[11];
  assign o[2858] = i[11];
  assign o[2859] = i[11];
  assign o[2860] = i[11];
  assign o[2861] = i[11];
  assign o[2862] = i[11];
  assign o[2863] = i[11];
  assign o[2864] = i[11];
  assign o[2865] = i[11];
  assign o[2866] = i[11];
  assign o[2867] = i[11];
  assign o[2868] = i[11];
  assign o[2869] = i[11];
  assign o[2870] = i[11];
  assign o[2871] = i[11];
  assign o[2872] = i[11];
  assign o[2873] = i[11];
  assign o[2874] = i[11];
  assign o[2875] = i[11];
  assign o[2876] = i[11];
  assign o[2877] = i[11];
  assign o[2878] = i[11];
  assign o[2879] = i[11];
  assign o[2880] = i[11];
  assign o[2881] = i[11];
  assign o[2882] = i[11];
  assign o[2883] = i[11];
  assign o[2884] = i[11];
  assign o[2885] = i[11];
  assign o[2886] = i[11];
  assign o[2887] = i[11];
  assign o[2888] = i[11];
  assign o[2889] = i[11];
  assign o[2890] = i[11];
  assign o[2891] = i[11];
  assign o[2892] = i[11];
  assign o[2893] = i[11];
  assign o[2894] = i[11];
  assign o[2895] = i[11];
  assign o[2896] = i[11];
  assign o[2897] = i[11];
  assign o[2898] = i[11];
  assign o[2899] = i[11];
  assign o[2900] = i[11];
  assign o[2901] = i[11];
  assign o[2902] = i[11];
  assign o[2903] = i[11];
  assign o[2904] = i[11];
  assign o[2905] = i[11];
  assign o[2906] = i[11];
  assign o[2907] = i[11];
  assign o[2908] = i[11];
  assign o[2909] = i[11];
  assign o[2910] = i[11];
  assign o[2911] = i[11];
  assign o[2912] = i[11];
  assign o[2913] = i[11];
  assign o[2914] = i[11];
  assign o[2915] = i[11];
  assign o[2916] = i[11];
  assign o[2917] = i[11];
  assign o[2918] = i[11];
  assign o[2919] = i[11];
  assign o[2920] = i[11];
  assign o[2921] = i[11];
  assign o[2922] = i[11];
  assign o[2923] = i[11];
  assign o[2924] = i[11];
  assign o[2925] = i[11];
  assign o[2926] = i[11];
  assign o[2927] = i[11];
  assign o[2928] = i[11];
  assign o[2929] = i[11];
  assign o[2930] = i[11];
  assign o[2931] = i[11];
  assign o[2932] = i[11];
  assign o[2933] = i[11];
  assign o[2934] = i[11];
  assign o[2935] = i[11];
  assign o[2936] = i[11];
  assign o[2937] = i[11];
  assign o[2938] = i[11];
  assign o[2939] = i[11];
  assign o[2940] = i[11];
  assign o[2941] = i[11];
  assign o[2942] = i[11];
  assign o[2943] = i[11];
  assign o[2944] = i[11];
  assign o[2945] = i[11];
  assign o[2946] = i[11];
  assign o[2947] = i[11];
  assign o[2948] = i[11];
  assign o[2949] = i[11];
  assign o[2950] = i[11];
  assign o[2951] = i[11];
  assign o[2952] = i[11];
  assign o[2953] = i[11];
  assign o[2954] = i[11];
  assign o[2955] = i[11];
  assign o[2956] = i[11];
  assign o[2957] = i[11];
  assign o[2958] = i[11];
  assign o[2959] = i[11];
  assign o[2960] = i[11];
  assign o[2961] = i[11];
  assign o[2962] = i[11];
  assign o[2963] = i[11];
  assign o[2964] = i[11];
  assign o[2965] = i[11];
  assign o[2966] = i[11];
  assign o[2967] = i[11];
  assign o[2968] = i[11];
  assign o[2969] = i[11];
  assign o[2970] = i[11];
  assign o[2971] = i[11];
  assign o[2972] = i[11];
  assign o[2973] = i[11];
  assign o[2974] = i[11];
  assign o[2975] = i[11];
  assign o[2976] = i[11];
  assign o[2977] = i[11];
  assign o[2978] = i[11];
  assign o[2979] = i[11];
  assign o[2980] = i[11];
  assign o[2981] = i[11];
  assign o[2982] = i[11];
  assign o[2983] = i[11];
  assign o[2984] = i[11];
  assign o[2985] = i[11];
  assign o[2986] = i[11];
  assign o[2987] = i[11];
  assign o[2988] = i[11];
  assign o[2989] = i[11];
  assign o[2990] = i[11];
  assign o[2991] = i[11];
  assign o[2992] = i[11];
  assign o[2993] = i[11];
  assign o[2994] = i[11];
  assign o[2995] = i[11];
  assign o[2996] = i[11];
  assign o[2997] = i[11];
  assign o[2998] = i[11];
  assign o[2999] = i[11];
  assign o[3000] = i[11];
  assign o[3001] = i[11];
  assign o[3002] = i[11];
  assign o[3003] = i[11];
  assign o[3004] = i[11];
  assign o[3005] = i[11];
  assign o[3006] = i[11];
  assign o[3007] = i[11];
  assign o[3008] = i[11];
  assign o[3009] = i[11];
  assign o[3010] = i[11];
  assign o[3011] = i[11];
  assign o[3012] = i[11];
  assign o[3013] = i[11];
  assign o[3014] = i[11];
  assign o[3015] = i[11];
  assign o[3016] = i[11];
  assign o[3017] = i[11];
  assign o[3018] = i[11];
  assign o[3019] = i[11];
  assign o[3020] = i[11];
  assign o[3021] = i[11];
  assign o[3022] = i[11];
  assign o[3023] = i[11];
  assign o[3024] = i[11];
  assign o[3025] = i[11];
  assign o[3026] = i[11];
  assign o[3027] = i[11];
  assign o[3028] = i[11];
  assign o[3029] = i[11];
  assign o[3030] = i[11];
  assign o[3031] = i[11];
  assign o[3032] = i[11];
  assign o[3033] = i[11];
  assign o[3034] = i[11];
  assign o[3035] = i[11];
  assign o[3036] = i[11];
  assign o[3037] = i[11];
  assign o[3038] = i[11];
  assign o[3039] = i[11];
  assign o[3040] = i[11];
  assign o[3041] = i[11];
  assign o[3042] = i[11];
  assign o[3043] = i[11];
  assign o[3044] = i[11];
  assign o[3045] = i[11];
  assign o[3046] = i[11];
  assign o[3047] = i[11];
  assign o[3048] = i[11];
  assign o[3049] = i[11];
  assign o[3050] = i[11];
  assign o[3051] = i[11];
  assign o[3052] = i[11];
  assign o[3053] = i[11];
  assign o[3054] = i[11];
  assign o[3055] = i[11];
  assign o[3056] = i[11];
  assign o[3057] = i[11];
  assign o[3058] = i[11];
  assign o[3059] = i[11];
  assign o[3060] = i[11];
  assign o[3061] = i[11];
  assign o[3062] = i[11];
  assign o[3063] = i[11];
  assign o[3064] = i[11];
  assign o[3065] = i[11];
  assign o[3066] = i[11];
  assign o[3067] = i[11];
  assign o[3068] = i[11];
  assign o[3069] = i[11];
  assign o[3070] = i[11];
  assign o[3071] = i[11];
  assign o[2560] = i[10];
  assign o[2561] = i[10];
  assign o[2562] = i[10];
  assign o[2563] = i[10];
  assign o[2564] = i[10];
  assign o[2565] = i[10];
  assign o[2566] = i[10];
  assign o[2567] = i[10];
  assign o[2568] = i[10];
  assign o[2569] = i[10];
  assign o[2570] = i[10];
  assign o[2571] = i[10];
  assign o[2572] = i[10];
  assign o[2573] = i[10];
  assign o[2574] = i[10];
  assign o[2575] = i[10];
  assign o[2576] = i[10];
  assign o[2577] = i[10];
  assign o[2578] = i[10];
  assign o[2579] = i[10];
  assign o[2580] = i[10];
  assign o[2581] = i[10];
  assign o[2582] = i[10];
  assign o[2583] = i[10];
  assign o[2584] = i[10];
  assign o[2585] = i[10];
  assign o[2586] = i[10];
  assign o[2587] = i[10];
  assign o[2588] = i[10];
  assign o[2589] = i[10];
  assign o[2590] = i[10];
  assign o[2591] = i[10];
  assign o[2592] = i[10];
  assign o[2593] = i[10];
  assign o[2594] = i[10];
  assign o[2595] = i[10];
  assign o[2596] = i[10];
  assign o[2597] = i[10];
  assign o[2598] = i[10];
  assign o[2599] = i[10];
  assign o[2600] = i[10];
  assign o[2601] = i[10];
  assign o[2602] = i[10];
  assign o[2603] = i[10];
  assign o[2604] = i[10];
  assign o[2605] = i[10];
  assign o[2606] = i[10];
  assign o[2607] = i[10];
  assign o[2608] = i[10];
  assign o[2609] = i[10];
  assign o[2610] = i[10];
  assign o[2611] = i[10];
  assign o[2612] = i[10];
  assign o[2613] = i[10];
  assign o[2614] = i[10];
  assign o[2615] = i[10];
  assign o[2616] = i[10];
  assign o[2617] = i[10];
  assign o[2618] = i[10];
  assign o[2619] = i[10];
  assign o[2620] = i[10];
  assign o[2621] = i[10];
  assign o[2622] = i[10];
  assign o[2623] = i[10];
  assign o[2624] = i[10];
  assign o[2625] = i[10];
  assign o[2626] = i[10];
  assign o[2627] = i[10];
  assign o[2628] = i[10];
  assign o[2629] = i[10];
  assign o[2630] = i[10];
  assign o[2631] = i[10];
  assign o[2632] = i[10];
  assign o[2633] = i[10];
  assign o[2634] = i[10];
  assign o[2635] = i[10];
  assign o[2636] = i[10];
  assign o[2637] = i[10];
  assign o[2638] = i[10];
  assign o[2639] = i[10];
  assign o[2640] = i[10];
  assign o[2641] = i[10];
  assign o[2642] = i[10];
  assign o[2643] = i[10];
  assign o[2644] = i[10];
  assign o[2645] = i[10];
  assign o[2646] = i[10];
  assign o[2647] = i[10];
  assign o[2648] = i[10];
  assign o[2649] = i[10];
  assign o[2650] = i[10];
  assign o[2651] = i[10];
  assign o[2652] = i[10];
  assign o[2653] = i[10];
  assign o[2654] = i[10];
  assign o[2655] = i[10];
  assign o[2656] = i[10];
  assign o[2657] = i[10];
  assign o[2658] = i[10];
  assign o[2659] = i[10];
  assign o[2660] = i[10];
  assign o[2661] = i[10];
  assign o[2662] = i[10];
  assign o[2663] = i[10];
  assign o[2664] = i[10];
  assign o[2665] = i[10];
  assign o[2666] = i[10];
  assign o[2667] = i[10];
  assign o[2668] = i[10];
  assign o[2669] = i[10];
  assign o[2670] = i[10];
  assign o[2671] = i[10];
  assign o[2672] = i[10];
  assign o[2673] = i[10];
  assign o[2674] = i[10];
  assign o[2675] = i[10];
  assign o[2676] = i[10];
  assign o[2677] = i[10];
  assign o[2678] = i[10];
  assign o[2679] = i[10];
  assign o[2680] = i[10];
  assign o[2681] = i[10];
  assign o[2682] = i[10];
  assign o[2683] = i[10];
  assign o[2684] = i[10];
  assign o[2685] = i[10];
  assign o[2686] = i[10];
  assign o[2687] = i[10];
  assign o[2688] = i[10];
  assign o[2689] = i[10];
  assign o[2690] = i[10];
  assign o[2691] = i[10];
  assign o[2692] = i[10];
  assign o[2693] = i[10];
  assign o[2694] = i[10];
  assign o[2695] = i[10];
  assign o[2696] = i[10];
  assign o[2697] = i[10];
  assign o[2698] = i[10];
  assign o[2699] = i[10];
  assign o[2700] = i[10];
  assign o[2701] = i[10];
  assign o[2702] = i[10];
  assign o[2703] = i[10];
  assign o[2704] = i[10];
  assign o[2705] = i[10];
  assign o[2706] = i[10];
  assign o[2707] = i[10];
  assign o[2708] = i[10];
  assign o[2709] = i[10];
  assign o[2710] = i[10];
  assign o[2711] = i[10];
  assign o[2712] = i[10];
  assign o[2713] = i[10];
  assign o[2714] = i[10];
  assign o[2715] = i[10];
  assign o[2716] = i[10];
  assign o[2717] = i[10];
  assign o[2718] = i[10];
  assign o[2719] = i[10];
  assign o[2720] = i[10];
  assign o[2721] = i[10];
  assign o[2722] = i[10];
  assign o[2723] = i[10];
  assign o[2724] = i[10];
  assign o[2725] = i[10];
  assign o[2726] = i[10];
  assign o[2727] = i[10];
  assign o[2728] = i[10];
  assign o[2729] = i[10];
  assign o[2730] = i[10];
  assign o[2731] = i[10];
  assign o[2732] = i[10];
  assign o[2733] = i[10];
  assign o[2734] = i[10];
  assign o[2735] = i[10];
  assign o[2736] = i[10];
  assign o[2737] = i[10];
  assign o[2738] = i[10];
  assign o[2739] = i[10];
  assign o[2740] = i[10];
  assign o[2741] = i[10];
  assign o[2742] = i[10];
  assign o[2743] = i[10];
  assign o[2744] = i[10];
  assign o[2745] = i[10];
  assign o[2746] = i[10];
  assign o[2747] = i[10];
  assign o[2748] = i[10];
  assign o[2749] = i[10];
  assign o[2750] = i[10];
  assign o[2751] = i[10];
  assign o[2752] = i[10];
  assign o[2753] = i[10];
  assign o[2754] = i[10];
  assign o[2755] = i[10];
  assign o[2756] = i[10];
  assign o[2757] = i[10];
  assign o[2758] = i[10];
  assign o[2759] = i[10];
  assign o[2760] = i[10];
  assign o[2761] = i[10];
  assign o[2762] = i[10];
  assign o[2763] = i[10];
  assign o[2764] = i[10];
  assign o[2765] = i[10];
  assign o[2766] = i[10];
  assign o[2767] = i[10];
  assign o[2768] = i[10];
  assign o[2769] = i[10];
  assign o[2770] = i[10];
  assign o[2771] = i[10];
  assign o[2772] = i[10];
  assign o[2773] = i[10];
  assign o[2774] = i[10];
  assign o[2775] = i[10];
  assign o[2776] = i[10];
  assign o[2777] = i[10];
  assign o[2778] = i[10];
  assign o[2779] = i[10];
  assign o[2780] = i[10];
  assign o[2781] = i[10];
  assign o[2782] = i[10];
  assign o[2783] = i[10];
  assign o[2784] = i[10];
  assign o[2785] = i[10];
  assign o[2786] = i[10];
  assign o[2787] = i[10];
  assign o[2788] = i[10];
  assign o[2789] = i[10];
  assign o[2790] = i[10];
  assign o[2791] = i[10];
  assign o[2792] = i[10];
  assign o[2793] = i[10];
  assign o[2794] = i[10];
  assign o[2795] = i[10];
  assign o[2796] = i[10];
  assign o[2797] = i[10];
  assign o[2798] = i[10];
  assign o[2799] = i[10];
  assign o[2800] = i[10];
  assign o[2801] = i[10];
  assign o[2802] = i[10];
  assign o[2803] = i[10];
  assign o[2804] = i[10];
  assign o[2805] = i[10];
  assign o[2806] = i[10];
  assign o[2807] = i[10];
  assign o[2808] = i[10];
  assign o[2809] = i[10];
  assign o[2810] = i[10];
  assign o[2811] = i[10];
  assign o[2812] = i[10];
  assign o[2813] = i[10];
  assign o[2814] = i[10];
  assign o[2815] = i[10];
  assign o[2304] = i[9];
  assign o[2305] = i[9];
  assign o[2306] = i[9];
  assign o[2307] = i[9];
  assign o[2308] = i[9];
  assign o[2309] = i[9];
  assign o[2310] = i[9];
  assign o[2311] = i[9];
  assign o[2312] = i[9];
  assign o[2313] = i[9];
  assign o[2314] = i[9];
  assign o[2315] = i[9];
  assign o[2316] = i[9];
  assign o[2317] = i[9];
  assign o[2318] = i[9];
  assign o[2319] = i[9];
  assign o[2320] = i[9];
  assign o[2321] = i[9];
  assign o[2322] = i[9];
  assign o[2323] = i[9];
  assign o[2324] = i[9];
  assign o[2325] = i[9];
  assign o[2326] = i[9];
  assign o[2327] = i[9];
  assign o[2328] = i[9];
  assign o[2329] = i[9];
  assign o[2330] = i[9];
  assign o[2331] = i[9];
  assign o[2332] = i[9];
  assign o[2333] = i[9];
  assign o[2334] = i[9];
  assign o[2335] = i[9];
  assign o[2336] = i[9];
  assign o[2337] = i[9];
  assign o[2338] = i[9];
  assign o[2339] = i[9];
  assign o[2340] = i[9];
  assign o[2341] = i[9];
  assign o[2342] = i[9];
  assign o[2343] = i[9];
  assign o[2344] = i[9];
  assign o[2345] = i[9];
  assign o[2346] = i[9];
  assign o[2347] = i[9];
  assign o[2348] = i[9];
  assign o[2349] = i[9];
  assign o[2350] = i[9];
  assign o[2351] = i[9];
  assign o[2352] = i[9];
  assign o[2353] = i[9];
  assign o[2354] = i[9];
  assign o[2355] = i[9];
  assign o[2356] = i[9];
  assign o[2357] = i[9];
  assign o[2358] = i[9];
  assign o[2359] = i[9];
  assign o[2360] = i[9];
  assign o[2361] = i[9];
  assign o[2362] = i[9];
  assign o[2363] = i[9];
  assign o[2364] = i[9];
  assign o[2365] = i[9];
  assign o[2366] = i[9];
  assign o[2367] = i[9];
  assign o[2368] = i[9];
  assign o[2369] = i[9];
  assign o[2370] = i[9];
  assign o[2371] = i[9];
  assign o[2372] = i[9];
  assign o[2373] = i[9];
  assign o[2374] = i[9];
  assign o[2375] = i[9];
  assign o[2376] = i[9];
  assign o[2377] = i[9];
  assign o[2378] = i[9];
  assign o[2379] = i[9];
  assign o[2380] = i[9];
  assign o[2381] = i[9];
  assign o[2382] = i[9];
  assign o[2383] = i[9];
  assign o[2384] = i[9];
  assign o[2385] = i[9];
  assign o[2386] = i[9];
  assign o[2387] = i[9];
  assign o[2388] = i[9];
  assign o[2389] = i[9];
  assign o[2390] = i[9];
  assign o[2391] = i[9];
  assign o[2392] = i[9];
  assign o[2393] = i[9];
  assign o[2394] = i[9];
  assign o[2395] = i[9];
  assign o[2396] = i[9];
  assign o[2397] = i[9];
  assign o[2398] = i[9];
  assign o[2399] = i[9];
  assign o[2400] = i[9];
  assign o[2401] = i[9];
  assign o[2402] = i[9];
  assign o[2403] = i[9];
  assign o[2404] = i[9];
  assign o[2405] = i[9];
  assign o[2406] = i[9];
  assign o[2407] = i[9];
  assign o[2408] = i[9];
  assign o[2409] = i[9];
  assign o[2410] = i[9];
  assign o[2411] = i[9];
  assign o[2412] = i[9];
  assign o[2413] = i[9];
  assign o[2414] = i[9];
  assign o[2415] = i[9];
  assign o[2416] = i[9];
  assign o[2417] = i[9];
  assign o[2418] = i[9];
  assign o[2419] = i[9];
  assign o[2420] = i[9];
  assign o[2421] = i[9];
  assign o[2422] = i[9];
  assign o[2423] = i[9];
  assign o[2424] = i[9];
  assign o[2425] = i[9];
  assign o[2426] = i[9];
  assign o[2427] = i[9];
  assign o[2428] = i[9];
  assign o[2429] = i[9];
  assign o[2430] = i[9];
  assign o[2431] = i[9];
  assign o[2432] = i[9];
  assign o[2433] = i[9];
  assign o[2434] = i[9];
  assign o[2435] = i[9];
  assign o[2436] = i[9];
  assign o[2437] = i[9];
  assign o[2438] = i[9];
  assign o[2439] = i[9];
  assign o[2440] = i[9];
  assign o[2441] = i[9];
  assign o[2442] = i[9];
  assign o[2443] = i[9];
  assign o[2444] = i[9];
  assign o[2445] = i[9];
  assign o[2446] = i[9];
  assign o[2447] = i[9];
  assign o[2448] = i[9];
  assign o[2449] = i[9];
  assign o[2450] = i[9];
  assign o[2451] = i[9];
  assign o[2452] = i[9];
  assign o[2453] = i[9];
  assign o[2454] = i[9];
  assign o[2455] = i[9];
  assign o[2456] = i[9];
  assign o[2457] = i[9];
  assign o[2458] = i[9];
  assign o[2459] = i[9];
  assign o[2460] = i[9];
  assign o[2461] = i[9];
  assign o[2462] = i[9];
  assign o[2463] = i[9];
  assign o[2464] = i[9];
  assign o[2465] = i[9];
  assign o[2466] = i[9];
  assign o[2467] = i[9];
  assign o[2468] = i[9];
  assign o[2469] = i[9];
  assign o[2470] = i[9];
  assign o[2471] = i[9];
  assign o[2472] = i[9];
  assign o[2473] = i[9];
  assign o[2474] = i[9];
  assign o[2475] = i[9];
  assign o[2476] = i[9];
  assign o[2477] = i[9];
  assign o[2478] = i[9];
  assign o[2479] = i[9];
  assign o[2480] = i[9];
  assign o[2481] = i[9];
  assign o[2482] = i[9];
  assign o[2483] = i[9];
  assign o[2484] = i[9];
  assign o[2485] = i[9];
  assign o[2486] = i[9];
  assign o[2487] = i[9];
  assign o[2488] = i[9];
  assign o[2489] = i[9];
  assign o[2490] = i[9];
  assign o[2491] = i[9];
  assign o[2492] = i[9];
  assign o[2493] = i[9];
  assign o[2494] = i[9];
  assign o[2495] = i[9];
  assign o[2496] = i[9];
  assign o[2497] = i[9];
  assign o[2498] = i[9];
  assign o[2499] = i[9];
  assign o[2500] = i[9];
  assign o[2501] = i[9];
  assign o[2502] = i[9];
  assign o[2503] = i[9];
  assign o[2504] = i[9];
  assign o[2505] = i[9];
  assign o[2506] = i[9];
  assign o[2507] = i[9];
  assign o[2508] = i[9];
  assign o[2509] = i[9];
  assign o[2510] = i[9];
  assign o[2511] = i[9];
  assign o[2512] = i[9];
  assign o[2513] = i[9];
  assign o[2514] = i[9];
  assign o[2515] = i[9];
  assign o[2516] = i[9];
  assign o[2517] = i[9];
  assign o[2518] = i[9];
  assign o[2519] = i[9];
  assign o[2520] = i[9];
  assign o[2521] = i[9];
  assign o[2522] = i[9];
  assign o[2523] = i[9];
  assign o[2524] = i[9];
  assign o[2525] = i[9];
  assign o[2526] = i[9];
  assign o[2527] = i[9];
  assign o[2528] = i[9];
  assign o[2529] = i[9];
  assign o[2530] = i[9];
  assign o[2531] = i[9];
  assign o[2532] = i[9];
  assign o[2533] = i[9];
  assign o[2534] = i[9];
  assign o[2535] = i[9];
  assign o[2536] = i[9];
  assign o[2537] = i[9];
  assign o[2538] = i[9];
  assign o[2539] = i[9];
  assign o[2540] = i[9];
  assign o[2541] = i[9];
  assign o[2542] = i[9];
  assign o[2543] = i[9];
  assign o[2544] = i[9];
  assign o[2545] = i[9];
  assign o[2546] = i[9];
  assign o[2547] = i[9];
  assign o[2548] = i[9];
  assign o[2549] = i[9];
  assign o[2550] = i[9];
  assign o[2551] = i[9];
  assign o[2552] = i[9];
  assign o[2553] = i[9];
  assign o[2554] = i[9];
  assign o[2555] = i[9];
  assign o[2556] = i[9];
  assign o[2557] = i[9];
  assign o[2558] = i[9];
  assign o[2559] = i[9];
  assign o[2048] = i[8];
  assign o[2049] = i[8];
  assign o[2050] = i[8];
  assign o[2051] = i[8];
  assign o[2052] = i[8];
  assign o[2053] = i[8];
  assign o[2054] = i[8];
  assign o[2055] = i[8];
  assign o[2056] = i[8];
  assign o[2057] = i[8];
  assign o[2058] = i[8];
  assign o[2059] = i[8];
  assign o[2060] = i[8];
  assign o[2061] = i[8];
  assign o[2062] = i[8];
  assign o[2063] = i[8];
  assign o[2064] = i[8];
  assign o[2065] = i[8];
  assign o[2066] = i[8];
  assign o[2067] = i[8];
  assign o[2068] = i[8];
  assign o[2069] = i[8];
  assign o[2070] = i[8];
  assign o[2071] = i[8];
  assign o[2072] = i[8];
  assign o[2073] = i[8];
  assign o[2074] = i[8];
  assign o[2075] = i[8];
  assign o[2076] = i[8];
  assign o[2077] = i[8];
  assign o[2078] = i[8];
  assign o[2079] = i[8];
  assign o[2080] = i[8];
  assign o[2081] = i[8];
  assign o[2082] = i[8];
  assign o[2083] = i[8];
  assign o[2084] = i[8];
  assign o[2085] = i[8];
  assign o[2086] = i[8];
  assign o[2087] = i[8];
  assign o[2088] = i[8];
  assign o[2089] = i[8];
  assign o[2090] = i[8];
  assign o[2091] = i[8];
  assign o[2092] = i[8];
  assign o[2093] = i[8];
  assign o[2094] = i[8];
  assign o[2095] = i[8];
  assign o[2096] = i[8];
  assign o[2097] = i[8];
  assign o[2098] = i[8];
  assign o[2099] = i[8];
  assign o[2100] = i[8];
  assign o[2101] = i[8];
  assign o[2102] = i[8];
  assign o[2103] = i[8];
  assign o[2104] = i[8];
  assign o[2105] = i[8];
  assign o[2106] = i[8];
  assign o[2107] = i[8];
  assign o[2108] = i[8];
  assign o[2109] = i[8];
  assign o[2110] = i[8];
  assign o[2111] = i[8];
  assign o[2112] = i[8];
  assign o[2113] = i[8];
  assign o[2114] = i[8];
  assign o[2115] = i[8];
  assign o[2116] = i[8];
  assign o[2117] = i[8];
  assign o[2118] = i[8];
  assign o[2119] = i[8];
  assign o[2120] = i[8];
  assign o[2121] = i[8];
  assign o[2122] = i[8];
  assign o[2123] = i[8];
  assign o[2124] = i[8];
  assign o[2125] = i[8];
  assign o[2126] = i[8];
  assign o[2127] = i[8];
  assign o[2128] = i[8];
  assign o[2129] = i[8];
  assign o[2130] = i[8];
  assign o[2131] = i[8];
  assign o[2132] = i[8];
  assign o[2133] = i[8];
  assign o[2134] = i[8];
  assign o[2135] = i[8];
  assign o[2136] = i[8];
  assign o[2137] = i[8];
  assign o[2138] = i[8];
  assign o[2139] = i[8];
  assign o[2140] = i[8];
  assign o[2141] = i[8];
  assign o[2142] = i[8];
  assign o[2143] = i[8];
  assign o[2144] = i[8];
  assign o[2145] = i[8];
  assign o[2146] = i[8];
  assign o[2147] = i[8];
  assign o[2148] = i[8];
  assign o[2149] = i[8];
  assign o[2150] = i[8];
  assign o[2151] = i[8];
  assign o[2152] = i[8];
  assign o[2153] = i[8];
  assign o[2154] = i[8];
  assign o[2155] = i[8];
  assign o[2156] = i[8];
  assign o[2157] = i[8];
  assign o[2158] = i[8];
  assign o[2159] = i[8];
  assign o[2160] = i[8];
  assign o[2161] = i[8];
  assign o[2162] = i[8];
  assign o[2163] = i[8];
  assign o[2164] = i[8];
  assign o[2165] = i[8];
  assign o[2166] = i[8];
  assign o[2167] = i[8];
  assign o[2168] = i[8];
  assign o[2169] = i[8];
  assign o[2170] = i[8];
  assign o[2171] = i[8];
  assign o[2172] = i[8];
  assign o[2173] = i[8];
  assign o[2174] = i[8];
  assign o[2175] = i[8];
  assign o[2176] = i[8];
  assign o[2177] = i[8];
  assign o[2178] = i[8];
  assign o[2179] = i[8];
  assign o[2180] = i[8];
  assign o[2181] = i[8];
  assign o[2182] = i[8];
  assign o[2183] = i[8];
  assign o[2184] = i[8];
  assign o[2185] = i[8];
  assign o[2186] = i[8];
  assign o[2187] = i[8];
  assign o[2188] = i[8];
  assign o[2189] = i[8];
  assign o[2190] = i[8];
  assign o[2191] = i[8];
  assign o[2192] = i[8];
  assign o[2193] = i[8];
  assign o[2194] = i[8];
  assign o[2195] = i[8];
  assign o[2196] = i[8];
  assign o[2197] = i[8];
  assign o[2198] = i[8];
  assign o[2199] = i[8];
  assign o[2200] = i[8];
  assign o[2201] = i[8];
  assign o[2202] = i[8];
  assign o[2203] = i[8];
  assign o[2204] = i[8];
  assign o[2205] = i[8];
  assign o[2206] = i[8];
  assign o[2207] = i[8];
  assign o[2208] = i[8];
  assign o[2209] = i[8];
  assign o[2210] = i[8];
  assign o[2211] = i[8];
  assign o[2212] = i[8];
  assign o[2213] = i[8];
  assign o[2214] = i[8];
  assign o[2215] = i[8];
  assign o[2216] = i[8];
  assign o[2217] = i[8];
  assign o[2218] = i[8];
  assign o[2219] = i[8];
  assign o[2220] = i[8];
  assign o[2221] = i[8];
  assign o[2222] = i[8];
  assign o[2223] = i[8];
  assign o[2224] = i[8];
  assign o[2225] = i[8];
  assign o[2226] = i[8];
  assign o[2227] = i[8];
  assign o[2228] = i[8];
  assign o[2229] = i[8];
  assign o[2230] = i[8];
  assign o[2231] = i[8];
  assign o[2232] = i[8];
  assign o[2233] = i[8];
  assign o[2234] = i[8];
  assign o[2235] = i[8];
  assign o[2236] = i[8];
  assign o[2237] = i[8];
  assign o[2238] = i[8];
  assign o[2239] = i[8];
  assign o[2240] = i[8];
  assign o[2241] = i[8];
  assign o[2242] = i[8];
  assign o[2243] = i[8];
  assign o[2244] = i[8];
  assign o[2245] = i[8];
  assign o[2246] = i[8];
  assign o[2247] = i[8];
  assign o[2248] = i[8];
  assign o[2249] = i[8];
  assign o[2250] = i[8];
  assign o[2251] = i[8];
  assign o[2252] = i[8];
  assign o[2253] = i[8];
  assign o[2254] = i[8];
  assign o[2255] = i[8];
  assign o[2256] = i[8];
  assign o[2257] = i[8];
  assign o[2258] = i[8];
  assign o[2259] = i[8];
  assign o[2260] = i[8];
  assign o[2261] = i[8];
  assign o[2262] = i[8];
  assign o[2263] = i[8];
  assign o[2264] = i[8];
  assign o[2265] = i[8];
  assign o[2266] = i[8];
  assign o[2267] = i[8];
  assign o[2268] = i[8];
  assign o[2269] = i[8];
  assign o[2270] = i[8];
  assign o[2271] = i[8];
  assign o[2272] = i[8];
  assign o[2273] = i[8];
  assign o[2274] = i[8];
  assign o[2275] = i[8];
  assign o[2276] = i[8];
  assign o[2277] = i[8];
  assign o[2278] = i[8];
  assign o[2279] = i[8];
  assign o[2280] = i[8];
  assign o[2281] = i[8];
  assign o[2282] = i[8];
  assign o[2283] = i[8];
  assign o[2284] = i[8];
  assign o[2285] = i[8];
  assign o[2286] = i[8];
  assign o[2287] = i[8];
  assign o[2288] = i[8];
  assign o[2289] = i[8];
  assign o[2290] = i[8];
  assign o[2291] = i[8];
  assign o[2292] = i[8];
  assign o[2293] = i[8];
  assign o[2294] = i[8];
  assign o[2295] = i[8];
  assign o[2296] = i[8];
  assign o[2297] = i[8];
  assign o[2298] = i[8];
  assign o[2299] = i[8];
  assign o[2300] = i[8];
  assign o[2301] = i[8];
  assign o[2302] = i[8];
  assign o[2303] = i[8];
  assign o[1792] = i[7];
  assign o[1793] = i[7];
  assign o[1794] = i[7];
  assign o[1795] = i[7];
  assign o[1796] = i[7];
  assign o[1797] = i[7];
  assign o[1798] = i[7];
  assign o[1799] = i[7];
  assign o[1800] = i[7];
  assign o[1801] = i[7];
  assign o[1802] = i[7];
  assign o[1803] = i[7];
  assign o[1804] = i[7];
  assign o[1805] = i[7];
  assign o[1806] = i[7];
  assign o[1807] = i[7];
  assign o[1808] = i[7];
  assign o[1809] = i[7];
  assign o[1810] = i[7];
  assign o[1811] = i[7];
  assign o[1812] = i[7];
  assign o[1813] = i[7];
  assign o[1814] = i[7];
  assign o[1815] = i[7];
  assign o[1816] = i[7];
  assign o[1817] = i[7];
  assign o[1818] = i[7];
  assign o[1819] = i[7];
  assign o[1820] = i[7];
  assign o[1821] = i[7];
  assign o[1822] = i[7];
  assign o[1823] = i[7];
  assign o[1824] = i[7];
  assign o[1825] = i[7];
  assign o[1826] = i[7];
  assign o[1827] = i[7];
  assign o[1828] = i[7];
  assign o[1829] = i[7];
  assign o[1830] = i[7];
  assign o[1831] = i[7];
  assign o[1832] = i[7];
  assign o[1833] = i[7];
  assign o[1834] = i[7];
  assign o[1835] = i[7];
  assign o[1836] = i[7];
  assign o[1837] = i[7];
  assign o[1838] = i[7];
  assign o[1839] = i[7];
  assign o[1840] = i[7];
  assign o[1841] = i[7];
  assign o[1842] = i[7];
  assign o[1843] = i[7];
  assign o[1844] = i[7];
  assign o[1845] = i[7];
  assign o[1846] = i[7];
  assign o[1847] = i[7];
  assign o[1848] = i[7];
  assign o[1849] = i[7];
  assign o[1850] = i[7];
  assign o[1851] = i[7];
  assign o[1852] = i[7];
  assign o[1853] = i[7];
  assign o[1854] = i[7];
  assign o[1855] = i[7];
  assign o[1856] = i[7];
  assign o[1857] = i[7];
  assign o[1858] = i[7];
  assign o[1859] = i[7];
  assign o[1860] = i[7];
  assign o[1861] = i[7];
  assign o[1862] = i[7];
  assign o[1863] = i[7];
  assign o[1864] = i[7];
  assign o[1865] = i[7];
  assign o[1866] = i[7];
  assign o[1867] = i[7];
  assign o[1868] = i[7];
  assign o[1869] = i[7];
  assign o[1870] = i[7];
  assign o[1871] = i[7];
  assign o[1872] = i[7];
  assign o[1873] = i[7];
  assign o[1874] = i[7];
  assign o[1875] = i[7];
  assign o[1876] = i[7];
  assign o[1877] = i[7];
  assign o[1878] = i[7];
  assign o[1879] = i[7];
  assign o[1880] = i[7];
  assign o[1881] = i[7];
  assign o[1882] = i[7];
  assign o[1883] = i[7];
  assign o[1884] = i[7];
  assign o[1885] = i[7];
  assign o[1886] = i[7];
  assign o[1887] = i[7];
  assign o[1888] = i[7];
  assign o[1889] = i[7];
  assign o[1890] = i[7];
  assign o[1891] = i[7];
  assign o[1892] = i[7];
  assign o[1893] = i[7];
  assign o[1894] = i[7];
  assign o[1895] = i[7];
  assign o[1896] = i[7];
  assign o[1897] = i[7];
  assign o[1898] = i[7];
  assign o[1899] = i[7];
  assign o[1900] = i[7];
  assign o[1901] = i[7];
  assign o[1902] = i[7];
  assign o[1903] = i[7];
  assign o[1904] = i[7];
  assign o[1905] = i[7];
  assign o[1906] = i[7];
  assign o[1907] = i[7];
  assign o[1908] = i[7];
  assign o[1909] = i[7];
  assign o[1910] = i[7];
  assign o[1911] = i[7];
  assign o[1912] = i[7];
  assign o[1913] = i[7];
  assign o[1914] = i[7];
  assign o[1915] = i[7];
  assign o[1916] = i[7];
  assign o[1917] = i[7];
  assign o[1918] = i[7];
  assign o[1919] = i[7];
  assign o[1920] = i[7];
  assign o[1921] = i[7];
  assign o[1922] = i[7];
  assign o[1923] = i[7];
  assign o[1924] = i[7];
  assign o[1925] = i[7];
  assign o[1926] = i[7];
  assign o[1927] = i[7];
  assign o[1928] = i[7];
  assign o[1929] = i[7];
  assign o[1930] = i[7];
  assign o[1931] = i[7];
  assign o[1932] = i[7];
  assign o[1933] = i[7];
  assign o[1934] = i[7];
  assign o[1935] = i[7];
  assign o[1936] = i[7];
  assign o[1937] = i[7];
  assign o[1938] = i[7];
  assign o[1939] = i[7];
  assign o[1940] = i[7];
  assign o[1941] = i[7];
  assign o[1942] = i[7];
  assign o[1943] = i[7];
  assign o[1944] = i[7];
  assign o[1945] = i[7];
  assign o[1946] = i[7];
  assign o[1947] = i[7];
  assign o[1948] = i[7];
  assign o[1949] = i[7];
  assign o[1950] = i[7];
  assign o[1951] = i[7];
  assign o[1952] = i[7];
  assign o[1953] = i[7];
  assign o[1954] = i[7];
  assign o[1955] = i[7];
  assign o[1956] = i[7];
  assign o[1957] = i[7];
  assign o[1958] = i[7];
  assign o[1959] = i[7];
  assign o[1960] = i[7];
  assign o[1961] = i[7];
  assign o[1962] = i[7];
  assign o[1963] = i[7];
  assign o[1964] = i[7];
  assign o[1965] = i[7];
  assign o[1966] = i[7];
  assign o[1967] = i[7];
  assign o[1968] = i[7];
  assign o[1969] = i[7];
  assign o[1970] = i[7];
  assign o[1971] = i[7];
  assign o[1972] = i[7];
  assign o[1973] = i[7];
  assign o[1974] = i[7];
  assign o[1975] = i[7];
  assign o[1976] = i[7];
  assign o[1977] = i[7];
  assign o[1978] = i[7];
  assign o[1979] = i[7];
  assign o[1980] = i[7];
  assign o[1981] = i[7];
  assign o[1982] = i[7];
  assign o[1983] = i[7];
  assign o[1984] = i[7];
  assign o[1985] = i[7];
  assign o[1986] = i[7];
  assign o[1987] = i[7];
  assign o[1988] = i[7];
  assign o[1989] = i[7];
  assign o[1990] = i[7];
  assign o[1991] = i[7];
  assign o[1992] = i[7];
  assign o[1993] = i[7];
  assign o[1994] = i[7];
  assign o[1995] = i[7];
  assign o[1996] = i[7];
  assign o[1997] = i[7];
  assign o[1998] = i[7];
  assign o[1999] = i[7];
  assign o[2000] = i[7];
  assign o[2001] = i[7];
  assign o[2002] = i[7];
  assign o[2003] = i[7];
  assign o[2004] = i[7];
  assign o[2005] = i[7];
  assign o[2006] = i[7];
  assign o[2007] = i[7];
  assign o[2008] = i[7];
  assign o[2009] = i[7];
  assign o[2010] = i[7];
  assign o[2011] = i[7];
  assign o[2012] = i[7];
  assign o[2013] = i[7];
  assign o[2014] = i[7];
  assign o[2015] = i[7];
  assign o[2016] = i[7];
  assign o[2017] = i[7];
  assign o[2018] = i[7];
  assign o[2019] = i[7];
  assign o[2020] = i[7];
  assign o[2021] = i[7];
  assign o[2022] = i[7];
  assign o[2023] = i[7];
  assign o[2024] = i[7];
  assign o[2025] = i[7];
  assign o[2026] = i[7];
  assign o[2027] = i[7];
  assign o[2028] = i[7];
  assign o[2029] = i[7];
  assign o[2030] = i[7];
  assign o[2031] = i[7];
  assign o[2032] = i[7];
  assign o[2033] = i[7];
  assign o[2034] = i[7];
  assign o[2035] = i[7];
  assign o[2036] = i[7];
  assign o[2037] = i[7];
  assign o[2038] = i[7];
  assign o[2039] = i[7];
  assign o[2040] = i[7];
  assign o[2041] = i[7];
  assign o[2042] = i[7];
  assign o[2043] = i[7];
  assign o[2044] = i[7];
  assign o[2045] = i[7];
  assign o[2046] = i[7];
  assign o[2047] = i[7];
  assign o[1536] = i[6];
  assign o[1537] = i[6];
  assign o[1538] = i[6];
  assign o[1539] = i[6];
  assign o[1540] = i[6];
  assign o[1541] = i[6];
  assign o[1542] = i[6];
  assign o[1543] = i[6];
  assign o[1544] = i[6];
  assign o[1545] = i[6];
  assign o[1546] = i[6];
  assign o[1547] = i[6];
  assign o[1548] = i[6];
  assign o[1549] = i[6];
  assign o[1550] = i[6];
  assign o[1551] = i[6];
  assign o[1552] = i[6];
  assign o[1553] = i[6];
  assign o[1554] = i[6];
  assign o[1555] = i[6];
  assign o[1556] = i[6];
  assign o[1557] = i[6];
  assign o[1558] = i[6];
  assign o[1559] = i[6];
  assign o[1560] = i[6];
  assign o[1561] = i[6];
  assign o[1562] = i[6];
  assign o[1563] = i[6];
  assign o[1564] = i[6];
  assign o[1565] = i[6];
  assign o[1566] = i[6];
  assign o[1567] = i[6];
  assign o[1568] = i[6];
  assign o[1569] = i[6];
  assign o[1570] = i[6];
  assign o[1571] = i[6];
  assign o[1572] = i[6];
  assign o[1573] = i[6];
  assign o[1574] = i[6];
  assign o[1575] = i[6];
  assign o[1576] = i[6];
  assign o[1577] = i[6];
  assign o[1578] = i[6];
  assign o[1579] = i[6];
  assign o[1580] = i[6];
  assign o[1581] = i[6];
  assign o[1582] = i[6];
  assign o[1583] = i[6];
  assign o[1584] = i[6];
  assign o[1585] = i[6];
  assign o[1586] = i[6];
  assign o[1587] = i[6];
  assign o[1588] = i[6];
  assign o[1589] = i[6];
  assign o[1590] = i[6];
  assign o[1591] = i[6];
  assign o[1592] = i[6];
  assign o[1593] = i[6];
  assign o[1594] = i[6];
  assign o[1595] = i[6];
  assign o[1596] = i[6];
  assign o[1597] = i[6];
  assign o[1598] = i[6];
  assign o[1599] = i[6];
  assign o[1600] = i[6];
  assign o[1601] = i[6];
  assign o[1602] = i[6];
  assign o[1603] = i[6];
  assign o[1604] = i[6];
  assign o[1605] = i[6];
  assign o[1606] = i[6];
  assign o[1607] = i[6];
  assign o[1608] = i[6];
  assign o[1609] = i[6];
  assign o[1610] = i[6];
  assign o[1611] = i[6];
  assign o[1612] = i[6];
  assign o[1613] = i[6];
  assign o[1614] = i[6];
  assign o[1615] = i[6];
  assign o[1616] = i[6];
  assign o[1617] = i[6];
  assign o[1618] = i[6];
  assign o[1619] = i[6];
  assign o[1620] = i[6];
  assign o[1621] = i[6];
  assign o[1622] = i[6];
  assign o[1623] = i[6];
  assign o[1624] = i[6];
  assign o[1625] = i[6];
  assign o[1626] = i[6];
  assign o[1627] = i[6];
  assign o[1628] = i[6];
  assign o[1629] = i[6];
  assign o[1630] = i[6];
  assign o[1631] = i[6];
  assign o[1632] = i[6];
  assign o[1633] = i[6];
  assign o[1634] = i[6];
  assign o[1635] = i[6];
  assign o[1636] = i[6];
  assign o[1637] = i[6];
  assign o[1638] = i[6];
  assign o[1639] = i[6];
  assign o[1640] = i[6];
  assign o[1641] = i[6];
  assign o[1642] = i[6];
  assign o[1643] = i[6];
  assign o[1644] = i[6];
  assign o[1645] = i[6];
  assign o[1646] = i[6];
  assign o[1647] = i[6];
  assign o[1648] = i[6];
  assign o[1649] = i[6];
  assign o[1650] = i[6];
  assign o[1651] = i[6];
  assign o[1652] = i[6];
  assign o[1653] = i[6];
  assign o[1654] = i[6];
  assign o[1655] = i[6];
  assign o[1656] = i[6];
  assign o[1657] = i[6];
  assign o[1658] = i[6];
  assign o[1659] = i[6];
  assign o[1660] = i[6];
  assign o[1661] = i[6];
  assign o[1662] = i[6];
  assign o[1663] = i[6];
  assign o[1664] = i[6];
  assign o[1665] = i[6];
  assign o[1666] = i[6];
  assign o[1667] = i[6];
  assign o[1668] = i[6];
  assign o[1669] = i[6];
  assign o[1670] = i[6];
  assign o[1671] = i[6];
  assign o[1672] = i[6];
  assign o[1673] = i[6];
  assign o[1674] = i[6];
  assign o[1675] = i[6];
  assign o[1676] = i[6];
  assign o[1677] = i[6];
  assign o[1678] = i[6];
  assign o[1679] = i[6];
  assign o[1680] = i[6];
  assign o[1681] = i[6];
  assign o[1682] = i[6];
  assign o[1683] = i[6];
  assign o[1684] = i[6];
  assign o[1685] = i[6];
  assign o[1686] = i[6];
  assign o[1687] = i[6];
  assign o[1688] = i[6];
  assign o[1689] = i[6];
  assign o[1690] = i[6];
  assign o[1691] = i[6];
  assign o[1692] = i[6];
  assign o[1693] = i[6];
  assign o[1694] = i[6];
  assign o[1695] = i[6];
  assign o[1696] = i[6];
  assign o[1697] = i[6];
  assign o[1698] = i[6];
  assign o[1699] = i[6];
  assign o[1700] = i[6];
  assign o[1701] = i[6];
  assign o[1702] = i[6];
  assign o[1703] = i[6];
  assign o[1704] = i[6];
  assign o[1705] = i[6];
  assign o[1706] = i[6];
  assign o[1707] = i[6];
  assign o[1708] = i[6];
  assign o[1709] = i[6];
  assign o[1710] = i[6];
  assign o[1711] = i[6];
  assign o[1712] = i[6];
  assign o[1713] = i[6];
  assign o[1714] = i[6];
  assign o[1715] = i[6];
  assign o[1716] = i[6];
  assign o[1717] = i[6];
  assign o[1718] = i[6];
  assign o[1719] = i[6];
  assign o[1720] = i[6];
  assign o[1721] = i[6];
  assign o[1722] = i[6];
  assign o[1723] = i[6];
  assign o[1724] = i[6];
  assign o[1725] = i[6];
  assign o[1726] = i[6];
  assign o[1727] = i[6];
  assign o[1728] = i[6];
  assign o[1729] = i[6];
  assign o[1730] = i[6];
  assign o[1731] = i[6];
  assign o[1732] = i[6];
  assign o[1733] = i[6];
  assign o[1734] = i[6];
  assign o[1735] = i[6];
  assign o[1736] = i[6];
  assign o[1737] = i[6];
  assign o[1738] = i[6];
  assign o[1739] = i[6];
  assign o[1740] = i[6];
  assign o[1741] = i[6];
  assign o[1742] = i[6];
  assign o[1743] = i[6];
  assign o[1744] = i[6];
  assign o[1745] = i[6];
  assign o[1746] = i[6];
  assign o[1747] = i[6];
  assign o[1748] = i[6];
  assign o[1749] = i[6];
  assign o[1750] = i[6];
  assign o[1751] = i[6];
  assign o[1752] = i[6];
  assign o[1753] = i[6];
  assign o[1754] = i[6];
  assign o[1755] = i[6];
  assign o[1756] = i[6];
  assign o[1757] = i[6];
  assign o[1758] = i[6];
  assign o[1759] = i[6];
  assign o[1760] = i[6];
  assign o[1761] = i[6];
  assign o[1762] = i[6];
  assign o[1763] = i[6];
  assign o[1764] = i[6];
  assign o[1765] = i[6];
  assign o[1766] = i[6];
  assign o[1767] = i[6];
  assign o[1768] = i[6];
  assign o[1769] = i[6];
  assign o[1770] = i[6];
  assign o[1771] = i[6];
  assign o[1772] = i[6];
  assign o[1773] = i[6];
  assign o[1774] = i[6];
  assign o[1775] = i[6];
  assign o[1776] = i[6];
  assign o[1777] = i[6];
  assign o[1778] = i[6];
  assign o[1779] = i[6];
  assign o[1780] = i[6];
  assign o[1781] = i[6];
  assign o[1782] = i[6];
  assign o[1783] = i[6];
  assign o[1784] = i[6];
  assign o[1785] = i[6];
  assign o[1786] = i[6];
  assign o[1787] = i[6];
  assign o[1788] = i[6];
  assign o[1789] = i[6];
  assign o[1790] = i[6];
  assign o[1791] = i[6];
  assign o[1280] = i[5];
  assign o[1281] = i[5];
  assign o[1282] = i[5];
  assign o[1283] = i[5];
  assign o[1284] = i[5];
  assign o[1285] = i[5];
  assign o[1286] = i[5];
  assign o[1287] = i[5];
  assign o[1288] = i[5];
  assign o[1289] = i[5];
  assign o[1290] = i[5];
  assign o[1291] = i[5];
  assign o[1292] = i[5];
  assign o[1293] = i[5];
  assign o[1294] = i[5];
  assign o[1295] = i[5];
  assign o[1296] = i[5];
  assign o[1297] = i[5];
  assign o[1298] = i[5];
  assign o[1299] = i[5];
  assign o[1300] = i[5];
  assign o[1301] = i[5];
  assign o[1302] = i[5];
  assign o[1303] = i[5];
  assign o[1304] = i[5];
  assign o[1305] = i[5];
  assign o[1306] = i[5];
  assign o[1307] = i[5];
  assign o[1308] = i[5];
  assign o[1309] = i[5];
  assign o[1310] = i[5];
  assign o[1311] = i[5];
  assign o[1312] = i[5];
  assign o[1313] = i[5];
  assign o[1314] = i[5];
  assign o[1315] = i[5];
  assign o[1316] = i[5];
  assign o[1317] = i[5];
  assign o[1318] = i[5];
  assign o[1319] = i[5];
  assign o[1320] = i[5];
  assign o[1321] = i[5];
  assign o[1322] = i[5];
  assign o[1323] = i[5];
  assign o[1324] = i[5];
  assign o[1325] = i[5];
  assign o[1326] = i[5];
  assign o[1327] = i[5];
  assign o[1328] = i[5];
  assign o[1329] = i[5];
  assign o[1330] = i[5];
  assign o[1331] = i[5];
  assign o[1332] = i[5];
  assign o[1333] = i[5];
  assign o[1334] = i[5];
  assign o[1335] = i[5];
  assign o[1336] = i[5];
  assign o[1337] = i[5];
  assign o[1338] = i[5];
  assign o[1339] = i[5];
  assign o[1340] = i[5];
  assign o[1341] = i[5];
  assign o[1342] = i[5];
  assign o[1343] = i[5];
  assign o[1344] = i[5];
  assign o[1345] = i[5];
  assign o[1346] = i[5];
  assign o[1347] = i[5];
  assign o[1348] = i[5];
  assign o[1349] = i[5];
  assign o[1350] = i[5];
  assign o[1351] = i[5];
  assign o[1352] = i[5];
  assign o[1353] = i[5];
  assign o[1354] = i[5];
  assign o[1355] = i[5];
  assign o[1356] = i[5];
  assign o[1357] = i[5];
  assign o[1358] = i[5];
  assign o[1359] = i[5];
  assign o[1360] = i[5];
  assign o[1361] = i[5];
  assign o[1362] = i[5];
  assign o[1363] = i[5];
  assign o[1364] = i[5];
  assign o[1365] = i[5];
  assign o[1366] = i[5];
  assign o[1367] = i[5];
  assign o[1368] = i[5];
  assign o[1369] = i[5];
  assign o[1370] = i[5];
  assign o[1371] = i[5];
  assign o[1372] = i[5];
  assign o[1373] = i[5];
  assign o[1374] = i[5];
  assign o[1375] = i[5];
  assign o[1376] = i[5];
  assign o[1377] = i[5];
  assign o[1378] = i[5];
  assign o[1379] = i[5];
  assign o[1380] = i[5];
  assign o[1381] = i[5];
  assign o[1382] = i[5];
  assign o[1383] = i[5];
  assign o[1384] = i[5];
  assign o[1385] = i[5];
  assign o[1386] = i[5];
  assign o[1387] = i[5];
  assign o[1388] = i[5];
  assign o[1389] = i[5];
  assign o[1390] = i[5];
  assign o[1391] = i[5];
  assign o[1392] = i[5];
  assign o[1393] = i[5];
  assign o[1394] = i[5];
  assign o[1395] = i[5];
  assign o[1396] = i[5];
  assign o[1397] = i[5];
  assign o[1398] = i[5];
  assign o[1399] = i[5];
  assign o[1400] = i[5];
  assign o[1401] = i[5];
  assign o[1402] = i[5];
  assign o[1403] = i[5];
  assign o[1404] = i[5];
  assign o[1405] = i[5];
  assign o[1406] = i[5];
  assign o[1407] = i[5];
  assign o[1408] = i[5];
  assign o[1409] = i[5];
  assign o[1410] = i[5];
  assign o[1411] = i[5];
  assign o[1412] = i[5];
  assign o[1413] = i[5];
  assign o[1414] = i[5];
  assign o[1415] = i[5];
  assign o[1416] = i[5];
  assign o[1417] = i[5];
  assign o[1418] = i[5];
  assign o[1419] = i[5];
  assign o[1420] = i[5];
  assign o[1421] = i[5];
  assign o[1422] = i[5];
  assign o[1423] = i[5];
  assign o[1424] = i[5];
  assign o[1425] = i[5];
  assign o[1426] = i[5];
  assign o[1427] = i[5];
  assign o[1428] = i[5];
  assign o[1429] = i[5];
  assign o[1430] = i[5];
  assign o[1431] = i[5];
  assign o[1432] = i[5];
  assign o[1433] = i[5];
  assign o[1434] = i[5];
  assign o[1435] = i[5];
  assign o[1436] = i[5];
  assign o[1437] = i[5];
  assign o[1438] = i[5];
  assign o[1439] = i[5];
  assign o[1440] = i[5];
  assign o[1441] = i[5];
  assign o[1442] = i[5];
  assign o[1443] = i[5];
  assign o[1444] = i[5];
  assign o[1445] = i[5];
  assign o[1446] = i[5];
  assign o[1447] = i[5];
  assign o[1448] = i[5];
  assign o[1449] = i[5];
  assign o[1450] = i[5];
  assign o[1451] = i[5];
  assign o[1452] = i[5];
  assign o[1453] = i[5];
  assign o[1454] = i[5];
  assign o[1455] = i[5];
  assign o[1456] = i[5];
  assign o[1457] = i[5];
  assign o[1458] = i[5];
  assign o[1459] = i[5];
  assign o[1460] = i[5];
  assign o[1461] = i[5];
  assign o[1462] = i[5];
  assign o[1463] = i[5];
  assign o[1464] = i[5];
  assign o[1465] = i[5];
  assign o[1466] = i[5];
  assign o[1467] = i[5];
  assign o[1468] = i[5];
  assign o[1469] = i[5];
  assign o[1470] = i[5];
  assign o[1471] = i[5];
  assign o[1472] = i[5];
  assign o[1473] = i[5];
  assign o[1474] = i[5];
  assign o[1475] = i[5];
  assign o[1476] = i[5];
  assign o[1477] = i[5];
  assign o[1478] = i[5];
  assign o[1479] = i[5];
  assign o[1480] = i[5];
  assign o[1481] = i[5];
  assign o[1482] = i[5];
  assign o[1483] = i[5];
  assign o[1484] = i[5];
  assign o[1485] = i[5];
  assign o[1486] = i[5];
  assign o[1487] = i[5];
  assign o[1488] = i[5];
  assign o[1489] = i[5];
  assign o[1490] = i[5];
  assign o[1491] = i[5];
  assign o[1492] = i[5];
  assign o[1493] = i[5];
  assign o[1494] = i[5];
  assign o[1495] = i[5];
  assign o[1496] = i[5];
  assign o[1497] = i[5];
  assign o[1498] = i[5];
  assign o[1499] = i[5];
  assign o[1500] = i[5];
  assign o[1501] = i[5];
  assign o[1502] = i[5];
  assign o[1503] = i[5];
  assign o[1504] = i[5];
  assign o[1505] = i[5];
  assign o[1506] = i[5];
  assign o[1507] = i[5];
  assign o[1508] = i[5];
  assign o[1509] = i[5];
  assign o[1510] = i[5];
  assign o[1511] = i[5];
  assign o[1512] = i[5];
  assign o[1513] = i[5];
  assign o[1514] = i[5];
  assign o[1515] = i[5];
  assign o[1516] = i[5];
  assign o[1517] = i[5];
  assign o[1518] = i[5];
  assign o[1519] = i[5];
  assign o[1520] = i[5];
  assign o[1521] = i[5];
  assign o[1522] = i[5];
  assign o[1523] = i[5];
  assign o[1524] = i[5];
  assign o[1525] = i[5];
  assign o[1526] = i[5];
  assign o[1527] = i[5];
  assign o[1528] = i[5];
  assign o[1529] = i[5];
  assign o[1530] = i[5];
  assign o[1531] = i[5];
  assign o[1532] = i[5];
  assign o[1533] = i[5];
  assign o[1534] = i[5];
  assign o[1535] = i[5];
  assign o[1024] = i[4];
  assign o[1025] = i[4];
  assign o[1026] = i[4];
  assign o[1027] = i[4];
  assign o[1028] = i[4];
  assign o[1029] = i[4];
  assign o[1030] = i[4];
  assign o[1031] = i[4];
  assign o[1032] = i[4];
  assign o[1033] = i[4];
  assign o[1034] = i[4];
  assign o[1035] = i[4];
  assign o[1036] = i[4];
  assign o[1037] = i[4];
  assign o[1038] = i[4];
  assign o[1039] = i[4];
  assign o[1040] = i[4];
  assign o[1041] = i[4];
  assign o[1042] = i[4];
  assign o[1043] = i[4];
  assign o[1044] = i[4];
  assign o[1045] = i[4];
  assign o[1046] = i[4];
  assign o[1047] = i[4];
  assign o[1048] = i[4];
  assign o[1049] = i[4];
  assign o[1050] = i[4];
  assign o[1051] = i[4];
  assign o[1052] = i[4];
  assign o[1053] = i[4];
  assign o[1054] = i[4];
  assign o[1055] = i[4];
  assign o[1056] = i[4];
  assign o[1057] = i[4];
  assign o[1058] = i[4];
  assign o[1059] = i[4];
  assign o[1060] = i[4];
  assign o[1061] = i[4];
  assign o[1062] = i[4];
  assign o[1063] = i[4];
  assign o[1064] = i[4];
  assign o[1065] = i[4];
  assign o[1066] = i[4];
  assign o[1067] = i[4];
  assign o[1068] = i[4];
  assign o[1069] = i[4];
  assign o[1070] = i[4];
  assign o[1071] = i[4];
  assign o[1072] = i[4];
  assign o[1073] = i[4];
  assign o[1074] = i[4];
  assign o[1075] = i[4];
  assign o[1076] = i[4];
  assign o[1077] = i[4];
  assign o[1078] = i[4];
  assign o[1079] = i[4];
  assign o[1080] = i[4];
  assign o[1081] = i[4];
  assign o[1082] = i[4];
  assign o[1083] = i[4];
  assign o[1084] = i[4];
  assign o[1085] = i[4];
  assign o[1086] = i[4];
  assign o[1087] = i[4];
  assign o[1088] = i[4];
  assign o[1089] = i[4];
  assign o[1090] = i[4];
  assign o[1091] = i[4];
  assign o[1092] = i[4];
  assign o[1093] = i[4];
  assign o[1094] = i[4];
  assign o[1095] = i[4];
  assign o[1096] = i[4];
  assign o[1097] = i[4];
  assign o[1098] = i[4];
  assign o[1099] = i[4];
  assign o[1100] = i[4];
  assign o[1101] = i[4];
  assign o[1102] = i[4];
  assign o[1103] = i[4];
  assign o[1104] = i[4];
  assign o[1105] = i[4];
  assign o[1106] = i[4];
  assign o[1107] = i[4];
  assign o[1108] = i[4];
  assign o[1109] = i[4];
  assign o[1110] = i[4];
  assign o[1111] = i[4];
  assign o[1112] = i[4];
  assign o[1113] = i[4];
  assign o[1114] = i[4];
  assign o[1115] = i[4];
  assign o[1116] = i[4];
  assign o[1117] = i[4];
  assign o[1118] = i[4];
  assign o[1119] = i[4];
  assign o[1120] = i[4];
  assign o[1121] = i[4];
  assign o[1122] = i[4];
  assign o[1123] = i[4];
  assign o[1124] = i[4];
  assign o[1125] = i[4];
  assign o[1126] = i[4];
  assign o[1127] = i[4];
  assign o[1128] = i[4];
  assign o[1129] = i[4];
  assign o[1130] = i[4];
  assign o[1131] = i[4];
  assign o[1132] = i[4];
  assign o[1133] = i[4];
  assign o[1134] = i[4];
  assign o[1135] = i[4];
  assign o[1136] = i[4];
  assign o[1137] = i[4];
  assign o[1138] = i[4];
  assign o[1139] = i[4];
  assign o[1140] = i[4];
  assign o[1141] = i[4];
  assign o[1142] = i[4];
  assign o[1143] = i[4];
  assign o[1144] = i[4];
  assign o[1145] = i[4];
  assign o[1146] = i[4];
  assign o[1147] = i[4];
  assign o[1148] = i[4];
  assign o[1149] = i[4];
  assign o[1150] = i[4];
  assign o[1151] = i[4];
  assign o[1152] = i[4];
  assign o[1153] = i[4];
  assign o[1154] = i[4];
  assign o[1155] = i[4];
  assign o[1156] = i[4];
  assign o[1157] = i[4];
  assign o[1158] = i[4];
  assign o[1159] = i[4];
  assign o[1160] = i[4];
  assign o[1161] = i[4];
  assign o[1162] = i[4];
  assign o[1163] = i[4];
  assign o[1164] = i[4];
  assign o[1165] = i[4];
  assign o[1166] = i[4];
  assign o[1167] = i[4];
  assign o[1168] = i[4];
  assign o[1169] = i[4];
  assign o[1170] = i[4];
  assign o[1171] = i[4];
  assign o[1172] = i[4];
  assign o[1173] = i[4];
  assign o[1174] = i[4];
  assign o[1175] = i[4];
  assign o[1176] = i[4];
  assign o[1177] = i[4];
  assign o[1178] = i[4];
  assign o[1179] = i[4];
  assign o[1180] = i[4];
  assign o[1181] = i[4];
  assign o[1182] = i[4];
  assign o[1183] = i[4];
  assign o[1184] = i[4];
  assign o[1185] = i[4];
  assign o[1186] = i[4];
  assign o[1187] = i[4];
  assign o[1188] = i[4];
  assign o[1189] = i[4];
  assign o[1190] = i[4];
  assign o[1191] = i[4];
  assign o[1192] = i[4];
  assign o[1193] = i[4];
  assign o[1194] = i[4];
  assign o[1195] = i[4];
  assign o[1196] = i[4];
  assign o[1197] = i[4];
  assign o[1198] = i[4];
  assign o[1199] = i[4];
  assign o[1200] = i[4];
  assign o[1201] = i[4];
  assign o[1202] = i[4];
  assign o[1203] = i[4];
  assign o[1204] = i[4];
  assign o[1205] = i[4];
  assign o[1206] = i[4];
  assign o[1207] = i[4];
  assign o[1208] = i[4];
  assign o[1209] = i[4];
  assign o[1210] = i[4];
  assign o[1211] = i[4];
  assign o[1212] = i[4];
  assign o[1213] = i[4];
  assign o[1214] = i[4];
  assign o[1215] = i[4];
  assign o[1216] = i[4];
  assign o[1217] = i[4];
  assign o[1218] = i[4];
  assign o[1219] = i[4];
  assign o[1220] = i[4];
  assign o[1221] = i[4];
  assign o[1222] = i[4];
  assign o[1223] = i[4];
  assign o[1224] = i[4];
  assign o[1225] = i[4];
  assign o[1226] = i[4];
  assign o[1227] = i[4];
  assign o[1228] = i[4];
  assign o[1229] = i[4];
  assign o[1230] = i[4];
  assign o[1231] = i[4];
  assign o[1232] = i[4];
  assign o[1233] = i[4];
  assign o[1234] = i[4];
  assign o[1235] = i[4];
  assign o[1236] = i[4];
  assign o[1237] = i[4];
  assign o[1238] = i[4];
  assign o[1239] = i[4];
  assign o[1240] = i[4];
  assign o[1241] = i[4];
  assign o[1242] = i[4];
  assign o[1243] = i[4];
  assign o[1244] = i[4];
  assign o[1245] = i[4];
  assign o[1246] = i[4];
  assign o[1247] = i[4];
  assign o[1248] = i[4];
  assign o[1249] = i[4];
  assign o[1250] = i[4];
  assign o[1251] = i[4];
  assign o[1252] = i[4];
  assign o[1253] = i[4];
  assign o[1254] = i[4];
  assign o[1255] = i[4];
  assign o[1256] = i[4];
  assign o[1257] = i[4];
  assign o[1258] = i[4];
  assign o[1259] = i[4];
  assign o[1260] = i[4];
  assign o[1261] = i[4];
  assign o[1262] = i[4];
  assign o[1263] = i[4];
  assign o[1264] = i[4];
  assign o[1265] = i[4];
  assign o[1266] = i[4];
  assign o[1267] = i[4];
  assign o[1268] = i[4];
  assign o[1269] = i[4];
  assign o[1270] = i[4];
  assign o[1271] = i[4];
  assign o[1272] = i[4];
  assign o[1273] = i[4];
  assign o[1274] = i[4];
  assign o[1275] = i[4];
  assign o[1276] = i[4];
  assign o[1277] = i[4];
  assign o[1278] = i[4];
  assign o[1279] = i[4];
  assign o[768] = i[3];
  assign o[769] = i[3];
  assign o[770] = i[3];
  assign o[771] = i[3];
  assign o[772] = i[3];
  assign o[773] = i[3];
  assign o[774] = i[3];
  assign o[775] = i[3];
  assign o[776] = i[3];
  assign o[777] = i[3];
  assign o[778] = i[3];
  assign o[779] = i[3];
  assign o[780] = i[3];
  assign o[781] = i[3];
  assign o[782] = i[3];
  assign o[783] = i[3];
  assign o[784] = i[3];
  assign o[785] = i[3];
  assign o[786] = i[3];
  assign o[787] = i[3];
  assign o[788] = i[3];
  assign o[789] = i[3];
  assign o[790] = i[3];
  assign o[791] = i[3];
  assign o[792] = i[3];
  assign o[793] = i[3];
  assign o[794] = i[3];
  assign o[795] = i[3];
  assign o[796] = i[3];
  assign o[797] = i[3];
  assign o[798] = i[3];
  assign o[799] = i[3];
  assign o[800] = i[3];
  assign o[801] = i[3];
  assign o[802] = i[3];
  assign o[803] = i[3];
  assign o[804] = i[3];
  assign o[805] = i[3];
  assign o[806] = i[3];
  assign o[807] = i[3];
  assign o[808] = i[3];
  assign o[809] = i[3];
  assign o[810] = i[3];
  assign o[811] = i[3];
  assign o[812] = i[3];
  assign o[813] = i[3];
  assign o[814] = i[3];
  assign o[815] = i[3];
  assign o[816] = i[3];
  assign o[817] = i[3];
  assign o[818] = i[3];
  assign o[819] = i[3];
  assign o[820] = i[3];
  assign o[821] = i[3];
  assign o[822] = i[3];
  assign o[823] = i[3];
  assign o[824] = i[3];
  assign o[825] = i[3];
  assign o[826] = i[3];
  assign o[827] = i[3];
  assign o[828] = i[3];
  assign o[829] = i[3];
  assign o[830] = i[3];
  assign o[831] = i[3];
  assign o[832] = i[3];
  assign o[833] = i[3];
  assign o[834] = i[3];
  assign o[835] = i[3];
  assign o[836] = i[3];
  assign o[837] = i[3];
  assign o[838] = i[3];
  assign o[839] = i[3];
  assign o[840] = i[3];
  assign o[841] = i[3];
  assign o[842] = i[3];
  assign o[843] = i[3];
  assign o[844] = i[3];
  assign o[845] = i[3];
  assign o[846] = i[3];
  assign o[847] = i[3];
  assign o[848] = i[3];
  assign o[849] = i[3];
  assign o[850] = i[3];
  assign o[851] = i[3];
  assign o[852] = i[3];
  assign o[853] = i[3];
  assign o[854] = i[3];
  assign o[855] = i[3];
  assign o[856] = i[3];
  assign o[857] = i[3];
  assign o[858] = i[3];
  assign o[859] = i[3];
  assign o[860] = i[3];
  assign o[861] = i[3];
  assign o[862] = i[3];
  assign o[863] = i[3];
  assign o[864] = i[3];
  assign o[865] = i[3];
  assign o[866] = i[3];
  assign o[867] = i[3];
  assign o[868] = i[3];
  assign o[869] = i[3];
  assign o[870] = i[3];
  assign o[871] = i[3];
  assign o[872] = i[3];
  assign o[873] = i[3];
  assign o[874] = i[3];
  assign o[875] = i[3];
  assign o[876] = i[3];
  assign o[877] = i[3];
  assign o[878] = i[3];
  assign o[879] = i[3];
  assign o[880] = i[3];
  assign o[881] = i[3];
  assign o[882] = i[3];
  assign o[883] = i[3];
  assign o[884] = i[3];
  assign o[885] = i[3];
  assign o[886] = i[3];
  assign o[887] = i[3];
  assign o[888] = i[3];
  assign o[889] = i[3];
  assign o[890] = i[3];
  assign o[891] = i[3];
  assign o[892] = i[3];
  assign o[893] = i[3];
  assign o[894] = i[3];
  assign o[895] = i[3];
  assign o[896] = i[3];
  assign o[897] = i[3];
  assign o[898] = i[3];
  assign o[899] = i[3];
  assign o[900] = i[3];
  assign o[901] = i[3];
  assign o[902] = i[3];
  assign o[903] = i[3];
  assign o[904] = i[3];
  assign o[905] = i[3];
  assign o[906] = i[3];
  assign o[907] = i[3];
  assign o[908] = i[3];
  assign o[909] = i[3];
  assign o[910] = i[3];
  assign o[911] = i[3];
  assign o[912] = i[3];
  assign o[913] = i[3];
  assign o[914] = i[3];
  assign o[915] = i[3];
  assign o[916] = i[3];
  assign o[917] = i[3];
  assign o[918] = i[3];
  assign o[919] = i[3];
  assign o[920] = i[3];
  assign o[921] = i[3];
  assign o[922] = i[3];
  assign o[923] = i[3];
  assign o[924] = i[3];
  assign o[925] = i[3];
  assign o[926] = i[3];
  assign o[927] = i[3];
  assign o[928] = i[3];
  assign o[929] = i[3];
  assign o[930] = i[3];
  assign o[931] = i[3];
  assign o[932] = i[3];
  assign o[933] = i[3];
  assign o[934] = i[3];
  assign o[935] = i[3];
  assign o[936] = i[3];
  assign o[937] = i[3];
  assign o[938] = i[3];
  assign o[939] = i[3];
  assign o[940] = i[3];
  assign o[941] = i[3];
  assign o[942] = i[3];
  assign o[943] = i[3];
  assign o[944] = i[3];
  assign o[945] = i[3];
  assign o[946] = i[3];
  assign o[947] = i[3];
  assign o[948] = i[3];
  assign o[949] = i[3];
  assign o[950] = i[3];
  assign o[951] = i[3];
  assign o[952] = i[3];
  assign o[953] = i[3];
  assign o[954] = i[3];
  assign o[955] = i[3];
  assign o[956] = i[3];
  assign o[957] = i[3];
  assign o[958] = i[3];
  assign o[959] = i[3];
  assign o[960] = i[3];
  assign o[961] = i[3];
  assign o[962] = i[3];
  assign o[963] = i[3];
  assign o[964] = i[3];
  assign o[965] = i[3];
  assign o[966] = i[3];
  assign o[967] = i[3];
  assign o[968] = i[3];
  assign o[969] = i[3];
  assign o[970] = i[3];
  assign o[971] = i[3];
  assign o[972] = i[3];
  assign o[973] = i[3];
  assign o[974] = i[3];
  assign o[975] = i[3];
  assign o[976] = i[3];
  assign o[977] = i[3];
  assign o[978] = i[3];
  assign o[979] = i[3];
  assign o[980] = i[3];
  assign o[981] = i[3];
  assign o[982] = i[3];
  assign o[983] = i[3];
  assign o[984] = i[3];
  assign o[985] = i[3];
  assign o[986] = i[3];
  assign o[987] = i[3];
  assign o[988] = i[3];
  assign o[989] = i[3];
  assign o[990] = i[3];
  assign o[991] = i[3];
  assign o[992] = i[3];
  assign o[993] = i[3];
  assign o[994] = i[3];
  assign o[995] = i[3];
  assign o[996] = i[3];
  assign o[997] = i[3];
  assign o[998] = i[3];
  assign o[999] = i[3];
  assign o[1000] = i[3];
  assign o[1001] = i[3];
  assign o[1002] = i[3];
  assign o[1003] = i[3];
  assign o[1004] = i[3];
  assign o[1005] = i[3];
  assign o[1006] = i[3];
  assign o[1007] = i[3];
  assign o[1008] = i[3];
  assign o[1009] = i[3];
  assign o[1010] = i[3];
  assign o[1011] = i[3];
  assign o[1012] = i[3];
  assign o[1013] = i[3];
  assign o[1014] = i[3];
  assign o[1015] = i[3];
  assign o[1016] = i[3];
  assign o[1017] = i[3];
  assign o[1018] = i[3];
  assign o[1019] = i[3];
  assign o[1020] = i[3];
  assign o[1021] = i[3];
  assign o[1022] = i[3];
  assign o[1023] = i[3];
  assign o[512] = i[2];
  assign o[513] = i[2];
  assign o[514] = i[2];
  assign o[515] = i[2];
  assign o[516] = i[2];
  assign o[517] = i[2];
  assign o[518] = i[2];
  assign o[519] = i[2];
  assign o[520] = i[2];
  assign o[521] = i[2];
  assign o[522] = i[2];
  assign o[523] = i[2];
  assign o[524] = i[2];
  assign o[525] = i[2];
  assign o[526] = i[2];
  assign o[527] = i[2];
  assign o[528] = i[2];
  assign o[529] = i[2];
  assign o[530] = i[2];
  assign o[531] = i[2];
  assign o[532] = i[2];
  assign o[533] = i[2];
  assign o[534] = i[2];
  assign o[535] = i[2];
  assign o[536] = i[2];
  assign o[537] = i[2];
  assign o[538] = i[2];
  assign o[539] = i[2];
  assign o[540] = i[2];
  assign o[541] = i[2];
  assign o[542] = i[2];
  assign o[543] = i[2];
  assign o[544] = i[2];
  assign o[545] = i[2];
  assign o[546] = i[2];
  assign o[547] = i[2];
  assign o[548] = i[2];
  assign o[549] = i[2];
  assign o[550] = i[2];
  assign o[551] = i[2];
  assign o[552] = i[2];
  assign o[553] = i[2];
  assign o[554] = i[2];
  assign o[555] = i[2];
  assign o[556] = i[2];
  assign o[557] = i[2];
  assign o[558] = i[2];
  assign o[559] = i[2];
  assign o[560] = i[2];
  assign o[561] = i[2];
  assign o[562] = i[2];
  assign o[563] = i[2];
  assign o[564] = i[2];
  assign o[565] = i[2];
  assign o[566] = i[2];
  assign o[567] = i[2];
  assign o[568] = i[2];
  assign o[569] = i[2];
  assign o[570] = i[2];
  assign o[571] = i[2];
  assign o[572] = i[2];
  assign o[573] = i[2];
  assign o[574] = i[2];
  assign o[575] = i[2];
  assign o[576] = i[2];
  assign o[577] = i[2];
  assign o[578] = i[2];
  assign o[579] = i[2];
  assign o[580] = i[2];
  assign o[581] = i[2];
  assign o[582] = i[2];
  assign o[583] = i[2];
  assign o[584] = i[2];
  assign o[585] = i[2];
  assign o[586] = i[2];
  assign o[587] = i[2];
  assign o[588] = i[2];
  assign o[589] = i[2];
  assign o[590] = i[2];
  assign o[591] = i[2];
  assign o[592] = i[2];
  assign o[593] = i[2];
  assign o[594] = i[2];
  assign o[595] = i[2];
  assign o[596] = i[2];
  assign o[597] = i[2];
  assign o[598] = i[2];
  assign o[599] = i[2];
  assign o[600] = i[2];
  assign o[601] = i[2];
  assign o[602] = i[2];
  assign o[603] = i[2];
  assign o[604] = i[2];
  assign o[605] = i[2];
  assign o[606] = i[2];
  assign o[607] = i[2];
  assign o[608] = i[2];
  assign o[609] = i[2];
  assign o[610] = i[2];
  assign o[611] = i[2];
  assign o[612] = i[2];
  assign o[613] = i[2];
  assign o[614] = i[2];
  assign o[615] = i[2];
  assign o[616] = i[2];
  assign o[617] = i[2];
  assign o[618] = i[2];
  assign o[619] = i[2];
  assign o[620] = i[2];
  assign o[621] = i[2];
  assign o[622] = i[2];
  assign o[623] = i[2];
  assign o[624] = i[2];
  assign o[625] = i[2];
  assign o[626] = i[2];
  assign o[627] = i[2];
  assign o[628] = i[2];
  assign o[629] = i[2];
  assign o[630] = i[2];
  assign o[631] = i[2];
  assign o[632] = i[2];
  assign o[633] = i[2];
  assign o[634] = i[2];
  assign o[635] = i[2];
  assign o[636] = i[2];
  assign o[637] = i[2];
  assign o[638] = i[2];
  assign o[639] = i[2];
  assign o[640] = i[2];
  assign o[641] = i[2];
  assign o[642] = i[2];
  assign o[643] = i[2];
  assign o[644] = i[2];
  assign o[645] = i[2];
  assign o[646] = i[2];
  assign o[647] = i[2];
  assign o[648] = i[2];
  assign o[649] = i[2];
  assign o[650] = i[2];
  assign o[651] = i[2];
  assign o[652] = i[2];
  assign o[653] = i[2];
  assign o[654] = i[2];
  assign o[655] = i[2];
  assign o[656] = i[2];
  assign o[657] = i[2];
  assign o[658] = i[2];
  assign o[659] = i[2];
  assign o[660] = i[2];
  assign o[661] = i[2];
  assign o[662] = i[2];
  assign o[663] = i[2];
  assign o[664] = i[2];
  assign o[665] = i[2];
  assign o[666] = i[2];
  assign o[667] = i[2];
  assign o[668] = i[2];
  assign o[669] = i[2];
  assign o[670] = i[2];
  assign o[671] = i[2];
  assign o[672] = i[2];
  assign o[673] = i[2];
  assign o[674] = i[2];
  assign o[675] = i[2];
  assign o[676] = i[2];
  assign o[677] = i[2];
  assign o[678] = i[2];
  assign o[679] = i[2];
  assign o[680] = i[2];
  assign o[681] = i[2];
  assign o[682] = i[2];
  assign o[683] = i[2];
  assign o[684] = i[2];
  assign o[685] = i[2];
  assign o[686] = i[2];
  assign o[687] = i[2];
  assign o[688] = i[2];
  assign o[689] = i[2];
  assign o[690] = i[2];
  assign o[691] = i[2];
  assign o[692] = i[2];
  assign o[693] = i[2];
  assign o[694] = i[2];
  assign o[695] = i[2];
  assign o[696] = i[2];
  assign o[697] = i[2];
  assign o[698] = i[2];
  assign o[699] = i[2];
  assign o[700] = i[2];
  assign o[701] = i[2];
  assign o[702] = i[2];
  assign o[703] = i[2];
  assign o[704] = i[2];
  assign o[705] = i[2];
  assign o[706] = i[2];
  assign o[707] = i[2];
  assign o[708] = i[2];
  assign o[709] = i[2];
  assign o[710] = i[2];
  assign o[711] = i[2];
  assign o[712] = i[2];
  assign o[713] = i[2];
  assign o[714] = i[2];
  assign o[715] = i[2];
  assign o[716] = i[2];
  assign o[717] = i[2];
  assign o[718] = i[2];
  assign o[719] = i[2];
  assign o[720] = i[2];
  assign o[721] = i[2];
  assign o[722] = i[2];
  assign o[723] = i[2];
  assign o[724] = i[2];
  assign o[725] = i[2];
  assign o[726] = i[2];
  assign o[727] = i[2];
  assign o[728] = i[2];
  assign o[729] = i[2];
  assign o[730] = i[2];
  assign o[731] = i[2];
  assign o[732] = i[2];
  assign o[733] = i[2];
  assign o[734] = i[2];
  assign o[735] = i[2];
  assign o[736] = i[2];
  assign o[737] = i[2];
  assign o[738] = i[2];
  assign o[739] = i[2];
  assign o[740] = i[2];
  assign o[741] = i[2];
  assign o[742] = i[2];
  assign o[743] = i[2];
  assign o[744] = i[2];
  assign o[745] = i[2];
  assign o[746] = i[2];
  assign o[747] = i[2];
  assign o[748] = i[2];
  assign o[749] = i[2];
  assign o[750] = i[2];
  assign o[751] = i[2];
  assign o[752] = i[2];
  assign o[753] = i[2];
  assign o[754] = i[2];
  assign o[755] = i[2];
  assign o[756] = i[2];
  assign o[757] = i[2];
  assign o[758] = i[2];
  assign o[759] = i[2];
  assign o[760] = i[2];
  assign o[761] = i[2];
  assign o[762] = i[2];
  assign o[763] = i[2];
  assign o[764] = i[2];
  assign o[765] = i[2];
  assign o[766] = i[2];
  assign o[767] = i[2];
  assign o[256] = i[1];
  assign o[257] = i[1];
  assign o[258] = i[1];
  assign o[259] = i[1];
  assign o[260] = i[1];
  assign o[261] = i[1];
  assign o[262] = i[1];
  assign o[263] = i[1];
  assign o[264] = i[1];
  assign o[265] = i[1];
  assign o[266] = i[1];
  assign o[267] = i[1];
  assign o[268] = i[1];
  assign o[269] = i[1];
  assign o[270] = i[1];
  assign o[271] = i[1];
  assign o[272] = i[1];
  assign o[273] = i[1];
  assign o[274] = i[1];
  assign o[275] = i[1];
  assign o[276] = i[1];
  assign o[277] = i[1];
  assign o[278] = i[1];
  assign o[279] = i[1];
  assign o[280] = i[1];
  assign o[281] = i[1];
  assign o[282] = i[1];
  assign o[283] = i[1];
  assign o[284] = i[1];
  assign o[285] = i[1];
  assign o[286] = i[1];
  assign o[287] = i[1];
  assign o[288] = i[1];
  assign o[289] = i[1];
  assign o[290] = i[1];
  assign o[291] = i[1];
  assign o[292] = i[1];
  assign o[293] = i[1];
  assign o[294] = i[1];
  assign o[295] = i[1];
  assign o[296] = i[1];
  assign o[297] = i[1];
  assign o[298] = i[1];
  assign o[299] = i[1];
  assign o[300] = i[1];
  assign o[301] = i[1];
  assign o[302] = i[1];
  assign o[303] = i[1];
  assign o[304] = i[1];
  assign o[305] = i[1];
  assign o[306] = i[1];
  assign o[307] = i[1];
  assign o[308] = i[1];
  assign o[309] = i[1];
  assign o[310] = i[1];
  assign o[311] = i[1];
  assign o[312] = i[1];
  assign o[313] = i[1];
  assign o[314] = i[1];
  assign o[315] = i[1];
  assign o[316] = i[1];
  assign o[317] = i[1];
  assign o[318] = i[1];
  assign o[319] = i[1];
  assign o[320] = i[1];
  assign o[321] = i[1];
  assign o[322] = i[1];
  assign o[323] = i[1];
  assign o[324] = i[1];
  assign o[325] = i[1];
  assign o[326] = i[1];
  assign o[327] = i[1];
  assign o[328] = i[1];
  assign o[329] = i[1];
  assign o[330] = i[1];
  assign o[331] = i[1];
  assign o[332] = i[1];
  assign o[333] = i[1];
  assign o[334] = i[1];
  assign o[335] = i[1];
  assign o[336] = i[1];
  assign o[337] = i[1];
  assign o[338] = i[1];
  assign o[339] = i[1];
  assign o[340] = i[1];
  assign o[341] = i[1];
  assign o[342] = i[1];
  assign o[343] = i[1];
  assign o[344] = i[1];
  assign o[345] = i[1];
  assign o[346] = i[1];
  assign o[347] = i[1];
  assign o[348] = i[1];
  assign o[349] = i[1];
  assign o[350] = i[1];
  assign o[351] = i[1];
  assign o[352] = i[1];
  assign o[353] = i[1];
  assign o[354] = i[1];
  assign o[355] = i[1];
  assign o[356] = i[1];
  assign o[357] = i[1];
  assign o[358] = i[1];
  assign o[359] = i[1];
  assign o[360] = i[1];
  assign o[361] = i[1];
  assign o[362] = i[1];
  assign o[363] = i[1];
  assign o[364] = i[1];
  assign o[365] = i[1];
  assign o[366] = i[1];
  assign o[367] = i[1];
  assign o[368] = i[1];
  assign o[369] = i[1];
  assign o[370] = i[1];
  assign o[371] = i[1];
  assign o[372] = i[1];
  assign o[373] = i[1];
  assign o[374] = i[1];
  assign o[375] = i[1];
  assign o[376] = i[1];
  assign o[377] = i[1];
  assign o[378] = i[1];
  assign o[379] = i[1];
  assign o[380] = i[1];
  assign o[381] = i[1];
  assign o[382] = i[1];
  assign o[383] = i[1];
  assign o[384] = i[1];
  assign o[385] = i[1];
  assign o[386] = i[1];
  assign o[387] = i[1];
  assign o[388] = i[1];
  assign o[389] = i[1];
  assign o[390] = i[1];
  assign o[391] = i[1];
  assign o[392] = i[1];
  assign o[393] = i[1];
  assign o[394] = i[1];
  assign o[395] = i[1];
  assign o[396] = i[1];
  assign o[397] = i[1];
  assign o[398] = i[1];
  assign o[399] = i[1];
  assign o[400] = i[1];
  assign o[401] = i[1];
  assign o[402] = i[1];
  assign o[403] = i[1];
  assign o[404] = i[1];
  assign o[405] = i[1];
  assign o[406] = i[1];
  assign o[407] = i[1];
  assign o[408] = i[1];
  assign o[409] = i[1];
  assign o[410] = i[1];
  assign o[411] = i[1];
  assign o[412] = i[1];
  assign o[413] = i[1];
  assign o[414] = i[1];
  assign o[415] = i[1];
  assign o[416] = i[1];
  assign o[417] = i[1];
  assign o[418] = i[1];
  assign o[419] = i[1];
  assign o[420] = i[1];
  assign o[421] = i[1];
  assign o[422] = i[1];
  assign o[423] = i[1];
  assign o[424] = i[1];
  assign o[425] = i[1];
  assign o[426] = i[1];
  assign o[427] = i[1];
  assign o[428] = i[1];
  assign o[429] = i[1];
  assign o[430] = i[1];
  assign o[431] = i[1];
  assign o[432] = i[1];
  assign o[433] = i[1];
  assign o[434] = i[1];
  assign o[435] = i[1];
  assign o[436] = i[1];
  assign o[437] = i[1];
  assign o[438] = i[1];
  assign o[439] = i[1];
  assign o[440] = i[1];
  assign o[441] = i[1];
  assign o[442] = i[1];
  assign o[443] = i[1];
  assign o[444] = i[1];
  assign o[445] = i[1];
  assign o[446] = i[1];
  assign o[447] = i[1];
  assign o[448] = i[1];
  assign o[449] = i[1];
  assign o[450] = i[1];
  assign o[451] = i[1];
  assign o[452] = i[1];
  assign o[453] = i[1];
  assign o[454] = i[1];
  assign o[455] = i[1];
  assign o[456] = i[1];
  assign o[457] = i[1];
  assign o[458] = i[1];
  assign o[459] = i[1];
  assign o[460] = i[1];
  assign o[461] = i[1];
  assign o[462] = i[1];
  assign o[463] = i[1];
  assign o[464] = i[1];
  assign o[465] = i[1];
  assign o[466] = i[1];
  assign o[467] = i[1];
  assign o[468] = i[1];
  assign o[469] = i[1];
  assign o[470] = i[1];
  assign o[471] = i[1];
  assign o[472] = i[1];
  assign o[473] = i[1];
  assign o[474] = i[1];
  assign o[475] = i[1];
  assign o[476] = i[1];
  assign o[477] = i[1];
  assign o[478] = i[1];
  assign o[479] = i[1];
  assign o[480] = i[1];
  assign o[481] = i[1];
  assign o[482] = i[1];
  assign o[483] = i[1];
  assign o[484] = i[1];
  assign o[485] = i[1];
  assign o[486] = i[1];
  assign o[487] = i[1];
  assign o[488] = i[1];
  assign o[489] = i[1];
  assign o[490] = i[1];
  assign o[491] = i[1];
  assign o[492] = i[1];
  assign o[493] = i[1];
  assign o[494] = i[1];
  assign o[495] = i[1];
  assign o[496] = i[1];
  assign o[497] = i[1];
  assign o[498] = i[1];
  assign o[499] = i[1];
  assign o[500] = i[1];
  assign o[501] = i[1];
  assign o[502] = i[1];
  assign o[503] = i[1];
  assign o[504] = i[1];
  assign o[505] = i[1];
  assign o[506] = i[1];
  assign o[507] = i[1];
  assign o[508] = i[1];
  assign o[509] = i[1];
  assign o[510] = i[1];
  assign o[511] = i[1];
  assign o[0] = i[0];
  assign o[1] = i[0];
  assign o[2] = i[0];
  assign o[3] = i[0];
  assign o[4] = i[0];
  assign o[5] = i[0];
  assign o[6] = i[0];
  assign o[7] = i[0];
  assign o[8] = i[0];
  assign o[9] = i[0];
  assign o[10] = i[0];
  assign o[11] = i[0];
  assign o[12] = i[0];
  assign o[13] = i[0];
  assign o[14] = i[0];
  assign o[15] = i[0];
  assign o[16] = i[0];
  assign o[17] = i[0];
  assign o[18] = i[0];
  assign o[19] = i[0];
  assign o[20] = i[0];
  assign o[21] = i[0];
  assign o[22] = i[0];
  assign o[23] = i[0];
  assign o[24] = i[0];
  assign o[25] = i[0];
  assign o[26] = i[0];
  assign o[27] = i[0];
  assign o[28] = i[0];
  assign o[29] = i[0];
  assign o[30] = i[0];
  assign o[31] = i[0];
  assign o[32] = i[0];
  assign o[33] = i[0];
  assign o[34] = i[0];
  assign o[35] = i[0];
  assign o[36] = i[0];
  assign o[37] = i[0];
  assign o[38] = i[0];
  assign o[39] = i[0];
  assign o[40] = i[0];
  assign o[41] = i[0];
  assign o[42] = i[0];
  assign o[43] = i[0];
  assign o[44] = i[0];
  assign o[45] = i[0];
  assign o[46] = i[0];
  assign o[47] = i[0];
  assign o[48] = i[0];
  assign o[49] = i[0];
  assign o[50] = i[0];
  assign o[51] = i[0];
  assign o[52] = i[0];
  assign o[53] = i[0];
  assign o[54] = i[0];
  assign o[55] = i[0];
  assign o[56] = i[0];
  assign o[57] = i[0];
  assign o[58] = i[0];
  assign o[59] = i[0];
  assign o[60] = i[0];
  assign o[61] = i[0];
  assign o[62] = i[0];
  assign o[63] = i[0];
  assign o[64] = i[0];
  assign o[65] = i[0];
  assign o[66] = i[0];
  assign o[67] = i[0];
  assign o[68] = i[0];
  assign o[69] = i[0];
  assign o[70] = i[0];
  assign o[71] = i[0];
  assign o[72] = i[0];
  assign o[73] = i[0];
  assign o[74] = i[0];
  assign o[75] = i[0];
  assign o[76] = i[0];
  assign o[77] = i[0];
  assign o[78] = i[0];
  assign o[79] = i[0];
  assign o[80] = i[0];
  assign o[81] = i[0];
  assign o[82] = i[0];
  assign o[83] = i[0];
  assign o[84] = i[0];
  assign o[85] = i[0];
  assign o[86] = i[0];
  assign o[87] = i[0];
  assign o[88] = i[0];
  assign o[89] = i[0];
  assign o[90] = i[0];
  assign o[91] = i[0];
  assign o[92] = i[0];
  assign o[93] = i[0];
  assign o[94] = i[0];
  assign o[95] = i[0];
  assign o[96] = i[0];
  assign o[97] = i[0];
  assign o[98] = i[0];
  assign o[99] = i[0];
  assign o[100] = i[0];
  assign o[101] = i[0];
  assign o[102] = i[0];
  assign o[103] = i[0];
  assign o[104] = i[0];
  assign o[105] = i[0];
  assign o[106] = i[0];
  assign o[107] = i[0];
  assign o[108] = i[0];
  assign o[109] = i[0];
  assign o[110] = i[0];
  assign o[111] = i[0];
  assign o[112] = i[0];
  assign o[113] = i[0];
  assign o[114] = i[0];
  assign o[115] = i[0];
  assign o[116] = i[0];
  assign o[117] = i[0];
  assign o[118] = i[0];
  assign o[119] = i[0];
  assign o[120] = i[0];
  assign o[121] = i[0];
  assign o[122] = i[0];
  assign o[123] = i[0];
  assign o[124] = i[0];
  assign o[125] = i[0];
  assign o[126] = i[0];
  assign o[127] = i[0];
  assign o[128] = i[0];
  assign o[129] = i[0];
  assign o[130] = i[0];
  assign o[131] = i[0];
  assign o[132] = i[0];
  assign o[133] = i[0];
  assign o[134] = i[0];
  assign o[135] = i[0];
  assign o[136] = i[0];
  assign o[137] = i[0];
  assign o[138] = i[0];
  assign o[139] = i[0];
  assign o[140] = i[0];
  assign o[141] = i[0];
  assign o[142] = i[0];
  assign o[143] = i[0];
  assign o[144] = i[0];
  assign o[145] = i[0];
  assign o[146] = i[0];
  assign o[147] = i[0];
  assign o[148] = i[0];
  assign o[149] = i[0];
  assign o[150] = i[0];
  assign o[151] = i[0];
  assign o[152] = i[0];
  assign o[153] = i[0];
  assign o[154] = i[0];
  assign o[155] = i[0];
  assign o[156] = i[0];
  assign o[157] = i[0];
  assign o[158] = i[0];
  assign o[159] = i[0];
  assign o[160] = i[0];
  assign o[161] = i[0];
  assign o[162] = i[0];
  assign o[163] = i[0];
  assign o[164] = i[0];
  assign o[165] = i[0];
  assign o[166] = i[0];
  assign o[167] = i[0];
  assign o[168] = i[0];
  assign o[169] = i[0];
  assign o[170] = i[0];
  assign o[171] = i[0];
  assign o[172] = i[0];
  assign o[173] = i[0];
  assign o[174] = i[0];
  assign o[175] = i[0];
  assign o[176] = i[0];
  assign o[177] = i[0];
  assign o[178] = i[0];
  assign o[179] = i[0];
  assign o[180] = i[0];
  assign o[181] = i[0];
  assign o[182] = i[0];
  assign o[183] = i[0];
  assign o[184] = i[0];
  assign o[185] = i[0];
  assign o[186] = i[0];
  assign o[187] = i[0];
  assign o[188] = i[0];
  assign o[189] = i[0];
  assign o[190] = i[0];
  assign o[191] = i[0];
  assign o[192] = i[0];
  assign o[193] = i[0];
  assign o[194] = i[0];
  assign o[195] = i[0];
  assign o[196] = i[0];
  assign o[197] = i[0];
  assign o[198] = i[0];
  assign o[199] = i[0];
  assign o[200] = i[0];
  assign o[201] = i[0];
  assign o[202] = i[0];
  assign o[203] = i[0];
  assign o[204] = i[0];
  assign o[205] = i[0];
  assign o[206] = i[0];
  assign o[207] = i[0];
  assign o[208] = i[0];
  assign o[209] = i[0];
  assign o[210] = i[0];
  assign o[211] = i[0];
  assign o[212] = i[0];
  assign o[213] = i[0];
  assign o[214] = i[0];
  assign o[215] = i[0];
  assign o[216] = i[0];
  assign o[217] = i[0];
  assign o[218] = i[0];
  assign o[219] = i[0];
  assign o[220] = i[0];
  assign o[221] = i[0];
  assign o[222] = i[0];
  assign o[223] = i[0];
  assign o[224] = i[0];
  assign o[225] = i[0];
  assign o[226] = i[0];
  assign o[227] = i[0];
  assign o[228] = i[0];
  assign o[229] = i[0];
  assign o[230] = i[0];
  assign o[231] = i[0];
  assign o[232] = i[0];
  assign o[233] = i[0];
  assign o[234] = i[0];
  assign o[235] = i[0];
  assign o[236] = i[0];
  assign o[237] = i[0];
  assign o[238] = i[0];
  assign o[239] = i[0];
  assign o[240] = i[0];
  assign o[241] = i[0];
  assign o[242] = i[0];
  assign o[243] = i[0];
  assign o[244] = i[0];
  assign o[245] = i[0];
  assign o[246] = i[0];
  assign o[247] = i[0];
  assign o[248] = i[0];
  assign o[249] = i[0];
  assign o[250] = i[0];
  assign o[251] = i[0];
  assign o[252] = i[0];
  assign o[253] = i[0];
  assign o[254] = i[0];
  assign o[255] = i[0];

endmodule

