

module top
(
  en_ls_i,
  clk_i,
  reset_i,
  clk_o,
  reset_o,
  fsb_v_i_o,
  fsb_data_i_o,
  fsb_yumi_o_i,
  fsb_v_o_i,
  fsb_data_o_i,
  fsb_ready_i_o,
  node_v_i_o,
  node_data_i_o,
  node_ready_o_i,
  node_v_o_i,
  node_data_o_i,
  node_yumi_i_o
);

  output [499:0] fsb_data_i_o;
  input [499:0] fsb_data_o_i;
  output [499:0] node_data_i_o;
  input [499:0] node_data_o_i;
  input en_ls_i;
  input clk_i;
  input reset_i;
  input fsb_yumi_o_i;
  input fsb_v_o_i;
  input node_ready_o_i;
  input node_v_o_i;
  output clk_o;
  output reset_o;
  output fsb_v_i_o;
  output fsb_ready_i_o;
  output node_v_i_o;
  output node_yumi_i_o;

  bsg_fsb_node_level_shift_fsb_domain
  wrapper
  (
    .fsb_data_i_o(fsb_data_i_o),
    .fsb_data_o_i(fsb_data_o_i),
    .node_data_i_o(node_data_i_o),
    .node_data_o_i(node_data_o_i),
    .en_ls_i(en_ls_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fsb_yumi_o_i(fsb_yumi_o_i),
    .fsb_v_o_i(fsb_v_o_i),
    .node_ready_o_i(node_ready_o_i),
    .node_v_o_i(node_v_o_i),
    .clk_o(clk_o),
    .reset_o(reset_o),
    .fsb_v_i_o(fsb_v_i_o),
    .fsb_ready_i_o(fsb_ready_i_o),
    .node_v_i_o(node_v_i_o),
    .node_yumi_i_o(node_yumi_i_o)
  );


endmodule



module bsg_level_shift_up_down_source_width_p1
(
  v0_en_i,
  v0_data_i,
  v1_data_o
);

  input [0:0] v0_data_i;
  output [0:0] v1_data_o;
  input v0_en_i;
  wire [0:0] v1_data_o;
  assign v1_data_o[0] = v0_data_i[0] & v0_en_i;

endmodule



module bsg_level_shift_up_down_sink_width_p1
(
  v0_data_i,
  v1_en_i,
  v1_data_o
);

  input [0:0] v0_data_i;
  output [0:0] v1_data_o;
  input v1_en_i;
  wire [0:0] v1_data_o;
  assign v1_data_o[0] = v0_data_i[0] & v1_en_i;

endmodule



module bsg_level_shift_up_down_sink_width_p500
(
  v0_data_i,
  v1_en_i,
  v1_data_o
);

  input [499:0] v0_data_i;
  output [499:0] v1_data_o;
  input v1_en_i;
  wire [499:0] v1_data_o;
  assign v1_data_o[499] = v0_data_i[499] & v1_en_i;
  assign v1_data_o[498] = v0_data_i[498] & v1_en_i;
  assign v1_data_o[497] = v0_data_i[497] & v1_en_i;
  assign v1_data_o[496] = v0_data_i[496] & v1_en_i;
  assign v1_data_o[495] = v0_data_i[495] & v1_en_i;
  assign v1_data_o[494] = v0_data_i[494] & v1_en_i;
  assign v1_data_o[493] = v0_data_i[493] & v1_en_i;
  assign v1_data_o[492] = v0_data_i[492] & v1_en_i;
  assign v1_data_o[491] = v0_data_i[491] & v1_en_i;
  assign v1_data_o[490] = v0_data_i[490] & v1_en_i;
  assign v1_data_o[489] = v0_data_i[489] & v1_en_i;
  assign v1_data_o[488] = v0_data_i[488] & v1_en_i;
  assign v1_data_o[487] = v0_data_i[487] & v1_en_i;
  assign v1_data_o[486] = v0_data_i[486] & v1_en_i;
  assign v1_data_o[485] = v0_data_i[485] & v1_en_i;
  assign v1_data_o[484] = v0_data_i[484] & v1_en_i;
  assign v1_data_o[483] = v0_data_i[483] & v1_en_i;
  assign v1_data_o[482] = v0_data_i[482] & v1_en_i;
  assign v1_data_o[481] = v0_data_i[481] & v1_en_i;
  assign v1_data_o[480] = v0_data_i[480] & v1_en_i;
  assign v1_data_o[479] = v0_data_i[479] & v1_en_i;
  assign v1_data_o[478] = v0_data_i[478] & v1_en_i;
  assign v1_data_o[477] = v0_data_i[477] & v1_en_i;
  assign v1_data_o[476] = v0_data_i[476] & v1_en_i;
  assign v1_data_o[475] = v0_data_i[475] & v1_en_i;
  assign v1_data_o[474] = v0_data_i[474] & v1_en_i;
  assign v1_data_o[473] = v0_data_i[473] & v1_en_i;
  assign v1_data_o[472] = v0_data_i[472] & v1_en_i;
  assign v1_data_o[471] = v0_data_i[471] & v1_en_i;
  assign v1_data_o[470] = v0_data_i[470] & v1_en_i;
  assign v1_data_o[469] = v0_data_i[469] & v1_en_i;
  assign v1_data_o[468] = v0_data_i[468] & v1_en_i;
  assign v1_data_o[467] = v0_data_i[467] & v1_en_i;
  assign v1_data_o[466] = v0_data_i[466] & v1_en_i;
  assign v1_data_o[465] = v0_data_i[465] & v1_en_i;
  assign v1_data_o[464] = v0_data_i[464] & v1_en_i;
  assign v1_data_o[463] = v0_data_i[463] & v1_en_i;
  assign v1_data_o[462] = v0_data_i[462] & v1_en_i;
  assign v1_data_o[461] = v0_data_i[461] & v1_en_i;
  assign v1_data_o[460] = v0_data_i[460] & v1_en_i;
  assign v1_data_o[459] = v0_data_i[459] & v1_en_i;
  assign v1_data_o[458] = v0_data_i[458] & v1_en_i;
  assign v1_data_o[457] = v0_data_i[457] & v1_en_i;
  assign v1_data_o[456] = v0_data_i[456] & v1_en_i;
  assign v1_data_o[455] = v0_data_i[455] & v1_en_i;
  assign v1_data_o[454] = v0_data_i[454] & v1_en_i;
  assign v1_data_o[453] = v0_data_i[453] & v1_en_i;
  assign v1_data_o[452] = v0_data_i[452] & v1_en_i;
  assign v1_data_o[451] = v0_data_i[451] & v1_en_i;
  assign v1_data_o[450] = v0_data_i[450] & v1_en_i;
  assign v1_data_o[449] = v0_data_i[449] & v1_en_i;
  assign v1_data_o[448] = v0_data_i[448] & v1_en_i;
  assign v1_data_o[447] = v0_data_i[447] & v1_en_i;
  assign v1_data_o[446] = v0_data_i[446] & v1_en_i;
  assign v1_data_o[445] = v0_data_i[445] & v1_en_i;
  assign v1_data_o[444] = v0_data_i[444] & v1_en_i;
  assign v1_data_o[443] = v0_data_i[443] & v1_en_i;
  assign v1_data_o[442] = v0_data_i[442] & v1_en_i;
  assign v1_data_o[441] = v0_data_i[441] & v1_en_i;
  assign v1_data_o[440] = v0_data_i[440] & v1_en_i;
  assign v1_data_o[439] = v0_data_i[439] & v1_en_i;
  assign v1_data_o[438] = v0_data_i[438] & v1_en_i;
  assign v1_data_o[437] = v0_data_i[437] & v1_en_i;
  assign v1_data_o[436] = v0_data_i[436] & v1_en_i;
  assign v1_data_o[435] = v0_data_i[435] & v1_en_i;
  assign v1_data_o[434] = v0_data_i[434] & v1_en_i;
  assign v1_data_o[433] = v0_data_i[433] & v1_en_i;
  assign v1_data_o[432] = v0_data_i[432] & v1_en_i;
  assign v1_data_o[431] = v0_data_i[431] & v1_en_i;
  assign v1_data_o[430] = v0_data_i[430] & v1_en_i;
  assign v1_data_o[429] = v0_data_i[429] & v1_en_i;
  assign v1_data_o[428] = v0_data_i[428] & v1_en_i;
  assign v1_data_o[427] = v0_data_i[427] & v1_en_i;
  assign v1_data_o[426] = v0_data_i[426] & v1_en_i;
  assign v1_data_o[425] = v0_data_i[425] & v1_en_i;
  assign v1_data_o[424] = v0_data_i[424] & v1_en_i;
  assign v1_data_o[423] = v0_data_i[423] & v1_en_i;
  assign v1_data_o[422] = v0_data_i[422] & v1_en_i;
  assign v1_data_o[421] = v0_data_i[421] & v1_en_i;
  assign v1_data_o[420] = v0_data_i[420] & v1_en_i;
  assign v1_data_o[419] = v0_data_i[419] & v1_en_i;
  assign v1_data_o[418] = v0_data_i[418] & v1_en_i;
  assign v1_data_o[417] = v0_data_i[417] & v1_en_i;
  assign v1_data_o[416] = v0_data_i[416] & v1_en_i;
  assign v1_data_o[415] = v0_data_i[415] & v1_en_i;
  assign v1_data_o[414] = v0_data_i[414] & v1_en_i;
  assign v1_data_o[413] = v0_data_i[413] & v1_en_i;
  assign v1_data_o[412] = v0_data_i[412] & v1_en_i;
  assign v1_data_o[411] = v0_data_i[411] & v1_en_i;
  assign v1_data_o[410] = v0_data_i[410] & v1_en_i;
  assign v1_data_o[409] = v0_data_i[409] & v1_en_i;
  assign v1_data_o[408] = v0_data_i[408] & v1_en_i;
  assign v1_data_o[407] = v0_data_i[407] & v1_en_i;
  assign v1_data_o[406] = v0_data_i[406] & v1_en_i;
  assign v1_data_o[405] = v0_data_i[405] & v1_en_i;
  assign v1_data_o[404] = v0_data_i[404] & v1_en_i;
  assign v1_data_o[403] = v0_data_i[403] & v1_en_i;
  assign v1_data_o[402] = v0_data_i[402] & v1_en_i;
  assign v1_data_o[401] = v0_data_i[401] & v1_en_i;
  assign v1_data_o[400] = v0_data_i[400] & v1_en_i;
  assign v1_data_o[399] = v0_data_i[399] & v1_en_i;
  assign v1_data_o[398] = v0_data_i[398] & v1_en_i;
  assign v1_data_o[397] = v0_data_i[397] & v1_en_i;
  assign v1_data_o[396] = v0_data_i[396] & v1_en_i;
  assign v1_data_o[395] = v0_data_i[395] & v1_en_i;
  assign v1_data_o[394] = v0_data_i[394] & v1_en_i;
  assign v1_data_o[393] = v0_data_i[393] & v1_en_i;
  assign v1_data_o[392] = v0_data_i[392] & v1_en_i;
  assign v1_data_o[391] = v0_data_i[391] & v1_en_i;
  assign v1_data_o[390] = v0_data_i[390] & v1_en_i;
  assign v1_data_o[389] = v0_data_i[389] & v1_en_i;
  assign v1_data_o[388] = v0_data_i[388] & v1_en_i;
  assign v1_data_o[387] = v0_data_i[387] & v1_en_i;
  assign v1_data_o[386] = v0_data_i[386] & v1_en_i;
  assign v1_data_o[385] = v0_data_i[385] & v1_en_i;
  assign v1_data_o[384] = v0_data_i[384] & v1_en_i;
  assign v1_data_o[383] = v0_data_i[383] & v1_en_i;
  assign v1_data_o[382] = v0_data_i[382] & v1_en_i;
  assign v1_data_o[381] = v0_data_i[381] & v1_en_i;
  assign v1_data_o[380] = v0_data_i[380] & v1_en_i;
  assign v1_data_o[379] = v0_data_i[379] & v1_en_i;
  assign v1_data_o[378] = v0_data_i[378] & v1_en_i;
  assign v1_data_o[377] = v0_data_i[377] & v1_en_i;
  assign v1_data_o[376] = v0_data_i[376] & v1_en_i;
  assign v1_data_o[375] = v0_data_i[375] & v1_en_i;
  assign v1_data_o[374] = v0_data_i[374] & v1_en_i;
  assign v1_data_o[373] = v0_data_i[373] & v1_en_i;
  assign v1_data_o[372] = v0_data_i[372] & v1_en_i;
  assign v1_data_o[371] = v0_data_i[371] & v1_en_i;
  assign v1_data_o[370] = v0_data_i[370] & v1_en_i;
  assign v1_data_o[369] = v0_data_i[369] & v1_en_i;
  assign v1_data_o[368] = v0_data_i[368] & v1_en_i;
  assign v1_data_o[367] = v0_data_i[367] & v1_en_i;
  assign v1_data_o[366] = v0_data_i[366] & v1_en_i;
  assign v1_data_o[365] = v0_data_i[365] & v1_en_i;
  assign v1_data_o[364] = v0_data_i[364] & v1_en_i;
  assign v1_data_o[363] = v0_data_i[363] & v1_en_i;
  assign v1_data_o[362] = v0_data_i[362] & v1_en_i;
  assign v1_data_o[361] = v0_data_i[361] & v1_en_i;
  assign v1_data_o[360] = v0_data_i[360] & v1_en_i;
  assign v1_data_o[359] = v0_data_i[359] & v1_en_i;
  assign v1_data_o[358] = v0_data_i[358] & v1_en_i;
  assign v1_data_o[357] = v0_data_i[357] & v1_en_i;
  assign v1_data_o[356] = v0_data_i[356] & v1_en_i;
  assign v1_data_o[355] = v0_data_i[355] & v1_en_i;
  assign v1_data_o[354] = v0_data_i[354] & v1_en_i;
  assign v1_data_o[353] = v0_data_i[353] & v1_en_i;
  assign v1_data_o[352] = v0_data_i[352] & v1_en_i;
  assign v1_data_o[351] = v0_data_i[351] & v1_en_i;
  assign v1_data_o[350] = v0_data_i[350] & v1_en_i;
  assign v1_data_o[349] = v0_data_i[349] & v1_en_i;
  assign v1_data_o[348] = v0_data_i[348] & v1_en_i;
  assign v1_data_o[347] = v0_data_i[347] & v1_en_i;
  assign v1_data_o[346] = v0_data_i[346] & v1_en_i;
  assign v1_data_o[345] = v0_data_i[345] & v1_en_i;
  assign v1_data_o[344] = v0_data_i[344] & v1_en_i;
  assign v1_data_o[343] = v0_data_i[343] & v1_en_i;
  assign v1_data_o[342] = v0_data_i[342] & v1_en_i;
  assign v1_data_o[341] = v0_data_i[341] & v1_en_i;
  assign v1_data_o[340] = v0_data_i[340] & v1_en_i;
  assign v1_data_o[339] = v0_data_i[339] & v1_en_i;
  assign v1_data_o[338] = v0_data_i[338] & v1_en_i;
  assign v1_data_o[337] = v0_data_i[337] & v1_en_i;
  assign v1_data_o[336] = v0_data_i[336] & v1_en_i;
  assign v1_data_o[335] = v0_data_i[335] & v1_en_i;
  assign v1_data_o[334] = v0_data_i[334] & v1_en_i;
  assign v1_data_o[333] = v0_data_i[333] & v1_en_i;
  assign v1_data_o[332] = v0_data_i[332] & v1_en_i;
  assign v1_data_o[331] = v0_data_i[331] & v1_en_i;
  assign v1_data_o[330] = v0_data_i[330] & v1_en_i;
  assign v1_data_o[329] = v0_data_i[329] & v1_en_i;
  assign v1_data_o[328] = v0_data_i[328] & v1_en_i;
  assign v1_data_o[327] = v0_data_i[327] & v1_en_i;
  assign v1_data_o[326] = v0_data_i[326] & v1_en_i;
  assign v1_data_o[325] = v0_data_i[325] & v1_en_i;
  assign v1_data_o[324] = v0_data_i[324] & v1_en_i;
  assign v1_data_o[323] = v0_data_i[323] & v1_en_i;
  assign v1_data_o[322] = v0_data_i[322] & v1_en_i;
  assign v1_data_o[321] = v0_data_i[321] & v1_en_i;
  assign v1_data_o[320] = v0_data_i[320] & v1_en_i;
  assign v1_data_o[319] = v0_data_i[319] & v1_en_i;
  assign v1_data_o[318] = v0_data_i[318] & v1_en_i;
  assign v1_data_o[317] = v0_data_i[317] & v1_en_i;
  assign v1_data_o[316] = v0_data_i[316] & v1_en_i;
  assign v1_data_o[315] = v0_data_i[315] & v1_en_i;
  assign v1_data_o[314] = v0_data_i[314] & v1_en_i;
  assign v1_data_o[313] = v0_data_i[313] & v1_en_i;
  assign v1_data_o[312] = v0_data_i[312] & v1_en_i;
  assign v1_data_o[311] = v0_data_i[311] & v1_en_i;
  assign v1_data_o[310] = v0_data_i[310] & v1_en_i;
  assign v1_data_o[309] = v0_data_i[309] & v1_en_i;
  assign v1_data_o[308] = v0_data_i[308] & v1_en_i;
  assign v1_data_o[307] = v0_data_i[307] & v1_en_i;
  assign v1_data_o[306] = v0_data_i[306] & v1_en_i;
  assign v1_data_o[305] = v0_data_i[305] & v1_en_i;
  assign v1_data_o[304] = v0_data_i[304] & v1_en_i;
  assign v1_data_o[303] = v0_data_i[303] & v1_en_i;
  assign v1_data_o[302] = v0_data_i[302] & v1_en_i;
  assign v1_data_o[301] = v0_data_i[301] & v1_en_i;
  assign v1_data_o[300] = v0_data_i[300] & v1_en_i;
  assign v1_data_o[299] = v0_data_i[299] & v1_en_i;
  assign v1_data_o[298] = v0_data_i[298] & v1_en_i;
  assign v1_data_o[297] = v0_data_i[297] & v1_en_i;
  assign v1_data_o[296] = v0_data_i[296] & v1_en_i;
  assign v1_data_o[295] = v0_data_i[295] & v1_en_i;
  assign v1_data_o[294] = v0_data_i[294] & v1_en_i;
  assign v1_data_o[293] = v0_data_i[293] & v1_en_i;
  assign v1_data_o[292] = v0_data_i[292] & v1_en_i;
  assign v1_data_o[291] = v0_data_i[291] & v1_en_i;
  assign v1_data_o[290] = v0_data_i[290] & v1_en_i;
  assign v1_data_o[289] = v0_data_i[289] & v1_en_i;
  assign v1_data_o[288] = v0_data_i[288] & v1_en_i;
  assign v1_data_o[287] = v0_data_i[287] & v1_en_i;
  assign v1_data_o[286] = v0_data_i[286] & v1_en_i;
  assign v1_data_o[285] = v0_data_i[285] & v1_en_i;
  assign v1_data_o[284] = v0_data_i[284] & v1_en_i;
  assign v1_data_o[283] = v0_data_i[283] & v1_en_i;
  assign v1_data_o[282] = v0_data_i[282] & v1_en_i;
  assign v1_data_o[281] = v0_data_i[281] & v1_en_i;
  assign v1_data_o[280] = v0_data_i[280] & v1_en_i;
  assign v1_data_o[279] = v0_data_i[279] & v1_en_i;
  assign v1_data_o[278] = v0_data_i[278] & v1_en_i;
  assign v1_data_o[277] = v0_data_i[277] & v1_en_i;
  assign v1_data_o[276] = v0_data_i[276] & v1_en_i;
  assign v1_data_o[275] = v0_data_i[275] & v1_en_i;
  assign v1_data_o[274] = v0_data_i[274] & v1_en_i;
  assign v1_data_o[273] = v0_data_i[273] & v1_en_i;
  assign v1_data_o[272] = v0_data_i[272] & v1_en_i;
  assign v1_data_o[271] = v0_data_i[271] & v1_en_i;
  assign v1_data_o[270] = v0_data_i[270] & v1_en_i;
  assign v1_data_o[269] = v0_data_i[269] & v1_en_i;
  assign v1_data_o[268] = v0_data_i[268] & v1_en_i;
  assign v1_data_o[267] = v0_data_i[267] & v1_en_i;
  assign v1_data_o[266] = v0_data_i[266] & v1_en_i;
  assign v1_data_o[265] = v0_data_i[265] & v1_en_i;
  assign v1_data_o[264] = v0_data_i[264] & v1_en_i;
  assign v1_data_o[263] = v0_data_i[263] & v1_en_i;
  assign v1_data_o[262] = v0_data_i[262] & v1_en_i;
  assign v1_data_o[261] = v0_data_i[261] & v1_en_i;
  assign v1_data_o[260] = v0_data_i[260] & v1_en_i;
  assign v1_data_o[259] = v0_data_i[259] & v1_en_i;
  assign v1_data_o[258] = v0_data_i[258] & v1_en_i;
  assign v1_data_o[257] = v0_data_i[257] & v1_en_i;
  assign v1_data_o[256] = v0_data_i[256] & v1_en_i;
  assign v1_data_o[255] = v0_data_i[255] & v1_en_i;
  assign v1_data_o[254] = v0_data_i[254] & v1_en_i;
  assign v1_data_o[253] = v0_data_i[253] & v1_en_i;
  assign v1_data_o[252] = v0_data_i[252] & v1_en_i;
  assign v1_data_o[251] = v0_data_i[251] & v1_en_i;
  assign v1_data_o[250] = v0_data_i[250] & v1_en_i;
  assign v1_data_o[249] = v0_data_i[249] & v1_en_i;
  assign v1_data_o[248] = v0_data_i[248] & v1_en_i;
  assign v1_data_o[247] = v0_data_i[247] & v1_en_i;
  assign v1_data_o[246] = v0_data_i[246] & v1_en_i;
  assign v1_data_o[245] = v0_data_i[245] & v1_en_i;
  assign v1_data_o[244] = v0_data_i[244] & v1_en_i;
  assign v1_data_o[243] = v0_data_i[243] & v1_en_i;
  assign v1_data_o[242] = v0_data_i[242] & v1_en_i;
  assign v1_data_o[241] = v0_data_i[241] & v1_en_i;
  assign v1_data_o[240] = v0_data_i[240] & v1_en_i;
  assign v1_data_o[239] = v0_data_i[239] & v1_en_i;
  assign v1_data_o[238] = v0_data_i[238] & v1_en_i;
  assign v1_data_o[237] = v0_data_i[237] & v1_en_i;
  assign v1_data_o[236] = v0_data_i[236] & v1_en_i;
  assign v1_data_o[235] = v0_data_i[235] & v1_en_i;
  assign v1_data_o[234] = v0_data_i[234] & v1_en_i;
  assign v1_data_o[233] = v0_data_i[233] & v1_en_i;
  assign v1_data_o[232] = v0_data_i[232] & v1_en_i;
  assign v1_data_o[231] = v0_data_i[231] & v1_en_i;
  assign v1_data_o[230] = v0_data_i[230] & v1_en_i;
  assign v1_data_o[229] = v0_data_i[229] & v1_en_i;
  assign v1_data_o[228] = v0_data_i[228] & v1_en_i;
  assign v1_data_o[227] = v0_data_i[227] & v1_en_i;
  assign v1_data_o[226] = v0_data_i[226] & v1_en_i;
  assign v1_data_o[225] = v0_data_i[225] & v1_en_i;
  assign v1_data_o[224] = v0_data_i[224] & v1_en_i;
  assign v1_data_o[223] = v0_data_i[223] & v1_en_i;
  assign v1_data_o[222] = v0_data_i[222] & v1_en_i;
  assign v1_data_o[221] = v0_data_i[221] & v1_en_i;
  assign v1_data_o[220] = v0_data_i[220] & v1_en_i;
  assign v1_data_o[219] = v0_data_i[219] & v1_en_i;
  assign v1_data_o[218] = v0_data_i[218] & v1_en_i;
  assign v1_data_o[217] = v0_data_i[217] & v1_en_i;
  assign v1_data_o[216] = v0_data_i[216] & v1_en_i;
  assign v1_data_o[215] = v0_data_i[215] & v1_en_i;
  assign v1_data_o[214] = v0_data_i[214] & v1_en_i;
  assign v1_data_o[213] = v0_data_i[213] & v1_en_i;
  assign v1_data_o[212] = v0_data_i[212] & v1_en_i;
  assign v1_data_o[211] = v0_data_i[211] & v1_en_i;
  assign v1_data_o[210] = v0_data_i[210] & v1_en_i;
  assign v1_data_o[209] = v0_data_i[209] & v1_en_i;
  assign v1_data_o[208] = v0_data_i[208] & v1_en_i;
  assign v1_data_o[207] = v0_data_i[207] & v1_en_i;
  assign v1_data_o[206] = v0_data_i[206] & v1_en_i;
  assign v1_data_o[205] = v0_data_i[205] & v1_en_i;
  assign v1_data_o[204] = v0_data_i[204] & v1_en_i;
  assign v1_data_o[203] = v0_data_i[203] & v1_en_i;
  assign v1_data_o[202] = v0_data_i[202] & v1_en_i;
  assign v1_data_o[201] = v0_data_i[201] & v1_en_i;
  assign v1_data_o[200] = v0_data_i[200] & v1_en_i;
  assign v1_data_o[199] = v0_data_i[199] & v1_en_i;
  assign v1_data_o[198] = v0_data_i[198] & v1_en_i;
  assign v1_data_o[197] = v0_data_i[197] & v1_en_i;
  assign v1_data_o[196] = v0_data_i[196] & v1_en_i;
  assign v1_data_o[195] = v0_data_i[195] & v1_en_i;
  assign v1_data_o[194] = v0_data_i[194] & v1_en_i;
  assign v1_data_o[193] = v0_data_i[193] & v1_en_i;
  assign v1_data_o[192] = v0_data_i[192] & v1_en_i;
  assign v1_data_o[191] = v0_data_i[191] & v1_en_i;
  assign v1_data_o[190] = v0_data_i[190] & v1_en_i;
  assign v1_data_o[189] = v0_data_i[189] & v1_en_i;
  assign v1_data_o[188] = v0_data_i[188] & v1_en_i;
  assign v1_data_o[187] = v0_data_i[187] & v1_en_i;
  assign v1_data_o[186] = v0_data_i[186] & v1_en_i;
  assign v1_data_o[185] = v0_data_i[185] & v1_en_i;
  assign v1_data_o[184] = v0_data_i[184] & v1_en_i;
  assign v1_data_o[183] = v0_data_i[183] & v1_en_i;
  assign v1_data_o[182] = v0_data_i[182] & v1_en_i;
  assign v1_data_o[181] = v0_data_i[181] & v1_en_i;
  assign v1_data_o[180] = v0_data_i[180] & v1_en_i;
  assign v1_data_o[179] = v0_data_i[179] & v1_en_i;
  assign v1_data_o[178] = v0_data_i[178] & v1_en_i;
  assign v1_data_o[177] = v0_data_i[177] & v1_en_i;
  assign v1_data_o[176] = v0_data_i[176] & v1_en_i;
  assign v1_data_o[175] = v0_data_i[175] & v1_en_i;
  assign v1_data_o[174] = v0_data_i[174] & v1_en_i;
  assign v1_data_o[173] = v0_data_i[173] & v1_en_i;
  assign v1_data_o[172] = v0_data_i[172] & v1_en_i;
  assign v1_data_o[171] = v0_data_i[171] & v1_en_i;
  assign v1_data_o[170] = v0_data_i[170] & v1_en_i;
  assign v1_data_o[169] = v0_data_i[169] & v1_en_i;
  assign v1_data_o[168] = v0_data_i[168] & v1_en_i;
  assign v1_data_o[167] = v0_data_i[167] & v1_en_i;
  assign v1_data_o[166] = v0_data_i[166] & v1_en_i;
  assign v1_data_o[165] = v0_data_i[165] & v1_en_i;
  assign v1_data_o[164] = v0_data_i[164] & v1_en_i;
  assign v1_data_o[163] = v0_data_i[163] & v1_en_i;
  assign v1_data_o[162] = v0_data_i[162] & v1_en_i;
  assign v1_data_o[161] = v0_data_i[161] & v1_en_i;
  assign v1_data_o[160] = v0_data_i[160] & v1_en_i;
  assign v1_data_o[159] = v0_data_i[159] & v1_en_i;
  assign v1_data_o[158] = v0_data_i[158] & v1_en_i;
  assign v1_data_o[157] = v0_data_i[157] & v1_en_i;
  assign v1_data_o[156] = v0_data_i[156] & v1_en_i;
  assign v1_data_o[155] = v0_data_i[155] & v1_en_i;
  assign v1_data_o[154] = v0_data_i[154] & v1_en_i;
  assign v1_data_o[153] = v0_data_i[153] & v1_en_i;
  assign v1_data_o[152] = v0_data_i[152] & v1_en_i;
  assign v1_data_o[151] = v0_data_i[151] & v1_en_i;
  assign v1_data_o[150] = v0_data_i[150] & v1_en_i;
  assign v1_data_o[149] = v0_data_i[149] & v1_en_i;
  assign v1_data_o[148] = v0_data_i[148] & v1_en_i;
  assign v1_data_o[147] = v0_data_i[147] & v1_en_i;
  assign v1_data_o[146] = v0_data_i[146] & v1_en_i;
  assign v1_data_o[145] = v0_data_i[145] & v1_en_i;
  assign v1_data_o[144] = v0_data_i[144] & v1_en_i;
  assign v1_data_o[143] = v0_data_i[143] & v1_en_i;
  assign v1_data_o[142] = v0_data_i[142] & v1_en_i;
  assign v1_data_o[141] = v0_data_i[141] & v1_en_i;
  assign v1_data_o[140] = v0_data_i[140] & v1_en_i;
  assign v1_data_o[139] = v0_data_i[139] & v1_en_i;
  assign v1_data_o[138] = v0_data_i[138] & v1_en_i;
  assign v1_data_o[137] = v0_data_i[137] & v1_en_i;
  assign v1_data_o[136] = v0_data_i[136] & v1_en_i;
  assign v1_data_o[135] = v0_data_i[135] & v1_en_i;
  assign v1_data_o[134] = v0_data_i[134] & v1_en_i;
  assign v1_data_o[133] = v0_data_i[133] & v1_en_i;
  assign v1_data_o[132] = v0_data_i[132] & v1_en_i;
  assign v1_data_o[131] = v0_data_i[131] & v1_en_i;
  assign v1_data_o[130] = v0_data_i[130] & v1_en_i;
  assign v1_data_o[129] = v0_data_i[129] & v1_en_i;
  assign v1_data_o[128] = v0_data_i[128] & v1_en_i;
  assign v1_data_o[127] = v0_data_i[127] & v1_en_i;
  assign v1_data_o[126] = v0_data_i[126] & v1_en_i;
  assign v1_data_o[125] = v0_data_i[125] & v1_en_i;
  assign v1_data_o[124] = v0_data_i[124] & v1_en_i;
  assign v1_data_o[123] = v0_data_i[123] & v1_en_i;
  assign v1_data_o[122] = v0_data_i[122] & v1_en_i;
  assign v1_data_o[121] = v0_data_i[121] & v1_en_i;
  assign v1_data_o[120] = v0_data_i[120] & v1_en_i;
  assign v1_data_o[119] = v0_data_i[119] & v1_en_i;
  assign v1_data_o[118] = v0_data_i[118] & v1_en_i;
  assign v1_data_o[117] = v0_data_i[117] & v1_en_i;
  assign v1_data_o[116] = v0_data_i[116] & v1_en_i;
  assign v1_data_o[115] = v0_data_i[115] & v1_en_i;
  assign v1_data_o[114] = v0_data_i[114] & v1_en_i;
  assign v1_data_o[113] = v0_data_i[113] & v1_en_i;
  assign v1_data_o[112] = v0_data_i[112] & v1_en_i;
  assign v1_data_o[111] = v0_data_i[111] & v1_en_i;
  assign v1_data_o[110] = v0_data_i[110] & v1_en_i;
  assign v1_data_o[109] = v0_data_i[109] & v1_en_i;
  assign v1_data_o[108] = v0_data_i[108] & v1_en_i;
  assign v1_data_o[107] = v0_data_i[107] & v1_en_i;
  assign v1_data_o[106] = v0_data_i[106] & v1_en_i;
  assign v1_data_o[105] = v0_data_i[105] & v1_en_i;
  assign v1_data_o[104] = v0_data_i[104] & v1_en_i;
  assign v1_data_o[103] = v0_data_i[103] & v1_en_i;
  assign v1_data_o[102] = v0_data_i[102] & v1_en_i;
  assign v1_data_o[101] = v0_data_i[101] & v1_en_i;
  assign v1_data_o[100] = v0_data_i[100] & v1_en_i;
  assign v1_data_o[99] = v0_data_i[99] & v1_en_i;
  assign v1_data_o[98] = v0_data_i[98] & v1_en_i;
  assign v1_data_o[97] = v0_data_i[97] & v1_en_i;
  assign v1_data_o[96] = v0_data_i[96] & v1_en_i;
  assign v1_data_o[95] = v0_data_i[95] & v1_en_i;
  assign v1_data_o[94] = v0_data_i[94] & v1_en_i;
  assign v1_data_o[93] = v0_data_i[93] & v1_en_i;
  assign v1_data_o[92] = v0_data_i[92] & v1_en_i;
  assign v1_data_o[91] = v0_data_i[91] & v1_en_i;
  assign v1_data_o[90] = v0_data_i[90] & v1_en_i;
  assign v1_data_o[89] = v0_data_i[89] & v1_en_i;
  assign v1_data_o[88] = v0_data_i[88] & v1_en_i;
  assign v1_data_o[87] = v0_data_i[87] & v1_en_i;
  assign v1_data_o[86] = v0_data_i[86] & v1_en_i;
  assign v1_data_o[85] = v0_data_i[85] & v1_en_i;
  assign v1_data_o[84] = v0_data_i[84] & v1_en_i;
  assign v1_data_o[83] = v0_data_i[83] & v1_en_i;
  assign v1_data_o[82] = v0_data_i[82] & v1_en_i;
  assign v1_data_o[81] = v0_data_i[81] & v1_en_i;
  assign v1_data_o[80] = v0_data_i[80] & v1_en_i;
  assign v1_data_o[79] = v0_data_i[79] & v1_en_i;
  assign v1_data_o[78] = v0_data_i[78] & v1_en_i;
  assign v1_data_o[77] = v0_data_i[77] & v1_en_i;
  assign v1_data_o[76] = v0_data_i[76] & v1_en_i;
  assign v1_data_o[75] = v0_data_i[75] & v1_en_i;
  assign v1_data_o[74] = v0_data_i[74] & v1_en_i;
  assign v1_data_o[73] = v0_data_i[73] & v1_en_i;
  assign v1_data_o[72] = v0_data_i[72] & v1_en_i;
  assign v1_data_o[71] = v0_data_i[71] & v1_en_i;
  assign v1_data_o[70] = v0_data_i[70] & v1_en_i;
  assign v1_data_o[69] = v0_data_i[69] & v1_en_i;
  assign v1_data_o[68] = v0_data_i[68] & v1_en_i;
  assign v1_data_o[67] = v0_data_i[67] & v1_en_i;
  assign v1_data_o[66] = v0_data_i[66] & v1_en_i;
  assign v1_data_o[65] = v0_data_i[65] & v1_en_i;
  assign v1_data_o[64] = v0_data_i[64] & v1_en_i;
  assign v1_data_o[63] = v0_data_i[63] & v1_en_i;
  assign v1_data_o[62] = v0_data_i[62] & v1_en_i;
  assign v1_data_o[61] = v0_data_i[61] & v1_en_i;
  assign v1_data_o[60] = v0_data_i[60] & v1_en_i;
  assign v1_data_o[59] = v0_data_i[59] & v1_en_i;
  assign v1_data_o[58] = v0_data_i[58] & v1_en_i;
  assign v1_data_o[57] = v0_data_i[57] & v1_en_i;
  assign v1_data_o[56] = v0_data_i[56] & v1_en_i;
  assign v1_data_o[55] = v0_data_i[55] & v1_en_i;
  assign v1_data_o[54] = v0_data_i[54] & v1_en_i;
  assign v1_data_o[53] = v0_data_i[53] & v1_en_i;
  assign v1_data_o[52] = v0_data_i[52] & v1_en_i;
  assign v1_data_o[51] = v0_data_i[51] & v1_en_i;
  assign v1_data_o[50] = v0_data_i[50] & v1_en_i;
  assign v1_data_o[49] = v0_data_i[49] & v1_en_i;
  assign v1_data_o[48] = v0_data_i[48] & v1_en_i;
  assign v1_data_o[47] = v0_data_i[47] & v1_en_i;
  assign v1_data_o[46] = v0_data_i[46] & v1_en_i;
  assign v1_data_o[45] = v0_data_i[45] & v1_en_i;
  assign v1_data_o[44] = v0_data_i[44] & v1_en_i;
  assign v1_data_o[43] = v0_data_i[43] & v1_en_i;
  assign v1_data_o[42] = v0_data_i[42] & v1_en_i;
  assign v1_data_o[41] = v0_data_i[41] & v1_en_i;
  assign v1_data_o[40] = v0_data_i[40] & v1_en_i;
  assign v1_data_o[39] = v0_data_i[39] & v1_en_i;
  assign v1_data_o[38] = v0_data_i[38] & v1_en_i;
  assign v1_data_o[37] = v0_data_i[37] & v1_en_i;
  assign v1_data_o[36] = v0_data_i[36] & v1_en_i;
  assign v1_data_o[35] = v0_data_i[35] & v1_en_i;
  assign v1_data_o[34] = v0_data_i[34] & v1_en_i;
  assign v1_data_o[33] = v0_data_i[33] & v1_en_i;
  assign v1_data_o[32] = v0_data_i[32] & v1_en_i;
  assign v1_data_o[31] = v0_data_i[31] & v1_en_i;
  assign v1_data_o[30] = v0_data_i[30] & v1_en_i;
  assign v1_data_o[29] = v0_data_i[29] & v1_en_i;
  assign v1_data_o[28] = v0_data_i[28] & v1_en_i;
  assign v1_data_o[27] = v0_data_i[27] & v1_en_i;
  assign v1_data_o[26] = v0_data_i[26] & v1_en_i;
  assign v1_data_o[25] = v0_data_i[25] & v1_en_i;
  assign v1_data_o[24] = v0_data_i[24] & v1_en_i;
  assign v1_data_o[23] = v0_data_i[23] & v1_en_i;
  assign v1_data_o[22] = v0_data_i[22] & v1_en_i;
  assign v1_data_o[21] = v0_data_i[21] & v1_en_i;
  assign v1_data_o[20] = v0_data_i[20] & v1_en_i;
  assign v1_data_o[19] = v0_data_i[19] & v1_en_i;
  assign v1_data_o[18] = v0_data_i[18] & v1_en_i;
  assign v1_data_o[17] = v0_data_i[17] & v1_en_i;
  assign v1_data_o[16] = v0_data_i[16] & v1_en_i;
  assign v1_data_o[15] = v0_data_i[15] & v1_en_i;
  assign v1_data_o[14] = v0_data_i[14] & v1_en_i;
  assign v1_data_o[13] = v0_data_i[13] & v1_en_i;
  assign v1_data_o[12] = v0_data_i[12] & v1_en_i;
  assign v1_data_o[11] = v0_data_i[11] & v1_en_i;
  assign v1_data_o[10] = v0_data_i[10] & v1_en_i;
  assign v1_data_o[9] = v0_data_i[9] & v1_en_i;
  assign v1_data_o[8] = v0_data_i[8] & v1_en_i;
  assign v1_data_o[7] = v0_data_i[7] & v1_en_i;
  assign v1_data_o[6] = v0_data_i[6] & v1_en_i;
  assign v1_data_o[5] = v0_data_i[5] & v1_en_i;
  assign v1_data_o[4] = v0_data_i[4] & v1_en_i;
  assign v1_data_o[3] = v0_data_i[3] & v1_en_i;
  assign v1_data_o[2] = v0_data_i[2] & v1_en_i;
  assign v1_data_o[1] = v0_data_i[1] & v1_en_i;
  assign v1_data_o[0] = v0_data_i[0] & v1_en_i;

endmodule



module bsg_level_shift_up_down_source_width_p500
(
  v0_en_i,
  v0_data_i,
  v1_data_o
);

  input [499:0] v0_data_i;
  output [499:0] v1_data_o;
  input v0_en_i;
  wire [499:0] v1_data_o;
  assign v1_data_o[499] = v0_data_i[499] & v0_en_i;
  assign v1_data_o[498] = v0_data_i[498] & v0_en_i;
  assign v1_data_o[497] = v0_data_i[497] & v0_en_i;
  assign v1_data_o[496] = v0_data_i[496] & v0_en_i;
  assign v1_data_o[495] = v0_data_i[495] & v0_en_i;
  assign v1_data_o[494] = v0_data_i[494] & v0_en_i;
  assign v1_data_o[493] = v0_data_i[493] & v0_en_i;
  assign v1_data_o[492] = v0_data_i[492] & v0_en_i;
  assign v1_data_o[491] = v0_data_i[491] & v0_en_i;
  assign v1_data_o[490] = v0_data_i[490] & v0_en_i;
  assign v1_data_o[489] = v0_data_i[489] & v0_en_i;
  assign v1_data_o[488] = v0_data_i[488] & v0_en_i;
  assign v1_data_o[487] = v0_data_i[487] & v0_en_i;
  assign v1_data_o[486] = v0_data_i[486] & v0_en_i;
  assign v1_data_o[485] = v0_data_i[485] & v0_en_i;
  assign v1_data_o[484] = v0_data_i[484] & v0_en_i;
  assign v1_data_o[483] = v0_data_i[483] & v0_en_i;
  assign v1_data_o[482] = v0_data_i[482] & v0_en_i;
  assign v1_data_o[481] = v0_data_i[481] & v0_en_i;
  assign v1_data_o[480] = v0_data_i[480] & v0_en_i;
  assign v1_data_o[479] = v0_data_i[479] & v0_en_i;
  assign v1_data_o[478] = v0_data_i[478] & v0_en_i;
  assign v1_data_o[477] = v0_data_i[477] & v0_en_i;
  assign v1_data_o[476] = v0_data_i[476] & v0_en_i;
  assign v1_data_o[475] = v0_data_i[475] & v0_en_i;
  assign v1_data_o[474] = v0_data_i[474] & v0_en_i;
  assign v1_data_o[473] = v0_data_i[473] & v0_en_i;
  assign v1_data_o[472] = v0_data_i[472] & v0_en_i;
  assign v1_data_o[471] = v0_data_i[471] & v0_en_i;
  assign v1_data_o[470] = v0_data_i[470] & v0_en_i;
  assign v1_data_o[469] = v0_data_i[469] & v0_en_i;
  assign v1_data_o[468] = v0_data_i[468] & v0_en_i;
  assign v1_data_o[467] = v0_data_i[467] & v0_en_i;
  assign v1_data_o[466] = v0_data_i[466] & v0_en_i;
  assign v1_data_o[465] = v0_data_i[465] & v0_en_i;
  assign v1_data_o[464] = v0_data_i[464] & v0_en_i;
  assign v1_data_o[463] = v0_data_i[463] & v0_en_i;
  assign v1_data_o[462] = v0_data_i[462] & v0_en_i;
  assign v1_data_o[461] = v0_data_i[461] & v0_en_i;
  assign v1_data_o[460] = v0_data_i[460] & v0_en_i;
  assign v1_data_o[459] = v0_data_i[459] & v0_en_i;
  assign v1_data_o[458] = v0_data_i[458] & v0_en_i;
  assign v1_data_o[457] = v0_data_i[457] & v0_en_i;
  assign v1_data_o[456] = v0_data_i[456] & v0_en_i;
  assign v1_data_o[455] = v0_data_i[455] & v0_en_i;
  assign v1_data_o[454] = v0_data_i[454] & v0_en_i;
  assign v1_data_o[453] = v0_data_i[453] & v0_en_i;
  assign v1_data_o[452] = v0_data_i[452] & v0_en_i;
  assign v1_data_o[451] = v0_data_i[451] & v0_en_i;
  assign v1_data_o[450] = v0_data_i[450] & v0_en_i;
  assign v1_data_o[449] = v0_data_i[449] & v0_en_i;
  assign v1_data_o[448] = v0_data_i[448] & v0_en_i;
  assign v1_data_o[447] = v0_data_i[447] & v0_en_i;
  assign v1_data_o[446] = v0_data_i[446] & v0_en_i;
  assign v1_data_o[445] = v0_data_i[445] & v0_en_i;
  assign v1_data_o[444] = v0_data_i[444] & v0_en_i;
  assign v1_data_o[443] = v0_data_i[443] & v0_en_i;
  assign v1_data_o[442] = v0_data_i[442] & v0_en_i;
  assign v1_data_o[441] = v0_data_i[441] & v0_en_i;
  assign v1_data_o[440] = v0_data_i[440] & v0_en_i;
  assign v1_data_o[439] = v0_data_i[439] & v0_en_i;
  assign v1_data_o[438] = v0_data_i[438] & v0_en_i;
  assign v1_data_o[437] = v0_data_i[437] & v0_en_i;
  assign v1_data_o[436] = v0_data_i[436] & v0_en_i;
  assign v1_data_o[435] = v0_data_i[435] & v0_en_i;
  assign v1_data_o[434] = v0_data_i[434] & v0_en_i;
  assign v1_data_o[433] = v0_data_i[433] & v0_en_i;
  assign v1_data_o[432] = v0_data_i[432] & v0_en_i;
  assign v1_data_o[431] = v0_data_i[431] & v0_en_i;
  assign v1_data_o[430] = v0_data_i[430] & v0_en_i;
  assign v1_data_o[429] = v0_data_i[429] & v0_en_i;
  assign v1_data_o[428] = v0_data_i[428] & v0_en_i;
  assign v1_data_o[427] = v0_data_i[427] & v0_en_i;
  assign v1_data_o[426] = v0_data_i[426] & v0_en_i;
  assign v1_data_o[425] = v0_data_i[425] & v0_en_i;
  assign v1_data_o[424] = v0_data_i[424] & v0_en_i;
  assign v1_data_o[423] = v0_data_i[423] & v0_en_i;
  assign v1_data_o[422] = v0_data_i[422] & v0_en_i;
  assign v1_data_o[421] = v0_data_i[421] & v0_en_i;
  assign v1_data_o[420] = v0_data_i[420] & v0_en_i;
  assign v1_data_o[419] = v0_data_i[419] & v0_en_i;
  assign v1_data_o[418] = v0_data_i[418] & v0_en_i;
  assign v1_data_o[417] = v0_data_i[417] & v0_en_i;
  assign v1_data_o[416] = v0_data_i[416] & v0_en_i;
  assign v1_data_o[415] = v0_data_i[415] & v0_en_i;
  assign v1_data_o[414] = v0_data_i[414] & v0_en_i;
  assign v1_data_o[413] = v0_data_i[413] & v0_en_i;
  assign v1_data_o[412] = v0_data_i[412] & v0_en_i;
  assign v1_data_o[411] = v0_data_i[411] & v0_en_i;
  assign v1_data_o[410] = v0_data_i[410] & v0_en_i;
  assign v1_data_o[409] = v0_data_i[409] & v0_en_i;
  assign v1_data_o[408] = v0_data_i[408] & v0_en_i;
  assign v1_data_o[407] = v0_data_i[407] & v0_en_i;
  assign v1_data_o[406] = v0_data_i[406] & v0_en_i;
  assign v1_data_o[405] = v0_data_i[405] & v0_en_i;
  assign v1_data_o[404] = v0_data_i[404] & v0_en_i;
  assign v1_data_o[403] = v0_data_i[403] & v0_en_i;
  assign v1_data_o[402] = v0_data_i[402] & v0_en_i;
  assign v1_data_o[401] = v0_data_i[401] & v0_en_i;
  assign v1_data_o[400] = v0_data_i[400] & v0_en_i;
  assign v1_data_o[399] = v0_data_i[399] & v0_en_i;
  assign v1_data_o[398] = v0_data_i[398] & v0_en_i;
  assign v1_data_o[397] = v0_data_i[397] & v0_en_i;
  assign v1_data_o[396] = v0_data_i[396] & v0_en_i;
  assign v1_data_o[395] = v0_data_i[395] & v0_en_i;
  assign v1_data_o[394] = v0_data_i[394] & v0_en_i;
  assign v1_data_o[393] = v0_data_i[393] & v0_en_i;
  assign v1_data_o[392] = v0_data_i[392] & v0_en_i;
  assign v1_data_o[391] = v0_data_i[391] & v0_en_i;
  assign v1_data_o[390] = v0_data_i[390] & v0_en_i;
  assign v1_data_o[389] = v0_data_i[389] & v0_en_i;
  assign v1_data_o[388] = v0_data_i[388] & v0_en_i;
  assign v1_data_o[387] = v0_data_i[387] & v0_en_i;
  assign v1_data_o[386] = v0_data_i[386] & v0_en_i;
  assign v1_data_o[385] = v0_data_i[385] & v0_en_i;
  assign v1_data_o[384] = v0_data_i[384] & v0_en_i;
  assign v1_data_o[383] = v0_data_i[383] & v0_en_i;
  assign v1_data_o[382] = v0_data_i[382] & v0_en_i;
  assign v1_data_o[381] = v0_data_i[381] & v0_en_i;
  assign v1_data_o[380] = v0_data_i[380] & v0_en_i;
  assign v1_data_o[379] = v0_data_i[379] & v0_en_i;
  assign v1_data_o[378] = v0_data_i[378] & v0_en_i;
  assign v1_data_o[377] = v0_data_i[377] & v0_en_i;
  assign v1_data_o[376] = v0_data_i[376] & v0_en_i;
  assign v1_data_o[375] = v0_data_i[375] & v0_en_i;
  assign v1_data_o[374] = v0_data_i[374] & v0_en_i;
  assign v1_data_o[373] = v0_data_i[373] & v0_en_i;
  assign v1_data_o[372] = v0_data_i[372] & v0_en_i;
  assign v1_data_o[371] = v0_data_i[371] & v0_en_i;
  assign v1_data_o[370] = v0_data_i[370] & v0_en_i;
  assign v1_data_o[369] = v0_data_i[369] & v0_en_i;
  assign v1_data_o[368] = v0_data_i[368] & v0_en_i;
  assign v1_data_o[367] = v0_data_i[367] & v0_en_i;
  assign v1_data_o[366] = v0_data_i[366] & v0_en_i;
  assign v1_data_o[365] = v0_data_i[365] & v0_en_i;
  assign v1_data_o[364] = v0_data_i[364] & v0_en_i;
  assign v1_data_o[363] = v0_data_i[363] & v0_en_i;
  assign v1_data_o[362] = v0_data_i[362] & v0_en_i;
  assign v1_data_o[361] = v0_data_i[361] & v0_en_i;
  assign v1_data_o[360] = v0_data_i[360] & v0_en_i;
  assign v1_data_o[359] = v0_data_i[359] & v0_en_i;
  assign v1_data_o[358] = v0_data_i[358] & v0_en_i;
  assign v1_data_o[357] = v0_data_i[357] & v0_en_i;
  assign v1_data_o[356] = v0_data_i[356] & v0_en_i;
  assign v1_data_o[355] = v0_data_i[355] & v0_en_i;
  assign v1_data_o[354] = v0_data_i[354] & v0_en_i;
  assign v1_data_o[353] = v0_data_i[353] & v0_en_i;
  assign v1_data_o[352] = v0_data_i[352] & v0_en_i;
  assign v1_data_o[351] = v0_data_i[351] & v0_en_i;
  assign v1_data_o[350] = v0_data_i[350] & v0_en_i;
  assign v1_data_o[349] = v0_data_i[349] & v0_en_i;
  assign v1_data_o[348] = v0_data_i[348] & v0_en_i;
  assign v1_data_o[347] = v0_data_i[347] & v0_en_i;
  assign v1_data_o[346] = v0_data_i[346] & v0_en_i;
  assign v1_data_o[345] = v0_data_i[345] & v0_en_i;
  assign v1_data_o[344] = v0_data_i[344] & v0_en_i;
  assign v1_data_o[343] = v0_data_i[343] & v0_en_i;
  assign v1_data_o[342] = v0_data_i[342] & v0_en_i;
  assign v1_data_o[341] = v0_data_i[341] & v0_en_i;
  assign v1_data_o[340] = v0_data_i[340] & v0_en_i;
  assign v1_data_o[339] = v0_data_i[339] & v0_en_i;
  assign v1_data_o[338] = v0_data_i[338] & v0_en_i;
  assign v1_data_o[337] = v0_data_i[337] & v0_en_i;
  assign v1_data_o[336] = v0_data_i[336] & v0_en_i;
  assign v1_data_o[335] = v0_data_i[335] & v0_en_i;
  assign v1_data_o[334] = v0_data_i[334] & v0_en_i;
  assign v1_data_o[333] = v0_data_i[333] & v0_en_i;
  assign v1_data_o[332] = v0_data_i[332] & v0_en_i;
  assign v1_data_o[331] = v0_data_i[331] & v0_en_i;
  assign v1_data_o[330] = v0_data_i[330] & v0_en_i;
  assign v1_data_o[329] = v0_data_i[329] & v0_en_i;
  assign v1_data_o[328] = v0_data_i[328] & v0_en_i;
  assign v1_data_o[327] = v0_data_i[327] & v0_en_i;
  assign v1_data_o[326] = v0_data_i[326] & v0_en_i;
  assign v1_data_o[325] = v0_data_i[325] & v0_en_i;
  assign v1_data_o[324] = v0_data_i[324] & v0_en_i;
  assign v1_data_o[323] = v0_data_i[323] & v0_en_i;
  assign v1_data_o[322] = v0_data_i[322] & v0_en_i;
  assign v1_data_o[321] = v0_data_i[321] & v0_en_i;
  assign v1_data_o[320] = v0_data_i[320] & v0_en_i;
  assign v1_data_o[319] = v0_data_i[319] & v0_en_i;
  assign v1_data_o[318] = v0_data_i[318] & v0_en_i;
  assign v1_data_o[317] = v0_data_i[317] & v0_en_i;
  assign v1_data_o[316] = v0_data_i[316] & v0_en_i;
  assign v1_data_o[315] = v0_data_i[315] & v0_en_i;
  assign v1_data_o[314] = v0_data_i[314] & v0_en_i;
  assign v1_data_o[313] = v0_data_i[313] & v0_en_i;
  assign v1_data_o[312] = v0_data_i[312] & v0_en_i;
  assign v1_data_o[311] = v0_data_i[311] & v0_en_i;
  assign v1_data_o[310] = v0_data_i[310] & v0_en_i;
  assign v1_data_o[309] = v0_data_i[309] & v0_en_i;
  assign v1_data_o[308] = v0_data_i[308] & v0_en_i;
  assign v1_data_o[307] = v0_data_i[307] & v0_en_i;
  assign v1_data_o[306] = v0_data_i[306] & v0_en_i;
  assign v1_data_o[305] = v0_data_i[305] & v0_en_i;
  assign v1_data_o[304] = v0_data_i[304] & v0_en_i;
  assign v1_data_o[303] = v0_data_i[303] & v0_en_i;
  assign v1_data_o[302] = v0_data_i[302] & v0_en_i;
  assign v1_data_o[301] = v0_data_i[301] & v0_en_i;
  assign v1_data_o[300] = v0_data_i[300] & v0_en_i;
  assign v1_data_o[299] = v0_data_i[299] & v0_en_i;
  assign v1_data_o[298] = v0_data_i[298] & v0_en_i;
  assign v1_data_o[297] = v0_data_i[297] & v0_en_i;
  assign v1_data_o[296] = v0_data_i[296] & v0_en_i;
  assign v1_data_o[295] = v0_data_i[295] & v0_en_i;
  assign v1_data_o[294] = v0_data_i[294] & v0_en_i;
  assign v1_data_o[293] = v0_data_i[293] & v0_en_i;
  assign v1_data_o[292] = v0_data_i[292] & v0_en_i;
  assign v1_data_o[291] = v0_data_i[291] & v0_en_i;
  assign v1_data_o[290] = v0_data_i[290] & v0_en_i;
  assign v1_data_o[289] = v0_data_i[289] & v0_en_i;
  assign v1_data_o[288] = v0_data_i[288] & v0_en_i;
  assign v1_data_o[287] = v0_data_i[287] & v0_en_i;
  assign v1_data_o[286] = v0_data_i[286] & v0_en_i;
  assign v1_data_o[285] = v0_data_i[285] & v0_en_i;
  assign v1_data_o[284] = v0_data_i[284] & v0_en_i;
  assign v1_data_o[283] = v0_data_i[283] & v0_en_i;
  assign v1_data_o[282] = v0_data_i[282] & v0_en_i;
  assign v1_data_o[281] = v0_data_i[281] & v0_en_i;
  assign v1_data_o[280] = v0_data_i[280] & v0_en_i;
  assign v1_data_o[279] = v0_data_i[279] & v0_en_i;
  assign v1_data_o[278] = v0_data_i[278] & v0_en_i;
  assign v1_data_o[277] = v0_data_i[277] & v0_en_i;
  assign v1_data_o[276] = v0_data_i[276] & v0_en_i;
  assign v1_data_o[275] = v0_data_i[275] & v0_en_i;
  assign v1_data_o[274] = v0_data_i[274] & v0_en_i;
  assign v1_data_o[273] = v0_data_i[273] & v0_en_i;
  assign v1_data_o[272] = v0_data_i[272] & v0_en_i;
  assign v1_data_o[271] = v0_data_i[271] & v0_en_i;
  assign v1_data_o[270] = v0_data_i[270] & v0_en_i;
  assign v1_data_o[269] = v0_data_i[269] & v0_en_i;
  assign v1_data_o[268] = v0_data_i[268] & v0_en_i;
  assign v1_data_o[267] = v0_data_i[267] & v0_en_i;
  assign v1_data_o[266] = v0_data_i[266] & v0_en_i;
  assign v1_data_o[265] = v0_data_i[265] & v0_en_i;
  assign v1_data_o[264] = v0_data_i[264] & v0_en_i;
  assign v1_data_o[263] = v0_data_i[263] & v0_en_i;
  assign v1_data_o[262] = v0_data_i[262] & v0_en_i;
  assign v1_data_o[261] = v0_data_i[261] & v0_en_i;
  assign v1_data_o[260] = v0_data_i[260] & v0_en_i;
  assign v1_data_o[259] = v0_data_i[259] & v0_en_i;
  assign v1_data_o[258] = v0_data_i[258] & v0_en_i;
  assign v1_data_o[257] = v0_data_i[257] & v0_en_i;
  assign v1_data_o[256] = v0_data_i[256] & v0_en_i;
  assign v1_data_o[255] = v0_data_i[255] & v0_en_i;
  assign v1_data_o[254] = v0_data_i[254] & v0_en_i;
  assign v1_data_o[253] = v0_data_i[253] & v0_en_i;
  assign v1_data_o[252] = v0_data_i[252] & v0_en_i;
  assign v1_data_o[251] = v0_data_i[251] & v0_en_i;
  assign v1_data_o[250] = v0_data_i[250] & v0_en_i;
  assign v1_data_o[249] = v0_data_i[249] & v0_en_i;
  assign v1_data_o[248] = v0_data_i[248] & v0_en_i;
  assign v1_data_o[247] = v0_data_i[247] & v0_en_i;
  assign v1_data_o[246] = v0_data_i[246] & v0_en_i;
  assign v1_data_o[245] = v0_data_i[245] & v0_en_i;
  assign v1_data_o[244] = v0_data_i[244] & v0_en_i;
  assign v1_data_o[243] = v0_data_i[243] & v0_en_i;
  assign v1_data_o[242] = v0_data_i[242] & v0_en_i;
  assign v1_data_o[241] = v0_data_i[241] & v0_en_i;
  assign v1_data_o[240] = v0_data_i[240] & v0_en_i;
  assign v1_data_o[239] = v0_data_i[239] & v0_en_i;
  assign v1_data_o[238] = v0_data_i[238] & v0_en_i;
  assign v1_data_o[237] = v0_data_i[237] & v0_en_i;
  assign v1_data_o[236] = v0_data_i[236] & v0_en_i;
  assign v1_data_o[235] = v0_data_i[235] & v0_en_i;
  assign v1_data_o[234] = v0_data_i[234] & v0_en_i;
  assign v1_data_o[233] = v0_data_i[233] & v0_en_i;
  assign v1_data_o[232] = v0_data_i[232] & v0_en_i;
  assign v1_data_o[231] = v0_data_i[231] & v0_en_i;
  assign v1_data_o[230] = v0_data_i[230] & v0_en_i;
  assign v1_data_o[229] = v0_data_i[229] & v0_en_i;
  assign v1_data_o[228] = v0_data_i[228] & v0_en_i;
  assign v1_data_o[227] = v0_data_i[227] & v0_en_i;
  assign v1_data_o[226] = v0_data_i[226] & v0_en_i;
  assign v1_data_o[225] = v0_data_i[225] & v0_en_i;
  assign v1_data_o[224] = v0_data_i[224] & v0_en_i;
  assign v1_data_o[223] = v0_data_i[223] & v0_en_i;
  assign v1_data_o[222] = v0_data_i[222] & v0_en_i;
  assign v1_data_o[221] = v0_data_i[221] & v0_en_i;
  assign v1_data_o[220] = v0_data_i[220] & v0_en_i;
  assign v1_data_o[219] = v0_data_i[219] & v0_en_i;
  assign v1_data_o[218] = v0_data_i[218] & v0_en_i;
  assign v1_data_o[217] = v0_data_i[217] & v0_en_i;
  assign v1_data_o[216] = v0_data_i[216] & v0_en_i;
  assign v1_data_o[215] = v0_data_i[215] & v0_en_i;
  assign v1_data_o[214] = v0_data_i[214] & v0_en_i;
  assign v1_data_o[213] = v0_data_i[213] & v0_en_i;
  assign v1_data_o[212] = v0_data_i[212] & v0_en_i;
  assign v1_data_o[211] = v0_data_i[211] & v0_en_i;
  assign v1_data_o[210] = v0_data_i[210] & v0_en_i;
  assign v1_data_o[209] = v0_data_i[209] & v0_en_i;
  assign v1_data_o[208] = v0_data_i[208] & v0_en_i;
  assign v1_data_o[207] = v0_data_i[207] & v0_en_i;
  assign v1_data_o[206] = v0_data_i[206] & v0_en_i;
  assign v1_data_o[205] = v0_data_i[205] & v0_en_i;
  assign v1_data_o[204] = v0_data_i[204] & v0_en_i;
  assign v1_data_o[203] = v0_data_i[203] & v0_en_i;
  assign v1_data_o[202] = v0_data_i[202] & v0_en_i;
  assign v1_data_o[201] = v0_data_i[201] & v0_en_i;
  assign v1_data_o[200] = v0_data_i[200] & v0_en_i;
  assign v1_data_o[199] = v0_data_i[199] & v0_en_i;
  assign v1_data_o[198] = v0_data_i[198] & v0_en_i;
  assign v1_data_o[197] = v0_data_i[197] & v0_en_i;
  assign v1_data_o[196] = v0_data_i[196] & v0_en_i;
  assign v1_data_o[195] = v0_data_i[195] & v0_en_i;
  assign v1_data_o[194] = v0_data_i[194] & v0_en_i;
  assign v1_data_o[193] = v0_data_i[193] & v0_en_i;
  assign v1_data_o[192] = v0_data_i[192] & v0_en_i;
  assign v1_data_o[191] = v0_data_i[191] & v0_en_i;
  assign v1_data_o[190] = v0_data_i[190] & v0_en_i;
  assign v1_data_o[189] = v0_data_i[189] & v0_en_i;
  assign v1_data_o[188] = v0_data_i[188] & v0_en_i;
  assign v1_data_o[187] = v0_data_i[187] & v0_en_i;
  assign v1_data_o[186] = v0_data_i[186] & v0_en_i;
  assign v1_data_o[185] = v0_data_i[185] & v0_en_i;
  assign v1_data_o[184] = v0_data_i[184] & v0_en_i;
  assign v1_data_o[183] = v0_data_i[183] & v0_en_i;
  assign v1_data_o[182] = v0_data_i[182] & v0_en_i;
  assign v1_data_o[181] = v0_data_i[181] & v0_en_i;
  assign v1_data_o[180] = v0_data_i[180] & v0_en_i;
  assign v1_data_o[179] = v0_data_i[179] & v0_en_i;
  assign v1_data_o[178] = v0_data_i[178] & v0_en_i;
  assign v1_data_o[177] = v0_data_i[177] & v0_en_i;
  assign v1_data_o[176] = v0_data_i[176] & v0_en_i;
  assign v1_data_o[175] = v0_data_i[175] & v0_en_i;
  assign v1_data_o[174] = v0_data_i[174] & v0_en_i;
  assign v1_data_o[173] = v0_data_i[173] & v0_en_i;
  assign v1_data_o[172] = v0_data_i[172] & v0_en_i;
  assign v1_data_o[171] = v0_data_i[171] & v0_en_i;
  assign v1_data_o[170] = v0_data_i[170] & v0_en_i;
  assign v1_data_o[169] = v0_data_i[169] & v0_en_i;
  assign v1_data_o[168] = v0_data_i[168] & v0_en_i;
  assign v1_data_o[167] = v0_data_i[167] & v0_en_i;
  assign v1_data_o[166] = v0_data_i[166] & v0_en_i;
  assign v1_data_o[165] = v0_data_i[165] & v0_en_i;
  assign v1_data_o[164] = v0_data_i[164] & v0_en_i;
  assign v1_data_o[163] = v0_data_i[163] & v0_en_i;
  assign v1_data_o[162] = v0_data_i[162] & v0_en_i;
  assign v1_data_o[161] = v0_data_i[161] & v0_en_i;
  assign v1_data_o[160] = v0_data_i[160] & v0_en_i;
  assign v1_data_o[159] = v0_data_i[159] & v0_en_i;
  assign v1_data_o[158] = v0_data_i[158] & v0_en_i;
  assign v1_data_o[157] = v0_data_i[157] & v0_en_i;
  assign v1_data_o[156] = v0_data_i[156] & v0_en_i;
  assign v1_data_o[155] = v0_data_i[155] & v0_en_i;
  assign v1_data_o[154] = v0_data_i[154] & v0_en_i;
  assign v1_data_o[153] = v0_data_i[153] & v0_en_i;
  assign v1_data_o[152] = v0_data_i[152] & v0_en_i;
  assign v1_data_o[151] = v0_data_i[151] & v0_en_i;
  assign v1_data_o[150] = v0_data_i[150] & v0_en_i;
  assign v1_data_o[149] = v0_data_i[149] & v0_en_i;
  assign v1_data_o[148] = v0_data_i[148] & v0_en_i;
  assign v1_data_o[147] = v0_data_i[147] & v0_en_i;
  assign v1_data_o[146] = v0_data_i[146] & v0_en_i;
  assign v1_data_o[145] = v0_data_i[145] & v0_en_i;
  assign v1_data_o[144] = v0_data_i[144] & v0_en_i;
  assign v1_data_o[143] = v0_data_i[143] & v0_en_i;
  assign v1_data_o[142] = v0_data_i[142] & v0_en_i;
  assign v1_data_o[141] = v0_data_i[141] & v0_en_i;
  assign v1_data_o[140] = v0_data_i[140] & v0_en_i;
  assign v1_data_o[139] = v0_data_i[139] & v0_en_i;
  assign v1_data_o[138] = v0_data_i[138] & v0_en_i;
  assign v1_data_o[137] = v0_data_i[137] & v0_en_i;
  assign v1_data_o[136] = v0_data_i[136] & v0_en_i;
  assign v1_data_o[135] = v0_data_i[135] & v0_en_i;
  assign v1_data_o[134] = v0_data_i[134] & v0_en_i;
  assign v1_data_o[133] = v0_data_i[133] & v0_en_i;
  assign v1_data_o[132] = v0_data_i[132] & v0_en_i;
  assign v1_data_o[131] = v0_data_i[131] & v0_en_i;
  assign v1_data_o[130] = v0_data_i[130] & v0_en_i;
  assign v1_data_o[129] = v0_data_i[129] & v0_en_i;
  assign v1_data_o[128] = v0_data_i[128] & v0_en_i;
  assign v1_data_o[127] = v0_data_i[127] & v0_en_i;
  assign v1_data_o[126] = v0_data_i[126] & v0_en_i;
  assign v1_data_o[125] = v0_data_i[125] & v0_en_i;
  assign v1_data_o[124] = v0_data_i[124] & v0_en_i;
  assign v1_data_o[123] = v0_data_i[123] & v0_en_i;
  assign v1_data_o[122] = v0_data_i[122] & v0_en_i;
  assign v1_data_o[121] = v0_data_i[121] & v0_en_i;
  assign v1_data_o[120] = v0_data_i[120] & v0_en_i;
  assign v1_data_o[119] = v0_data_i[119] & v0_en_i;
  assign v1_data_o[118] = v0_data_i[118] & v0_en_i;
  assign v1_data_o[117] = v0_data_i[117] & v0_en_i;
  assign v1_data_o[116] = v0_data_i[116] & v0_en_i;
  assign v1_data_o[115] = v0_data_i[115] & v0_en_i;
  assign v1_data_o[114] = v0_data_i[114] & v0_en_i;
  assign v1_data_o[113] = v0_data_i[113] & v0_en_i;
  assign v1_data_o[112] = v0_data_i[112] & v0_en_i;
  assign v1_data_o[111] = v0_data_i[111] & v0_en_i;
  assign v1_data_o[110] = v0_data_i[110] & v0_en_i;
  assign v1_data_o[109] = v0_data_i[109] & v0_en_i;
  assign v1_data_o[108] = v0_data_i[108] & v0_en_i;
  assign v1_data_o[107] = v0_data_i[107] & v0_en_i;
  assign v1_data_o[106] = v0_data_i[106] & v0_en_i;
  assign v1_data_o[105] = v0_data_i[105] & v0_en_i;
  assign v1_data_o[104] = v0_data_i[104] & v0_en_i;
  assign v1_data_o[103] = v0_data_i[103] & v0_en_i;
  assign v1_data_o[102] = v0_data_i[102] & v0_en_i;
  assign v1_data_o[101] = v0_data_i[101] & v0_en_i;
  assign v1_data_o[100] = v0_data_i[100] & v0_en_i;
  assign v1_data_o[99] = v0_data_i[99] & v0_en_i;
  assign v1_data_o[98] = v0_data_i[98] & v0_en_i;
  assign v1_data_o[97] = v0_data_i[97] & v0_en_i;
  assign v1_data_o[96] = v0_data_i[96] & v0_en_i;
  assign v1_data_o[95] = v0_data_i[95] & v0_en_i;
  assign v1_data_o[94] = v0_data_i[94] & v0_en_i;
  assign v1_data_o[93] = v0_data_i[93] & v0_en_i;
  assign v1_data_o[92] = v0_data_i[92] & v0_en_i;
  assign v1_data_o[91] = v0_data_i[91] & v0_en_i;
  assign v1_data_o[90] = v0_data_i[90] & v0_en_i;
  assign v1_data_o[89] = v0_data_i[89] & v0_en_i;
  assign v1_data_o[88] = v0_data_i[88] & v0_en_i;
  assign v1_data_o[87] = v0_data_i[87] & v0_en_i;
  assign v1_data_o[86] = v0_data_i[86] & v0_en_i;
  assign v1_data_o[85] = v0_data_i[85] & v0_en_i;
  assign v1_data_o[84] = v0_data_i[84] & v0_en_i;
  assign v1_data_o[83] = v0_data_i[83] & v0_en_i;
  assign v1_data_o[82] = v0_data_i[82] & v0_en_i;
  assign v1_data_o[81] = v0_data_i[81] & v0_en_i;
  assign v1_data_o[80] = v0_data_i[80] & v0_en_i;
  assign v1_data_o[79] = v0_data_i[79] & v0_en_i;
  assign v1_data_o[78] = v0_data_i[78] & v0_en_i;
  assign v1_data_o[77] = v0_data_i[77] & v0_en_i;
  assign v1_data_o[76] = v0_data_i[76] & v0_en_i;
  assign v1_data_o[75] = v0_data_i[75] & v0_en_i;
  assign v1_data_o[74] = v0_data_i[74] & v0_en_i;
  assign v1_data_o[73] = v0_data_i[73] & v0_en_i;
  assign v1_data_o[72] = v0_data_i[72] & v0_en_i;
  assign v1_data_o[71] = v0_data_i[71] & v0_en_i;
  assign v1_data_o[70] = v0_data_i[70] & v0_en_i;
  assign v1_data_o[69] = v0_data_i[69] & v0_en_i;
  assign v1_data_o[68] = v0_data_i[68] & v0_en_i;
  assign v1_data_o[67] = v0_data_i[67] & v0_en_i;
  assign v1_data_o[66] = v0_data_i[66] & v0_en_i;
  assign v1_data_o[65] = v0_data_i[65] & v0_en_i;
  assign v1_data_o[64] = v0_data_i[64] & v0_en_i;
  assign v1_data_o[63] = v0_data_i[63] & v0_en_i;
  assign v1_data_o[62] = v0_data_i[62] & v0_en_i;
  assign v1_data_o[61] = v0_data_i[61] & v0_en_i;
  assign v1_data_o[60] = v0_data_i[60] & v0_en_i;
  assign v1_data_o[59] = v0_data_i[59] & v0_en_i;
  assign v1_data_o[58] = v0_data_i[58] & v0_en_i;
  assign v1_data_o[57] = v0_data_i[57] & v0_en_i;
  assign v1_data_o[56] = v0_data_i[56] & v0_en_i;
  assign v1_data_o[55] = v0_data_i[55] & v0_en_i;
  assign v1_data_o[54] = v0_data_i[54] & v0_en_i;
  assign v1_data_o[53] = v0_data_i[53] & v0_en_i;
  assign v1_data_o[52] = v0_data_i[52] & v0_en_i;
  assign v1_data_o[51] = v0_data_i[51] & v0_en_i;
  assign v1_data_o[50] = v0_data_i[50] & v0_en_i;
  assign v1_data_o[49] = v0_data_i[49] & v0_en_i;
  assign v1_data_o[48] = v0_data_i[48] & v0_en_i;
  assign v1_data_o[47] = v0_data_i[47] & v0_en_i;
  assign v1_data_o[46] = v0_data_i[46] & v0_en_i;
  assign v1_data_o[45] = v0_data_i[45] & v0_en_i;
  assign v1_data_o[44] = v0_data_i[44] & v0_en_i;
  assign v1_data_o[43] = v0_data_i[43] & v0_en_i;
  assign v1_data_o[42] = v0_data_i[42] & v0_en_i;
  assign v1_data_o[41] = v0_data_i[41] & v0_en_i;
  assign v1_data_o[40] = v0_data_i[40] & v0_en_i;
  assign v1_data_o[39] = v0_data_i[39] & v0_en_i;
  assign v1_data_o[38] = v0_data_i[38] & v0_en_i;
  assign v1_data_o[37] = v0_data_i[37] & v0_en_i;
  assign v1_data_o[36] = v0_data_i[36] & v0_en_i;
  assign v1_data_o[35] = v0_data_i[35] & v0_en_i;
  assign v1_data_o[34] = v0_data_i[34] & v0_en_i;
  assign v1_data_o[33] = v0_data_i[33] & v0_en_i;
  assign v1_data_o[32] = v0_data_i[32] & v0_en_i;
  assign v1_data_o[31] = v0_data_i[31] & v0_en_i;
  assign v1_data_o[30] = v0_data_i[30] & v0_en_i;
  assign v1_data_o[29] = v0_data_i[29] & v0_en_i;
  assign v1_data_o[28] = v0_data_i[28] & v0_en_i;
  assign v1_data_o[27] = v0_data_i[27] & v0_en_i;
  assign v1_data_o[26] = v0_data_i[26] & v0_en_i;
  assign v1_data_o[25] = v0_data_i[25] & v0_en_i;
  assign v1_data_o[24] = v0_data_i[24] & v0_en_i;
  assign v1_data_o[23] = v0_data_i[23] & v0_en_i;
  assign v1_data_o[22] = v0_data_i[22] & v0_en_i;
  assign v1_data_o[21] = v0_data_i[21] & v0_en_i;
  assign v1_data_o[20] = v0_data_i[20] & v0_en_i;
  assign v1_data_o[19] = v0_data_i[19] & v0_en_i;
  assign v1_data_o[18] = v0_data_i[18] & v0_en_i;
  assign v1_data_o[17] = v0_data_i[17] & v0_en_i;
  assign v1_data_o[16] = v0_data_i[16] & v0_en_i;
  assign v1_data_o[15] = v0_data_i[15] & v0_en_i;
  assign v1_data_o[14] = v0_data_i[14] & v0_en_i;
  assign v1_data_o[13] = v0_data_i[13] & v0_en_i;
  assign v1_data_o[12] = v0_data_i[12] & v0_en_i;
  assign v1_data_o[11] = v0_data_i[11] & v0_en_i;
  assign v1_data_o[10] = v0_data_i[10] & v0_en_i;
  assign v1_data_o[9] = v0_data_i[9] & v0_en_i;
  assign v1_data_o[8] = v0_data_i[8] & v0_en_i;
  assign v1_data_o[7] = v0_data_i[7] & v0_en_i;
  assign v1_data_o[6] = v0_data_i[6] & v0_en_i;
  assign v1_data_o[5] = v0_data_i[5] & v0_en_i;
  assign v1_data_o[4] = v0_data_i[4] & v0_en_i;
  assign v1_data_o[3] = v0_data_i[3] & v0_en_i;
  assign v1_data_o[2] = v0_data_i[2] & v0_en_i;
  assign v1_data_o[1] = v0_data_i[1] & v0_en_i;
  assign v1_data_o[0] = v0_data_i[0] & v0_en_i;

endmodule



module bsg_fsb_node_level_shift_fsb_domain
(
  en_ls_i,
  clk_i,
  reset_i,
  clk_o,
  reset_o,
  fsb_v_i_o,
  fsb_data_i_o,
  fsb_yumi_o_i,
  fsb_v_o_i,
  fsb_data_o_i,
  fsb_ready_i_o,
  node_v_i_o,
  node_data_i_o,
  node_ready_o_i,
  node_v_o_i,
  node_data_o_i,
  node_yumi_i_o
);

  output [499:0] fsb_data_i_o;
  input [499:0] fsb_data_o_i;
  output [499:0] node_data_i_o;
  input [499:0] node_data_o_i;
  input en_ls_i;
  input clk_i;
  input reset_i;
  input fsb_yumi_o_i;
  input fsb_v_o_i;
  input node_ready_o_i;
  input node_v_o_i;
  output clk_o;
  output reset_o;
  output fsb_v_i_o;
  output fsb_ready_i_o;
  output node_v_i_o;
  output node_yumi_i_o;
  wire [499:0] fsb_data_i_o,node_data_i_o;
  wire clk_o,reset_o,fsb_v_i_o,fsb_ready_i_o,node_v_i_o,node_yumi_i_o;

  bsg_level_shift_up_down_source_width_p1
  clk_ls_inst
  (
    .v0_en_i(1'b1),
    .v0_data_i(clk_i),
    .v1_data_o(clk_o)
  );


  bsg_level_shift_up_down_source_width_p1
  reset_ls_inst
  (
    .v0_en_i(1'b1),
    .v0_data_i(reset_i),
    .v1_data_o(reset_o)
  );


  bsg_level_shift_up_down_sink_width_p1
  n2f_v_ls_inst
  (
    .v0_data_i(node_v_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(fsb_v_i_o)
  );


  bsg_level_shift_up_down_sink_width_p500
  n2f_data_ls_inst
  (
    .v0_data_i(node_data_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(fsb_data_i_o)
  );


  bsg_level_shift_up_down_source_width_p1
  f2n_yumi_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(fsb_yumi_o_i),
    .v1_data_o(node_yumi_i_o)
  );


  bsg_level_shift_up_down_source_width_p1
  f2n_v_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(fsb_v_o_i),
    .v1_data_o(node_v_i_o)
  );


  bsg_level_shift_up_down_source_width_p500
  f2n_data_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(fsb_data_o_i),
    .v1_data_o(node_data_i_o)
  );


  bsg_level_shift_up_down_sink_width_p1
  n2f_ready_ls_inst
  (
    .v0_data_i(node_ready_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(fsb_ready_i_o)
  );


endmodule

