

module top
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_i
);

  input [2047:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_o;
  output valid_o;

  bsg_parallel_in_serial_out
  wrapper
  (
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .valid_i(valid_i),
    .yumi_i(yumi_i),
    .ready_o(ready_o),
    .valid_o(valid_o)
  );


endmodule



module bsg_array_reverse_width_p32_els_p64
(
  i,
  o
);

  input [2047:0] i;
  output [2047:0] o;
  wire [2047:0] o;
  assign o[2047] = i[31];
  assign o[2046] = i[30];
  assign o[2045] = i[29];
  assign o[2044] = i[28];
  assign o[2043] = i[27];
  assign o[2042] = i[26];
  assign o[2041] = i[25];
  assign o[2040] = i[24];
  assign o[2039] = i[23];
  assign o[2038] = i[22];
  assign o[2037] = i[21];
  assign o[2036] = i[20];
  assign o[2035] = i[19];
  assign o[2034] = i[18];
  assign o[2033] = i[17];
  assign o[2032] = i[16];
  assign o[2031] = i[15];
  assign o[2030] = i[14];
  assign o[2029] = i[13];
  assign o[2028] = i[12];
  assign o[2027] = i[11];
  assign o[2026] = i[10];
  assign o[2025] = i[9];
  assign o[2024] = i[8];
  assign o[2023] = i[7];
  assign o[2022] = i[6];
  assign o[2021] = i[5];
  assign o[2020] = i[4];
  assign o[2019] = i[3];
  assign o[2018] = i[2];
  assign o[2017] = i[1];
  assign o[2016] = i[0];
  assign o[2015] = i[63];
  assign o[2014] = i[62];
  assign o[2013] = i[61];
  assign o[2012] = i[60];
  assign o[2011] = i[59];
  assign o[2010] = i[58];
  assign o[2009] = i[57];
  assign o[2008] = i[56];
  assign o[2007] = i[55];
  assign o[2006] = i[54];
  assign o[2005] = i[53];
  assign o[2004] = i[52];
  assign o[2003] = i[51];
  assign o[2002] = i[50];
  assign o[2001] = i[49];
  assign o[2000] = i[48];
  assign o[1999] = i[47];
  assign o[1998] = i[46];
  assign o[1997] = i[45];
  assign o[1996] = i[44];
  assign o[1995] = i[43];
  assign o[1994] = i[42];
  assign o[1993] = i[41];
  assign o[1992] = i[40];
  assign o[1991] = i[39];
  assign o[1990] = i[38];
  assign o[1989] = i[37];
  assign o[1988] = i[36];
  assign o[1987] = i[35];
  assign o[1986] = i[34];
  assign o[1985] = i[33];
  assign o[1984] = i[32];
  assign o[1983] = i[95];
  assign o[1982] = i[94];
  assign o[1981] = i[93];
  assign o[1980] = i[92];
  assign o[1979] = i[91];
  assign o[1978] = i[90];
  assign o[1977] = i[89];
  assign o[1976] = i[88];
  assign o[1975] = i[87];
  assign o[1974] = i[86];
  assign o[1973] = i[85];
  assign o[1972] = i[84];
  assign o[1971] = i[83];
  assign o[1970] = i[82];
  assign o[1969] = i[81];
  assign o[1968] = i[80];
  assign o[1967] = i[79];
  assign o[1966] = i[78];
  assign o[1965] = i[77];
  assign o[1964] = i[76];
  assign o[1963] = i[75];
  assign o[1962] = i[74];
  assign o[1961] = i[73];
  assign o[1960] = i[72];
  assign o[1959] = i[71];
  assign o[1958] = i[70];
  assign o[1957] = i[69];
  assign o[1956] = i[68];
  assign o[1955] = i[67];
  assign o[1954] = i[66];
  assign o[1953] = i[65];
  assign o[1952] = i[64];
  assign o[1951] = i[127];
  assign o[1950] = i[126];
  assign o[1949] = i[125];
  assign o[1948] = i[124];
  assign o[1947] = i[123];
  assign o[1946] = i[122];
  assign o[1945] = i[121];
  assign o[1944] = i[120];
  assign o[1943] = i[119];
  assign o[1942] = i[118];
  assign o[1941] = i[117];
  assign o[1940] = i[116];
  assign o[1939] = i[115];
  assign o[1938] = i[114];
  assign o[1937] = i[113];
  assign o[1936] = i[112];
  assign o[1935] = i[111];
  assign o[1934] = i[110];
  assign o[1933] = i[109];
  assign o[1932] = i[108];
  assign o[1931] = i[107];
  assign o[1930] = i[106];
  assign o[1929] = i[105];
  assign o[1928] = i[104];
  assign o[1927] = i[103];
  assign o[1926] = i[102];
  assign o[1925] = i[101];
  assign o[1924] = i[100];
  assign o[1923] = i[99];
  assign o[1922] = i[98];
  assign o[1921] = i[97];
  assign o[1920] = i[96];
  assign o[1919] = i[159];
  assign o[1918] = i[158];
  assign o[1917] = i[157];
  assign o[1916] = i[156];
  assign o[1915] = i[155];
  assign o[1914] = i[154];
  assign o[1913] = i[153];
  assign o[1912] = i[152];
  assign o[1911] = i[151];
  assign o[1910] = i[150];
  assign o[1909] = i[149];
  assign o[1908] = i[148];
  assign o[1907] = i[147];
  assign o[1906] = i[146];
  assign o[1905] = i[145];
  assign o[1904] = i[144];
  assign o[1903] = i[143];
  assign o[1902] = i[142];
  assign o[1901] = i[141];
  assign o[1900] = i[140];
  assign o[1899] = i[139];
  assign o[1898] = i[138];
  assign o[1897] = i[137];
  assign o[1896] = i[136];
  assign o[1895] = i[135];
  assign o[1894] = i[134];
  assign o[1893] = i[133];
  assign o[1892] = i[132];
  assign o[1891] = i[131];
  assign o[1890] = i[130];
  assign o[1889] = i[129];
  assign o[1888] = i[128];
  assign o[1887] = i[191];
  assign o[1886] = i[190];
  assign o[1885] = i[189];
  assign o[1884] = i[188];
  assign o[1883] = i[187];
  assign o[1882] = i[186];
  assign o[1881] = i[185];
  assign o[1880] = i[184];
  assign o[1879] = i[183];
  assign o[1878] = i[182];
  assign o[1877] = i[181];
  assign o[1876] = i[180];
  assign o[1875] = i[179];
  assign o[1874] = i[178];
  assign o[1873] = i[177];
  assign o[1872] = i[176];
  assign o[1871] = i[175];
  assign o[1870] = i[174];
  assign o[1869] = i[173];
  assign o[1868] = i[172];
  assign o[1867] = i[171];
  assign o[1866] = i[170];
  assign o[1865] = i[169];
  assign o[1864] = i[168];
  assign o[1863] = i[167];
  assign o[1862] = i[166];
  assign o[1861] = i[165];
  assign o[1860] = i[164];
  assign o[1859] = i[163];
  assign o[1858] = i[162];
  assign o[1857] = i[161];
  assign o[1856] = i[160];
  assign o[1855] = i[223];
  assign o[1854] = i[222];
  assign o[1853] = i[221];
  assign o[1852] = i[220];
  assign o[1851] = i[219];
  assign o[1850] = i[218];
  assign o[1849] = i[217];
  assign o[1848] = i[216];
  assign o[1847] = i[215];
  assign o[1846] = i[214];
  assign o[1845] = i[213];
  assign o[1844] = i[212];
  assign o[1843] = i[211];
  assign o[1842] = i[210];
  assign o[1841] = i[209];
  assign o[1840] = i[208];
  assign o[1839] = i[207];
  assign o[1838] = i[206];
  assign o[1837] = i[205];
  assign o[1836] = i[204];
  assign o[1835] = i[203];
  assign o[1834] = i[202];
  assign o[1833] = i[201];
  assign o[1832] = i[200];
  assign o[1831] = i[199];
  assign o[1830] = i[198];
  assign o[1829] = i[197];
  assign o[1828] = i[196];
  assign o[1827] = i[195];
  assign o[1826] = i[194];
  assign o[1825] = i[193];
  assign o[1824] = i[192];
  assign o[1823] = i[255];
  assign o[1822] = i[254];
  assign o[1821] = i[253];
  assign o[1820] = i[252];
  assign o[1819] = i[251];
  assign o[1818] = i[250];
  assign o[1817] = i[249];
  assign o[1816] = i[248];
  assign o[1815] = i[247];
  assign o[1814] = i[246];
  assign o[1813] = i[245];
  assign o[1812] = i[244];
  assign o[1811] = i[243];
  assign o[1810] = i[242];
  assign o[1809] = i[241];
  assign o[1808] = i[240];
  assign o[1807] = i[239];
  assign o[1806] = i[238];
  assign o[1805] = i[237];
  assign o[1804] = i[236];
  assign o[1803] = i[235];
  assign o[1802] = i[234];
  assign o[1801] = i[233];
  assign o[1800] = i[232];
  assign o[1799] = i[231];
  assign o[1798] = i[230];
  assign o[1797] = i[229];
  assign o[1796] = i[228];
  assign o[1795] = i[227];
  assign o[1794] = i[226];
  assign o[1793] = i[225];
  assign o[1792] = i[224];
  assign o[1791] = i[287];
  assign o[1790] = i[286];
  assign o[1789] = i[285];
  assign o[1788] = i[284];
  assign o[1787] = i[283];
  assign o[1786] = i[282];
  assign o[1785] = i[281];
  assign o[1784] = i[280];
  assign o[1783] = i[279];
  assign o[1782] = i[278];
  assign o[1781] = i[277];
  assign o[1780] = i[276];
  assign o[1779] = i[275];
  assign o[1778] = i[274];
  assign o[1777] = i[273];
  assign o[1776] = i[272];
  assign o[1775] = i[271];
  assign o[1774] = i[270];
  assign o[1773] = i[269];
  assign o[1772] = i[268];
  assign o[1771] = i[267];
  assign o[1770] = i[266];
  assign o[1769] = i[265];
  assign o[1768] = i[264];
  assign o[1767] = i[263];
  assign o[1766] = i[262];
  assign o[1765] = i[261];
  assign o[1764] = i[260];
  assign o[1763] = i[259];
  assign o[1762] = i[258];
  assign o[1761] = i[257];
  assign o[1760] = i[256];
  assign o[1759] = i[319];
  assign o[1758] = i[318];
  assign o[1757] = i[317];
  assign o[1756] = i[316];
  assign o[1755] = i[315];
  assign o[1754] = i[314];
  assign o[1753] = i[313];
  assign o[1752] = i[312];
  assign o[1751] = i[311];
  assign o[1750] = i[310];
  assign o[1749] = i[309];
  assign o[1748] = i[308];
  assign o[1747] = i[307];
  assign o[1746] = i[306];
  assign o[1745] = i[305];
  assign o[1744] = i[304];
  assign o[1743] = i[303];
  assign o[1742] = i[302];
  assign o[1741] = i[301];
  assign o[1740] = i[300];
  assign o[1739] = i[299];
  assign o[1738] = i[298];
  assign o[1737] = i[297];
  assign o[1736] = i[296];
  assign o[1735] = i[295];
  assign o[1734] = i[294];
  assign o[1733] = i[293];
  assign o[1732] = i[292];
  assign o[1731] = i[291];
  assign o[1730] = i[290];
  assign o[1729] = i[289];
  assign o[1728] = i[288];
  assign o[1727] = i[351];
  assign o[1726] = i[350];
  assign o[1725] = i[349];
  assign o[1724] = i[348];
  assign o[1723] = i[347];
  assign o[1722] = i[346];
  assign o[1721] = i[345];
  assign o[1720] = i[344];
  assign o[1719] = i[343];
  assign o[1718] = i[342];
  assign o[1717] = i[341];
  assign o[1716] = i[340];
  assign o[1715] = i[339];
  assign o[1714] = i[338];
  assign o[1713] = i[337];
  assign o[1712] = i[336];
  assign o[1711] = i[335];
  assign o[1710] = i[334];
  assign o[1709] = i[333];
  assign o[1708] = i[332];
  assign o[1707] = i[331];
  assign o[1706] = i[330];
  assign o[1705] = i[329];
  assign o[1704] = i[328];
  assign o[1703] = i[327];
  assign o[1702] = i[326];
  assign o[1701] = i[325];
  assign o[1700] = i[324];
  assign o[1699] = i[323];
  assign o[1698] = i[322];
  assign o[1697] = i[321];
  assign o[1696] = i[320];
  assign o[1695] = i[383];
  assign o[1694] = i[382];
  assign o[1693] = i[381];
  assign o[1692] = i[380];
  assign o[1691] = i[379];
  assign o[1690] = i[378];
  assign o[1689] = i[377];
  assign o[1688] = i[376];
  assign o[1687] = i[375];
  assign o[1686] = i[374];
  assign o[1685] = i[373];
  assign o[1684] = i[372];
  assign o[1683] = i[371];
  assign o[1682] = i[370];
  assign o[1681] = i[369];
  assign o[1680] = i[368];
  assign o[1679] = i[367];
  assign o[1678] = i[366];
  assign o[1677] = i[365];
  assign o[1676] = i[364];
  assign o[1675] = i[363];
  assign o[1674] = i[362];
  assign o[1673] = i[361];
  assign o[1672] = i[360];
  assign o[1671] = i[359];
  assign o[1670] = i[358];
  assign o[1669] = i[357];
  assign o[1668] = i[356];
  assign o[1667] = i[355];
  assign o[1666] = i[354];
  assign o[1665] = i[353];
  assign o[1664] = i[352];
  assign o[1663] = i[415];
  assign o[1662] = i[414];
  assign o[1661] = i[413];
  assign o[1660] = i[412];
  assign o[1659] = i[411];
  assign o[1658] = i[410];
  assign o[1657] = i[409];
  assign o[1656] = i[408];
  assign o[1655] = i[407];
  assign o[1654] = i[406];
  assign o[1653] = i[405];
  assign o[1652] = i[404];
  assign o[1651] = i[403];
  assign o[1650] = i[402];
  assign o[1649] = i[401];
  assign o[1648] = i[400];
  assign o[1647] = i[399];
  assign o[1646] = i[398];
  assign o[1645] = i[397];
  assign o[1644] = i[396];
  assign o[1643] = i[395];
  assign o[1642] = i[394];
  assign o[1641] = i[393];
  assign o[1640] = i[392];
  assign o[1639] = i[391];
  assign o[1638] = i[390];
  assign o[1637] = i[389];
  assign o[1636] = i[388];
  assign o[1635] = i[387];
  assign o[1634] = i[386];
  assign o[1633] = i[385];
  assign o[1632] = i[384];
  assign o[1631] = i[447];
  assign o[1630] = i[446];
  assign o[1629] = i[445];
  assign o[1628] = i[444];
  assign o[1627] = i[443];
  assign o[1626] = i[442];
  assign o[1625] = i[441];
  assign o[1624] = i[440];
  assign o[1623] = i[439];
  assign o[1622] = i[438];
  assign o[1621] = i[437];
  assign o[1620] = i[436];
  assign o[1619] = i[435];
  assign o[1618] = i[434];
  assign o[1617] = i[433];
  assign o[1616] = i[432];
  assign o[1615] = i[431];
  assign o[1614] = i[430];
  assign o[1613] = i[429];
  assign o[1612] = i[428];
  assign o[1611] = i[427];
  assign o[1610] = i[426];
  assign o[1609] = i[425];
  assign o[1608] = i[424];
  assign o[1607] = i[423];
  assign o[1606] = i[422];
  assign o[1605] = i[421];
  assign o[1604] = i[420];
  assign o[1603] = i[419];
  assign o[1602] = i[418];
  assign o[1601] = i[417];
  assign o[1600] = i[416];
  assign o[1599] = i[479];
  assign o[1598] = i[478];
  assign o[1597] = i[477];
  assign o[1596] = i[476];
  assign o[1595] = i[475];
  assign o[1594] = i[474];
  assign o[1593] = i[473];
  assign o[1592] = i[472];
  assign o[1591] = i[471];
  assign o[1590] = i[470];
  assign o[1589] = i[469];
  assign o[1588] = i[468];
  assign o[1587] = i[467];
  assign o[1586] = i[466];
  assign o[1585] = i[465];
  assign o[1584] = i[464];
  assign o[1583] = i[463];
  assign o[1582] = i[462];
  assign o[1581] = i[461];
  assign o[1580] = i[460];
  assign o[1579] = i[459];
  assign o[1578] = i[458];
  assign o[1577] = i[457];
  assign o[1576] = i[456];
  assign o[1575] = i[455];
  assign o[1574] = i[454];
  assign o[1573] = i[453];
  assign o[1572] = i[452];
  assign o[1571] = i[451];
  assign o[1570] = i[450];
  assign o[1569] = i[449];
  assign o[1568] = i[448];
  assign o[1567] = i[511];
  assign o[1566] = i[510];
  assign o[1565] = i[509];
  assign o[1564] = i[508];
  assign o[1563] = i[507];
  assign o[1562] = i[506];
  assign o[1561] = i[505];
  assign o[1560] = i[504];
  assign o[1559] = i[503];
  assign o[1558] = i[502];
  assign o[1557] = i[501];
  assign o[1556] = i[500];
  assign o[1555] = i[499];
  assign o[1554] = i[498];
  assign o[1553] = i[497];
  assign o[1552] = i[496];
  assign o[1551] = i[495];
  assign o[1550] = i[494];
  assign o[1549] = i[493];
  assign o[1548] = i[492];
  assign o[1547] = i[491];
  assign o[1546] = i[490];
  assign o[1545] = i[489];
  assign o[1544] = i[488];
  assign o[1543] = i[487];
  assign o[1542] = i[486];
  assign o[1541] = i[485];
  assign o[1540] = i[484];
  assign o[1539] = i[483];
  assign o[1538] = i[482];
  assign o[1537] = i[481];
  assign o[1536] = i[480];
  assign o[1535] = i[543];
  assign o[1534] = i[542];
  assign o[1533] = i[541];
  assign o[1532] = i[540];
  assign o[1531] = i[539];
  assign o[1530] = i[538];
  assign o[1529] = i[537];
  assign o[1528] = i[536];
  assign o[1527] = i[535];
  assign o[1526] = i[534];
  assign o[1525] = i[533];
  assign o[1524] = i[532];
  assign o[1523] = i[531];
  assign o[1522] = i[530];
  assign o[1521] = i[529];
  assign o[1520] = i[528];
  assign o[1519] = i[527];
  assign o[1518] = i[526];
  assign o[1517] = i[525];
  assign o[1516] = i[524];
  assign o[1515] = i[523];
  assign o[1514] = i[522];
  assign o[1513] = i[521];
  assign o[1512] = i[520];
  assign o[1511] = i[519];
  assign o[1510] = i[518];
  assign o[1509] = i[517];
  assign o[1508] = i[516];
  assign o[1507] = i[515];
  assign o[1506] = i[514];
  assign o[1505] = i[513];
  assign o[1504] = i[512];
  assign o[1503] = i[575];
  assign o[1502] = i[574];
  assign o[1501] = i[573];
  assign o[1500] = i[572];
  assign o[1499] = i[571];
  assign o[1498] = i[570];
  assign o[1497] = i[569];
  assign o[1496] = i[568];
  assign o[1495] = i[567];
  assign o[1494] = i[566];
  assign o[1493] = i[565];
  assign o[1492] = i[564];
  assign o[1491] = i[563];
  assign o[1490] = i[562];
  assign o[1489] = i[561];
  assign o[1488] = i[560];
  assign o[1487] = i[559];
  assign o[1486] = i[558];
  assign o[1485] = i[557];
  assign o[1484] = i[556];
  assign o[1483] = i[555];
  assign o[1482] = i[554];
  assign o[1481] = i[553];
  assign o[1480] = i[552];
  assign o[1479] = i[551];
  assign o[1478] = i[550];
  assign o[1477] = i[549];
  assign o[1476] = i[548];
  assign o[1475] = i[547];
  assign o[1474] = i[546];
  assign o[1473] = i[545];
  assign o[1472] = i[544];
  assign o[1471] = i[607];
  assign o[1470] = i[606];
  assign o[1469] = i[605];
  assign o[1468] = i[604];
  assign o[1467] = i[603];
  assign o[1466] = i[602];
  assign o[1465] = i[601];
  assign o[1464] = i[600];
  assign o[1463] = i[599];
  assign o[1462] = i[598];
  assign o[1461] = i[597];
  assign o[1460] = i[596];
  assign o[1459] = i[595];
  assign o[1458] = i[594];
  assign o[1457] = i[593];
  assign o[1456] = i[592];
  assign o[1455] = i[591];
  assign o[1454] = i[590];
  assign o[1453] = i[589];
  assign o[1452] = i[588];
  assign o[1451] = i[587];
  assign o[1450] = i[586];
  assign o[1449] = i[585];
  assign o[1448] = i[584];
  assign o[1447] = i[583];
  assign o[1446] = i[582];
  assign o[1445] = i[581];
  assign o[1444] = i[580];
  assign o[1443] = i[579];
  assign o[1442] = i[578];
  assign o[1441] = i[577];
  assign o[1440] = i[576];
  assign o[1439] = i[639];
  assign o[1438] = i[638];
  assign o[1437] = i[637];
  assign o[1436] = i[636];
  assign o[1435] = i[635];
  assign o[1434] = i[634];
  assign o[1433] = i[633];
  assign o[1432] = i[632];
  assign o[1431] = i[631];
  assign o[1430] = i[630];
  assign o[1429] = i[629];
  assign o[1428] = i[628];
  assign o[1427] = i[627];
  assign o[1426] = i[626];
  assign o[1425] = i[625];
  assign o[1424] = i[624];
  assign o[1423] = i[623];
  assign o[1422] = i[622];
  assign o[1421] = i[621];
  assign o[1420] = i[620];
  assign o[1419] = i[619];
  assign o[1418] = i[618];
  assign o[1417] = i[617];
  assign o[1416] = i[616];
  assign o[1415] = i[615];
  assign o[1414] = i[614];
  assign o[1413] = i[613];
  assign o[1412] = i[612];
  assign o[1411] = i[611];
  assign o[1410] = i[610];
  assign o[1409] = i[609];
  assign o[1408] = i[608];
  assign o[1407] = i[671];
  assign o[1406] = i[670];
  assign o[1405] = i[669];
  assign o[1404] = i[668];
  assign o[1403] = i[667];
  assign o[1402] = i[666];
  assign o[1401] = i[665];
  assign o[1400] = i[664];
  assign o[1399] = i[663];
  assign o[1398] = i[662];
  assign o[1397] = i[661];
  assign o[1396] = i[660];
  assign o[1395] = i[659];
  assign o[1394] = i[658];
  assign o[1393] = i[657];
  assign o[1392] = i[656];
  assign o[1391] = i[655];
  assign o[1390] = i[654];
  assign o[1389] = i[653];
  assign o[1388] = i[652];
  assign o[1387] = i[651];
  assign o[1386] = i[650];
  assign o[1385] = i[649];
  assign o[1384] = i[648];
  assign o[1383] = i[647];
  assign o[1382] = i[646];
  assign o[1381] = i[645];
  assign o[1380] = i[644];
  assign o[1379] = i[643];
  assign o[1378] = i[642];
  assign o[1377] = i[641];
  assign o[1376] = i[640];
  assign o[1375] = i[703];
  assign o[1374] = i[702];
  assign o[1373] = i[701];
  assign o[1372] = i[700];
  assign o[1371] = i[699];
  assign o[1370] = i[698];
  assign o[1369] = i[697];
  assign o[1368] = i[696];
  assign o[1367] = i[695];
  assign o[1366] = i[694];
  assign o[1365] = i[693];
  assign o[1364] = i[692];
  assign o[1363] = i[691];
  assign o[1362] = i[690];
  assign o[1361] = i[689];
  assign o[1360] = i[688];
  assign o[1359] = i[687];
  assign o[1358] = i[686];
  assign o[1357] = i[685];
  assign o[1356] = i[684];
  assign o[1355] = i[683];
  assign o[1354] = i[682];
  assign o[1353] = i[681];
  assign o[1352] = i[680];
  assign o[1351] = i[679];
  assign o[1350] = i[678];
  assign o[1349] = i[677];
  assign o[1348] = i[676];
  assign o[1347] = i[675];
  assign o[1346] = i[674];
  assign o[1345] = i[673];
  assign o[1344] = i[672];
  assign o[1343] = i[735];
  assign o[1342] = i[734];
  assign o[1341] = i[733];
  assign o[1340] = i[732];
  assign o[1339] = i[731];
  assign o[1338] = i[730];
  assign o[1337] = i[729];
  assign o[1336] = i[728];
  assign o[1335] = i[727];
  assign o[1334] = i[726];
  assign o[1333] = i[725];
  assign o[1332] = i[724];
  assign o[1331] = i[723];
  assign o[1330] = i[722];
  assign o[1329] = i[721];
  assign o[1328] = i[720];
  assign o[1327] = i[719];
  assign o[1326] = i[718];
  assign o[1325] = i[717];
  assign o[1324] = i[716];
  assign o[1323] = i[715];
  assign o[1322] = i[714];
  assign o[1321] = i[713];
  assign o[1320] = i[712];
  assign o[1319] = i[711];
  assign o[1318] = i[710];
  assign o[1317] = i[709];
  assign o[1316] = i[708];
  assign o[1315] = i[707];
  assign o[1314] = i[706];
  assign o[1313] = i[705];
  assign o[1312] = i[704];
  assign o[1311] = i[767];
  assign o[1310] = i[766];
  assign o[1309] = i[765];
  assign o[1308] = i[764];
  assign o[1307] = i[763];
  assign o[1306] = i[762];
  assign o[1305] = i[761];
  assign o[1304] = i[760];
  assign o[1303] = i[759];
  assign o[1302] = i[758];
  assign o[1301] = i[757];
  assign o[1300] = i[756];
  assign o[1299] = i[755];
  assign o[1298] = i[754];
  assign o[1297] = i[753];
  assign o[1296] = i[752];
  assign o[1295] = i[751];
  assign o[1294] = i[750];
  assign o[1293] = i[749];
  assign o[1292] = i[748];
  assign o[1291] = i[747];
  assign o[1290] = i[746];
  assign o[1289] = i[745];
  assign o[1288] = i[744];
  assign o[1287] = i[743];
  assign o[1286] = i[742];
  assign o[1285] = i[741];
  assign o[1284] = i[740];
  assign o[1283] = i[739];
  assign o[1282] = i[738];
  assign o[1281] = i[737];
  assign o[1280] = i[736];
  assign o[1279] = i[799];
  assign o[1278] = i[798];
  assign o[1277] = i[797];
  assign o[1276] = i[796];
  assign o[1275] = i[795];
  assign o[1274] = i[794];
  assign o[1273] = i[793];
  assign o[1272] = i[792];
  assign o[1271] = i[791];
  assign o[1270] = i[790];
  assign o[1269] = i[789];
  assign o[1268] = i[788];
  assign o[1267] = i[787];
  assign o[1266] = i[786];
  assign o[1265] = i[785];
  assign o[1264] = i[784];
  assign o[1263] = i[783];
  assign o[1262] = i[782];
  assign o[1261] = i[781];
  assign o[1260] = i[780];
  assign o[1259] = i[779];
  assign o[1258] = i[778];
  assign o[1257] = i[777];
  assign o[1256] = i[776];
  assign o[1255] = i[775];
  assign o[1254] = i[774];
  assign o[1253] = i[773];
  assign o[1252] = i[772];
  assign o[1251] = i[771];
  assign o[1250] = i[770];
  assign o[1249] = i[769];
  assign o[1248] = i[768];
  assign o[1247] = i[831];
  assign o[1246] = i[830];
  assign o[1245] = i[829];
  assign o[1244] = i[828];
  assign o[1243] = i[827];
  assign o[1242] = i[826];
  assign o[1241] = i[825];
  assign o[1240] = i[824];
  assign o[1239] = i[823];
  assign o[1238] = i[822];
  assign o[1237] = i[821];
  assign o[1236] = i[820];
  assign o[1235] = i[819];
  assign o[1234] = i[818];
  assign o[1233] = i[817];
  assign o[1232] = i[816];
  assign o[1231] = i[815];
  assign o[1230] = i[814];
  assign o[1229] = i[813];
  assign o[1228] = i[812];
  assign o[1227] = i[811];
  assign o[1226] = i[810];
  assign o[1225] = i[809];
  assign o[1224] = i[808];
  assign o[1223] = i[807];
  assign o[1222] = i[806];
  assign o[1221] = i[805];
  assign o[1220] = i[804];
  assign o[1219] = i[803];
  assign o[1218] = i[802];
  assign o[1217] = i[801];
  assign o[1216] = i[800];
  assign o[1215] = i[863];
  assign o[1214] = i[862];
  assign o[1213] = i[861];
  assign o[1212] = i[860];
  assign o[1211] = i[859];
  assign o[1210] = i[858];
  assign o[1209] = i[857];
  assign o[1208] = i[856];
  assign o[1207] = i[855];
  assign o[1206] = i[854];
  assign o[1205] = i[853];
  assign o[1204] = i[852];
  assign o[1203] = i[851];
  assign o[1202] = i[850];
  assign o[1201] = i[849];
  assign o[1200] = i[848];
  assign o[1199] = i[847];
  assign o[1198] = i[846];
  assign o[1197] = i[845];
  assign o[1196] = i[844];
  assign o[1195] = i[843];
  assign o[1194] = i[842];
  assign o[1193] = i[841];
  assign o[1192] = i[840];
  assign o[1191] = i[839];
  assign o[1190] = i[838];
  assign o[1189] = i[837];
  assign o[1188] = i[836];
  assign o[1187] = i[835];
  assign o[1186] = i[834];
  assign o[1185] = i[833];
  assign o[1184] = i[832];
  assign o[1183] = i[895];
  assign o[1182] = i[894];
  assign o[1181] = i[893];
  assign o[1180] = i[892];
  assign o[1179] = i[891];
  assign o[1178] = i[890];
  assign o[1177] = i[889];
  assign o[1176] = i[888];
  assign o[1175] = i[887];
  assign o[1174] = i[886];
  assign o[1173] = i[885];
  assign o[1172] = i[884];
  assign o[1171] = i[883];
  assign o[1170] = i[882];
  assign o[1169] = i[881];
  assign o[1168] = i[880];
  assign o[1167] = i[879];
  assign o[1166] = i[878];
  assign o[1165] = i[877];
  assign o[1164] = i[876];
  assign o[1163] = i[875];
  assign o[1162] = i[874];
  assign o[1161] = i[873];
  assign o[1160] = i[872];
  assign o[1159] = i[871];
  assign o[1158] = i[870];
  assign o[1157] = i[869];
  assign o[1156] = i[868];
  assign o[1155] = i[867];
  assign o[1154] = i[866];
  assign o[1153] = i[865];
  assign o[1152] = i[864];
  assign o[1151] = i[927];
  assign o[1150] = i[926];
  assign o[1149] = i[925];
  assign o[1148] = i[924];
  assign o[1147] = i[923];
  assign o[1146] = i[922];
  assign o[1145] = i[921];
  assign o[1144] = i[920];
  assign o[1143] = i[919];
  assign o[1142] = i[918];
  assign o[1141] = i[917];
  assign o[1140] = i[916];
  assign o[1139] = i[915];
  assign o[1138] = i[914];
  assign o[1137] = i[913];
  assign o[1136] = i[912];
  assign o[1135] = i[911];
  assign o[1134] = i[910];
  assign o[1133] = i[909];
  assign o[1132] = i[908];
  assign o[1131] = i[907];
  assign o[1130] = i[906];
  assign o[1129] = i[905];
  assign o[1128] = i[904];
  assign o[1127] = i[903];
  assign o[1126] = i[902];
  assign o[1125] = i[901];
  assign o[1124] = i[900];
  assign o[1123] = i[899];
  assign o[1122] = i[898];
  assign o[1121] = i[897];
  assign o[1120] = i[896];
  assign o[1119] = i[959];
  assign o[1118] = i[958];
  assign o[1117] = i[957];
  assign o[1116] = i[956];
  assign o[1115] = i[955];
  assign o[1114] = i[954];
  assign o[1113] = i[953];
  assign o[1112] = i[952];
  assign o[1111] = i[951];
  assign o[1110] = i[950];
  assign o[1109] = i[949];
  assign o[1108] = i[948];
  assign o[1107] = i[947];
  assign o[1106] = i[946];
  assign o[1105] = i[945];
  assign o[1104] = i[944];
  assign o[1103] = i[943];
  assign o[1102] = i[942];
  assign o[1101] = i[941];
  assign o[1100] = i[940];
  assign o[1099] = i[939];
  assign o[1098] = i[938];
  assign o[1097] = i[937];
  assign o[1096] = i[936];
  assign o[1095] = i[935];
  assign o[1094] = i[934];
  assign o[1093] = i[933];
  assign o[1092] = i[932];
  assign o[1091] = i[931];
  assign o[1090] = i[930];
  assign o[1089] = i[929];
  assign o[1088] = i[928];
  assign o[1087] = i[991];
  assign o[1086] = i[990];
  assign o[1085] = i[989];
  assign o[1084] = i[988];
  assign o[1083] = i[987];
  assign o[1082] = i[986];
  assign o[1081] = i[985];
  assign o[1080] = i[984];
  assign o[1079] = i[983];
  assign o[1078] = i[982];
  assign o[1077] = i[981];
  assign o[1076] = i[980];
  assign o[1075] = i[979];
  assign o[1074] = i[978];
  assign o[1073] = i[977];
  assign o[1072] = i[976];
  assign o[1071] = i[975];
  assign o[1070] = i[974];
  assign o[1069] = i[973];
  assign o[1068] = i[972];
  assign o[1067] = i[971];
  assign o[1066] = i[970];
  assign o[1065] = i[969];
  assign o[1064] = i[968];
  assign o[1063] = i[967];
  assign o[1062] = i[966];
  assign o[1061] = i[965];
  assign o[1060] = i[964];
  assign o[1059] = i[963];
  assign o[1058] = i[962];
  assign o[1057] = i[961];
  assign o[1056] = i[960];
  assign o[1055] = i[1023];
  assign o[1054] = i[1022];
  assign o[1053] = i[1021];
  assign o[1052] = i[1020];
  assign o[1051] = i[1019];
  assign o[1050] = i[1018];
  assign o[1049] = i[1017];
  assign o[1048] = i[1016];
  assign o[1047] = i[1015];
  assign o[1046] = i[1014];
  assign o[1045] = i[1013];
  assign o[1044] = i[1012];
  assign o[1043] = i[1011];
  assign o[1042] = i[1010];
  assign o[1041] = i[1009];
  assign o[1040] = i[1008];
  assign o[1039] = i[1007];
  assign o[1038] = i[1006];
  assign o[1037] = i[1005];
  assign o[1036] = i[1004];
  assign o[1035] = i[1003];
  assign o[1034] = i[1002];
  assign o[1033] = i[1001];
  assign o[1032] = i[1000];
  assign o[1031] = i[999];
  assign o[1030] = i[998];
  assign o[1029] = i[997];
  assign o[1028] = i[996];
  assign o[1027] = i[995];
  assign o[1026] = i[994];
  assign o[1025] = i[993];
  assign o[1024] = i[992];
  assign o[1023] = i[1055];
  assign o[1022] = i[1054];
  assign o[1021] = i[1053];
  assign o[1020] = i[1052];
  assign o[1019] = i[1051];
  assign o[1018] = i[1050];
  assign o[1017] = i[1049];
  assign o[1016] = i[1048];
  assign o[1015] = i[1047];
  assign o[1014] = i[1046];
  assign o[1013] = i[1045];
  assign o[1012] = i[1044];
  assign o[1011] = i[1043];
  assign o[1010] = i[1042];
  assign o[1009] = i[1041];
  assign o[1008] = i[1040];
  assign o[1007] = i[1039];
  assign o[1006] = i[1038];
  assign o[1005] = i[1037];
  assign o[1004] = i[1036];
  assign o[1003] = i[1035];
  assign o[1002] = i[1034];
  assign o[1001] = i[1033];
  assign o[1000] = i[1032];
  assign o[999] = i[1031];
  assign o[998] = i[1030];
  assign o[997] = i[1029];
  assign o[996] = i[1028];
  assign o[995] = i[1027];
  assign o[994] = i[1026];
  assign o[993] = i[1025];
  assign o[992] = i[1024];
  assign o[991] = i[1087];
  assign o[990] = i[1086];
  assign o[989] = i[1085];
  assign o[988] = i[1084];
  assign o[987] = i[1083];
  assign o[986] = i[1082];
  assign o[985] = i[1081];
  assign o[984] = i[1080];
  assign o[983] = i[1079];
  assign o[982] = i[1078];
  assign o[981] = i[1077];
  assign o[980] = i[1076];
  assign o[979] = i[1075];
  assign o[978] = i[1074];
  assign o[977] = i[1073];
  assign o[976] = i[1072];
  assign o[975] = i[1071];
  assign o[974] = i[1070];
  assign o[973] = i[1069];
  assign o[972] = i[1068];
  assign o[971] = i[1067];
  assign o[970] = i[1066];
  assign o[969] = i[1065];
  assign o[968] = i[1064];
  assign o[967] = i[1063];
  assign o[966] = i[1062];
  assign o[965] = i[1061];
  assign o[964] = i[1060];
  assign o[963] = i[1059];
  assign o[962] = i[1058];
  assign o[961] = i[1057];
  assign o[960] = i[1056];
  assign o[959] = i[1119];
  assign o[958] = i[1118];
  assign o[957] = i[1117];
  assign o[956] = i[1116];
  assign o[955] = i[1115];
  assign o[954] = i[1114];
  assign o[953] = i[1113];
  assign o[952] = i[1112];
  assign o[951] = i[1111];
  assign o[950] = i[1110];
  assign o[949] = i[1109];
  assign o[948] = i[1108];
  assign o[947] = i[1107];
  assign o[946] = i[1106];
  assign o[945] = i[1105];
  assign o[944] = i[1104];
  assign o[943] = i[1103];
  assign o[942] = i[1102];
  assign o[941] = i[1101];
  assign o[940] = i[1100];
  assign o[939] = i[1099];
  assign o[938] = i[1098];
  assign o[937] = i[1097];
  assign o[936] = i[1096];
  assign o[935] = i[1095];
  assign o[934] = i[1094];
  assign o[933] = i[1093];
  assign o[932] = i[1092];
  assign o[931] = i[1091];
  assign o[930] = i[1090];
  assign o[929] = i[1089];
  assign o[928] = i[1088];
  assign o[927] = i[1151];
  assign o[926] = i[1150];
  assign o[925] = i[1149];
  assign o[924] = i[1148];
  assign o[923] = i[1147];
  assign o[922] = i[1146];
  assign o[921] = i[1145];
  assign o[920] = i[1144];
  assign o[919] = i[1143];
  assign o[918] = i[1142];
  assign o[917] = i[1141];
  assign o[916] = i[1140];
  assign o[915] = i[1139];
  assign o[914] = i[1138];
  assign o[913] = i[1137];
  assign o[912] = i[1136];
  assign o[911] = i[1135];
  assign o[910] = i[1134];
  assign o[909] = i[1133];
  assign o[908] = i[1132];
  assign o[907] = i[1131];
  assign o[906] = i[1130];
  assign o[905] = i[1129];
  assign o[904] = i[1128];
  assign o[903] = i[1127];
  assign o[902] = i[1126];
  assign o[901] = i[1125];
  assign o[900] = i[1124];
  assign o[899] = i[1123];
  assign o[898] = i[1122];
  assign o[897] = i[1121];
  assign o[896] = i[1120];
  assign o[895] = i[1183];
  assign o[894] = i[1182];
  assign o[893] = i[1181];
  assign o[892] = i[1180];
  assign o[891] = i[1179];
  assign o[890] = i[1178];
  assign o[889] = i[1177];
  assign o[888] = i[1176];
  assign o[887] = i[1175];
  assign o[886] = i[1174];
  assign o[885] = i[1173];
  assign o[884] = i[1172];
  assign o[883] = i[1171];
  assign o[882] = i[1170];
  assign o[881] = i[1169];
  assign o[880] = i[1168];
  assign o[879] = i[1167];
  assign o[878] = i[1166];
  assign o[877] = i[1165];
  assign o[876] = i[1164];
  assign o[875] = i[1163];
  assign o[874] = i[1162];
  assign o[873] = i[1161];
  assign o[872] = i[1160];
  assign o[871] = i[1159];
  assign o[870] = i[1158];
  assign o[869] = i[1157];
  assign o[868] = i[1156];
  assign o[867] = i[1155];
  assign o[866] = i[1154];
  assign o[865] = i[1153];
  assign o[864] = i[1152];
  assign o[863] = i[1215];
  assign o[862] = i[1214];
  assign o[861] = i[1213];
  assign o[860] = i[1212];
  assign o[859] = i[1211];
  assign o[858] = i[1210];
  assign o[857] = i[1209];
  assign o[856] = i[1208];
  assign o[855] = i[1207];
  assign o[854] = i[1206];
  assign o[853] = i[1205];
  assign o[852] = i[1204];
  assign o[851] = i[1203];
  assign o[850] = i[1202];
  assign o[849] = i[1201];
  assign o[848] = i[1200];
  assign o[847] = i[1199];
  assign o[846] = i[1198];
  assign o[845] = i[1197];
  assign o[844] = i[1196];
  assign o[843] = i[1195];
  assign o[842] = i[1194];
  assign o[841] = i[1193];
  assign o[840] = i[1192];
  assign o[839] = i[1191];
  assign o[838] = i[1190];
  assign o[837] = i[1189];
  assign o[836] = i[1188];
  assign o[835] = i[1187];
  assign o[834] = i[1186];
  assign o[833] = i[1185];
  assign o[832] = i[1184];
  assign o[831] = i[1247];
  assign o[830] = i[1246];
  assign o[829] = i[1245];
  assign o[828] = i[1244];
  assign o[827] = i[1243];
  assign o[826] = i[1242];
  assign o[825] = i[1241];
  assign o[824] = i[1240];
  assign o[823] = i[1239];
  assign o[822] = i[1238];
  assign o[821] = i[1237];
  assign o[820] = i[1236];
  assign o[819] = i[1235];
  assign o[818] = i[1234];
  assign o[817] = i[1233];
  assign o[816] = i[1232];
  assign o[815] = i[1231];
  assign o[814] = i[1230];
  assign o[813] = i[1229];
  assign o[812] = i[1228];
  assign o[811] = i[1227];
  assign o[810] = i[1226];
  assign o[809] = i[1225];
  assign o[808] = i[1224];
  assign o[807] = i[1223];
  assign o[806] = i[1222];
  assign o[805] = i[1221];
  assign o[804] = i[1220];
  assign o[803] = i[1219];
  assign o[802] = i[1218];
  assign o[801] = i[1217];
  assign o[800] = i[1216];
  assign o[799] = i[1279];
  assign o[798] = i[1278];
  assign o[797] = i[1277];
  assign o[796] = i[1276];
  assign o[795] = i[1275];
  assign o[794] = i[1274];
  assign o[793] = i[1273];
  assign o[792] = i[1272];
  assign o[791] = i[1271];
  assign o[790] = i[1270];
  assign o[789] = i[1269];
  assign o[788] = i[1268];
  assign o[787] = i[1267];
  assign o[786] = i[1266];
  assign o[785] = i[1265];
  assign o[784] = i[1264];
  assign o[783] = i[1263];
  assign o[782] = i[1262];
  assign o[781] = i[1261];
  assign o[780] = i[1260];
  assign o[779] = i[1259];
  assign o[778] = i[1258];
  assign o[777] = i[1257];
  assign o[776] = i[1256];
  assign o[775] = i[1255];
  assign o[774] = i[1254];
  assign o[773] = i[1253];
  assign o[772] = i[1252];
  assign o[771] = i[1251];
  assign o[770] = i[1250];
  assign o[769] = i[1249];
  assign o[768] = i[1248];
  assign o[767] = i[1311];
  assign o[766] = i[1310];
  assign o[765] = i[1309];
  assign o[764] = i[1308];
  assign o[763] = i[1307];
  assign o[762] = i[1306];
  assign o[761] = i[1305];
  assign o[760] = i[1304];
  assign o[759] = i[1303];
  assign o[758] = i[1302];
  assign o[757] = i[1301];
  assign o[756] = i[1300];
  assign o[755] = i[1299];
  assign o[754] = i[1298];
  assign o[753] = i[1297];
  assign o[752] = i[1296];
  assign o[751] = i[1295];
  assign o[750] = i[1294];
  assign o[749] = i[1293];
  assign o[748] = i[1292];
  assign o[747] = i[1291];
  assign o[746] = i[1290];
  assign o[745] = i[1289];
  assign o[744] = i[1288];
  assign o[743] = i[1287];
  assign o[742] = i[1286];
  assign o[741] = i[1285];
  assign o[740] = i[1284];
  assign o[739] = i[1283];
  assign o[738] = i[1282];
  assign o[737] = i[1281];
  assign o[736] = i[1280];
  assign o[735] = i[1343];
  assign o[734] = i[1342];
  assign o[733] = i[1341];
  assign o[732] = i[1340];
  assign o[731] = i[1339];
  assign o[730] = i[1338];
  assign o[729] = i[1337];
  assign o[728] = i[1336];
  assign o[727] = i[1335];
  assign o[726] = i[1334];
  assign o[725] = i[1333];
  assign o[724] = i[1332];
  assign o[723] = i[1331];
  assign o[722] = i[1330];
  assign o[721] = i[1329];
  assign o[720] = i[1328];
  assign o[719] = i[1327];
  assign o[718] = i[1326];
  assign o[717] = i[1325];
  assign o[716] = i[1324];
  assign o[715] = i[1323];
  assign o[714] = i[1322];
  assign o[713] = i[1321];
  assign o[712] = i[1320];
  assign o[711] = i[1319];
  assign o[710] = i[1318];
  assign o[709] = i[1317];
  assign o[708] = i[1316];
  assign o[707] = i[1315];
  assign o[706] = i[1314];
  assign o[705] = i[1313];
  assign o[704] = i[1312];
  assign o[703] = i[1375];
  assign o[702] = i[1374];
  assign o[701] = i[1373];
  assign o[700] = i[1372];
  assign o[699] = i[1371];
  assign o[698] = i[1370];
  assign o[697] = i[1369];
  assign o[696] = i[1368];
  assign o[695] = i[1367];
  assign o[694] = i[1366];
  assign o[693] = i[1365];
  assign o[692] = i[1364];
  assign o[691] = i[1363];
  assign o[690] = i[1362];
  assign o[689] = i[1361];
  assign o[688] = i[1360];
  assign o[687] = i[1359];
  assign o[686] = i[1358];
  assign o[685] = i[1357];
  assign o[684] = i[1356];
  assign o[683] = i[1355];
  assign o[682] = i[1354];
  assign o[681] = i[1353];
  assign o[680] = i[1352];
  assign o[679] = i[1351];
  assign o[678] = i[1350];
  assign o[677] = i[1349];
  assign o[676] = i[1348];
  assign o[675] = i[1347];
  assign o[674] = i[1346];
  assign o[673] = i[1345];
  assign o[672] = i[1344];
  assign o[671] = i[1407];
  assign o[670] = i[1406];
  assign o[669] = i[1405];
  assign o[668] = i[1404];
  assign o[667] = i[1403];
  assign o[666] = i[1402];
  assign o[665] = i[1401];
  assign o[664] = i[1400];
  assign o[663] = i[1399];
  assign o[662] = i[1398];
  assign o[661] = i[1397];
  assign o[660] = i[1396];
  assign o[659] = i[1395];
  assign o[658] = i[1394];
  assign o[657] = i[1393];
  assign o[656] = i[1392];
  assign o[655] = i[1391];
  assign o[654] = i[1390];
  assign o[653] = i[1389];
  assign o[652] = i[1388];
  assign o[651] = i[1387];
  assign o[650] = i[1386];
  assign o[649] = i[1385];
  assign o[648] = i[1384];
  assign o[647] = i[1383];
  assign o[646] = i[1382];
  assign o[645] = i[1381];
  assign o[644] = i[1380];
  assign o[643] = i[1379];
  assign o[642] = i[1378];
  assign o[641] = i[1377];
  assign o[640] = i[1376];
  assign o[639] = i[1439];
  assign o[638] = i[1438];
  assign o[637] = i[1437];
  assign o[636] = i[1436];
  assign o[635] = i[1435];
  assign o[634] = i[1434];
  assign o[633] = i[1433];
  assign o[632] = i[1432];
  assign o[631] = i[1431];
  assign o[630] = i[1430];
  assign o[629] = i[1429];
  assign o[628] = i[1428];
  assign o[627] = i[1427];
  assign o[626] = i[1426];
  assign o[625] = i[1425];
  assign o[624] = i[1424];
  assign o[623] = i[1423];
  assign o[622] = i[1422];
  assign o[621] = i[1421];
  assign o[620] = i[1420];
  assign o[619] = i[1419];
  assign o[618] = i[1418];
  assign o[617] = i[1417];
  assign o[616] = i[1416];
  assign o[615] = i[1415];
  assign o[614] = i[1414];
  assign o[613] = i[1413];
  assign o[612] = i[1412];
  assign o[611] = i[1411];
  assign o[610] = i[1410];
  assign o[609] = i[1409];
  assign o[608] = i[1408];
  assign o[607] = i[1471];
  assign o[606] = i[1470];
  assign o[605] = i[1469];
  assign o[604] = i[1468];
  assign o[603] = i[1467];
  assign o[602] = i[1466];
  assign o[601] = i[1465];
  assign o[600] = i[1464];
  assign o[599] = i[1463];
  assign o[598] = i[1462];
  assign o[597] = i[1461];
  assign o[596] = i[1460];
  assign o[595] = i[1459];
  assign o[594] = i[1458];
  assign o[593] = i[1457];
  assign o[592] = i[1456];
  assign o[591] = i[1455];
  assign o[590] = i[1454];
  assign o[589] = i[1453];
  assign o[588] = i[1452];
  assign o[587] = i[1451];
  assign o[586] = i[1450];
  assign o[585] = i[1449];
  assign o[584] = i[1448];
  assign o[583] = i[1447];
  assign o[582] = i[1446];
  assign o[581] = i[1445];
  assign o[580] = i[1444];
  assign o[579] = i[1443];
  assign o[578] = i[1442];
  assign o[577] = i[1441];
  assign o[576] = i[1440];
  assign o[575] = i[1503];
  assign o[574] = i[1502];
  assign o[573] = i[1501];
  assign o[572] = i[1500];
  assign o[571] = i[1499];
  assign o[570] = i[1498];
  assign o[569] = i[1497];
  assign o[568] = i[1496];
  assign o[567] = i[1495];
  assign o[566] = i[1494];
  assign o[565] = i[1493];
  assign o[564] = i[1492];
  assign o[563] = i[1491];
  assign o[562] = i[1490];
  assign o[561] = i[1489];
  assign o[560] = i[1488];
  assign o[559] = i[1487];
  assign o[558] = i[1486];
  assign o[557] = i[1485];
  assign o[556] = i[1484];
  assign o[555] = i[1483];
  assign o[554] = i[1482];
  assign o[553] = i[1481];
  assign o[552] = i[1480];
  assign o[551] = i[1479];
  assign o[550] = i[1478];
  assign o[549] = i[1477];
  assign o[548] = i[1476];
  assign o[547] = i[1475];
  assign o[546] = i[1474];
  assign o[545] = i[1473];
  assign o[544] = i[1472];
  assign o[543] = i[1535];
  assign o[542] = i[1534];
  assign o[541] = i[1533];
  assign o[540] = i[1532];
  assign o[539] = i[1531];
  assign o[538] = i[1530];
  assign o[537] = i[1529];
  assign o[536] = i[1528];
  assign o[535] = i[1527];
  assign o[534] = i[1526];
  assign o[533] = i[1525];
  assign o[532] = i[1524];
  assign o[531] = i[1523];
  assign o[530] = i[1522];
  assign o[529] = i[1521];
  assign o[528] = i[1520];
  assign o[527] = i[1519];
  assign o[526] = i[1518];
  assign o[525] = i[1517];
  assign o[524] = i[1516];
  assign o[523] = i[1515];
  assign o[522] = i[1514];
  assign o[521] = i[1513];
  assign o[520] = i[1512];
  assign o[519] = i[1511];
  assign o[518] = i[1510];
  assign o[517] = i[1509];
  assign o[516] = i[1508];
  assign o[515] = i[1507];
  assign o[514] = i[1506];
  assign o[513] = i[1505];
  assign o[512] = i[1504];
  assign o[511] = i[1567];
  assign o[510] = i[1566];
  assign o[509] = i[1565];
  assign o[508] = i[1564];
  assign o[507] = i[1563];
  assign o[506] = i[1562];
  assign o[505] = i[1561];
  assign o[504] = i[1560];
  assign o[503] = i[1559];
  assign o[502] = i[1558];
  assign o[501] = i[1557];
  assign o[500] = i[1556];
  assign o[499] = i[1555];
  assign o[498] = i[1554];
  assign o[497] = i[1553];
  assign o[496] = i[1552];
  assign o[495] = i[1551];
  assign o[494] = i[1550];
  assign o[493] = i[1549];
  assign o[492] = i[1548];
  assign o[491] = i[1547];
  assign o[490] = i[1546];
  assign o[489] = i[1545];
  assign o[488] = i[1544];
  assign o[487] = i[1543];
  assign o[486] = i[1542];
  assign o[485] = i[1541];
  assign o[484] = i[1540];
  assign o[483] = i[1539];
  assign o[482] = i[1538];
  assign o[481] = i[1537];
  assign o[480] = i[1536];
  assign o[479] = i[1599];
  assign o[478] = i[1598];
  assign o[477] = i[1597];
  assign o[476] = i[1596];
  assign o[475] = i[1595];
  assign o[474] = i[1594];
  assign o[473] = i[1593];
  assign o[472] = i[1592];
  assign o[471] = i[1591];
  assign o[470] = i[1590];
  assign o[469] = i[1589];
  assign o[468] = i[1588];
  assign o[467] = i[1587];
  assign o[466] = i[1586];
  assign o[465] = i[1585];
  assign o[464] = i[1584];
  assign o[463] = i[1583];
  assign o[462] = i[1582];
  assign o[461] = i[1581];
  assign o[460] = i[1580];
  assign o[459] = i[1579];
  assign o[458] = i[1578];
  assign o[457] = i[1577];
  assign o[456] = i[1576];
  assign o[455] = i[1575];
  assign o[454] = i[1574];
  assign o[453] = i[1573];
  assign o[452] = i[1572];
  assign o[451] = i[1571];
  assign o[450] = i[1570];
  assign o[449] = i[1569];
  assign o[448] = i[1568];
  assign o[447] = i[1631];
  assign o[446] = i[1630];
  assign o[445] = i[1629];
  assign o[444] = i[1628];
  assign o[443] = i[1627];
  assign o[442] = i[1626];
  assign o[441] = i[1625];
  assign o[440] = i[1624];
  assign o[439] = i[1623];
  assign o[438] = i[1622];
  assign o[437] = i[1621];
  assign o[436] = i[1620];
  assign o[435] = i[1619];
  assign o[434] = i[1618];
  assign o[433] = i[1617];
  assign o[432] = i[1616];
  assign o[431] = i[1615];
  assign o[430] = i[1614];
  assign o[429] = i[1613];
  assign o[428] = i[1612];
  assign o[427] = i[1611];
  assign o[426] = i[1610];
  assign o[425] = i[1609];
  assign o[424] = i[1608];
  assign o[423] = i[1607];
  assign o[422] = i[1606];
  assign o[421] = i[1605];
  assign o[420] = i[1604];
  assign o[419] = i[1603];
  assign o[418] = i[1602];
  assign o[417] = i[1601];
  assign o[416] = i[1600];
  assign o[415] = i[1663];
  assign o[414] = i[1662];
  assign o[413] = i[1661];
  assign o[412] = i[1660];
  assign o[411] = i[1659];
  assign o[410] = i[1658];
  assign o[409] = i[1657];
  assign o[408] = i[1656];
  assign o[407] = i[1655];
  assign o[406] = i[1654];
  assign o[405] = i[1653];
  assign o[404] = i[1652];
  assign o[403] = i[1651];
  assign o[402] = i[1650];
  assign o[401] = i[1649];
  assign o[400] = i[1648];
  assign o[399] = i[1647];
  assign o[398] = i[1646];
  assign o[397] = i[1645];
  assign o[396] = i[1644];
  assign o[395] = i[1643];
  assign o[394] = i[1642];
  assign o[393] = i[1641];
  assign o[392] = i[1640];
  assign o[391] = i[1639];
  assign o[390] = i[1638];
  assign o[389] = i[1637];
  assign o[388] = i[1636];
  assign o[387] = i[1635];
  assign o[386] = i[1634];
  assign o[385] = i[1633];
  assign o[384] = i[1632];
  assign o[383] = i[1695];
  assign o[382] = i[1694];
  assign o[381] = i[1693];
  assign o[380] = i[1692];
  assign o[379] = i[1691];
  assign o[378] = i[1690];
  assign o[377] = i[1689];
  assign o[376] = i[1688];
  assign o[375] = i[1687];
  assign o[374] = i[1686];
  assign o[373] = i[1685];
  assign o[372] = i[1684];
  assign o[371] = i[1683];
  assign o[370] = i[1682];
  assign o[369] = i[1681];
  assign o[368] = i[1680];
  assign o[367] = i[1679];
  assign o[366] = i[1678];
  assign o[365] = i[1677];
  assign o[364] = i[1676];
  assign o[363] = i[1675];
  assign o[362] = i[1674];
  assign o[361] = i[1673];
  assign o[360] = i[1672];
  assign o[359] = i[1671];
  assign o[358] = i[1670];
  assign o[357] = i[1669];
  assign o[356] = i[1668];
  assign o[355] = i[1667];
  assign o[354] = i[1666];
  assign o[353] = i[1665];
  assign o[352] = i[1664];
  assign o[351] = i[1727];
  assign o[350] = i[1726];
  assign o[349] = i[1725];
  assign o[348] = i[1724];
  assign o[347] = i[1723];
  assign o[346] = i[1722];
  assign o[345] = i[1721];
  assign o[344] = i[1720];
  assign o[343] = i[1719];
  assign o[342] = i[1718];
  assign o[341] = i[1717];
  assign o[340] = i[1716];
  assign o[339] = i[1715];
  assign o[338] = i[1714];
  assign o[337] = i[1713];
  assign o[336] = i[1712];
  assign o[335] = i[1711];
  assign o[334] = i[1710];
  assign o[333] = i[1709];
  assign o[332] = i[1708];
  assign o[331] = i[1707];
  assign o[330] = i[1706];
  assign o[329] = i[1705];
  assign o[328] = i[1704];
  assign o[327] = i[1703];
  assign o[326] = i[1702];
  assign o[325] = i[1701];
  assign o[324] = i[1700];
  assign o[323] = i[1699];
  assign o[322] = i[1698];
  assign o[321] = i[1697];
  assign o[320] = i[1696];
  assign o[319] = i[1759];
  assign o[318] = i[1758];
  assign o[317] = i[1757];
  assign o[316] = i[1756];
  assign o[315] = i[1755];
  assign o[314] = i[1754];
  assign o[313] = i[1753];
  assign o[312] = i[1752];
  assign o[311] = i[1751];
  assign o[310] = i[1750];
  assign o[309] = i[1749];
  assign o[308] = i[1748];
  assign o[307] = i[1747];
  assign o[306] = i[1746];
  assign o[305] = i[1745];
  assign o[304] = i[1744];
  assign o[303] = i[1743];
  assign o[302] = i[1742];
  assign o[301] = i[1741];
  assign o[300] = i[1740];
  assign o[299] = i[1739];
  assign o[298] = i[1738];
  assign o[297] = i[1737];
  assign o[296] = i[1736];
  assign o[295] = i[1735];
  assign o[294] = i[1734];
  assign o[293] = i[1733];
  assign o[292] = i[1732];
  assign o[291] = i[1731];
  assign o[290] = i[1730];
  assign o[289] = i[1729];
  assign o[288] = i[1728];
  assign o[287] = i[1791];
  assign o[286] = i[1790];
  assign o[285] = i[1789];
  assign o[284] = i[1788];
  assign o[283] = i[1787];
  assign o[282] = i[1786];
  assign o[281] = i[1785];
  assign o[280] = i[1784];
  assign o[279] = i[1783];
  assign o[278] = i[1782];
  assign o[277] = i[1781];
  assign o[276] = i[1780];
  assign o[275] = i[1779];
  assign o[274] = i[1778];
  assign o[273] = i[1777];
  assign o[272] = i[1776];
  assign o[271] = i[1775];
  assign o[270] = i[1774];
  assign o[269] = i[1773];
  assign o[268] = i[1772];
  assign o[267] = i[1771];
  assign o[266] = i[1770];
  assign o[265] = i[1769];
  assign o[264] = i[1768];
  assign o[263] = i[1767];
  assign o[262] = i[1766];
  assign o[261] = i[1765];
  assign o[260] = i[1764];
  assign o[259] = i[1763];
  assign o[258] = i[1762];
  assign o[257] = i[1761];
  assign o[256] = i[1760];
  assign o[255] = i[1823];
  assign o[254] = i[1822];
  assign o[253] = i[1821];
  assign o[252] = i[1820];
  assign o[251] = i[1819];
  assign o[250] = i[1818];
  assign o[249] = i[1817];
  assign o[248] = i[1816];
  assign o[247] = i[1815];
  assign o[246] = i[1814];
  assign o[245] = i[1813];
  assign o[244] = i[1812];
  assign o[243] = i[1811];
  assign o[242] = i[1810];
  assign o[241] = i[1809];
  assign o[240] = i[1808];
  assign o[239] = i[1807];
  assign o[238] = i[1806];
  assign o[237] = i[1805];
  assign o[236] = i[1804];
  assign o[235] = i[1803];
  assign o[234] = i[1802];
  assign o[233] = i[1801];
  assign o[232] = i[1800];
  assign o[231] = i[1799];
  assign o[230] = i[1798];
  assign o[229] = i[1797];
  assign o[228] = i[1796];
  assign o[227] = i[1795];
  assign o[226] = i[1794];
  assign o[225] = i[1793];
  assign o[224] = i[1792];
  assign o[223] = i[1855];
  assign o[222] = i[1854];
  assign o[221] = i[1853];
  assign o[220] = i[1852];
  assign o[219] = i[1851];
  assign o[218] = i[1850];
  assign o[217] = i[1849];
  assign o[216] = i[1848];
  assign o[215] = i[1847];
  assign o[214] = i[1846];
  assign o[213] = i[1845];
  assign o[212] = i[1844];
  assign o[211] = i[1843];
  assign o[210] = i[1842];
  assign o[209] = i[1841];
  assign o[208] = i[1840];
  assign o[207] = i[1839];
  assign o[206] = i[1838];
  assign o[205] = i[1837];
  assign o[204] = i[1836];
  assign o[203] = i[1835];
  assign o[202] = i[1834];
  assign o[201] = i[1833];
  assign o[200] = i[1832];
  assign o[199] = i[1831];
  assign o[198] = i[1830];
  assign o[197] = i[1829];
  assign o[196] = i[1828];
  assign o[195] = i[1827];
  assign o[194] = i[1826];
  assign o[193] = i[1825];
  assign o[192] = i[1824];
  assign o[191] = i[1887];
  assign o[190] = i[1886];
  assign o[189] = i[1885];
  assign o[188] = i[1884];
  assign o[187] = i[1883];
  assign o[186] = i[1882];
  assign o[185] = i[1881];
  assign o[184] = i[1880];
  assign o[183] = i[1879];
  assign o[182] = i[1878];
  assign o[181] = i[1877];
  assign o[180] = i[1876];
  assign o[179] = i[1875];
  assign o[178] = i[1874];
  assign o[177] = i[1873];
  assign o[176] = i[1872];
  assign o[175] = i[1871];
  assign o[174] = i[1870];
  assign o[173] = i[1869];
  assign o[172] = i[1868];
  assign o[171] = i[1867];
  assign o[170] = i[1866];
  assign o[169] = i[1865];
  assign o[168] = i[1864];
  assign o[167] = i[1863];
  assign o[166] = i[1862];
  assign o[165] = i[1861];
  assign o[164] = i[1860];
  assign o[163] = i[1859];
  assign o[162] = i[1858];
  assign o[161] = i[1857];
  assign o[160] = i[1856];
  assign o[159] = i[1919];
  assign o[158] = i[1918];
  assign o[157] = i[1917];
  assign o[156] = i[1916];
  assign o[155] = i[1915];
  assign o[154] = i[1914];
  assign o[153] = i[1913];
  assign o[152] = i[1912];
  assign o[151] = i[1911];
  assign o[150] = i[1910];
  assign o[149] = i[1909];
  assign o[148] = i[1908];
  assign o[147] = i[1907];
  assign o[146] = i[1906];
  assign o[145] = i[1905];
  assign o[144] = i[1904];
  assign o[143] = i[1903];
  assign o[142] = i[1902];
  assign o[141] = i[1901];
  assign o[140] = i[1900];
  assign o[139] = i[1899];
  assign o[138] = i[1898];
  assign o[137] = i[1897];
  assign o[136] = i[1896];
  assign o[135] = i[1895];
  assign o[134] = i[1894];
  assign o[133] = i[1893];
  assign o[132] = i[1892];
  assign o[131] = i[1891];
  assign o[130] = i[1890];
  assign o[129] = i[1889];
  assign o[128] = i[1888];
  assign o[127] = i[1951];
  assign o[126] = i[1950];
  assign o[125] = i[1949];
  assign o[124] = i[1948];
  assign o[123] = i[1947];
  assign o[122] = i[1946];
  assign o[121] = i[1945];
  assign o[120] = i[1944];
  assign o[119] = i[1943];
  assign o[118] = i[1942];
  assign o[117] = i[1941];
  assign o[116] = i[1940];
  assign o[115] = i[1939];
  assign o[114] = i[1938];
  assign o[113] = i[1937];
  assign o[112] = i[1936];
  assign o[111] = i[1935];
  assign o[110] = i[1934];
  assign o[109] = i[1933];
  assign o[108] = i[1932];
  assign o[107] = i[1931];
  assign o[106] = i[1930];
  assign o[105] = i[1929];
  assign o[104] = i[1928];
  assign o[103] = i[1927];
  assign o[102] = i[1926];
  assign o[101] = i[1925];
  assign o[100] = i[1924];
  assign o[99] = i[1923];
  assign o[98] = i[1922];
  assign o[97] = i[1921];
  assign o[96] = i[1920];
  assign o[95] = i[1983];
  assign o[94] = i[1982];
  assign o[93] = i[1981];
  assign o[92] = i[1980];
  assign o[91] = i[1979];
  assign o[90] = i[1978];
  assign o[89] = i[1977];
  assign o[88] = i[1976];
  assign o[87] = i[1975];
  assign o[86] = i[1974];
  assign o[85] = i[1973];
  assign o[84] = i[1972];
  assign o[83] = i[1971];
  assign o[82] = i[1970];
  assign o[81] = i[1969];
  assign o[80] = i[1968];
  assign o[79] = i[1967];
  assign o[78] = i[1966];
  assign o[77] = i[1965];
  assign o[76] = i[1964];
  assign o[75] = i[1963];
  assign o[74] = i[1962];
  assign o[73] = i[1961];
  assign o[72] = i[1960];
  assign o[71] = i[1959];
  assign o[70] = i[1958];
  assign o[69] = i[1957];
  assign o[68] = i[1956];
  assign o[67] = i[1955];
  assign o[66] = i[1954];
  assign o[65] = i[1953];
  assign o[64] = i[1952];
  assign o[63] = i[2015];
  assign o[62] = i[2014];
  assign o[61] = i[2013];
  assign o[60] = i[2012];
  assign o[59] = i[2011];
  assign o[58] = i[2010];
  assign o[57] = i[2009];
  assign o[56] = i[2008];
  assign o[55] = i[2007];
  assign o[54] = i[2006];
  assign o[53] = i[2005];
  assign o[52] = i[2004];
  assign o[51] = i[2003];
  assign o[50] = i[2002];
  assign o[49] = i[2001];
  assign o[48] = i[2000];
  assign o[47] = i[1999];
  assign o[46] = i[1998];
  assign o[45] = i[1997];
  assign o[44] = i[1996];
  assign o[43] = i[1995];
  assign o[42] = i[1994];
  assign o[41] = i[1993];
  assign o[40] = i[1992];
  assign o[39] = i[1991];
  assign o[38] = i[1990];
  assign o[37] = i[1989];
  assign o[36] = i[1988];
  assign o[35] = i[1987];
  assign o[34] = i[1986];
  assign o[33] = i[1985];
  assign o[32] = i[1984];
  assign o[31] = i[2047];
  assign o[30] = i[2046];
  assign o[29] = i[2045];
  assign o[28] = i[2044];
  assign o[27] = i[2043];
  assign o[26] = i[2042];
  assign o[25] = i[2041];
  assign o[24] = i[2040];
  assign o[23] = i[2039];
  assign o[22] = i[2038];
  assign o[21] = i[2037];
  assign o[20] = i[2036];
  assign o[19] = i[2035];
  assign o[18] = i[2034];
  assign o[17] = i[2033];
  assign o[16] = i[2032];
  assign o[15] = i[2031];
  assign o[14] = i[2030];
  assign o[13] = i[2029];
  assign o[12] = i[2028];
  assign o[11] = i[2027];
  assign o[10] = i[2026];
  assign o[9] = i[2025];
  assign o[8] = i[2024];
  assign o[7] = i[2023];
  assign o[6] = i[2022];
  assign o[5] = i[2021];
  assign o[4] = i[2020];
  assign o[3] = i[2019];
  assign o[2] = i[2018];
  assign o[1] = i[2017];
  assign o[0] = i[2016];

endmodule



module bsg_parallel_in_serial_out
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_i
);

  input [2047:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_o;
  output valid_o;
  wire [31:0] data_o;
  wire ready_o,valid_o,N0,N1,\piso.done_tx_n ,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,
  N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163;
  wire [5:0] \piso.shift_ctr_r ;
  wire [0:0] \piso.state_n ;
  wire [2047:0] \piso.data_li ,\piso.data_r ;
  reg valid_o_sv2v_reg,\piso.data_r_2047_sv2v_reg ,\piso.data_r_2046_sv2v_reg ,
  \piso.data_r_2045_sv2v_reg ,\piso.data_r_2044_sv2v_reg ,\piso.data_r_2043_sv2v_reg ,
  \piso.data_r_2042_sv2v_reg ,\piso.data_r_2041_sv2v_reg ,
  \piso.data_r_2040_sv2v_reg ,\piso.data_r_2039_sv2v_reg ,\piso.data_r_2038_sv2v_reg ,
  \piso.data_r_2037_sv2v_reg ,\piso.data_r_2036_sv2v_reg ,\piso.data_r_2035_sv2v_reg ,
  \piso.data_r_2034_sv2v_reg ,\piso.data_r_2033_sv2v_reg ,\piso.data_r_2032_sv2v_reg ,
  \piso.data_r_2031_sv2v_reg ,\piso.data_r_2030_sv2v_reg ,\piso.data_r_2029_sv2v_reg ,
  \piso.data_r_2028_sv2v_reg ,\piso.data_r_2027_sv2v_reg ,\piso.data_r_2026_sv2v_reg ,
  \piso.data_r_2025_sv2v_reg ,\piso.data_r_2024_sv2v_reg ,\piso.data_r_2023_sv2v_reg ,
  \piso.data_r_2022_sv2v_reg ,\piso.data_r_2021_sv2v_reg ,
  \piso.data_r_2020_sv2v_reg ,\piso.data_r_2019_sv2v_reg ,\piso.data_r_2018_sv2v_reg ,
  \piso.data_r_2017_sv2v_reg ,\piso.data_r_2016_sv2v_reg ,\piso.data_r_2015_sv2v_reg ,
  \piso.data_r_2014_sv2v_reg ,\piso.data_r_2013_sv2v_reg ,\piso.data_r_2012_sv2v_reg ,
  \piso.data_r_2011_sv2v_reg ,\piso.data_r_2010_sv2v_reg ,\piso.data_r_2009_sv2v_reg ,
  \piso.data_r_2008_sv2v_reg ,\piso.data_r_2007_sv2v_reg ,\piso.data_r_2006_sv2v_reg ,
  \piso.data_r_2005_sv2v_reg ,\piso.data_r_2004_sv2v_reg ,\piso.data_r_2003_sv2v_reg ,
  \piso.data_r_2002_sv2v_reg ,\piso.data_r_2001_sv2v_reg ,
  \piso.data_r_2000_sv2v_reg ,\piso.data_r_1999_sv2v_reg ,\piso.data_r_1998_sv2v_reg ,
  \piso.data_r_1997_sv2v_reg ,\piso.data_r_1996_sv2v_reg ,\piso.data_r_1995_sv2v_reg ,
  \piso.data_r_1994_sv2v_reg ,\piso.data_r_1993_sv2v_reg ,\piso.data_r_1992_sv2v_reg ,
  \piso.data_r_1991_sv2v_reg ,\piso.data_r_1990_sv2v_reg ,\piso.data_r_1989_sv2v_reg ,
  \piso.data_r_1988_sv2v_reg ,\piso.data_r_1987_sv2v_reg ,\piso.data_r_1986_sv2v_reg ,
  \piso.data_r_1985_sv2v_reg ,\piso.data_r_1984_sv2v_reg ,\piso.data_r_1983_sv2v_reg ,
  \piso.data_r_1982_sv2v_reg ,\piso.data_r_1981_sv2v_reg ,
  \piso.data_r_1980_sv2v_reg ,\piso.data_r_1979_sv2v_reg ,\piso.data_r_1978_sv2v_reg ,
  \piso.data_r_1977_sv2v_reg ,\piso.data_r_1976_sv2v_reg ,\piso.data_r_1975_sv2v_reg ,
  \piso.data_r_1974_sv2v_reg ,\piso.data_r_1973_sv2v_reg ,\piso.data_r_1972_sv2v_reg ,
  \piso.data_r_1971_sv2v_reg ,\piso.data_r_1970_sv2v_reg ,\piso.data_r_1969_sv2v_reg ,
  \piso.data_r_1968_sv2v_reg ,\piso.data_r_1967_sv2v_reg ,\piso.data_r_1966_sv2v_reg ,
  \piso.data_r_1965_sv2v_reg ,\piso.data_r_1964_sv2v_reg ,\piso.data_r_1963_sv2v_reg ,
  \piso.data_r_1962_sv2v_reg ,\piso.data_r_1961_sv2v_reg ,
  \piso.data_r_1960_sv2v_reg ,\piso.data_r_1959_sv2v_reg ,\piso.data_r_1958_sv2v_reg ,
  \piso.data_r_1957_sv2v_reg ,\piso.data_r_1956_sv2v_reg ,\piso.data_r_1955_sv2v_reg ,
  \piso.data_r_1954_sv2v_reg ,\piso.data_r_1953_sv2v_reg ,\piso.data_r_1952_sv2v_reg ,
  \piso.data_r_1951_sv2v_reg ,\piso.data_r_1950_sv2v_reg ,\piso.data_r_1949_sv2v_reg ,
  \piso.data_r_1948_sv2v_reg ,\piso.data_r_1947_sv2v_reg ,\piso.data_r_1946_sv2v_reg ,
  \piso.data_r_1945_sv2v_reg ,\piso.data_r_1944_sv2v_reg ,\piso.data_r_1943_sv2v_reg ,
  \piso.data_r_1942_sv2v_reg ,\piso.data_r_1941_sv2v_reg ,
  \piso.data_r_1940_sv2v_reg ,\piso.data_r_1939_sv2v_reg ,\piso.data_r_1938_sv2v_reg ,
  \piso.data_r_1937_sv2v_reg ,\piso.data_r_1936_sv2v_reg ,\piso.data_r_1935_sv2v_reg ,
  \piso.data_r_1934_sv2v_reg ,\piso.data_r_1933_sv2v_reg ,\piso.data_r_1932_sv2v_reg ,
  \piso.data_r_1931_sv2v_reg ,\piso.data_r_1930_sv2v_reg ,\piso.data_r_1929_sv2v_reg ,
  \piso.data_r_1928_sv2v_reg ,\piso.data_r_1927_sv2v_reg ,\piso.data_r_1926_sv2v_reg ,
  \piso.data_r_1925_sv2v_reg ,\piso.data_r_1924_sv2v_reg ,\piso.data_r_1923_sv2v_reg ,
  \piso.data_r_1922_sv2v_reg ,\piso.data_r_1921_sv2v_reg ,
  \piso.data_r_1920_sv2v_reg ,\piso.data_r_1919_sv2v_reg ,\piso.data_r_1918_sv2v_reg ,
  \piso.data_r_1917_sv2v_reg ,\piso.data_r_1916_sv2v_reg ,\piso.data_r_1915_sv2v_reg ,
  \piso.data_r_1914_sv2v_reg ,\piso.data_r_1913_sv2v_reg ,\piso.data_r_1912_sv2v_reg ,
  \piso.data_r_1911_sv2v_reg ,\piso.data_r_1910_sv2v_reg ,\piso.data_r_1909_sv2v_reg ,
  \piso.data_r_1908_sv2v_reg ,\piso.data_r_1907_sv2v_reg ,\piso.data_r_1906_sv2v_reg ,
  \piso.data_r_1905_sv2v_reg ,\piso.data_r_1904_sv2v_reg ,\piso.data_r_1903_sv2v_reg ,
  \piso.data_r_1902_sv2v_reg ,\piso.data_r_1901_sv2v_reg ,
  \piso.data_r_1900_sv2v_reg ,\piso.data_r_1899_sv2v_reg ,\piso.data_r_1898_sv2v_reg ,
  \piso.data_r_1897_sv2v_reg ,\piso.data_r_1896_sv2v_reg ,\piso.data_r_1895_sv2v_reg ,
  \piso.data_r_1894_sv2v_reg ,\piso.data_r_1893_sv2v_reg ,\piso.data_r_1892_sv2v_reg ,
  \piso.data_r_1891_sv2v_reg ,\piso.data_r_1890_sv2v_reg ,\piso.data_r_1889_sv2v_reg ,
  \piso.data_r_1888_sv2v_reg ,\piso.data_r_1887_sv2v_reg ,\piso.data_r_1886_sv2v_reg ,
  \piso.data_r_1885_sv2v_reg ,\piso.data_r_1884_sv2v_reg ,\piso.data_r_1883_sv2v_reg ,
  \piso.data_r_1882_sv2v_reg ,\piso.data_r_1881_sv2v_reg ,
  \piso.data_r_1880_sv2v_reg ,\piso.data_r_1879_sv2v_reg ,\piso.data_r_1878_sv2v_reg ,
  \piso.data_r_1877_sv2v_reg ,\piso.data_r_1876_sv2v_reg ,\piso.data_r_1875_sv2v_reg ,
  \piso.data_r_1874_sv2v_reg ,\piso.data_r_1873_sv2v_reg ,\piso.data_r_1872_sv2v_reg ,
  \piso.data_r_1871_sv2v_reg ,\piso.data_r_1870_sv2v_reg ,\piso.data_r_1869_sv2v_reg ,
  \piso.data_r_1868_sv2v_reg ,\piso.data_r_1867_sv2v_reg ,\piso.data_r_1866_sv2v_reg ,
  \piso.data_r_1865_sv2v_reg ,\piso.data_r_1864_sv2v_reg ,\piso.data_r_1863_sv2v_reg ,
  \piso.data_r_1862_sv2v_reg ,\piso.data_r_1861_sv2v_reg ,
  \piso.data_r_1860_sv2v_reg ,\piso.data_r_1859_sv2v_reg ,\piso.data_r_1858_sv2v_reg ,
  \piso.data_r_1857_sv2v_reg ,\piso.data_r_1856_sv2v_reg ,\piso.data_r_1855_sv2v_reg ,
  \piso.data_r_1854_sv2v_reg ,\piso.data_r_1853_sv2v_reg ,\piso.data_r_1852_sv2v_reg ,
  \piso.data_r_1851_sv2v_reg ,\piso.data_r_1850_sv2v_reg ,\piso.data_r_1849_sv2v_reg ,
  \piso.data_r_1848_sv2v_reg ,\piso.data_r_1847_sv2v_reg ,\piso.data_r_1846_sv2v_reg ,
  \piso.data_r_1845_sv2v_reg ,\piso.data_r_1844_sv2v_reg ,\piso.data_r_1843_sv2v_reg ,
  \piso.data_r_1842_sv2v_reg ,\piso.data_r_1841_sv2v_reg ,
  \piso.data_r_1840_sv2v_reg ,\piso.data_r_1839_sv2v_reg ,\piso.data_r_1838_sv2v_reg ,
  \piso.data_r_1837_sv2v_reg ,\piso.data_r_1836_sv2v_reg ,\piso.data_r_1835_sv2v_reg ,
  \piso.data_r_1834_sv2v_reg ,\piso.data_r_1833_sv2v_reg ,\piso.data_r_1832_sv2v_reg ,
  \piso.data_r_1831_sv2v_reg ,\piso.data_r_1830_sv2v_reg ,\piso.data_r_1829_sv2v_reg ,
  \piso.data_r_1828_sv2v_reg ,\piso.data_r_1827_sv2v_reg ,\piso.data_r_1826_sv2v_reg ,
  \piso.data_r_1825_sv2v_reg ,\piso.data_r_1824_sv2v_reg ,\piso.data_r_1823_sv2v_reg ,
  \piso.data_r_1822_sv2v_reg ,\piso.data_r_1821_sv2v_reg ,
  \piso.data_r_1820_sv2v_reg ,\piso.data_r_1819_sv2v_reg ,\piso.data_r_1818_sv2v_reg ,
  \piso.data_r_1817_sv2v_reg ,\piso.data_r_1816_sv2v_reg ,\piso.data_r_1815_sv2v_reg ,
  \piso.data_r_1814_sv2v_reg ,\piso.data_r_1813_sv2v_reg ,\piso.data_r_1812_sv2v_reg ,
  \piso.data_r_1811_sv2v_reg ,\piso.data_r_1810_sv2v_reg ,\piso.data_r_1809_sv2v_reg ,
  \piso.data_r_1808_sv2v_reg ,\piso.data_r_1807_sv2v_reg ,\piso.data_r_1806_sv2v_reg ,
  \piso.data_r_1805_sv2v_reg ,\piso.data_r_1804_sv2v_reg ,\piso.data_r_1803_sv2v_reg ,
  \piso.data_r_1802_sv2v_reg ,\piso.data_r_1801_sv2v_reg ,
  \piso.data_r_1800_sv2v_reg ,\piso.data_r_1799_sv2v_reg ,\piso.data_r_1798_sv2v_reg ,
  \piso.data_r_1797_sv2v_reg ,\piso.data_r_1796_sv2v_reg ,\piso.data_r_1795_sv2v_reg ,
  \piso.data_r_1794_sv2v_reg ,\piso.data_r_1793_sv2v_reg ,\piso.data_r_1792_sv2v_reg ,
  \piso.data_r_1791_sv2v_reg ,\piso.data_r_1790_sv2v_reg ,\piso.data_r_1789_sv2v_reg ,
  \piso.data_r_1788_sv2v_reg ,\piso.data_r_1787_sv2v_reg ,\piso.data_r_1786_sv2v_reg ,
  \piso.data_r_1785_sv2v_reg ,\piso.data_r_1784_sv2v_reg ,\piso.data_r_1783_sv2v_reg ,
  \piso.data_r_1782_sv2v_reg ,\piso.data_r_1781_sv2v_reg ,
  \piso.data_r_1780_sv2v_reg ,\piso.data_r_1779_sv2v_reg ,\piso.data_r_1778_sv2v_reg ,
  \piso.data_r_1777_sv2v_reg ,\piso.data_r_1776_sv2v_reg ,\piso.data_r_1775_sv2v_reg ,
  \piso.data_r_1774_sv2v_reg ,\piso.data_r_1773_sv2v_reg ,\piso.data_r_1772_sv2v_reg ,
  \piso.data_r_1771_sv2v_reg ,\piso.data_r_1770_sv2v_reg ,\piso.data_r_1769_sv2v_reg ,
  \piso.data_r_1768_sv2v_reg ,\piso.data_r_1767_sv2v_reg ,\piso.data_r_1766_sv2v_reg ,
  \piso.data_r_1765_sv2v_reg ,\piso.data_r_1764_sv2v_reg ,\piso.data_r_1763_sv2v_reg ,
  \piso.data_r_1762_sv2v_reg ,\piso.data_r_1761_sv2v_reg ,
  \piso.data_r_1760_sv2v_reg ,\piso.data_r_1759_sv2v_reg ,\piso.data_r_1758_sv2v_reg ,
  \piso.data_r_1757_sv2v_reg ,\piso.data_r_1756_sv2v_reg ,\piso.data_r_1755_sv2v_reg ,
  \piso.data_r_1754_sv2v_reg ,\piso.data_r_1753_sv2v_reg ,\piso.data_r_1752_sv2v_reg ,
  \piso.data_r_1751_sv2v_reg ,\piso.data_r_1750_sv2v_reg ,\piso.data_r_1749_sv2v_reg ,
  \piso.data_r_1748_sv2v_reg ,\piso.data_r_1747_sv2v_reg ,\piso.data_r_1746_sv2v_reg ,
  \piso.data_r_1745_sv2v_reg ,\piso.data_r_1744_sv2v_reg ,\piso.data_r_1743_sv2v_reg ,
  \piso.data_r_1742_sv2v_reg ,\piso.data_r_1741_sv2v_reg ,
  \piso.data_r_1740_sv2v_reg ,\piso.data_r_1739_sv2v_reg ,\piso.data_r_1738_sv2v_reg ,
  \piso.data_r_1737_sv2v_reg ,\piso.data_r_1736_sv2v_reg ,\piso.data_r_1735_sv2v_reg ,
  \piso.data_r_1734_sv2v_reg ,\piso.data_r_1733_sv2v_reg ,\piso.data_r_1732_sv2v_reg ,
  \piso.data_r_1731_sv2v_reg ,\piso.data_r_1730_sv2v_reg ,\piso.data_r_1729_sv2v_reg ,
  \piso.data_r_1728_sv2v_reg ,\piso.data_r_1727_sv2v_reg ,\piso.data_r_1726_sv2v_reg ,
  \piso.data_r_1725_sv2v_reg ,\piso.data_r_1724_sv2v_reg ,\piso.data_r_1723_sv2v_reg ,
  \piso.data_r_1722_sv2v_reg ,\piso.data_r_1721_sv2v_reg ,
  \piso.data_r_1720_sv2v_reg ,\piso.data_r_1719_sv2v_reg ,\piso.data_r_1718_sv2v_reg ,
  \piso.data_r_1717_sv2v_reg ,\piso.data_r_1716_sv2v_reg ,\piso.data_r_1715_sv2v_reg ,
  \piso.data_r_1714_sv2v_reg ,\piso.data_r_1713_sv2v_reg ,\piso.data_r_1712_sv2v_reg ,
  \piso.data_r_1711_sv2v_reg ,\piso.data_r_1710_sv2v_reg ,\piso.data_r_1709_sv2v_reg ,
  \piso.data_r_1708_sv2v_reg ,\piso.data_r_1707_sv2v_reg ,\piso.data_r_1706_sv2v_reg ,
  \piso.data_r_1705_sv2v_reg ,\piso.data_r_1704_sv2v_reg ,\piso.data_r_1703_sv2v_reg ,
  \piso.data_r_1702_sv2v_reg ,\piso.data_r_1701_sv2v_reg ,
  \piso.data_r_1700_sv2v_reg ,\piso.data_r_1699_sv2v_reg ,\piso.data_r_1698_sv2v_reg ,
  \piso.data_r_1697_sv2v_reg ,\piso.data_r_1696_sv2v_reg ,\piso.data_r_1695_sv2v_reg ,
  \piso.data_r_1694_sv2v_reg ,\piso.data_r_1693_sv2v_reg ,\piso.data_r_1692_sv2v_reg ,
  \piso.data_r_1691_sv2v_reg ,\piso.data_r_1690_sv2v_reg ,\piso.data_r_1689_sv2v_reg ,
  \piso.data_r_1688_sv2v_reg ,\piso.data_r_1687_sv2v_reg ,\piso.data_r_1686_sv2v_reg ,
  \piso.data_r_1685_sv2v_reg ,\piso.data_r_1684_sv2v_reg ,\piso.data_r_1683_sv2v_reg ,
  \piso.data_r_1682_sv2v_reg ,\piso.data_r_1681_sv2v_reg ,
  \piso.data_r_1680_sv2v_reg ,\piso.data_r_1679_sv2v_reg ,\piso.data_r_1678_sv2v_reg ,
  \piso.data_r_1677_sv2v_reg ,\piso.data_r_1676_sv2v_reg ,\piso.data_r_1675_sv2v_reg ,
  \piso.data_r_1674_sv2v_reg ,\piso.data_r_1673_sv2v_reg ,\piso.data_r_1672_sv2v_reg ,
  \piso.data_r_1671_sv2v_reg ,\piso.data_r_1670_sv2v_reg ,\piso.data_r_1669_sv2v_reg ,
  \piso.data_r_1668_sv2v_reg ,\piso.data_r_1667_sv2v_reg ,\piso.data_r_1666_sv2v_reg ,
  \piso.data_r_1665_sv2v_reg ,\piso.data_r_1664_sv2v_reg ,\piso.data_r_1663_sv2v_reg ,
  \piso.data_r_1662_sv2v_reg ,\piso.data_r_1661_sv2v_reg ,
  \piso.data_r_1660_sv2v_reg ,\piso.data_r_1659_sv2v_reg ,\piso.data_r_1658_sv2v_reg ,
  \piso.data_r_1657_sv2v_reg ,\piso.data_r_1656_sv2v_reg ,\piso.data_r_1655_sv2v_reg ,
  \piso.data_r_1654_sv2v_reg ,\piso.data_r_1653_sv2v_reg ,\piso.data_r_1652_sv2v_reg ,
  \piso.data_r_1651_sv2v_reg ,\piso.data_r_1650_sv2v_reg ,\piso.data_r_1649_sv2v_reg ,
  \piso.data_r_1648_sv2v_reg ,\piso.data_r_1647_sv2v_reg ,\piso.data_r_1646_sv2v_reg ,
  \piso.data_r_1645_sv2v_reg ,\piso.data_r_1644_sv2v_reg ,\piso.data_r_1643_sv2v_reg ,
  \piso.data_r_1642_sv2v_reg ,\piso.data_r_1641_sv2v_reg ,
  \piso.data_r_1640_sv2v_reg ,\piso.data_r_1639_sv2v_reg ,\piso.data_r_1638_sv2v_reg ,
  \piso.data_r_1637_sv2v_reg ,\piso.data_r_1636_sv2v_reg ,\piso.data_r_1635_sv2v_reg ,
  \piso.data_r_1634_sv2v_reg ,\piso.data_r_1633_sv2v_reg ,\piso.data_r_1632_sv2v_reg ,
  \piso.data_r_1631_sv2v_reg ,\piso.data_r_1630_sv2v_reg ,\piso.data_r_1629_sv2v_reg ,
  \piso.data_r_1628_sv2v_reg ,\piso.data_r_1627_sv2v_reg ,\piso.data_r_1626_sv2v_reg ,
  \piso.data_r_1625_sv2v_reg ,\piso.data_r_1624_sv2v_reg ,\piso.data_r_1623_sv2v_reg ,
  \piso.data_r_1622_sv2v_reg ,\piso.data_r_1621_sv2v_reg ,
  \piso.data_r_1620_sv2v_reg ,\piso.data_r_1619_sv2v_reg ,\piso.data_r_1618_sv2v_reg ,
  \piso.data_r_1617_sv2v_reg ,\piso.data_r_1616_sv2v_reg ,\piso.data_r_1615_sv2v_reg ,
  \piso.data_r_1614_sv2v_reg ,\piso.data_r_1613_sv2v_reg ,\piso.data_r_1612_sv2v_reg ,
  \piso.data_r_1611_sv2v_reg ,\piso.data_r_1610_sv2v_reg ,\piso.data_r_1609_sv2v_reg ,
  \piso.data_r_1608_sv2v_reg ,\piso.data_r_1607_sv2v_reg ,\piso.data_r_1606_sv2v_reg ,
  \piso.data_r_1605_sv2v_reg ,\piso.data_r_1604_sv2v_reg ,\piso.data_r_1603_sv2v_reg ,
  \piso.data_r_1602_sv2v_reg ,\piso.data_r_1601_sv2v_reg ,
  \piso.data_r_1600_sv2v_reg ,\piso.data_r_1599_sv2v_reg ,\piso.data_r_1598_sv2v_reg ,
  \piso.data_r_1597_sv2v_reg ,\piso.data_r_1596_sv2v_reg ,\piso.data_r_1595_sv2v_reg ,
  \piso.data_r_1594_sv2v_reg ,\piso.data_r_1593_sv2v_reg ,\piso.data_r_1592_sv2v_reg ,
  \piso.data_r_1591_sv2v_reg ,\piso.data_r_1590_sv2v_reg ,\piso.data_r_1589_sv2v_reg ,
  \piso.data_r_1588_sv2v_reg ,\piso.data_r_1587_sv2v_reg ,\piso.data_r_1586_sv2v_reg ,
  \piso.data_r_1585_sv2v_reg ,\piso.data_r_1584_sv2v_reg ,\piso.data_r_1583_sv2v_reg ,
  \piso.data_r_1582_sv2v_reg ,\piso.data_r_1581_sv2v_reg ,
  \piso.data_r_1580_sv2v_reg ,\piso.data_r_1579_sv2v_reg ,\piso.data_r_1578_sv2v_reg ,
  \piso.data_r_1577_sv2v_reg ,\piso.data_r_1576_sv2v_reg ,\piso.data_r_1575_sv2v_reg ,
  \piso.data_r_1574_sv2v_reg ,\piso.data_r_1573_sv2v_reg ,\piso.data_r_1572_sv2v_reg ,
  \piso.data_r_1571_sv2v_reg ,\piso.data_r_1570_sv2v_reg ,\piso.data_r_1569_sv2v_reg ,
  \piso.data_r_1568_sv2v_reg ,\piso.data_r_1567_sv2v_reg ,\piso.data_r_1566_sv2v_reg ,
  \piso.data_r_1565_sv2v_reg ,\piso.data_r_1564_sv2v_reg ,\piso.data_r_1563_sv2v_reg ,
  \piso.data_r_1562_sv2v_reg ,\piso.data_r_1561_sv2v_reg ,
  \piso.data_r_1560_sv2v_reg ,\piso.data_r_1559_sv2v_reg ,\piso.data_r_1558_sv2v_reg ,
  \piso.data_r_1557_sv2v_reg ,\piso.data_r_1556_sv2v_reg ,\piso.data_r_1555_sv2v_reg ,
  \piso.data_r_1554_sv2v_reg ,\piso.data_r_1553_sv2v_reg ,\piso.data_r_1552_sv2v_reg ,
  \piso.data_r_1551_sv2v_reg ,\piso.data_r_1550_sv2v_reg ,\piso.data_r_1549_sv2v_reg ,
  \piso.data_r_1548_sv2v_reg ,\piso.data_r_1547_sv2v_reg ,\piso.data_r_1546_sv2v_reg ,
  \piso.data_r_1545_sv2v_reg ,\piso.data_r_1544_sv2v_reg ,\piso.data_r_1543_sv2v_reg ,
  \piso.data_r_1542_sv2v_reg ,\piso.data_r_1541_sv2v_reg ,
  \piso.data_r_1540_sv2v_reg ,\piso.data_r_1539_sv2v_reg ,\piso.data_r_1538_sv2v_reg ,
  \piso.data_r_1537_sv2v_reg ,\piso.data_r_1536_sv2v_reg ,\piso.data_r_1535_sv2v_reg ,
  \piso.data_r_1534_sv2v_reg ,\piso.data_r_1533_sv2v_reg ,\piso.data_r_1532_sv2v_reg ,
  \piso.data_r_1531_sv2v_reg ,\piso.data_r_1530_sv2v_reg ,\piso.data_r_1529_sv2v_reg ,
  \piso.data_r_1528_sv2v_reg ,\piso.data_r_1527_sv2v_reg ,\piso.data_r_1526_sv2v_reg ,
  \piso.data_r_1525_sv2v_reg ,\piso.data_r_1524_sv2v_reg ,\piso.data_r_1523_sv2v_reg ,
  \piso.data_r_1522_sv2v_reg ,\piso.data_r_1521_sv2v_reg ,
  \piso.data_r_1520_sv2v_reg ,\piso.data_r_1519_sv2v_reg ,\piso.data_r_1518_sv2v_reg ,
  \piso.data_r_1517_sv2v_reg ,\piso.data_r_1516_sv2v_reg ,\piso.data_r_1515_sv2v_reg ,
  \piso.data_r_1514_sv2v_reg ,\piso.data_r_1513_sv2v_reg ,\piso.data_r_1512_sv2v_reg ,
  \piso.data_r_1511_sv2v_reg ,\piso.data_r_1510_sv2v_reg ,\piso.data_r_1509_sv2v_reg ,
  \piso.data_r_1508_sv2v_reg ,\piso.data_r_1507_sv2v_reg ,\piso.data_r_1506_sv2v_reg ,
  \piso.data_r_1505_sv2v_reg ,\piso.data_r_1504_sv2v_reg ,\piso.data_r_1503_sv2v_reg ,
  \piso.data_r_1502_sv2v_reg ,\piso.data_r_1501_sv2v_reg ,
  \piso.data_r_1500_sv2v_reg ,\piso.data_r_1499_sv2v_reg ,\piso.data_r_1498_sv2v_reg ,
  \piso.data_r_1497_sv2v_reg ,\piso.data_r_1496_sv2v_reg ,\piso.data_r_1495_sv2v_reg ,
  \piso.data_r_1494_sv2v_reg ,\piso.data_r_1493_sv2v_reg ,\piso.data_r_1492_sv2v_reg ,
  \piso.data_r_1491_sv2v_reg ,\piso.data_r_1490_sv2v_reg ,\piso.data_r_1489_sv2v_reg ,
  \piso.data_r_1488_sv2v_reg ,\piso.data_r_1487_sv2v_reg ,\piso.data_r_1486_sv2v_reg ,
  \piso.data_r_1485_sv2v_reg ,\piso.data_r_1484_sv2v_reg ,\piso.data_r_1483_sv2v_reg ,
  \piso.data_r_1482_sv2v_reg ,\piso.data_r_1481_sv2v_reg ,
  \piso.data_r_1480_sv2v_reg ,\piso.data_r_1479_sv2v_reg ,\piso.data_r_1478_sv2v_reg ,
  \piso.data_r_1477_sv2v_reg ,\piso.data_r_1476_sv2v_reg ,\piso.data_r_1475_sv2v_reg ,
  \piso.data_r_1474_sv2v_reg ,\piso.data_r_1473_sv2v_reg ,\piso.data_r_1472_sv2v_reg ,
  \piso.data_r_1471_sv2v_reg ,\piso.data_r_1470_sv2v_reg ,\piso.data_r_1469_sv2v_reg ,
  \piso.data_r_1468_sv2v_reg ,\piso.data_r_1467_sv2v_reg ,\piso.data_r_1466_sv2v_reg ,
  \piso.data_r_1465_sv2v_reg ,\piso.data_r_1464_sv2v_reg ,\piso.data_r_1463_sv2v_reg ,
  \piso.data_r_1462_sv2v_reg ,\piso.data_r_1461_sv2v_reg ,
  \piso.data_r_1460_sv2v_reg ,\piso.data_r_1459_sv2v_reg ,\piso.data_r_1458_sv2v_reg ,
  \piso.data_r_1457_sv2v_reg ,\piso.data_r_1456_sv2v_reg ,\piso.data_r_1455_sv2v_reg ,
  \piso.data_r_1454_sv2v_reg ,\piso.data_r_1453_sv2v_reg ,\piso.data_r_1452_sv2v_reg ,
  \piso.data_r_1451_sv2v_reg ,\piso.data_r_1450_sv2v_reg ,\piso.data_r_1449_sv2v_reg ,
  \piso.data_r_1448_sv2v_reg ,\piso.data_r_1447_sv2v_reg ,\piso.data_r_1446_sv2v_reg ,
  \piso.data_r_1445_sv2v_reg ,\piso.data_r_1444_sv2v_reg ,\piso.data_r_1443_sv2v_reg ,
  \piso.data_r_1442_sv2v_reg ,\piso.data_r_1441_sv2v_reg ,
  \piso.data_r_1440_sv2v_reg ,\piso.data_r_1439_sv2v_reg ,\piso.data_r_1438_sv2v_reg ,
  \piso.data_r_1437_sv2v_reg ,\piso.data_r_1436_sv2v_reg ,\piso.data_r_1435_sv2v_reg ,
  \piso.data_r_1434_sv2v_reg ,\piso.data_r_1433_sv2v_reg ,\piso.data_r_1432_sv2v_reg ,
  \piso.data_r_1431_sv2v_reg ,\piso.data_r_1430_sv2v_reg ,\piso.data_r_1429_sv2v_reg ,
  \piso.data_r_1428_sv2v_reg ,\piso.data_r_1427_sv2v_reg ,\piso.data_r_1426_sv2v_reg ,
  \piso.data_r_1425_sv2v_reg ,\piso.data_r_1424_sv2v_reg ,\piso.data_r_1423_sv2v_reg ,
  \piso.data_r_1422_sv2v_reg ,\piso.data_r_1421_sv2v_reg ,
  \piso.data_r_1420_sv2v_reg ,\piso.data_r_1419_sv2v_reg ,\piso.data_r_1418_sv2v_reg ,
  \piso.data_r_1417_sv2v_reg ,\piso.data_r_1416_sv2v_reg ,\piso.data_r_1415_sv2v_reg ,
  \piso.data_r_1414_sv2v_reg ,\piso.data_r_1413_sv2v_reg ,\piso.data_r_1412_sv2v_reg ,
  \piso.data_r_1411_sv2v_reg ,\piso.data_r_1410_sv2v_reg ,\piso.data_r_1409_sv2v_reg ,
  \piso.data_r_1408_sv2v_reg ,\piso.data_r_1407_sv2v_reg ,\piso.data_r_1406_sv2v_reg ,
  \piso.data_r_1405_sv2v_reg ,\piso.data_r_1404_sv2v_reg ,\piso.data_r_1403_sv2v_reg ,
  \piso.data_r_1402_sv2v_reg ,\piso.data_r_1401_sv2v_reg ,
  \piso.data_r_1400_sv2v_reg ,\piso.data_r_1399_sv2v_reg ,\piso.data_r_1398_sv2v_reg ,
  \piso.data_r_1397_sv2v_reg ,\piso.data_r_1396_sv2v_reg ,\piso.data_r_1395_sv2v_reg ,
  \piso.data_r_1394_sv2v_reg ,\piso.data_r_1393_sv2v_reg ,\piso.data_r_1392_sv2v_reg ,
  \piso.data_r_1391_sv2v_reg ,\piso.data_r_1390_sv2v_reg ,\piso.data_r_1389_sv2v_reg ,
  \piso.data_r_1388_sv2v_reg ,\piso.data_r_1387_sv2v_reg ,\piso.data_r_1386_sv2v_reg ,
  \piso.data_r_1385_sv2v_reg ,\piso.data_r_1384_sv2v_reg ,\piso.data_r_1383_sv2v_reg ,
  \piso.data_r_1382_sv2v_reg ,\piso.data_r_1381_sv2v_reg ,
  \piso.data_r_1380_sv2v_reg ,\piso.data_r_1379_sv2v_reg ,\piso.data_r_1378_sv2v_reg ,
  \piso.data_r_1377_sv2v_reg ,\piso.data_r_1376_sv2v_reg ,\piso.data_r_1375_sv2v_reg ,
  \piso.data_r_1374_sv2v_reg ,\piso.data_r_1373_sv2v_reg ,\piso.data_r_1372_sv2v_reg ,
  \piso.data_r_1371_sv2v_reg ,\piso.data_r_1370_sv2v_reg ,\piso.data_r_1369_sv2v_reg ,
  \piso.data_r_1368_sv2v_reg ,\piso.data_r_1367_sv2v_reg ,\piso.data_r_1366_sv2v_reg ,
  \piso.data_r_1365_sv2v_reg ,\piso.data_r_1364_sv2v_reg ,\piso.data_r_1363_sv2v_reg ,
  \piso.data_r_1362_sv2v_reg ,\piso.data_r_1361_sv2v_reg ,
  \piso.data_r_1360_sv2v_reg ,\piso.data_r_1359_sv2v_reg ,\piso.data_r_1358_sv2v_reg ,
  \piso.data_r_1357_sv2v_reg ,\piso.data_r_1356_sv2v_reg ,\piso.data_r_1355_sv2v_reg ,
  \piso.data_r_1354_sv2v_reg ,\piso.data_r_1353_sv2v_reg ,\piso.data_r_1352_sv2v_reg ,
  \piso.data_r_1351_sv2v_reg ,\piso.data_r_1350_sv2v_reg ,\piso.data_r_1349_sv2v_reg ,
  \piso.data_r_1348_sv2v_reg ,\piso.data_r_1347_sv2v_reg ,\piso.data_r_1346_sv2v_reg ,
  \piso.data_r_1345_sv2v_reg ,\piso.data_r_1344_sv2v_reg ,\piso.data_r_1343_sv2v_reg ,
  \piso.data_r_1342_sv2v_reg ,\piso.data_r_1341_sv2v_reg ,
  \piso.data_r_1340_sv2v_reg ,\piso.data_r_1339_sv2v_reg ,\piso.data_r_1338_sv2v_reg ,
  \piso.data_r_1337_sv2v_reg ,\piso.data_r_1336_sv2v_reg ,\piso.data_r_1335_sv2v_reg ,
  \piso.data_r_1334_sv2v_reg ,\piso.data_r_1333_sv2v_reg ,\piso.data_r_1332_sv2v_reg ,
  \piso.data_r_1331_sv2v_reg ,\piso.data_r_1330_sv2v_reg ,\piso.data_r_1329_sv2v_reg ,
  \piso.data_r_1328_sv2v_reg ,\piso.data_r_1327_sv2v_reg ,\piso.data_r_1326_sv2v_reg ,
  \piso.data_r_1325_sv2v_reg ,\piso.data_r_1324_sv2v_reg ,\piso.data_r_1323_sv2v_reg ,
  \piso.data_r_1322_sv2v_reg ,\piso.data_r_1321_sv2v_reg ,
  \piso.data_r_1320_sv2v_reg ,\piso.data_r_1319_sv2v_reg ,\piso.data_r_1318_sv2v_reg ,
  \piso.data_r_1317_sv2v_reg ,\piso.data_r_1316_sv2v_reg ,\piso.data_r_1315_sv2v_reg ,
  \piso.data_r_1314_sv2v_reg ,\piso.data_r_1313_sv2v_reg ,\piso.data_r_1312_sv2v_reg ,
  \piso.data_r_1311_sv2v_reg ,\piso.data_r_1310_sv2v_reg ,\piso.data_r_1309_sv2v_reg ,
  \piso.data_r_1308_sv2v_reg ,\piso.data_r_1307_sv2v_reg ,\piso.data_r_1306_sv2v_reg ,
  \piso.data_r_1305_sv2v_reg ,\piso.data_r_1304_sv2v_reg ,\piso.data_r_1303_sv2v_reg ,
  \piso.data_r_1302_sv2v_reg ,\piso.data_r_1301_sv2v_reg ,
  \piso.data_r_1300_sv2v_reg ,\piso.data_r_1299_sv2v_reg ,\piso.data_r_1298_sv2v_reg ,
  \piso.data_r_1297_sv2v_reg ,\piso.data_r_1296_sv2v_reg ,\piso.data_r_1295_sv2v_reg ,
  \piso.data_r_1294_sv2v_reg ,\piso.data_r_1293_sv2v_reg ,\piso.data_r_1292_sv2v_reg ,
  \piso.data_r_1291_sv2v_reg ,\piso.data_r_1290_sv2v_reg ,\piso.data_r_1289_sv2v_reg ,
  \piso.data_r_1288_sv2v_reg ,\piso.data_r_1287_sv2v_reg ,\piso.data_r_1286_sv2v_reg ,
  \piso.data_r_1285_sv2v_reg ,\piso.data_r_1284_sv2v_reg ,\piso.data_r_1283_sv2v_reg ,
  \piso.data_r_1282_sv2v_reg ,\piso.data_r_1281_sv2v_reg ,
  \piso.data_r_1280_sv2v_reg ,\piso.data_r_1279_sv2v_reg ,\piso.data_r_1278_sv2v_reg ,
  \piso.data_r_1277_sv2v_reg ,\piso.data_r_1276_sv2v_reg ,\piso.data_r_1275_sv2v_reg ,
  \piso.data_r_1274_sv2v_reg ,\piso.data_r_1273_sv2v_reg ,\piso.data_r_1272_sv2v_reg ,
  \piso.data_r_1271_sv2v_reg ,\piso.data_r_1270_sv2v_reg ,\piso.data_r_1269_sv2v_reg ,
  \piso.data_r_1268_sv2v_reg ,\piso.data_r_1267_sv2v_reg ,\piso.data_r_1266_sv2v_reg ,
  \piso.data_r_1265_sv2v_reg ,\piso.data_r_1264_sv2v_reg ,\piso.data_r_1263_sv2v_reg ,
  \piso.data_r_1262_sv2v_reg ,\piso.data_r_1261_sv2v_reg ,
  \piso.data_r_1260_sv2v_reg ,\piso.data_r_1259_sv2v_reg ,\piso.data_r_1258_sv2v_reg ,
  \piso.data_r_1257_sv2v_reg ,\piso.data_r_1256_sv2v_reg ,\piso.data_r_1255_sv2v_reg ,
  \piso.data_r_1254_sv2v_reg ,\piso.data_r_1253_sv2v_reg ,\piso.data_r_1252_sv2v_reg ,
  \piso.data_r_1251_sv2v_reg ,\piso.data_r_1250_sv2v_reg ,\piso.data_r_1249_sv2v_reg ,
  \piso.data_r_1248_sv2v_reg ,\piso.data_r_1247_sv2v_reg ,\piso.data_r_1246_sv2v_reg ,
  \piso.data_r_1245_sv2v_reg ,\piso.data_r_1244_sv2v_reg ,\piso.data_r_1243_sv2v_reg ,
  \piso.data_r_1242_sv2v_reg ,\piso.data_r_1241_sv2v_reg ,
  \piso.data_r_1240_sv2v_reg ,\piso.data_r_1239_sv2v_reg ,\piso.data_r_1238_sv2v_reg ,
  \piso.data_r_1237_sv2v_reg ,\piso.data_r_1236_sv2v_reg ,\piso.data_r_1235_sv2v_reg ,
  \piso.data_r_1234_sv2v_reg ,\piso.data_r_1233_sv2v_reg ,\piso.data_r_1232_sv2v_reg ,
  \piso.data_r_1231_sv2v_reg ,\piso.data_r_1230_sv2v_reg ,\piso.data_r_1229_sv2v_reg ,
  \piso.data_r_1228_sv2v_reg ,\piso.data_r_1227_sv2v_reg ,\piso.data_r_1226_sv2v_reg ,
  \piso.data_r_1225_sv2v_reg ,\piso.data_r_1224_sv2v_reg ,\piso.data_r_1223_sv2v_reg ,
  \piso.data_r_1222_sv2v_reg ,\piso.data_r_1221_sv2v_reg ,
  \piso.data_r_1220_sv2v_reg ,\piso.data_r_1219_sv2v_reg ,\piso.data_r_1218_sv2v_reg ,
  \piso.data_r_1217_sv2v_reg ,\piso.data_r_1216_sv2v_reg ,\piso.data_r_1215_sv2v_reg ,
  \piso.data_r_1214_sv2v_reg ,\piso.data_r_1213_sv2v_reg ,\piso.data_r_1212_sv2v_reg ,
  \piso.data_r_1211_sv2v_reg ,\piso.data_r_1210_sv2v_reg ,\piso.data_r_1209_sv2v_reg ,
  \piso.data_r_1208_sv2v_reg ,\piso.data_r_1207_sv2v_reg ,\piso.data_r_1206_sv2v_reg ,
  \piso.data_r_1205_sv2v_reg ,\piso.data_r_1204_sv2v_reg ,\piso.data_r_1203_sv2v_reg ,
  \piso.data_r_1202_sv2v_reg ,\piso.data_r_1201_sv2v_reg ,
  \piso.data_r_1200_sv2v_reg ,\piso.data_r_1199_sv2v_reg ,\piso.data_r_1198_sv2v_reg ,
  \piso.data_r_1197_sv2v_reg ,\piso.data_r_1196_sv2v_reg ,\piso.data_r_1195_sv2v_reg ,
  \piso.data_r_1194_sv2v_reg ,\piso.data_r_1193_sv2v_reg ,\piso.data_r_1192_sv2v_reg ,
  \piso.data_r_1191_sv2v_reg ,\piso.data_r_1190_sv2v_reg ,\piso.data_r_1189_sv2v_reg ,
  \piso.data_r_1188_sv2v_reg ,\piso.data_r_1187_sv2v_reg ,\piso.data_r_1186_sv2v_reg ,
  \piso.data_r_1185_sv2v_reg ,\piso.data_r_1184_sv2v_reg ,\piso.data_r_1183_sv2v_reg ,
  \piso.data_r_1182_sv2v_reg ,\piso.data_r_1181_sv2v_reg ,
  \piso.data_r_1180_sv2v_reg ,\piso.data_r_1179_sv2v_reg ,\piso.data_r_1178_sv2v_reg ,
  \piso.data_r_1177_sv2v_reg ,\piso.data_r_1176_sv2v_reg ,\piso.data_r_1175_sv2v_reg ,
  \piso.data_r_1174_sv2v_reg ,\piso.data_r_1173_sv2v_reg ,\piso.data_r_1172_sv2v_reg ,
  \piso.data_r_1171_sv2v_reg ,\piso.data_r_1170_sv2v_reg ,\piso.data_r_1169_sv2v_reg ,
  \piso.data_r_1168_sv2v_reg ,\piso.data_r_1167_sv2v_reg ,\piso.data_r_1166_sv2v_reg ,
  \piso.data_r_1165_sv2v_reg ,\piso.data_r_1164_sv2v_reg ,\piso.data_r_1163_sv2v_reg ,
  \piso.data_r_1162_sv2v_reg ,\piso.data_r_1161_sv2v_reg ,
  \piso.data_r_1160_sv2v_reg ,\piso.data_r_1159_sv2v_reg ,\piso.data_r_1158_sv2v_reg ,
  \piso.data_r_1157_sv2v_reg ,\piso.data_r_1156_sv2v_reg ,\piso.data_r_1155_sv2v_reg ,
  \piso.data_r_1154_sv2v_reg ,\piso.data_r_1153_sv2v_reg ,\piso.data_r_1152_sv2v_reg ,
  \piso.data_r_1151_sv2v_reg ,\piso.data_r_1150_sv2v_reg ,\piso.data_r_1149_sv2v_reg ,
  \piso.data_r_1148_sv2v_reg ,\piso.data_r_1147_sv2v_reg ,\piso.data_r_1146_sv2v_reg ,
  \piso.data_r_1145_sv2v_reg ,\piso.data_r_1144_sv2v_reg ,\piso.data_r_1143_sv2v_reg ,
  \piso.data_r_1142_sv2v_reg ,\piso.data_r_1141_sv2v_reg ,
  \piso.data_r_1140_sv2v_reg ,\piso.data_r_1139_sv2v_reg ,\piso.data_r_1138_sv2v_reg ,
  \piso.data_r_1137_sv2v_reg ,\piso.data_r_1136_sv2v_reg ,\piso.data_r_1135_sv2v_reg ,
  \piso.data_r_1134_sv2v_reg ,\piso.data_r_1133_sv2v_reg ,\piso.data_r_1132_sv2v_reg ,
  \piso.data_r_1131_sv2v_reg ,\piso.data_r_1130_sv2v_reg ,\piso.data_r_1129_sv2v_reg ,
  \piso.data_r_1128_sv2v_reg ,\piso.data_r_1127_sv2v_reg ,\piso.data_r_1126_sv2v_reg ,
  \piso.data_r_1125_sv2v_reg ,\piso.data_r_1124_sv2v_reg ,\piso.data_r_1123_sv2v_reg ,
  \piso.data_r_1122_sv2v_reg ,\piso.data_r_1121_sv2v_reg ,
  \piso.data_r_1120_sv2v_reg ,\piso.data_r_1119_sv2v_reg ,\piso.data_r_1118_sv2v_reg ,
  \piso.data_r_1117_sv2v_reg ,\piso.data_r_1116_sv2v_reg ,\piso.data_r_1115_sv2v_reg ,
  \piso.data_r_1114_sv2v_reg ,\piso.data_r_1113_sv2v_reg ,\piso.data_r_1112_sv2v_reg ,
  \piso.data_r_1111_sv2v_reg ,\piso.data_r_1110_sv2v_reg ,\piso.data_r_1109_sv2v_reg ,
  \piso.data_r_1108_sv2v_reg ,\piso.data_r_1107_sv2v_reg ,\piso.data_r_1106_sv2v_reg ,
  \piso.data_r_1105_sv2v_reg ,\piso.data_r_1104_sv2v_reg ,\piso.data_r_1103_sv2v_reg ,
  \piso.data_r_1102_sv2v_reg ,\piso.data_r_1101_sv2v_reg ,
  \piso.data_r_1100_sv2v_reg ,\piso.data_r_1099_sv2v_reg ,\piso.data_r_1098_sv2v_reg ,
  \piso.data_r_1097_sv2v_reg ,\piso.data_r_1096_sv2v_reg ,\piso.data_r_1095_sv2v_reg ,
  \piso.data_r_1094_sv2v_reg ,\piso.data_r_1093_sv2v_reg ,\piso.data_r_1092_sv2v_reg ,
  \piso.data_r_1091_sv2v_reg ,\piso.data_r_1090_sv2v_reg ,\piso.data_r_1089_sv2v_reg ,
  \piso.data_r_1088_sv2v_reg ,\piso.data_r_1087_sv2v_reg ,\piso.data_r_1086_sv2v_reg ,
  \piso.data_r_1085_sv2v_reg ,\piso.data_r_1084_sv2v_reg ,\piso.data_r_1083_sv2v_reg ,
  \piso.data_r_1082_sv2v_reg ,\piso.data_r_1081_sv2v_reg ,
  \piso.data_r_1080_sv2v_reg ,\piso.data_r_1079_sv2v_reg ,\piso.data_r_1078_sv2v_reg ,
  \piso.data_r_1077_sv2v_reg ,\piso.data_r_1076_sv2v_reg ,\piso.data_r_1075_sv2v_reg ,
  \piso.data_r_1074_sv2v_reg ,\piso.data_r_1073_sv2v_reg ,\piso.data_r_1072_sv2v_reg ,
  \piso.data_r_1071_sv2v_reg ,\piso.data_r_1070_sv2v_reg ,\piso.data_r_1069_sv2v_reg ,
  \piso.data_r_1068_sv2v_reg ,\piso.data_r_1067_sv2v_reg ,\piso.data_r_1066_sv2v_reg ,
  \piso.data_r_1065_sv2v_reg ,\piso.data_r_1064_sv2v_reg ,\piso.data_r_1063_sv2v_reg ,
  \piso.data_r_1062_sv2v_reg ,\piso.data_r_1061_sv2v_reg ,
  \piso.data_r_1060_sv2v_reg ,\piso.data_r_1059_sv2v_reg ,\piso.data_r_1058_sv2v_reg ,
  \piso.data_r_1057_sv2v_reg ,\piso.data_r_1056_sv2v_reg ,\piso.data_r_1055_sv2v_reg ,
  \piso.data_r_1054_sv2v_reg ,\piso.data_r_1053_sv2v_reg ,\piso.data_r_1052_sv2v_reg ,
  \piso.data_r_1051_sv2v_reg ,\piso.data_r_1050_sv2v_reg ,\piso.data_r_1049_sv2v_reg ,
  \piso.data_r_1048_sv2v_reg ,\piso.data_r_1047_sv2v_reg ,\piso.data_r_1046_sv2v_reg ,
  \piso.data_r_1045_sv2v_reg ,\piso.data_r_1044_sv2v_reg ,\piso.data_r_1043_sv2v_reg ,
  \piso.data_r_1042_sv2v_reg ,\piso.data_r_1041_sv2v_reg ,
  \piso.data_r_1040_sv2v_reg ,\piso.data_r_1039_sv2v_reg ,\piso.data_r_1038_sv2v_reg ,
  \piso.data_r_1037_sv2v_reg ,\piso.data_r_1036_sv2v_reg ,\piso.data_r_1035_sv2v_reg ,
  \piso.data_r_1034_sv2v_reg ,\piso.data_r_1033_sv2v_reg ,\piso.data_r_1032_sv2v_reg ,
  \piso.data_r_1031_sv2v_reg ,\piso.data_r_1030_sv2v_reg ,\piso.data_r_1029_sv2v_reg ,
  \piso.data_r_1028_sv2v_reg ,\piso.data_r_1027_sv2v_reg ,\piso.data_r_1026_sv2v_reg ,
  \piso.data_r_1025_sv2v_reg ,\piso.data_r_1024_sv2v_reg ,\piso.data_r_1023_sv2v_reg ,
  \piso.data_r_1022_sv2v_reg ,\piso.data_r_1021_sv2v_reg ,
  \piso.data_r_1020_sv2v_reg ,\piso.data_r_1019_sv2v_reg ,\piso.data_r_1018_sv2v_reg ,
  \piso.data_r_1017_sv2v_reg ,\piso.data_r_1016_sv2v_reg ,\piso.data_r_1015_sv2v_reg ,
  \piso.data_r_1014_sv2v_reg ,\piso.data_r_1013_sv2v_reg ,\piso.data_r_1012_sv2v_reg ,
  \piso.data_r_1011_sv2v_reg ,\piso.data_r_1010_sv2v_reg ,\piso.data_r_1009_sv2v_reg ,
  \piso.data_r_1008_sv2v_reg ,\piso.data_r_1007_sv2v_reg ,\piso.data_r_1006_sv2v_reg ,
  \piso.data_r_1005_sv2v_reg ,\piso.data_r_1004_sv2v_reg ,\piso.data_r_1003_sv2v_reg ,
  \piso.data_r_1002_sv2v_reg ,\piso.data_r_1001_sv2v_reg ,
  \piso.data_r_1000_sv2v_reg ,\piso.data_r_999_sv2v_reg ,\piso.data_r_998_sv2v_reg ,
  \piso.data_r_997_sv2v_reg ,\piso.data_r_996_sv2v_reg ,\piso.data_r_995_sv2v_reg ,
  \piso.data_r_994_sv2v_reg ,\piso.data_r_993_sv2v_reg ,\piso.data_r_992_sv2v_reg ,
  \piso.data_r_991_sv2v_reg ,\piso.data_r_990_sv2v_reg ,\piso.data_r_989_sv2v_reg ,
  \piso.data_r_988_sv2v_reg ,\piso.data_r_987_sv2v_reg ,\piso.data_r_986_sv2v_reg ,
  \piso.data_r_985_sv2v_reg ,\piso.data_r_984_sv2v_reg ,\piso.data_r_983_sv2v_reg ,
  \piso.data_r_982_sv2v_reg ,\piso.data_r_981_sv2v_reg ,\piso.data_r_980_sv2v_reg ,
  \piso.data_r_979_sv2v_reg ,\piso.data_r_978_sv2v_reg ,\piso.data_r_977_sv2v_reg ,
  \piso.data_r_976_sv2v_reg ,\piso.data_r_975_sv2v_reg ,\piso.data_r_974_sv2v_reg ,
  \piso.data_r_973_sv2v_reg ,\piso.data_r_972_sv2v_reg ,\piso.data_r_971_sv2v_reg ,
  \piso.data_r_970_sv2v_reg ,\piso.data_r_969_sv2v_reg ,\piso.data_r_968_sv2v_reg ,
  \piso.data_r_967_sv2v_reg ,\piso.data_r_966_sv2v_reg ,\piso.data_r_965_sv2v_reg ,
  \piso.data_r_964_sv2v_reg ,\piso.data_r_963_sv2v_reg ,\piso.data_r_962_sv2v_reg ,
  \piso.data_r_961_sv2v_reg ,\piso.data_r_960_sv2v_reg ,\piso.data_r_959_sv2v_reg ,
  \piso.data_r_958_sv2v_reg ,\piso.data_r_957_sv2v_reg ,\piso.data_r_956_sv2v_reg ,
  \piso.data_r_955_sv2v_reg ,\piso.data_r_954_sv2v_reg ,\piso.data_r_953_sv2v_reg ,
  \piso.data_r_952_sv2v_reg ,\piso.data_r_951_sv2v_reg ,\piso.data_r_950_sv2v_reg ,
  \piso.data_r_949_sv2v_reg ,\piso.data_r_948_sv2v_reg ,\piso.data_r_947_sv2v_reg ,
  \piso.data_r_946_sv2v_reg ,\piso.data_r_945_sv2v_reg ,\piso.data_r_944_sv2v_reg ,
  \piso.data_r_943_sv2v_reg ,\piso.data_r_942_sv2v_reg ,\piso.data_r_941_sv2v_reg ,
  \piso.data_r_940_sv2v_reg ,\piso.data_r_939_sv2v_reg ,\piso.data_r_938_sv2v_reg ,
  \piso.data_r_937_sv2v_reg ,\piso.data_r_936_sv2v_reg ,\piso.data_r_935_sv2v_reg ,
  \piso.data_r_934_sv2v_reg ,\piso.data_r_933_sv2v_reg ,\piso.data_r_932_sv2v_reg ,
  \piso.data_r_931_sv2v_reg ,\piso.data_r_930_sv2v_reg ,\piso.data_r_929_sv2v_reg ,
  \piso.data_r_928_sv2v_reg ,\piso.data_r_927_sv2v_reg ,\piso.data_r_926_sv2v_reg ,
  \piso.data_r_925_sv2v_reg ,\piso.data_r_924_sv2v_reg ,\piso.data_r_923_sv2v_reg ,
  \piso.data_r_922_sv2v_reg ,\piso.data_r_921_sv2v_reg ,
  \piso.data_r_920_sv2v_reg ,\piso.data_r_919_sv2v_reg ,\piso.data_r_918_sv2v_reg ,
  \piso.data_r_917_sv2v_reg ,\piso.data_r_916_sv2v_reg ,\piso.data_r_915_sv2v_reg ,
  \piso.data_r_914_sv2v_reg ,\piso.data_r_913_sv2v_reg ,\piso.data_r_912_sv2v_reg ,
  \piso.data_r_911_sv2v_reg ,\piso.data_r_910_sv2v_reg ,\piso.data_r_909_sv2v_reg ,
  \piso.data_r_908_sv2v_reg ,\piso.data_r_907_sv2v_reg ,\piso.data_r_906_sv2v_reg ,
  \piso.data_r_905_sv2v_reg ,\piso.data_r_904_sv2v_reg ,\piso.data_r_903_sv2v_reg ,
  \piso.data_r_902_sv2v_reg ,\piso.data_r_901_sv2v_reg ,\piso.data_r_900_sv2v_reg ,
  \piso.data_r_899_sv2v_reg ,\piso.data_r_898_sv2v_reg ,\piso.data_r_897_sv2v_reg ,
  \piso.data_r_896_sv2v_reg ,\piso.data_r_895_sv2v_reg ,\piso.data_r_894_sv2v_reg ,
  \piso.data_r_893_sv2v_reg ,\piso.data_r_892_sv2v_reg ,\piso.data_r_891_sv2v_reg ,
  \piso.data_r_890_sv2v_reg ,\piso.data_r_889_sv2v_reg ,\piso.data_r_888_sv2v_reg ,
  \piso.data_r_887_sv2v_reg ,\piso.data_r_886_sv2v_reg ,\piso.data_r_885_sv2v_reg ,
  \piso.data_r_884_sv2v_reg ,\piso.data_r_883_sv2v_reg ,\piso.data_r_882_sv2v_reg ,
  \piso.data_r_881_sv2v_reg ,\piso.data_r_880_sv2v_reg ,\piso.data_r_879_sv2v_reg ,
  \piso.data_r_878_sv2v_reg ,\piso.data_r_877_sv2v_reg ,\piso.data_r_876_sv2v_reg ,
  \piso.data_r_875_sv2v_reg ,\piso.data_r_874_sv2v_reg ,\piso.data_r_873_sv2v_reg ,
  \piso.data_r_872_sv2v_reg ,\piso.data_r_871_sv2v_reg ,\piso.data_r_870_sv2v_reg ,
  \piso.data_r_869_sv2v_reg ,\piso.data_r_868_sv2v_reg ,\piso.data_r_867_sv2v_reg ,
  \piso.data_r_866_sv2v_reg ,\piso.data_r_865_sv2v_reg ,\piso.data_r_864_sv2v_reg ,
  \piso.data_r_863_sv2v_reg ,\piso.data_r_862_sv2v_reg ,\piso.data_r_861_sv2v_reg ,
  \piso.data_r_860_sv2v_reg ,\piso.data_r_859_sv2v_reg ,\piso.data_r_858_sv2v_reg ,
  \piso.data_r_857_sv2v_reg ,\piso.data_r_856_sv2v_reg ,\piso.data_r_855_sv2v_reg ,
  \piso.data_r_854_sv2v_reg ,\piso.data_r_853_sv2v_reg ,\piso.data_r_852_sv2v_reg ,
  \piso.data_r_851_sv2v_reg ,\piso.data_r_850_sv2v_reg ,\piso.data_r_849_sv2v_reg ,
  \piso.data_r_848_sv2v_reg ,\piso.data_r_847_sv2v_reg ,\piso.data_r_846_sv2v_reg ,
  \piso.data_r_845_sv2v_reg ,\piso.data_r_844_sv2v_reg ,\piso.data_r_843_sv2v_reg ,
  \piso.data_r_842_sv2v_reg ,\piso.data_r_841_sv2v_reg ,
  \piso.data_r_840_sv2v_reg ,\piso.data_r_839_sv2v_reg ,\piso.data_r_838_sv2v_reg ,
  \piso.data_r_837_sv2v_reg ,\piso.data_r_836_sv2v_reg ,\piso.data_r_835_sv2v_reg ,
  \piso.data_r_834_sv2v_reg ,\piso.data_r_833_sv2v_reg ,\piso.data_r_832_sv2v_reg ,
  \piso.data_r_831_sv2v_reg ,\piso.data_r_830_sv2v_reg ,\piso.data_r_829_sv2v_reg ,
  \piso.data_r_828_sv2v_reg ,\piso.data_r_827_sv2v_reg ,\piso.data_r_826_sv2v_reg ,
  \piso.data_r_825_sv2v_reg ,\piso.data_r_824_sv2v_reg ,\piso.data_r_823_sv2v_reg ,
  \piso.data_r_822_sv2v_reg ,\piso.data_r_821_sv2v_reg ,\piso.data_r_820_sv2v_reg ,
  \piso.data_r_819_sv2v_reg ,\piso.data_r_818_sv2v_reg ,\piso.data_r_817_sv2v_reg ,
  \piso.data_r_816_sv2v_reg ,\piso.data_r_815_sv2v_reg ,\piso.data_r_814_sv2v_reg ,
  \piso.data_r_813_sv2v_reg ,\piso.data_r_812_sv2v_reg ,\piso.data_r_811_sv2v_reg ,
  \piso.data_r_810_sv2v_reg ,\piso.data_r_809_sv2v_reg ,\piso.data_r_808_sv2v_reg ,
  \piso.data_r_807_sv2v_reg ,\piso.data_r_806_sv2v_reg ,\piso.data_r_805_sv2v_reg ,
  \piso.data_r_804_sv2v_reg ,\piso.data_r_803_sv2v_reg ,\piso.data_r_802_sv2v_reg ,
  \piso.data_r_801_sv2v_reg ,\piso.data_r_800_sv2v_reg ,\piso.data_r_799_sv2v_reg ,
  \piso.data_r_798_sv2v_reg ,\piso.data_r_797_sv2v_reg ,\piso.data_r_796_sv2v_reg ,
  \piso.data_r_795_sv2v_reg ,\piso.data_r_794_sv2v_reg ,\piso.data_r_793_sv2v_reg ,
  \piso.data_r_792_sv2v_reg ,\piso.data_r_791_sv2v_reg ,\piso.data_r_790_sv2v_reg ,
  \piso.data_r_789_sv2v_reg ,\piso.data_r_788_sv2v_reg ,\piso.data_r_787_sv2v_reg ,
  \piso.data_r_786_sv2v_reg ,\piso.data_r_785_sv2v_reg ,\piso.data_r_784_sv2v_reg ,
  \piso.data_r_783_sv2v_reg ,\piso.data_r_782_sv2v_reg ,\piso.data_r_781_sv2v_reg ,
  \piso.data_r_780_sv2v_reg ,\piso.data_r_779_sv2v_reg ,\piso.data_r_778_sv2v_reg ,
  \piso.data_r_777_sv2v_reg ,\piso.data_r_776_sv2v_reg ,\piso.data_r_775_sv2v_reg ,
  \piso.data_r_774_sv2v_reg ,\piso.data_r_773_sv2v_reg ,\piso.data_r_772_sv2v_reg ,
  \piso.data_r_771_sv2v_reg ,\piso.data_r_770_sv2v_reg ,\piso.data_r_769_sv2v_reg ,
  \piso.data_r_768_sv2v_reg ,\piso.data_r_767_sv2v_reg ,\piso.data_r_766_sv2v_reg ,
  \piso.data_r_765_sv2v_reg ,\piso.data_r_764_sv2v_reg ,\piso.data_r_763_sv2v_reg ,
  \piso.data_r_762_sv2v_reg ,\piso.data_r_761_sv2v_reg ,
  \piso.data_r_760_sv2v_reg ,\piso.data_r_759_sv2v_reg ,\piso.data_r_758_sv2v_reg ,
  \piso.data_r_757_sv2v_reg ,\piso.data_r_756_sv2v_reg ,\piso.data_r_755_sv2v_reg ,
  \piso.data_r_754_sv2v_reg ,\piso.data_r_753_sv2v_reg ,\piso.data_r_752_sv2v_reg ,
  \piso.data_r_751_sv2v_reg ,\piso.data_r_750_sv2v_reg ,\piso.data_r_749_sv2v_reg ,
  \piso.data_r_748_sv2v_reg ,\piso.data_r_747_sv2v_reg ,\piso.data_r_746_sv2v_reg ,
  \piso.data_r_745_sv2v_reg ,\piso.data_r_744_sv2v_reg ,\piso.data_r_743_sv2v_reg ,
  \piso.data_r_742_sv2v_reg ,\piso.data_r_741_sv2v_reg ,\piso.data_r_740_sv2v_reg ,
  \piso.data_r_739_sv2v_reg ,\piso.data_r_738_sv2v_reg ,\piso.data_r_737_sv2v_reg ,
  \piso.data_r_736_sv2v_reg ,\piso.data_r_735_sv2v_reg ,\piso.data_r_734_sv2v_reg ,
  \piso.data_r_733_sv2v_reg ,\piso.data_r_732_sv2v_reg ,\piso.data_r_731_sv2v_reg ,
  \piso.data_r_730_sv2v_reg ,\piso.data_r_729_sv2v_reg ,\piso.data_r_728_sv2v_reg ,
  \piso.data_r_727_sv2v_reg ,\piso.data_r_726_sv2v_reg ,\piso.data_r_725_sv2v_reg ,
  \piso.data_r_724_sv2v_reg ,\piso.data_r_723_sv2v_reg ,\piso.data_r_722_sv2v_reg ,
  \piso.data_r_721_sv2v_reg ,\piso.data_r_720_sv2v_reg ,\piso.data_r_719_sv2v_reg ,
  \piso.data_r_718_sv2v_reg ,\piso.data_r_717_sv2v_reg ,\piso.data_r_716_sv2v_reg ,
  \piso.data_r_715_sv2v_reg ,\piso.data_r_714_sv2v_reg ,\piso.data_r_713_sv2v_reg ,
  \piso.data_r_712_sv2v_reg ,\piso.data_r_711_sv2v_reg ,\piso.data_r_710_sv2v_reg ,
  \piso.data_r_709_sv2v_reg ,\piso.data_r_708_sv2v_reg ,\piso.data_r_707_sv2v_reg ,
  \piso.data_r_706_sv2v_reg ,\piso.data_r_705_sv2v_reg ,\piso.data_r_704_sv2v_reg ,
  \piso.data_r_703_sv2v_reg ,\piso.data_r_702_sv2v_reg ,\piso.data_r_701_sv2v_reg ,
  \piso.data_r_700_sv2v_reg ,\piso.data_r_699_sv2v_reg ,\piso.data_r_698_sv2v_reg ,
  \piso.data_r_697_sv2v_reg ,\piso.data_r_696_sv2v_reg ,\piso.data_r_695_sv2v_reg ,
  \piso.data_r_694_sv2v_reg ,\piso.data_r_693_sv2v_reg ,\piso.data_r_692_sv2v_reg ,
  \piso.data_r_691_sv2v_reg ,\piso.data_r_690_sv2v_reg ,\piso.data_r_689_sv2v_reg ,
  \piso.data_r_688_sv2v_reg ,\piso.data_r_687_sv2v_reg ,\piso.data_r_686_sv2v_reg ,
  \piso.data_r_685_sv2v_reg ,\piso.data_r_684_sv2v_reg ,\piso.data_r_683_sv2v_reg ,
  \piso.data_r_682_sv2v_reg ,\piso.data_r_681_sv2v_reg ,
  \piso.data_r_680_sv2v_reg ,\piso.data_r_679_sv2v_reg ,\piso.data_r_678_sv2v_reg ,
  \piso.data_r_677_sv2v_reg ,\piso.data_r_676_sv2v_reg ,\piso.data_r_675_sv2v_reg ,
  \piso.data_r_674_sv2v_reg ,\piso.data_r_673_sv2v_reg ,\piso.data_r_672_sv2v_reg ,
  \piso.data_r_671_sv2v_reg ,\piso.data_r_670_sv2v_reg ,\piso.data_r_669_sv2v_reg ,
  \piso.data_r_668_sv2v_reg ,\piso.data_r_667_sv2v_reg ,\piso.data_r_666_sv2v_reg ,
  \piso.data_r_665_sv2v_reg ,\piso.data_r_664_sv2v_reg ,\piso.data_r_663_sv2v_reg ,
  \piso.data_r_662_sv2v_reg ,\piso.data_r_661_sv2v_reg ,\piso.data_r_660_sv2v_reg ,
  \piso.data_r_659_sv2v_reg ,\piso.data_r_658_sv2v_reg ,\piso.data_r_657_sv2v_reg ,
  \piso.data_r_656_sv2v_reg ,\piso.data_r_655_sv2v_reg ,\piso.data_r_654_sv2v_reg ,
  \piso.data_r_653_sv2v_reg ,\piso.data_r_652_sv2v_reg ,\piso.data_r_651_sv2v_reg ,
  \piso.data_r_650_sv2v_reg ,\piso.data_r_649_sv2v_reg ,\piso.data_r_648_sv2v_reg ,
  \piso.data_r_647_sv2v_reg ,\piso.data_r_646_sv2v_reg ,\piso.data_r_645_sv2v_reg ,
  \piso.data_r_644_sv2v_reg ,\piso.data_r_643_sv2v_reg ,\piso.data_r_642_sv2v_reg ,
  \piso.data_r_641_sv2v_reg ,\piso.data_r_640_sv2v_reg ,\piso.data_r_639_sv2v_reg ,
  \piso.data_r_638_sv2v_reg ,\piso.data_r_637_sv2v_reg ,\piso.data_r_636_sv2v_reg ,
  \piso.data_r_635_sv2v_reg ,\piso.data_r_634_sv2v_reg ,\piso.data_r_633_sv2v_reg ,
  \piso.data_r_632_sv2v_reg ,\piso.data_r_631_sv2v_reg ,\piso.data_r_630_sv2v_reg ,
  \piso.data_r_629_sv2v_reg ,\piso.data_r_628_sv2v_reg ,\piso.data_r_627_sv2v_reg ,
  \piso.data_r_626_sv2v_reg ,\piso.data_r_625_sv2v_reg ,\piso.data_r_624_sv2v_reg ,
  \piso.data_r_623_sv2v_reg ,\piso.data_r_622_sv2v_reg ,\piso.data_r_621_sv2v_reg ,
  \piso.data_r_620_sv2v_reg ,\piso.data_r_619_sv2v_reg ,\piso.data_r_618_sv2v_reg ,
  \piso.data_r_617_sv2v_reg ,\piso.data_r_616_sv2v_reg ,\piso.data_r_615_sv2v_reg ,
  \piso.data_r_614_sv2v_reg ,\piso.data_r_613_sv2v_reg ,\piso.data_r_612_sv2v_reg ,
  \piso.data_r_611_sv2v_reg ,\piso.data_r_610_sv2v_reg ,\piso.data_r_609_sv2v_reg ,
  \piso.data_r_608_sv2v_reg ,\piso.data_r_607_sv2v_reg ,\piso.data_r_606_sv2v_reg ,
  \piso.data_r_605_sv2v_reg ,\piso.data_r_604_sv2v_reg ,\piso.data_r_603_sv2v_reg ,
  \piso.data_r_602_sv2v_reg ,\piso.data_r_601_sv2v_reg ,
  \piso.data_r_600_sv2v_reg ,\piso.data_r_599_sv2v_reg ,\piso.data_r_598_sv2v_reg ,
  \piso.data_r_597_sv2v_reg ,\piso.data_r_596_sv2v_reg ,\piso.data_r_595_sv2v_reg ,
  \piso.data_r_594_sv2v_reg ,\piso.data_r_593_sv2v_reg ,\piso.data_r_592_sv2v_reg ,
  \piso.data_r_591_sv2v_reg ,\piso.data_r_590_sv2v_reg ,\piso.data_r_589_sv2v_reg ,
  \piso.data_r_588_sv2v_reg ,\piso.data_r_587_sv2v_reg ,\piso.data_r_586_sv2v_reg ,
  \piso.data_r_585_sv2v_reg ,\piso.data_r_584_sv2v_reg ,\piso.data_r_583_sv2v_reg ,
  \piso.data_r_582_sv2v_reg ,\piso.data_r_581_sv2v_reg ,\piso.data_r_580_sv2v_reg ,
  \piso.data_r_579_sv2v_reg ,\piso.data_r_578_sv2v_reg ,\piso.data_r_577_sv2v_reg ,
  \piso.data_r_576_sv2v_reg ,\piso.data_r_575_sv2v_reg ,\piso.data_r_574_sv2v_reg ,
  \piso.data_r_573_sv2v_reg ,\piso.data_r_572_sv2v_reg ,\piso.data_r_571_sv2v_reg ,
  \piso.data_r_570_sv2v_reg ,\piso.data_r_569_sv2v_reg ,\piso.data_r_568_sv2v_reg ,
  \piso.data_r_567_sv2v_reg ,\piso.data_r_566_sv2v_reg ,\piso.data_r_565_sv2v_reg ,
  \piso.data_r_564_sv2v_reg ,\piso.data_r_563_sv2v_reg ,\piso.data_r_562_sv2v_reg ,
  \piso.data_r_561_sv2v_reg ,\piso.data_r_560_sv2v_reg ,\piso.data_r_559_sv2v_reg ,
  \piso.data_r_558_sv2v_reg ,\piso.data_r_557_sv2v_reg ,\piso.data_r_556_sv2v_reg ,
  \piso.data_r_555_sv2v_reg ,\piso.data_r_554_sv2v_reg ,\piso.data_r_553_sv2v_reg ,
  \piso.data_r_552_sv2v_reg ,\piso.data_r_551_sv2v_reg ,\piso.data_r_550_sv2v_reg ,
  \piso.data_r_549_sv2v_reg ,\piso.data_r_548_sv2v_reg ,\piso.data_r_547_sv2v_reg ,
  \piso.data_r_546_sv2v_reg ,\piso.data_r_545_sv2v_reg ,\piso.data_r_544_sv2v_reg ,
  \piso.data_r_543_sv2v_reg ,\piso.data_r_542_sv2v_reg ,\piso.data_r_541_sv2v_reg ,
  \piso.data_r_540_sv2v_reg ,\piso.data_r_539_sv2v_reg ,\piso.data_r_538_sv2v_reg ,
  \piso.data_r_537_sv2v_reg ,\piso.data_r_536_sv2v_reg ,\piso.data_r_535_sv2v_reg ,
  \piso.data_r_534_sv2v_reg ,\piso.data_r_533_sv2v_reg ,\piso.data_r_532_sv2v_reg ,
  \piso.data_r_531_sv2v_reg ,\piso.data_r_530_sv2v_reg ,\piso.data_r_529_sv2v_reg ,
  \piso.data_r_528_sv2v_reg ,\piso.data_r_527_sv2v_reg ,\piso.data_r_526_sv2v_reg ,
  \piso.data_r_525_sv2v_reg ,\piso.data_r_524_sv2v_reg ,\piso.data_r_523_sv2v_reg ,
  \piso.data_r_522_sv2v_reg ,\piso.data_r_521_sv2v_reg ,
  \piso.data_r_520_sv2v_reg ,\piso.data_r_519_sv2v_reg ,\piso.data_r_518_sv2v_reg ,
  \piso.data_r_517_sv2v_reg ,\piso.data_r_516_sv2v_reg ,\piso.data_r_515_sv2v_reg ,
  \piso.data_r_514_sv2v_reg ,\piso.data_r_513_sv2v_reg ,\piso.data_r_512_sv2v_reg ,
  \piso.data_r_511_sv2v_reg ,\piso.data_r_510_sv2v_reg ,\piso.data_r_509_sv2v_reg ,
  \piso.data_r_508_sv2v_reg ,\piso.data_r_507_sv2v_reg ,\piso.data_r_506_sv2v_reg ,
  \piso.data_r_505_sv2v_reg ,\piso.data_r_504_sv2v_reg ,\piso.data_r_503_sv2v_reg ,
  \piso.data_r_502_sv2v_reg ,\piso.data_r_501_sv2v_reg ,\piso.data_r_500_sv2v_reg ,
  \piso.data_r_499_sv2v_reg ,\piso.data_r_498_sv2v_reg ,\piso.data_r_497_sv2v_reg ,
  \piso.data_r_496_sv2v_reg ,\piso.data_r_495_sv2v_reg ,\piso.data_r_494_sv2v_reg ,
  \piso.data_r_493_sv2v_reg ,\piso.data_r_492_sv2v_reg ,\piso.data_r_491_sv2v_reg ,
  \piso.data_r_490_sv2v_reg ,\piso.data_r_489_sv2v_reg ,\piso.data_r_488_sv2v_reg ,
  \piso.data_r_487_sv2v_reg ,\piso.data_r_486_sv2v_reg ,\piso.data_r_485_sv2v_reg ,
  \piso.data_r_484_sv2v_reg ,\piso.data_r_483_sv2v_reg ,\piso.data_r_482_sv2v_reg ,
  \piso.data_r_481_sv2v_reg ,\piso.data_r_480_sv2v_reg ,\piso.data_r_479_sv2v_reg ,
  \piso.data_r_478_sv2v_reg ,\piso.data_r_477_sv2v_reg ,\piso.data_r_476_sv2v_reg ,
  \piso.data_r_475_sv2v_reg ,\piso.data_r_474_sv2v_reg ,\piso.data_r_473_sv2v_reg ,
  \piso.data_r_472_sv2v_reg ,\piso.data_r_471_sv2v_reg ,\piso.data_r_470_sv2v_reg ,
  \piso.data_r_469_sv2v_reg ,\piso.data_r_468_sv2v_reg ,\piso.data_r_467_sv2v_reg ,
  \piso.data_r_466_sv2v_reg ,\piso.data_r_465_sv2v_reg ,\piso.data_r_464_sv2v_reg ,
  \piso.data_r_463_sv2v_reg ,\piso.data_r_462_sv2v_reg ,\piso.data_r_461_sv2v_reg ,
  \piso.data_r_460_sv2v_reg ,\piso.data_r_459_sv2v_reg ,\piso.data_r_458_sv2v_reg ,
  \piso.data_r_457_sv2v_reg ,\piso.data_r_456_sv2v_reg ,\piso.data_r_455_sv2v_reg ,
  \piso.data_r_454_sv2v_reg ,\piso.data_r_453_sv2v_reg ,\piso.data_r_452_sv2v_reg ,
  \piso.data_r_451_sv2v_reg ,\piso.data_r_450_sv2v_reg ,\piso.data_r_449_sv2v_reg ,
  \piso.data_r_448_sv2v_reg ,\piso.data_r_447_sv2v_reg ,\piso.data_r_446_sv2v_reg ,
  \piso.data_r_445_sv2v_reg ,\piso.data_r_444_sv2v_reg ,\piso.data_r_443_sv2v_reg ,
  \piso.data_r_442_sv2v_reg ,\piso.data_r_441_sv2v_reg ,
  \piso.data_r_440_sv2v_reg ,\piso.data_r_439_sv2v_reg ,\piso.data_r_438_sv2v_reg ,
  \piso.data_r_437_sv2v_reg ,\piso.data_r_436_sv2v_reg ,\piso.data_r_435_sv2v_reg ,
  \piso.data_r_434_sv2v_reg ,\piso.data_r_433_sv2v_reg ,\piso.data_r_432_sv2v_reg ,
  \piso.data_r_431_sv2v_reg ,\piso.data_r_430_sv2v_reg ,\piso.data_r_429_sv2v_reg ,
  \piso.data_r_428_sv2v_reg ,\piso.data_r_427_sv2v_reg ,\piso.data_r_426_sv2v_reg ,
  \piso.data_r_425_sv2v_reg ,\piso.data_r_424_sv2v_reg ,\piso.data_r_423_sv2v_reg ,
  \piso.data_r_422_sv2v_reg ,\piso.data_r_421_sv2v_reg ,\piso.data_r_420_sv2v_reg ,
  \piso.data_r_419_sv2v_reg ,\piso.data_r_418_sv2v_reg ,\piso.data_r_417_sv2v_reg ,
  \piso.data_r_416_sv2v_reg ,\piso.data_r_415_sv2v_reg ,\piso.data_r_414_sv2v_reg ,
  \piso.data_r_413_sv2v_reg ,\piso.data_r_412_sv2v_reg ,\piso.data_r_411_sv2v_reg ,
  \piso.data_r_410_sv2v_reg ,\piso.data_r_409_sv2v_reg ,\piso.data_r_408_sv2v_reg ,
  \piso.data_r_407_sv2v_reg ,\piso.data_r_406_sv2v_reg ,\piso.data_r_405_sv2v_reg ,
  \piso.data_r_404_sv2v_reg ,\piso.data_r_403_sv2v_reg ,\piso.data_r_402_sv2v_reg ,
  \piso.data_r_401_sv2v_reg ,\piso.data_r_400_sv2v_reg ,\piso.data_r_399_sv2v_reg ,
  \piso.data_r_398_sv2v_reg ,\piso.data_r_397_sv2v_reg ,\piso.data_r_396_sv2v_reg ,
  \piso.data_r_395_sv2v_reg ,\piso.data_r_394_sv2v_reg ,\piso.data_r_393_sv2v_reg ,
  \piso.data_r_392_sv2v_reg ,\piso.data_r_391_sv2v_reg ,\piso.data_r_390_sv2v_reg ,
  \piso.data_r_389_sv2v_reg ,\piso.data_r_388_sv2v_reg ,\piso.data_r_387_sv2v_reg ,
  \piso.data_r_386_sv2v_reg ,\piso.data_r_385_sv2v_reg ,\piso.data_r_384_sv2v_reg ,
  \piso.data_r_383_sv2v_reg ,\piso.data_r_382_sv2v_reg ,\piso.data_r_381_sv2v_reg ,
  \piso.data_r_380_sv2v_reg ,\piso.data_r_379_sv2v_reg ,\piso.data_r_378_sv2v_reg ,
  \piso.data_r_377_sv2v_reg ,\piso.data_r_376_sv2v_reg ,\piso.data_r_375_sv2v_reg ,
  \piso.data_r_374_sv2v_reg ,\piso.data_r_373_sv2v_reg ,\piso.data_r_372_sv2v_reg ,
  \piso.data_r_371_sv2v_reg ,\piso.data_r_370_sv2v_reg ,\piso.data_r_369_sv2v_reg ,
  \piso.data_r_368_sv2v_reg ,\piso.data_r_367_sv2v_reg ,\piso.data_r_366_sv2v_reg ,
  \piso.data_r_365_sv2v_reg ,\piso.data_r_364_sv2v_reg ,\piso.data_r_363_sv2v_reg ,
  \piso.data_r_362_sv2v_reg ,\piso.data_r_361_sv2v_reg ,
  \piso.data_r_360_sv2v_reg ,\piso.data_r_359_sv2v_reg ,\piso.data_r_358_sv2v_reg ,
  \piso.data_r_357_sv2v_reg ,\piso.data_r_356_sv2v_reg ,\piso.data_r_355_sv2v_reg ,
  \piso.data_r_354_sv2v_reg ,\piso.data_r_353_sv2v_reg ,\piso.data_r_352_sv2v_reg ,
  \piso.data_r_351_sv2v_reg ,\piso.data_r_350_sv2v_reg ,\piso.data_r_349_sv2v_reg ,
  \piso.data_r_348_sv2v_reg ,\piso.data_r_347_sv2v_reg ,\piso.data_r_346_sv2v_reg ,
  \piso.data_r_345_sv2v_reg ,\piso.data_r_344_sv2v_reg ,\piso.data_r_343_sv2v_reg ,
  \piso.data_r_342_sv2v_reg ,\piso.data_r_341_sv2v_reg ,\piso.data_r_340_sv2v_reg ,
  \piso.data_r_339_sv2v_reg ,\piso.data_r_338_sv2v_reg ,\piso.data_r_337_sv2v_reg ,
  \piso.data_r_336_sv2v_reg ,\piso.data_r_335_sv2v_reg ,\piso.data_r_334_sv2v_reg ,
  \piso.data_r_333_sv2v_reg ,\piso.data_r_332_sv2v_reg ,\piso.data_r_331_sv2v_reg ,
  \piso.data_r_330_sv2v_reg ,\piso.data_r_329_sv2v_reg ,\piso.data_r_328_sv2v_reg ,
  \piso.data_r_327_sv2v_reg ,\piso.data_r_326_sv2v_reg ,\piso.data_r_325_sv2v_reg ,
  \piso.data_r_324_sv2v_reg ,\piso.data_r_323_sv2v_reg ,\piso.data_r_322_sv2v_reg ,
  \piso.data_r_321_sv2v_reg ,\piso.data_r_320_sv2v_reg ,\piso.data_r_319_sv2v_reg ,
  \piso.data_r_318_sv2v_reg ,\piso.data_r_317_sv2v_reg ,\piso.data_r_316_sv2v_reg ,
  \piso.data_r_315_sv2v_reg ,\piso.data_r_314_sv2v_reg ,\piso.data_r_313_sv2v_reg ,
  \piso.data_r_312_sv2v_reg ,\piso.data_r_311_sv2v_reg ,\piso.data_r_310_sv2v_reg ,
  \piso.data_r_309_sv2v_reg ,\piso.data_r_308_sv2v_reg ,\piso.data_r_307_sv2v_reg ,
  \piso.data_r_306_sv2v_reg ,\piso.data_r_305_sv2v_reg ,\piso.data_r_304_sv2v_reg ,
  \piso.data_r_303_sv2v_reg ,\piso.data_r_302_sv2v_reg ,\piso.data_r_301_sv2v_reg ,
  \piso.data_r_300_sv2v_reg ,\piso.data_r_299_sv2v_reg ,\piso.data_r_298_sv2v_reg ,
  \piso.data_r_297_sv2v_reg ,\piso.data_r_296_sv2v_reg ,\piso.data_r_295_sv2v_reg ,
  \piso.data_r_294_sv2v_reg ,\piso.data_r_293_sv2v_reg ,\piso.data_r_292_sv2v_reg ,
  \piso.data_r_291_sv2v_reg ,\piso.data_r_290_sv2v_reg ,\piso.data_r_289_sv2v_reg ,
  \piso.data_r_288_sv2v_reg ,\piso.data_r_287_sv2v_reg ,\piso.data_r_286_sv2v_reg ,
  \piso.data_r_285_sv2v_reg ,\piso.data_r_284_sv2v_reg ,\piso.data_r_283_sv2v_reg ,
  \piso.data_r_282_sv2v_reg ,\piso.data_r_281_sv2v_reg ,
  \piso.data_r_280_sv2v_reg ,\piso.data_r_279_sv2v_reg ,\piso.data_r_278_sv2v_reg ,
  \piso.data_r_277_sv2v_reg ,\piso.data_r_276_sv2v_reg ,\piso.data_r_275_sv2v_reg ,
  \piso.data_r_274_sv2v_reg ,\piso.data_r_273_sv2v_reg ,\piso.data_r_272_sv2v_reg ,
  \piso.data_r_271_sv2v_reg ,\piso.data_r_270_sv2v_reg ,\piso.data_r_269_sv2v_reg ,
  \piso.data_r_268_sv2v_reg ,\piso.data_r_267_sv2v_reg ,\piso.data_r_266_sv2v_reg ,
  \piso.data_r_265_sv2v_reg ,\piso.data_r_264_sv2v_reg ,\piso.data_r_263_sv2v_reg ,
  \piso.data_r_262_sv2v_reg ,\piso.data_r_261_sv2v_reg ,\piso.data_r_260_sv2v_reg ,
  \piso.data_r_259_sv2v_reg ,\piso.data_r_258_sv2v_reg ,\piso.data_r_257_sv2v_reg ,
  \piso.data_r_256_sv2v_reg ,\piso.data_r_255_sv2v_reg ,\piso.data_r_254_sv2v_reg ,
  \piso.data_r_253_sv2v_reg ,\piso.data_r_252_sv2v_reg ,\piso.data_r_251_sv2v_reg ,
  \piso.data_r_250_sv2v_reg ,\piso.data_r_249_sv2v_reg ,\piso.data_r_248_sv2v_reg ,
  \piso.data_r_247_sv2v_reg ,\piso.data_r_246_sv2v_reg ,\piso.data_r_245_sv2v_reg ,
  \piso.data_r_244_sv2v_reg ,\piso.data_r_243_sv2v_reg ,\piso.data_r_242_sv2v_reg ,
  \piso.data_r_241_sv2v_reg ,\piso.data_r_240_sv2v_reg ,\piso.data_r_239_sv2v_reg ,
  \piso.data_r_238_sv2v_reg ,\piso.data_r_237_sv2v_reg ,\piso.data_r_236_sv2v_reg ,
  \piso.data_r_235_sv2v_reg ,\piso.data_r_234_sv2v_reg ,\piso.data_r_233_sv2v_reg ,
  \piso.data_r_232_sv2v_reg ,\piso.data_r_231_sv2v_reg ,\piso.data_r_230_sv2v_reg ,
  \piso.data_r_229_sv2v_reg ,\piso.data_r_228_sv2v_reg ,\piso.data_r_227_sv2v_reg ,
  \piso.data_r_226_sv2v_reg ,\piso.data_r_225_sv2v_reg ,\piso.data_r_224_sv2v_reg ,
  \piso.data_r_223_sv2v_reg ,\piso.data_r_222_sv2v_reg ,\piso.data_r_221_sv2v_reg ,
  \piso.data_r_220_sv2v_reg ,\piso.data_r_219_sv2v_reg ,\piso.data_r_218_sv2v_reg ,
  \piso.data_r_217_sv2v_reg ,\piso.data_r_216_sv2v_reg ,\piso.data_r_215_sv2v_reg ,
  \piso.data_r_214_sv2v_reg ,\piso.data_r_213_sv2v_reg ,\piso.data_r_212_sv2v_reg ,
  \piso.data_r_211_sv2v_reg ,\piso.data_r_210_sv2v_reg ,\piso.data_r_209_sv2v_reg ,
  \piso.data_r_208_sv2v_reg ,\piso.data_r_207_sv2v_reg ,\piso.data_r_206_sv2v_reg ,
  \piso.data_r_205_sv2v_reg ,\piso.data_r_204_sv2v_reg ,\piso.data_r_203_sv2v_reg ,
  \piso.data_r_202_sv2v_reg ,\piso.data_r_201_sv2v_reg ,
  \piso.data_r_200_sv2v_reg ,\piso.data_r_199_sv2v_reg ,\piso.data_r_198_sv2v_reg ,
  \piso.data_r_197_sv2v_reg ,\piso.data_r_196_sv2v_reg ,\piso.data_r_195_sv2v_reg ,
  \piso.data_r_194_sv2v_reg ,\piso.data_r_193_sv2v_reg ,\piso.data_r_192_sv2v_reg ,
  \piso.data_r_191_sv2v_reg ,\piso.data_r_190_sv2v_reg ,\piso.data_r_189_sv2v_reg ,
  \piso.data_r_188_sv2v_reg ,\piso.data_r_187_sv2v_reg ,\piso.data_r_186_sv2v_reg ,
  \piso.data_r_185_sv2v_reg ,\piso.data_r_184_sv2v_reg ,\piso.data_r_183_sv2v_reg ,
  \piso.data_r_182_sv2v_reg ,\piso.data_r_181_sv2v_reg ,\piso.data_r_180_sv2v_reg ,
  \piso.data_r_179_sv2v_reg ,\piso.data_r_178_sv2v_reg ,\piso.data_r_177_sv2v_reg ,
  \piso.data_r_176_sv2v_reg ,\piso.data_r_175_sv2v_reg ,\piso.data_r_174_sv2v_reg ,
  \piso.data_r_173_sv2v_reg ,\piso.data_r_172_sv2v_reg ,\piso.data_r_171_sv2v_reg ,
  \piso.data_r_170_sv2v_reg ,\piso.data_r_169_sv2v_reg ,\piso.data_r_168_sv2v_reg ,
  \piso.data_r_167_sv2v_reg ,\piso.data_r_166_sv2v_reg ,\piso.data_r_165_sv2v_reg ,
  \piso.data_r_164_sv2v_reg ,\piso.data_r_163_sv2v_reg ,\piso.data_r_162_sv2v_reg ,
  \piso.data_r_161_sv2v_reg ,\piso.data_r_160_sv2v_reg ,\piso.data_r_159_sv2v_reg ,
  \piso.data_r_158_sv2v_reg ,\piso.data_r_157_sv2v_reg ,\piso.data_r_156_sv2v_reg ,
  \piso.data_r_155_sv2v_reg ,\piso.data_r_154_sv2v_reg ,\piso.data_r_153_sv2v_reg ,
  \piso.data_r_152_sv2v_reg ,\piso.data_r_151_sv2v_reg ,\piso.data_r_150_sv2v_reg ,
  \piso.data_r_149_sv2v_reg ,\piso.data_r_148_sv2v_reg ,\piso.data_r_147_sv2v_reg ,
  \piso.data_r_146_sv2v_reg ,\piso.data_r_145_sv2v_reg ,\piso.data_r_144_sv2v_reg ,
  \piso.data_r_143_sv2v_reg ,\piso.data_r_142_sv2v_reg ,\piso.data_r_141_sv2v_reg ,
  \piso.data_r_140_sv2v_reg ,\piso.data_r_139_sv2v_reg ,\piso.data_r_138_sv2v_reg ,
  \piso.data_r_137_sv2v_reg ,\piso.data_r_136_sv2v_reg ,\piso.data_r_135_sv2v_reg ,
  \piso.data_r_134_sv2v_reg ,\piso.data_r_133_sv2v_reg ,\piso.data_r_132_sv2v_reg ,
  \piso.data_r_131_sv2v_reg ,\piso.data_r_130_sv2v_reg ,\piso.data_r_129_sv2v_reg ,
  \piso.data_r_128_sv2v_reg ,\piso.data_r_127_sv2v_reg ,\piso.data_r_126_sv2v_reg ,
  \piso.data_r_125_sv2v_reg ,\piso.data_r_124_sv2v_reg ,\piso.data_r_123_sv2v_reg ,
  \piso.data_r_122_sv2v_reg ,\piso.data_r_121_sv2v_reg ,
  \piso.data_r_120_sv2v_reg ,\piso.data_r_119_sv2v_reg ,\piso.data_r_118_sv2v_reg ,
  \piso.data_r_117_sv2v_reg ,\piso.data_r_116_sv2v_reg ,\piso.data_r_115_sv2v_reg ,
  \piso.data_r_114_sv2v_reg ,\piso.data_r_113_sv2v_reg ,\piso.data_r_112_sv2v_reg ,
  \piso.data_r_111_sv2v_reg ,\piso.data_r_110_sv2v_reg ,\piso.data_r_109_sv2v_reg ,
  \piso.data_r_108_sv2v_reg ,\piso.data_r_107_sv2v_reg ,\piso.data_r_106_sv2v_reg ,
  \piso.data_r_105_sv2v_reg ,\piso.data_r_104_sv2v_reg ,\piso.data_r_103_sv2v_reg ,
  \piso.data_r_102_sv2v_reg ,\piso.data_r_101_sv2v_reg ,\piso.data_r_100_sv2v_reg ,
  \piso.data_r_99_sv2v_reg ,\piso.data_r_98_sv2v_reg ,\piso.data_r_97_sv2v_reg ,
  \piso.data_r_96_sv2v_reg ,\piso.data_r_95_sv2v_reg ,\piso.data_r_94_sv2v_reg ,
  \piso.data_r_93_sv2v_reg ,\piso.data_r_92_sv2v_reg ,\piso.data_r_91_sv2v_reg ,
  \piso.data_r_90_sv2v_reg ,\piso.data_r_89_sv2v_reg ,\piso.data_r_88_sv2v_reg ,\piso.data_r_87_sv2v_reg ,
  \piso.data_r_86_sv2v_reg ,\piso.data_r_85_sv2v_reg ,\piso.data_r_84_sv2v_reg ,
  \piso.data_r_83_sv2v_reg ,\piso.data_r_82_sv2v_reg ,\piso.data_r_81_sv2v_reg ,
  \piso.data_r_80_sv2v_reg ,\piso.data_r_79_sv2v_reg ,\piso.data_r_78_sv2v_reg ,
  \piso.data_r_77_sv2v_reg ,\piso.data_r_76_sv2v_reg ,\piso.data_r_75_sv2v_reg ,
  \piso.data_r_74_sv2v_reg ,\piso.data_r_73_sv2v_reg ,\piso.data_r_72_sv2v_reg ,
  \piso.data_r_71_sv2v_reg ,\piso.data_r_70_sv2v_reg ,\piso.data_r_69_sv2v_reg ,
  \piso.data_r_68_sv2v_reg ,\piso.data_r_67_sv2v_reg ,\piso.data_r_66_sv2v_reg ,
  \piso.data_r_65_sv2v_reg ,\piso.data_r_64_sv2v_reg ,\piso.data_r_63_sv2v_reg ,
  \piso.data_r_62_sv2v_reg ,\piso.data_r_61_sv2v_reg ,\piso.data_r_60_sv2v_reg ,
  \piso.data_r_59_sv2v_reg ,\piso.data_r_58_sv2v_reg ,\piso.data_r_57_sv2v_reg ,
  \piso.data_r_56_sv2v_reg ,\piso.data_r_55_sv2v_reg ,\piso.data_r_54_sv2v_reg ,
  \piso.data_r_53_sv2v_reg ,\piso.data_r_52_sv2v_reg ,\piso.data_r_51_sv2v_reg ,
  \piso.data_r_50_sv2v_reg ,\piso.data_r_49_sv2v_reg ,\piso.data_r_48_sv2v_reg ,\piso.data_r_47_sv2v_reg ,
  \piso.data_r_46_sv2v_reg ,\piso.data_r_45_sv2v_reg ,\piso.data_r_44_sv2v_reg ,
  \piso.data_r_43_sv2v_reg ,\piso.data_r_42_sv2v_reg ,\piso.data_r_41_sv2v_reg ,
  \piso.data_r_40_sv2v_reg ,\piso.data_r_39_sv2v_reg ,\piso.data_r_38_sv2v_reg ,
  \piso.data_r_37_sv2v_reg ,\piso.data_r_36_sv2v_reg ,\piso.data_r_35_sv2v_reg ,
  \piso.data_r_34_sv2v_reg ,\piso.data_r_33_sv2v_reg ,\piso.data_r_32_sv2v_reg ,
  \piso.data_r_31_sv2v_reg ,\piso.data_r_30_sv2v_reg ,\piso.data_r_29_sv2v_reg ,
  \piso.data_r_28_sv2v_reg ,\piso.data_r_27_sv2v_reg ,\piso.data_r_26_sv2v_reg ,
  \piso.data_r_25_sv2v_reg ,\piso.data_r_24_sv2v_reg ,\piso.data_r_23_sv2v_reg ,
  \piso.data_r_22_sv2v_reg ,\piso.data_r_21_sv2v_reg ,\piso.data_r_20_sv2v_reg ,
  \piso.data_r_19_sv2v_reg ,\piso.data_r_18_sv2v_reg ,\piso.data_r_17_sv2v_reg ,
  \piso.data_r_16_sv2v_reg ,\piso.data_r_15_sv2v_reg ,\piso.data_r_14_sv2v_reg ,
  \piso.data_r_13_sv2v_reg ,\piso.data_r_12_sv2v_reg ,\piso.data_r_11_sv2v_reg ,
  \piso.data_r_10_sv2v_reg ,\piso.data_r_9_sv2v_reg ,\piso.data_r_8_sv2v_reg ,\piso.data_r_7_sv2v_reg ,
  \piso.data_r_6_sv2v_reg ,\piso.data_r_5_sv2v_reg ,\piso.data_r_4_sv2v_reg ,
  \piso.data_r_3_sv2v_reg ,\piso.data_r_2_sv2v_reg ,\piso.data_r_1_sv2v_reg ,
  \piso.data_r_0_sv2v_reg ,\piso.shift_ctr_r_5_sv2v_reg ,\piso.shift_ctr_r_4_sv2v_reg ,
  \piso.shift_ctr_r_3_sv2v_reg ,\piso.shift_ctr_r_2_sv2v_reg ,
  \piso.shift_ctr_r_1_sv2v_reg ,\piso.shift_ctr_r_0_sv2v_reg ;
  assign valid_o = valid_o_sv2v_reg;
  assign \piso.data_r [2047] = \piso.data_r_2047_sv2v_reg ;
  assign \piso.data_r [2046] = \piso.data_r_2046_sv2v_reg ;
  assign \piso.data_r [2045] = \piso.data_r_2045_sv2v_reg ;
  assign \piso.data_r [2044] = \piso.data_r_2044_sv2v_reg ;
  assign \piso.data_r [2043] = \piso.data_r_2043_sv2v_reg ;
  assign \piso.data_r [2042] = \piso.data_r_2042_sv2v_reg ;
  assign \piso.data_r [2041] = \piso.data_r_2041_sv2v_reg ;
  assign \piso.data_r [2040] = \piso.data_r_2040_sv2v_reg ;
  assign \piso.data_r [2039] = \piso.data_r_2039_sv2v_reg ;
  assign \piso.data_r [2038] = \piso.data_r_2038_sv2v_reg ;
  assign \piso.data_r [2037] = \piso.data_r_2037_sv2v_reg ;
  assign \piso.data_r [2036] = \piso.data_r_2036_sv2v_reg ;
  assign \piso.data_r [2035] = \piso.data_r_2035_sv2v_reg ;
  assign \piso.data_r [2034] = \piso.data_r_2034_sv2v_reg ;
  assign \piso.data_r [2033] = \piso.data_r_2033_sv2v_reg ;
  assign \piso.data_r [2032] = \piso.data_r_2032_sv2v_reg ;
  assign \piso.data_r [2031] = \piso.data_r_2031_sv2v_reg ;
  assign \piso.data_r [2030] = \piso.data_r_2030_sv2v_reg ;
  assign \piso.data_r [2029] = \piso.data_r_2029_sv2v_reg ;
  assign \piso.data_r [2028] = \piso.data_r_2028_sv2v_reg ;
  assign \piso.data_r [2027] = \piso.data_r_2027_sv2v_reg ;
  assign \piso.data_r [2026] = \piso.data_r_2026_sv2v_reg ;
  assign \piso.data_r [2025] = \piso.data_r_2025_sv2v_reg ;
  assign \piso.data_r [2024] = \piso.data_r_2024_sv2v_reg ;
  assign \piso.data_r [2023] = \piso.data_r_2023_sv2v_reg ;
  assign \piso.data_r [2022] = \piso.data_r_2022_sv2v_reg ;
  assign \piso.data_r [2021] = \piso.data_r_2021_sv2v_reg ;
  assign \piso.data_r [2020] = \piso.data_r_2020_sv2v_reg ;
  assign \piso.data_r [2019] = \piso.data_r_2019_sv2v_reg ;
  assign \piso.data_r [2018] = \piso.data_r_2018_sv2v_reg ;
  assign \piso.data_r [2017] = \piso.data_r_2017_sv2v_reg ;
  assign \piso.data_r [2016] = \piso.data_r_2016_sv2v_reg ;
  assign \piso.data_r [2015] = \piso.data_r_2015_sv2v_reg ;
  assign \piso.data_r [2014] = \piso.data_r_2014_sv2v_reg ;
  assign \piso.data_r [2013] = \piso.data_r_2013_sv2v_reg ;
  assign \piso.data_r [2012] = \piso.data_r_2012_sv2v_reg ;
  assign \piso.data_r [2011] = \piso.data_r_2011_sv2v_reg ;
  assign \piso.data_r [2010] = \piso.data_r_2010_sv2v_reg ;
  assign \piso.data_r [2009] = \piso.data_r_2009_sv2v_reg ;
  assign \piso.data_r [2008] = \piso.data_r_2008_sv2v_reg ;
  assign \piso.data_r [2007] = \piso.data_r_2007_sv2v_reg ;
  assign \piso.data_r [2006] = \piso.data_r_2006_sv2v_reg ;
  assign \piso.data_r [2005] = \piso.data_r_2005_sv2v_reg ;
  assign \piso.data_r [2004] = \piso.data_r_2004_sv2v_reg ;
  assign \piso.data_r [2003] = \piso.data_r_2003_sv2v_reg ;
  assign \piso.data_r [2002] = \piso.data_r_2002_sv2v_reg ;
  assign \piso.data_r [2001] = \piso.data_r_2001_sv2v_reg ;
  assign \piso.data_r [2000] = \piso.data_r_2000_sv2v_reg ;
  assign \piso.data_r [1999] = \piso.data_r_1999_sv2v_reg ;
  assign \piso.data_r [1998] = \piso.data_r_1998_sv2v_reg ;
  assign \piso.data_r [1997] = \piso.data_r_1997_sv2v_reg ;
  assign \piso.data_r [1996] = \piso.data_r_1996_sv2v_reg ;
  assign \piso.data_r [1995] = \piso.data_r_1995_sv2v_reg ;
  assign \piso.data_r [1994] = \piso.data_r_1994_sv2v_reg ;
  assign \piso.data_r [1993] = \piso.data_r_1993_sv2v_reg ;
  assign \piso.data_r [1992] = \piso.data_r_1992_sv2v_reg ;
  assign \piso.data_r [1991] = \piso.data_r_1991_sv2v_reg ;
  assign \piso.data_r [1990] = \piso.data_r_1990_sv2v_reg ;
  assign \piso.data_r [1989] = \piso.data_r_1989_sv2v_reg ;
  assign \piso.data_r [1988] = \piso.data_r_1988_sv2v_reg ;
  assign \piso.data_r [1987] = \piso.data_r_1987_sv2v_reg ;
  assign \piso.data_r [1986] = \piso.data_r_1986_sv2v_reg ;
  assign \piso.data_r [1985] = \piso.data_r_1985_sv2v_reg ;
  assign \piso.data_r [1984] = \piso.data_r_1984_sv2v_reg ;
  assign \piso.data_r [1983] = \piso.data_r_1983_sv2v_reg ;
  assign \piso.data_r [1982] = \piso.data_r_1982_sv2v_reg ;
  assign \piso.data_r [1981] = \piso.data_r_1981_sv2v_reg ;
  assign \piso.data_r [1980] = \piso.data_r_1980_sv2v_reg ;
  assign \piso.data_r [1979] = \piso.data_r_1979_sv2v_reg ;
  assign \piso.data_r [1978] = \piso.data_r_1978_sv2v_reg ;
  assign \piso.data_r [1977] = \piso.data_r_1977_sv2v_reg ;
  assign \piso.data_r [1976] = \piso.data_r_1976_sv2v_reg ;
  assign \piso.data_r [1975] = \piso.data_r_1975_sv2v_reg ;
  assign \piso.data_r [1974] = \piso.data_r_1974_sv2v_reg ;
  assign \piso.data_r [1973] = \piso.data_r_1973_sv2v_reg ;
  assign \piso.data_r [1972] = \piso.data_r_1972_sv2v_reg ;
  assign \piso.data_r [1971] = \piso.data_r_1971_sv2v_reg ;
  assign \piso.data_r [1970] = \piso.data_r_1970_sv2v_reg ;
  assign \piso.data_r [1969] = \piso.data_r_1969_sv2v_reg ;
  assign \piso.data_r [1968] = \piso.data_r_1968_sv2v_reg ;
  assign \piso.data_r [1967] = \piso.data_r_1967_sv2v_reg ;
  assign \piso.data_r [1966] = \piso.data_r_1966_sv2v_reg ;
  assign \piso.data_r [1965] = \piso.data_r_1965_sv2v_reg ;
  assign \piso.data_r [1964] = \piso.data_r_1964_sv2v_reg ;
  assign \piso.data_r [1963] = \piso.data_r_1963_sv2v_reg ;
  assign \piso.data_r [1962] = \piso.data_r_1962_sv2v_reg ;
  assign \piso.data_r [1961] = \piso.data_r_1961_sv2v_reg ;
  assign \piso.data_r [1960] = \piso.data_r_1960_sv2v_reg ;
  assign \piso.data_r [1959] = \piso.data_r_1959_sv2v_reg ;
  assign \piso.data_r [1958] = \piso.data_r_1958_sv2v_reg ;
  assign \piso.data_r [1957] = \piso.data_r_1957_sv2v_reg ;
  assign \piso.data_r [1956] = \piso.data_r_1956_sv2v_reg ;
  assign \piso.data_r [1955] = \piso.data_r_1955_sv2v_reg ;
  assign \piso.data_r [1954] = \piso.data_r_1954_sv2v_reg ;
  assign \piso.data_r [1953] = \piso.data_r_1953_sv2v_reg ;
  assign \piso.data_r [1952] = \piso.data_r_1952_sv2v_reg ;
  assign \piso.data_r [1951] = \piso.data_r_1951_sv2v_reg ;
  assign \piso.data_r [1950] = \piso.data_r_1950_sv2v_reg ;
  assign \piso.data_r [1949] = \piso.data_r_1949_sv2v_reg ;
  assign \piso.data_r [1948] = \piso.data_r_1948_sv2v_reg ;
  assign \piso.data_r [1947] = \piso.data_r_1947_sv2v_reg ;
  assign \piso.data_r [1946] = \piso.data_r_1946_sv2v_reg ;
  assign \piso.data_r [1945] = \piso.data_r_1945_sv2v_reg ;
  assign \piso.data_r [1944] = \piso.data_r_1944_sv2v_reg ;
  assign \piso.data_r [1943] = \piso.data_r_1943_sv2v_reg ;
  assign \piso.data_r [1942] = \piso.data_r_1942_sv2v_reg ;
  assign \piso.data_r [1941] = \piso.data_r_1941_sv2v_reg ;
  assign \piso.data_r [1940] = \piso.data_r_1940_sv2v_reg ;
  assign \piso.data_r [1939] = \piso.data_r_1939_sv2v_reg ;
  assign \piso.data_r [1938] = \piso.data_r_1938_sv2v_reg ;
  assign \piso.data_r [1937] = \piso.data_r_1937_sv2v_reg ;
  assign \piso.data_r [1936] = \piso.data_r_1936_sv2v_reg ;
  assign \piso.data_r [1935] = \piso.data_r_1935_sv2v_reg ;
  assign \piso.data_r [1934] = \piso.data_r_1934_sv2v_reg ;
  assign \piso.data_r [1933] = \piso.data_r_1933_sv2v_reg ;
  assign \piso.data_r [1932] = \piso.data_r_1932_sv2v_reg ;
  assign \piso.data_r [1931] = \piso.data_r_1931_sv2v_reg ;
  assign \piso.data_r [1930] = \piso.data_r_1930_sv2v_reg ;
  assign \piso.data_r [1929] = \piso.data_r_1929_sv2v_reg ;
  assign \piso.data_r [1928] = \piso.data_r_1928_sv2v_reg ;
  assign \piso.data_r [1927] = \piso.data_r_1927_sv2v_reg ;
  assign \piso.data_r [1926] = \piso.data_r_1926_sv2v_reg ;
  assign \piso.data_r [1925] = \piso.data_r_1925_sv2v_reg ;
  assign \piso.data_r [1924] = \piso.data_r_1924_sv2v_reg ;
  assign \piso.data_r [1923] = \piso.data_r_1923_sv2v_reg ;
  assign \piso.data_r [1922] = \piso.data_r_1922_sv2v_reg ;
  assign \piso.data_r [1921] = \piso.data_r_1921_sv2v_reg ;
  assign \piso.data_r [1920] = \piso.data_r_1920_sv2v_reg ;
  assign \piso.data_r [1919] = \piso.data_r_1919_sv2v_reg ;
  assign \piso.data_r [1918] = \piso.data_r_1918_sv2v_reg ;
  assign \piso.data_r [1917] = \piso.data_r_1917_sv2v_reg ;
  assign \piso.data_r [1916] = \piso.data_r_1916_sv2v_reg ;
  assign \piso.data_r [1915] = \piso.data_r_1915_sv2v_reg ;
  assign \piso.data_r [1914] = \piso.data_r_1914_sv2v_reg ;
  assign \piso.data_r [1913] = \piso.data_r_1913_sv2v_reg ;
  assign \piso.data_r [1912] = \piso.data_r_1912_sv2v_reg ;
  assign \piso.data_r [1911] = \piso.data_r_1911_sv2v_reg ;
  assign \piso.data_r [1910] = \piso.data_r_1910_sv2v_reg ;
  assign \piso.data_r [1909] = \piso.data_r_1909_sv2v_reg ;
  assign \piso.data_r [1908] = \piso.data_r_1908_sv2v_reg ;
  assign \piso.data_r [1907] = \piso.data_r_1907_sv2v_reg ;
  assign \piso.data_r [1906] = \piso.data_r_1906_sv2v_reg ;
  assign \piso.data_r [1905] = \piso.data_r_1905_sv2v_reg ;
  assign \piso.data_r [1904] = \piso.data_r_1904_sv2v_reg ;
  assign \piso.data_r [1903] = \piso.data_r_1903_sv2v_reg ;
  assign \piso.data_r [1902] = \piso.data_r_1902_sv2v_reg ;
  assign \piso.data_r [1901] = \piso.data_r_1901_sv2v_reg ;
  assign \piso.data_r [1900] = \piso.data_r_1900_sv2v_reg ;
  assign \piso.data_r [1899] = \piso.data_r_1899_sv2v_reg ;
  assign \piso.data_r [1898] = \piso.data_r_1898_sv2v_reg ;
  assign \piso.data_r [1897] = \piso.data_r_1897_sv2v_reg ;
  assign \piso.data_r [1896] = \piso.data_r_1896_sv2v_reg ;
  assign \piso.data_r [1895] = \piso.data_r_1895_sv2v_reg ;
  assign \piso.data_r [1894] = \piso.data_r_1894_sv2v_reg ;
  assign \piso.data_r [1893] = \piso.data_r_1893_sv2v_reg ;
  assign \piso.data_r [1892] = \piso.data_r_1892_sv2v_reg ;
  assign \piso.data_r [1891] = \piso.data_r_1891_sv2v_reg ;
  assign \piso.data_r [1890] = \piso.data_r_1890_sv2v_reg ;
  assign \piso.data_r [1889] = \piso.data_r_1889_sv2v_reg ;
  assign \piso.data_r [1888] = \piso.data_r_1888_sv2v_reg ;
  assign \piso.data_r [1887] = \piso.data_r_1887_sv2v_reg ;
  assign \piso.data_r [1886] = \piso.data_r_1886_sv2v_reg ;
  assign \piso.data_r [1885] = \piso.data_r_1885_sv2v_reg ;
  assign \piso.data_r [1884] = \piso.data_r_1884_sv2v_reg ;
  assign \piso.data_r [1883] = \piso.data_r_1883_sv2v_reg ;
  assign \piso.data_r [1882] = \piso.data_r_1882_sv2v_reg ;
  assign \piso.data_r [1881] = \piso.data_r_1881_sv2v_reg ;
  assign \piso.data_r [1880] = \piso.data_r_1880_sv2v_reg ;
  assign \piso.data_r [1879] = \piso.data_r_1879_sv2v_reg ;
  assign \piso.data_r [1878] = \piso.data_r_1878_sv2v_reg ;
  assign \piso.data_r [1877] = \piso.data_r_1877_sv2v_reg ;
  assign \piso.data_r [1876] = \piso.data_r_1876_sv2v_reg ;
  assign \piso.data_r [1875] = \piso.data_r_1875_sv2v_reg ;
  assign \piso.data_r [1874] = \piso.data_r_1874_sv2v_reg ;
  assign \piso.data_r [1873] = \piso.data_r_1873_sv2v_reg ;
  assign \piso.data_r [1872] = \piso.data_r_1872_sv2v_reg ;
  assign \piso.data_r [1871] = \piso.data_r_1871_sv2v_reg ;
  assign \piso.data_r [1870] = \piso.data_r_1870_sv2v_reg ;
  assign \piso.data_r [1869] = \piso.data_r_1869_sv2v_reg ;
  assign \piso.data_r [1868] = \piso.data_r_1868_sv2v_reg ;
  assign \piso.data_r [1867] = \piso.data_r_1867_sv2v_reg ;
  assign \piso.data_r [1866] = \piso.data_r_1866_sv2v_reg ;
  assign \piso.data_r [1865] = \piso.data_r_1865_sv2v_reg ;
  assign \piso.data_r [1864] = \piso.data_r_1864_sv2v_reg ;
  assign \piso.data_r [1863] = \piso.data_r_1863_sv2v_reg ;
  assign \piso.data_r [1862] = \piso.data_r_1862_sv2v_reg ;
  assign \piso.data_r [1861] = \piso.data_r_1861_sv2v_reg ;
  assign \piso.data_r [1860] = \piso.data_r_1860_sv2v_reg ;
  assign \piso.data_r [1859] = \piso.data_r_1859_sv2v_reg ;
  assign \piso.data_r [1858] = \piso.data_r_1858_sv2v_reg ;
  assign \piso.data_r [1857] = \piso.data_r_1857_sv2v_reg ;
  assign \piso.data_r [1856] = \piso.data_r_1856_sv2v_reg ;
  assign \piso.data_r [1855] = \piso.data_r_1855_sv2v_reg ;
  assign \piso.data_r [1854] = \piso.data_r_1854_sv2v_reg ;
  assign \piso.data_r [1853] = \piso.data_r_1853_sv2v_reg ;
  assign \piso.data_r [1852] = \piso.data_r_1852_sv2v_reg ;
  assign \piso.data_r [1851] = \piso.data_r_1851_sv2v_reg ;
  assign \piso.data_r [1850] = \piso.data_r_1850_sv2v_reg ;
  assign \piso.data_r [1849] = \piso.data_r_1849_sv2v_reg ;
  assign \piso.data_r [1848] = \piso.data_r_1848_sv2v_reg ;
  assign \piso.data_r [1847] = \piso.data_r_1847_sv2v_reg ;
  assign \piso.data_r [1846] = \piso.data_r_1846_sv2v_reg ;
  assign \piso.data_r [1845] = \piso.data_r_1845_sv2v_reg ;
  assign \piso.data_r [1844] = \piso.data_r_1844_sv2v_reg ;
  assign \piso.data_r [1843] = \piso.data_r_1843_sv2v_reg ;
  assign \piso.data_r [1842] = \piso.data_r_1842_sv2v_reg ;
  assign \piso.data_r [1841] = \piso.data_r_1841_sv2v_reg ;
  assign \piso.data_r [1840] = \piso.data_r_1840_sv2v_reg ;
  assign \piso.data_r [1839] = \piso.data_r_1839_sv2v_reg ;
  assign \piso.data_r [1838] = \piso.data_r_1838_sv2v_reg ;
  assign \piso.data_r [1837] = \piso.data_r_1837_sv2v_reg ;
  assign \piso.data_r [1836] = \piso.data_r_1836_sv2v_reg ;
  assign \piso.data_r [1835] = \piso.data_r_1835_sv2v_reg ;
  assign \piso.data_r [1834] = \piso.data_r_1834_sv2v_reg ;
  assign \piso.data_r [1833] = \piso.data_r_1833_sv2v_reg ;
  assign \piso.data_r [1832] = \piso.data_r_1832_sv2v_reg ;
  assign \piso.data_r [1831] = \piso.data_r_1831_sv2v_reg ;
  assign \piso.data_r [1830] = \piso.data_r_1830_sv2v_reg ;
  assign \piso.data_r [1829] = \piso.data_r_1829_sv2v_reg ;
  assign \piso.data_r [1828] = \piso.data_r_1828_sv2v_reg ;
  assign \piso.data_r [1827] = \piso.data_r_1827_sv2v_reg ;
  assign \piso.data_r [1826] = \piso.data_r_1826_sv2v_reg ;
  assign \piso.data_r [1825] = \piso.data_r_1825_sv2v_reg ;
  assign \piso.data_r [1824] = \piso.data_r_1824_sv2v_reg ;
  assign \piso.data_r [1823] = \piso.data_r_1823_sv2v_reg ;
  assign \piso.data_r [1822] = \piso.data_r_1822_sv2v_reg ;
  assign \piso.data_r [1821] = \piso.data_r_1821_sv2v_reg ;
  assign \piso.data_r [1820] = \piso.data_r_1820_sv2v_reg ;
  assign \piso.data_r [1819] = \piso.data_r_1819_sv2v_reg ;
  assign \piso.data_r [1818] = \piso.data_r_1818_sv2v_reg ;
  assign \piso.data_r [1817] = \piso.data_r_1817_sv2v_reg ;
  assign \piso.data_r [1816] = \piso.data_r_1816_sv2v_reg ;
  assign \piso.data_r [1815] = \piso.data_r_1815_sv2v_reg ;
  assign \piso.data_r [1814] = \piso.data_r_1814_sv2v_reg ;
  assign \piso.data_r [1813] = \piso.data_r_1813_sv2v_reg ;
  assign \piso.data_r [1812] = \piso.data_r_1812_sv2v_reg ;
  assign \piso.data_r [1811] = \piso.data_r_1811_sv2v_reg ;
  assign \piso.data_r [1810] = \piso.data_r_1810_sv2v_reg ;
  assign \piso.data_r [1809] = \piso.data_r_1809_sv2v_reg ;
  assign \piso.data_r [1808] = \piso.data_r_1808_sv2v_reg ;
  assign \piso.data_r [1807] = \piso.data_r_1807_sv2v_reg ;
  assign \piso.data_r [1806] = \piso.data_r_1806_sv2v_reg ;
  assign \piso.data_r [1805] = \piso.data_r_1805_sv2v_reg ;
  assign \piso.data_r [1804] = \piso.data_r_1804_sv2v_reg ;
  assign \piso.data_r [1803] = \piso.data_r_1803_sv2v_reg ;
  assign \piso.data_r [1802] = \piso.data_r_1802_sv2v_reg ;
  assign \piso.data_r [1801] = \piso.data_r_1801_sv2v_reg ;
  assign \piso.data_r [1800] = \piso.data_r_1800_sv2v_reg ;
  assign \piso.data_r [1799] = \piso.data_r_1799_sv2v_reg ;
  assign \piso.data_r [1798] = \piso.data_r_1798_sv2v_reg ;
  assign \piso.data_r [1797] = \piso.data_r_1797_sv2v_reg ;
  assign \piso.data_r [1796] = \piso.data_r_1796_sv2v_reg ;
  assign \piso.data_r [1795] = \piso.data_r_1795_sv2v_reg ;
  assign \piso.data_r [1794] = \piso.data_r_1794_sv2v_reg ;
  assign \piso.data_r [1793] = \piso.data_r_1793_sv2v_reg ;
  assign \piso.data_r [1792] = \piso.data_r_1792_sv2v_reg ;
  assign \piso.data_r [1791] = \piso.data_r_1791_sv2v_reg ;
  assign \piso.data_r [1790] = \piso.data_r_1790_sv2v_reg ;
  assign \piso.data_r [1789] = \piso.data_r_1789_sv2v_reg ;
  assign \piso.data_r [1788] = \piso.data_r_1788_sv2v_reg ;
  assign \piso.data_r [1787] = \piso.data_r_1787_sv2v_reg ;
  assign \piso.data_r [1786] = \piso.data_r_1786_sv2v_reg ;
  assign \piso.data_r [1785] = \piso.data_r_1785_sv2v_reg ;
  assign \piso.data_r [1784] = \piso.data_r_1784_sv2v_reg ;
  assign \piso.data_r [1783] = \piso.data_r_1783_sv2v_reg ;
  assign \piso.data_r [1782] = \piso.data_r_1782_sv2v_reg ;
  assign \piso.data_r [1781] = \piso.data_r_1781_sv2v_reg ;
  assign \piso.data_r [1780] = \piso.data_r_1780_sv2v_reg ;
  assign \piso.data_r [1779] = \piso.data_r_1779_sv2v_reg ;
  assign \piso.data_r [1778] = \piso.data_r_1778_sv2v_reg ;
  assign \piso.data_r [1777] = \piso.data_r_1777_sv2v_reg ;
  assign \piso.data_r [1776] = \piso.data_r_1776_sv2v_reg ;
  assign \piso.data_r [1775] = \piso.data_r_1775_sv2v_reg ;
  assign \piso.data_r [1774] = \piso.data_r_1774_sv2v_reg ;
  assign \piso.data_r [1773] = \piso.data_r_1773_sv2v_reg ;
  assign \piso.data_r [1772] = \piso.data_r_1772_sv2v_reg ;
  assign \piso.data_r [1771] = \piso.data_r_1771_sv2v_reg ;
  assign \piso.data_r [1770] = \piso.data_r_1770_sv2v_reg ;
  assign \piso.data_r [1769] = \piso.data_r_1769_sv2v_reg ;
  assign \piso.data_r [1768] = \piso.data_r_1768_sv2v_reg ;
  assign \piso.data_r [1767] = \piso.data_r_1767_sv2v_reg ;
  assign \piso.data_r [1766] = \piso.data_r_1766_sv2v_reg ;
  assign \piso.data_r [1765] = \piso.data_r_1765_sv2v_reg ;
  assign \piso.data_r [1764] = \piso.data_r_1764_sv2v_reg ;
  assign \piso.data_r [1763] = \piso.data_r_1763_sv2v_reg ;
  assign \piso.data_r [1762] = \piso.data_r_1762_sv2v_reg ;
  assign \piso.data_r [1761] = \piso.data_r_1761_sv2v_reg ;
  assign \piso.data_r [1760] = \piso.data_r_1760_sv2v_reg ;
  assign \piso.data_r [1759] = \piso.data_r_1759_sv2v_reg ;
  assign \piso.data_r [1758] = \piso.data_r_1758_sv2v_reg ;
  assign \piso.data_r [1757] = \piso.data_r_1757_sv2v_reg ;
  assign \piso.data_r [1756] = \piso.data_r_1756_sv2v_reg ;
  assign \piso.data_r [1755] = \piso.data_r_1755_sv2v_reg ;
  assign \piso.data_r [1754] = \piso.data_r_1754_sv2v_reg ;
  assign \piso.data_r [1753] = \piso.data_r_1753_sv2v_reg ;
  assign \piso.data_r [1752] = \piso.data_r_1752_sv2v_reg ;
  assign \piso.data_r [1751] = \piso.data_r_1751_sv2v_reg ;
  assign \piso.data_r [1750] = \piso.data_r_1750_sv2v_reg ;
  assign \piso.data_r [1749] = \piso.data_r_1749_sv2v_reg ;
  assign \piso.data_r [1748] = \piso.data_r_1748_sv2v_reg ;
  assign \piso.data_r [1747] = \piso.data_r_1747_sv2v_reg ;
  assign \piso.data_r [1746] = \piso.data_r_1746_sv2v_reg ;
  assign \piso.data_r [1745] = \piso.data_r_1745_sv2v_reg ;
  assign \piso.data_r [1744] = \piso.data_r_1744_sv2v_reg ;
  assign \piso.data_r [1743] = \piso.data_r_1743_sv2v_reg ;
  assign \piso.data_r [1742] = \piso.data_r_1742_sv2v_reg ;
  assign \piso.data_r [1741] = \piso.data_r_1741_sv2v_reg ;
  assign \piso.data_r [1740] = \piso.data_r_1740_sv2v_reg ;
  assign \piso.data_r [1739] = \piso.data_r_1739_sv2v_reg ;
  assign \piso.data_r [1738] = \piso.data_r_1738_sv2v_reg ;
  assign \piso.data_r [1737] = \piso.data_r_1737_sv2v_reg ;
  assign \piso.data_r [1736] = \piso.data_r_1736_sv2v_reg ;
  assign \piso.data_r [1735] = \piso.data_r_1735_sv2v_reg ;
  assign \piso.data_r [1734] = \piso.data_r_1734_sv2v_reg ;
  assign \piso.data_r [1733] = \piso.data_r_1733_sv2v_reg ;
  assign \piso.data_r [1732] = \piso.data_r_1732_sv2v_reg ;
  assign \piso.data_r [1731] = \piso.data_r_1731_sv2v_reg ;
  assign \piso.data_r [1730] = \piso.data_r_1730_sv2v_reg ;
  assign \piso.data_r [1729] = \piso.data_r_1729_sv2v_reg ;
  assign \piso.data_r [1728] = \piso.data_r_1728_sv2v_reg ;
  assign \piso.data_r [1727] = \piso.data_r_1727_sv2v_reg ;
  assign \piso.data_r [1726] = \piso.data_r_1726_sv2v_reg ;
  assign \piso.data_r [1725] = \piso.data_r_1725_sv2v_reg ;
  assign \piso.data_r [1724] = \piso.data_r_1724_sv2v_reg ;
  assign \piso.data_r [1723] = \piso.data_r_1723_sv2v_reg ;
  assign \piso.data_r [1722] = \piso.data_r_1722_sv2v_reg ;
  assign \piso.data_r [1721] = \piso.data_r_1721_sv2v_reg ;
  assign \piso.data_r [1720] = \piso.data_r_1720_sv2v_reg ;
  assign \piso.data_r [1719] = \piso.data_r_1719_sv2v_reg ;
  assign \piso.data_r [1718] = \piso.data_r_1718_sv2v_reg ;
  assign \piso.data_r [1717] = \piso.data_r_1717_sv2v_reg ;
  assign \piso.data_r [1716] = \piso.data_r_1716_sv2v_reg ;
  assign \piso.data_r [1715] = \piso.data_r_1715_sv2v_reg ;
  assign \piso.data_r [1714] = \piso.data_r_1714_sv2v_reg ;
  assign \piso.data_r [1713] = \piso.data_r_1713_sv2v_reg ;
  assign \piso.data_r [1712] = \piso.data_r_1712_sv2v_reg ;
  assign \piso.data_r [1711] = \piso.data_r_1711_sv2v_reg ;
  assign \piso.data_r [1710] = \piso.data_r_1710_sv2v_reg ;
  assign \piso.data_r [1709] = \piso.data_r_1709_sv2v_reg ;
  assign \piso.data_r [1708] = \piso.data_r_1708_sv2v_reg ;
  assign \piso.data_r [1707] = \piso.data_r_1707_sv2v_reg ;
  assign \piso.data_r [1706] = \piso.data_r_1706_sv2v_reg ;
  assign \piso.data_r [1705] = \piso.data_r_1705_sv2v_reg ;
  assign \piso.data_r [1704] = \piso.data_r_1704_sv2v_reg ;
  assign \piso.data_r [1703] = \piso.data_r_1703_sv2v_reg ;
  assign \piso.data_r [1702] = \piso.data_r_1702_sv2v_reg ;
  assign \piso.data_r [1701] = \piso.data_r_1701_sv2v_reg ;
  assign \piso.data_r [1700] = \piso.data_r_1700_sv2v_reg ;
  assign \piso.data_r [1699] = \piso.data_r_1699_sv2v_reg ;
  assign \piso.data_r [1698] = \piso.data_r_1698_sv2v_reg ;
  assign \piso.data_r [1697] = \piso.data_r_1697_sv2v_reg ;
  assign \piso.data_r [1696] = \piso.data_r_1696_sv2v_reg ;
  assign \piso.data_r [1695] = \piso.data_r_1695_sv2v_reg ;
  assign \piso.data_r [1694] = \piso.data_r_1694_sv2v_reg ;
  assign \piso.data_r [1693] = \piso.data_r_1693_sv2v_reg ;
  assign \piso.data_r [1692] = \piso.data_r_1692_sv2v_reg ;
  assign \piso.data_r [1691] = \piso.data_r_1691_sv2v_reg ;
  assign \piso.data_r [1690] = \piso.data_r_1690_sv2v_reg ;
  assign \piso.data_r [1689] = \piso.data_r_1689_sv2v_reg ;
  assign \piso.data_r [1688] = \piso.data_r_1688_sv2v_reg ;
  assign \piso.data_r [1687] = \piso.data_r_1687_sv2v_reg ;
  assign \piso.data_r [1686] = \piso.data_r_1686_sv2v_reg ;
  assign \piso.data_r [1685] = \piso.data_r_1685_sv2v_reg ;
  assign \piso.data_r [1684] = \piso.data_r_1684_sv2v_reg ;
  assign \piso.data_r [1683] = \piso.data_r_1683_sv2v_reg ;
  assign \piso.data_r [1682] = \piso.data_r_1682_sv2v_reg ;
  assign \piso.data_r [1681] = \piso.data_r_1681_sv2v_reg ;
  assign \piso.data_r [1680] = \piso.data_r_1680_sv2v_reg ;
  assign \piso.data_r [1679] = \piso.data_r_1679_sv2v_reg ;
  assign \piso.data_r [1678] = \piso.data_r_1678_sv2v_reg ;
  assign \piso.data_r [1677] = \piso.data_r_1677_sv2v_reg ;
  assign \piso.data_r [1676] = \piso.data_r_1676_sv2v_reg ;
  assign \piso.data_r [1675] = \piso.data_r_1675_sv2v_reg ;
  assign \piso.data_r [1674] = \piso.data_r_1674_sv2v_reg ;
  assign \piso.data_r [1673] = \piso.data_r_1673_sv2v_reg ;
  assign \piso.data_r [1672] = \piso.data_r_1672_sv2v_reg ;
  assign \piso.data_r [1671] = \piso.data_r_1671_sv2v_reg ;
  assign \piso.data_r [1670] = \piso.data_r_1670_sv2v_reg ;
  assign \piso.data_r [1669] = \piso.data_r_1669_sv2v_reg ;
  assign \piso.data_r [1668] = \piso.data_r_1668_sv2v_reg ;
  assign \piso.data_r [1667] = \piso.data_r_1667_sv2v_reg ;
  assign \piso.data_r [1666] = \piso.data_r_1666_sv2v_reg ;
  assign \piso.data_r [1665] = \piso.data_r_1665_sv2v_reg ;
  assign \piso.data_r [1664] = \piso.data_r_1664_sv2v_reg ;
  assign \piso.data_r [1663] = \piso.data_r_1663_sv2v_reg ;
  assign \piso.data_r [1662] = \piso.data_r_1662_sv2v_reg ;
  assign \piso.data_r [1661] = \piso.data_r_1661_sv2v_reg ;
  assign \piso.data_r [1660] = \piso.data_r_1660_sv2v_reg ;
  assign \piso.data_r [1659] = \piso.data_r_1659_sv2v_reg ;
  assign \piso.data_r [1658] = \piso.data_r_1658_sv2v_reg ;
  assign \piso.data_r [1657] = \piso.data_r_1657_sv2v_reg ;
  assign \piso.data_r [1656] = \piso.data_r_1656_sv2v_reg ;
  assign \piso.data_r [1655] = \piso.data_r_1655_sv2v_reg ;
  assign \piso.data_r [1654] = \piso.data_r_1654_sv2v_reg ;
  assign \piso.data_r [1653] = \piso.data_r_1653_sv2v_reg ;
  assign \piso.data_r [1652] = \piso.data_r_1652_sv2v_reg ;
  assign \piso.data_r [1651] = \piso.data_r_1651_sv2v_reg ;
  assign \piso.data_r [1650] = \piso.data_r_1650_sv2v_reg ;
  assign \piso.data_r [1649] = \piso.data_r_1649_sv2v_reg ;
  assign \piso.data_r [1648] = \piso.data_r_1648_sv2v_reg ;
  assign \piso.data_r [1647] = \piso.data_r_1647_sv2v_reg ;
  assign \piso.data_r [1646] = \piso.data_r_1646_sv2v_reg ;
  assign \piso.data_r [1645] = \piso.data_r_1645_sv2v_reg ;
  assign \piso.data_r [1644] = \piso.data_r_1644_sv2v_reg ;
  assign \piso.data_r [1643] = \piso.data_r_1643_sv2v_reg ;
  assign \piso.data_r [1642] = \piso.data_r_1642_sv2v_reg ;
  assign \piso.data_r [1641] = \piso.data_r_1641_sv2v_reg ;
  assign \piso.data_r [1640] = \piso.data_r_1640_sv2v_reg ;
  assign \piso.data_r [1639] = \piso.data_r_1639_sv2v_reg ;
  assign \piso.data_r [1638] = \piso.data_r_1638_sv2v_reg ;
  assign \piso.data_r [1637] = \piso.data_r_1637_sv2v_reg ;
  assign \piso.data_r [1636] = \piso.data_r_1636_sv2v_reg ;
  assign \piso.data_r [1635] = \piso.data_r_1635_sv2v_reg ;
  assign \piso.data_r [1634] = \piso.data_r_1634_sv2v_reg ;
  assign \piso.data_r [1633] = \piso.data_r_1633_sv2v_reg ;
  assign \piso.data_r [1632] = \piso.data_r_1632_sv2v_reg ;
  assign \piso.data_r [1631] = \piso.data_r_1631_sv2v_reg ;
  assign \piso.data_r [1630] = \piso.data_r_1630_sv2v_reg ;
  assign \piso.data_r [1629] = \piso.data_r_1629_sv2v_reg ;
  assign \piso.data_r [1628] = \piso.data_r_1628_sv2v_reg ;
  assign \piso.data_r [1627] = \piso.data_r_1627_sv2v_reg ;
  assign \piso.data_r [1626] = \piso.data_r_1626_sv2v_reg ;
  assign \piso.data_r [1625] = \piso.data_r_1625_sv2v_reg ;
  assign \piso.data_r [1624] = \piso.data_r_1624_sv2v_reg ;
  assign \piso.data_r [1623] = \piso.data_r_1623_sv2v_reg ;
  assign \piso.data_r [1622] = \piso.data_r_1622_sv2v_reg ;
  assign \piso.data_r [1621] = \piso.data_r_1621_sv2v_reg ;
  assign \piso.data_r [1620] = \piso.data_r_1620_sv2v_reg ;
  assign \piso.data_r [1619] = \piso.data_r_1619_sv2v_reg ;
  assign \piso.data_r [1618] = \piso.data_r_1618_sv2v_reg ;
  assign \piso.data_r [1617] = \piso.data_r_1617_sv2v_reg ;
  assign \piso.data_r [1616] = \piso.data_r_1616_sv2v_reg ;
  assign \piso.data_r [1615] = \piso.data_r_1615_sv2v_reg ;
  assign \piso.data_r [1614] = \piso.data_r_1614_sv2v_reg ;
  assign \piso.data_r [1613] = \piso.data_r_1613_sv2v_reg ;
  assign \piso.data_r [1612] = \piso.data_r_1612_sv2v_reg ;
  assign \piso.data_r [1611] = \piso.data_r_1611_sv2v_reg ;
  assign \piso.data_r [1610] = \piso.data_r_1610_sv2v_reg ;
  assign \piso.data_r [1609] = \piso.data_r_1609_sv2v_reg ;
  assign \piso.data_r [1608] = \piso.data_r_1608_sv2v_reg ;
  assign \piso.data_r [1607] = \piso.data_r_1607_sv2v_reg ;
  assign \piso.data_r [1606] = \piso.data_r_1606_sv2v_reg ;
  assign \piso.data_r [1605] = \piso.data_r_1605_sv2v_reg ;
  assign \piso.data_r [1604] = \piso.data_r_1604_sv2v_reg ;
  assign \piso.data_r [1603] = \piso.data_r_1603_sv2v_reg ;
  assign \piso.data_r [1602] = \piso.data_r_1602_sv2v_reg ;
  assign \piso.data_r [1601] = \piso.data_r_1601_sv2v_reg ;
  assign \piso.data_r [1600] = \piso.data_r_1600_sv2v_reg ;
  assign \piso.data_r [1599] = \piso.data_r_1599_sv2v_reg ;
  assign \piso.data_r [1598] = \piso.data_r_1598_sv2v_reg ;
  assign \piso.data_r [1597] = \piso.data_r_1597_sv2v_reg ;
  assign \piso.data_r [1596] = \piso.data_r_1596_sv2v_reg ;
  assign \piso.data_r [1595] = \piso.data_r_1595_sv2v_reg ;
  assign \piso.data_r [1594] = \piso.data_r_1594_sv2v_reg ;
  assign \piso.data_r [1593] = \piso.data_r_1593_sv2v_reg ;
  assign \piso.data_r [1592] = \piso.data_r_1592_sv2v_reg ;
  assign \piso.data_r [1591] = \piso.data_r_1591_sv2v_reg ;
  assign \piso.data_r [1590] = \piso.data_r_1590_sv2v_reg ;
  assign \piso.data_r [1589] = \piso.data_r_1589_sv2v_reg ;
  assign \piso.data_r [1588] = \piso.data_r_1588_sv2v_reg ;
  assign \piso.data_r [1587] = \piso.data_r_1587_sv2v_reg ;
  assign \piso.data_r [1586] = \piso.data_r_1586_sv2v_reg ;
  assign \piso.data_r [1585] = \piso.data_r_1585_sv2v_reg ;
  assign \piso.data_r [1584] = \piso.data_r_1584_sv2v_reg ;
  assign \piso.data_r [1583] = \piso.data_r_1583_sv2v_reg ;
  assign \piso.data_r [1582] = \piso.data_r_1582_sv2v_reg ;
  assign \piso.data_r [1581] = \piso.data_r_1581_sv2v_reg ;
  assign \piso.data_r [1580] = \piso.data_r_1580_sv2v_reg ;
  assign \piso.data_r [1579] = \piso.data_r_1579_sv2v_reg ;
  assign \piso.data_r [1578] = \piso.data_r_1578_sv2v_reg ;
  assign \piso.data_r [1577] = \piso.data_r_1577_sv2v_reg ;
  assign \piso.data_r [1576] = \piso.data_r_1576_sv2v_reg ;
  assign \piso.data_r [1575] = \piso.data_r_1575_sv2v_reg ;
  assign \piso.data_r [1574] = \piso.data_r_1574_sv2v_reg ;
  assign \piso.data_r [1573] = \piso.data_r_1573_sv2v_reg ;
  assign \piso.data_r [1572] = \piso.data_r_1572_sv2v_reg ;
  assign \piso.data_r [1571] = \piso.data_r_1571_sv2v_reg ;
  assign \piso.data_r [1570] = \piso.data_r_1570_sv2v_reg ;
  assign \piso.data_r [1569] = \piso.data_r_1569_sv2v_reg ;
  assign \piso.data_r [1568] = \piso.data_r_1568_sv2v_reg ;
  assign \piso.data_r [1567] = \piso.data_r_1567_sv2v_reg ;
  assign \piso.data_r [1566] = \piso.data_r_1566_sv2v_reg ;
  assign \piso.data_r [1565] = \piso.data_r_1565_sv2v_reg ;
  assign \piso.data_r [1564] = \piso.data_r_1564_sv2v_reg ;
  assign \piso.data_r [1563] = \piso.data_r_1563_sv2v_reg ;
  assign \piso.data_r [1562] = \piso.data_r_1562_sv2v_reg ;
  assign \piso.data_r [1561] = \piso.data_r_1561_sv2v_reg ;
  assign \piso.data_r [1560] = \piso.data_r_1560_sv2v_reg ;
  assign \piso.data_r [1559] = \piso.data_r_1559_sv2v_reg ;
  assign \piso.data_r [1558] = \piso.data_r_1558_sv2v_reg ;
  assign \piso.data_r [1557] = \piso.data_r_1557_sv2v_reg ;
  assign \piso.data_r [1556] = \piso.data_r_1556_sv2v_reg ;
  assign \piso.data_r [1555] = \piso.data_r_1555_sv2v_reg ;
  assign \piso.data_r [1554] = \piso.data_r_1554_sv2v_reg ;
  assign \piso.data_r [1553] = \piso.data_r_1553_sv2v_reg ;
  assign \piso.data_r [1552] = \piso.data_r_1552_sv2v_reg ;
  assign \piso.data_r [1551] = \piso.data_r_1551_sv2v_reg ;
  assign \piso.data_r [1550] = \piso.data_r_1550_sv2v_reg ;
  assign \piso.data_r [1549] = \piso.data_r_1549_sv2v_reg ;
  assign \piso.data_r [1548] = \piso.data_r_1548_sv2v_reg ;
  assign \piso.data_r [1547] = \piso.data_r_1547_sv2v_reg ;
  assign \piso.data_r [1546] = \piso.data_r_1546_sv2v_reg ;
  assign \piso.data_r [1545] = \piso.data_r_1545_sv2v_reg ;
  assign \piso.data_r [1544] = \piso.data_r_1544_sv2v_reg ;
  assign \piso.data_r [1543] = \piso.data_r_1543_sv2v_reg ;
  assign \piso.data_r [1542] = \piso.data_r_1542_sv2v_reg ;
  assign \piso.data_r [1541] = \piso.data_r_1541_sv2v_reg ;
  assign \piso.data_r [1540] = \piso.data_r_1540_sv2v_reg ;
  assign \piso.data_r [1539] = \piso.data_r_1539_sv2v_reg ;
  assign \piso.data_r [1538] = \piso.data_r_1538_sv2v_reg ;
  assign \piso.data_r [1537] = \piso.data_r_1537_sv2v_reg ;
  assign \piso.data_r [1536] = \piso.data_r_1536_sv2v_reg ;
  assign \piso.data_r [1535] = \piso.data_r_1535_sv2v_reg ;
  assign \piso.data_r [1534] = \piso.data_r_1534_sv2v_reg ;
  assign \piso.data_r [1533] = \piso.data_r_1533_sv2v_reg ;
  assign \piso.data_r [1532] = \piso.data_r_1532_sv2v_reg ;
  assign \piso.data_r [1531] = \piso.data_r_1531_sv2v_reg ;
  assign \piso.data_r [1530] = \piso.data_r_1530_sv2v_reg ;
  assign \piso.data_r [1529] = \piso.data_r_1529_sv2v_reg ;
  assign \piso.data_r [1528] = \piso.data_r_1528_sv2v_reg ;
  assign \piso.data_r [1527] = \piso.data_r_1527_sv2v_reg ;
  assign \piso.data_r [1526] = \piso.data_r_1526_sv2v_reg ;
  assign \piso.data_r [1525] = \piso.data_r_1525_sv2v_reg ;
  assign \piso.data_r [1524] = \piso.data_r_1524_sv2v_reg ;
  assign \piso.data_r [1523] = \piso.data_r_1523_sv2v_reg ;
  assign \piso.data_r [1522] = \piso.data_r_1522_sv2v_reg ;
  assign \piso.data_r [1521] = \piso.data_r_1521_sv2v_reg ;
  assign \piso.data_r [1520] = \piso.data_r_1520_sv2v_reg ;
  assign \piso.data_r [1519] = \piso.data_r_1519_sv2v_reg ;
  assign \piso.data_r [1518] = \piso.data_r_1518_sv2v_reg ;
  assign \piso.data_r [1517] = \piso.data_r_1517_sv2v_reg ;
  assign \piso.data_r [1516] = \piso.data_r_1516_sv2v_reg ;
  assign \piso.data_r [1515] = \piso.data_r_1515_sv2v_reg ;
  assign \piso.data_r [1514] = \piso.data_r_1514_sv2v_reg ;
  assign \piso.data_r [1513] = \piso.data_r_1513_sv2v_reg ;
  assign \piso.data_r [1512] = \piso.data_r_1512_sv2v_reg ;
  assign \piso.data_r [1511] = \piso.data_r_1511_sv2v_reg ;
  assign \piso.data_r [1510] = \piso.data_r_1510_sv2v_reg ;
  assign \piso.data_r [1509] = \piso.data_r_1509_sv2v_reg ;
  assign \piso.data_r [1508] = \piso.data_r_1508_sv2v_reg ;
  assign \piso.data_r [1507] = \piso.data_r_1507_sv2v_reg ;
  assign \piso.data_r [1506] = \piso.data_r_1506_sv2v_reg ;
  assign \piso.data_r [1505] = \piso.data_r_1505_sv2v_reg ;
  assign \piso.data_r [1504] = \piso.data_r_1504_sv2v_reg ;
  assign \piso.data_r [1503] = \piso.data_r_1503_sv2v_reg ;
  assign \piso.data_r [1502] = \piso.data_r_1502_sv2v_reg ;
  assign \piso.data_r [1501] = \piso.data_r_1501_sv2v_reg ;
  assign \piso.data_r [1500] = \piso.data_r_1500_sv2v_reg ;
  assign \piso.data_r [1499] = \piso.data_r_1499_sv2v_reg ;
  assign \piso.data_r [1498] = \piso.data_r_1498_sv2v_reg ;
  assign \piso.data_r [1497] = \piso.data_r_1497_sv2v_reg ;
  assign \piso.data_r [1496] = \piso.data_r_1496_sv2v_reg ;
  assign \piso.data_r [1495] = \piso.data_r_1495_sv2v_reg ;
  assign \piso.data_r [1494] = \piso.data_r_1494_sv2v_reg ;
  assign \piso.data_r [1493] = \piso.data_r_1493_sv2v_reg ;
  assign \piso.data_r [1492] = \piso.data_r_1492_sv2v_reg ;
  assign \piso.data_r [1491] = \piso.data_r_1491_sv2v_reg ;
  assign \piso.data_r [1490] = \piso.data_r_1490_sv2v_reg ;
  assign \piso.data_r [1489] = \piso.data_r_1489_sv2v_reg ;
  assign \piso.data_r [1488] = \piso.data_r_1488_sv2v_reg ;
  assign \piso.data_r [1487] = \piso.data_r_1487_sv2v_reg ;
  assign \piso.data_r [1486] = \piso.data_r_1486_sv2v_reg ;
  assign \piso.data_r [1485] = \piso.data_r_1485_sv2v_reg ;
  assign \piso.data_r [1484] = \piso.data_r_1484_sv2v_reg ;
  assign \piso.data_r [1483] = \piso.data_r_1483_sv2v_reg ;
  assign \piso.data_r [1482] = \piso.data_r_1482_sv2v_reg ;
  assign \piso.data_r [1481] = \piso.data_r_1481_sv2v_reg ;
  assign \piso.data_r [1480] = \piso.data_r_1480_sv2v_reg ;
  assign \piso.data_r [1479] = \piso.data_r_1479_sv2v_reg ;
  assign \piso.data_r [1478] = \piso.data_r_1478_sv2v_reg ;
  assign \piso.data_r [1477] = \piso.data_r_1477_sv2v_reg ;
  assign \piso.data_r [1476] = \piso.data_r_1476_sv2v_reg ;
  assign \piso.data_r [1475] = \piso.data_r_1475_sv2v_reg ;
  assign \piso.data_r [1474] = \piso.data_r_1474_sv2v_reg ;
  assign \piso.data_r [1473] = \piso.data_r_1473_sv2v_reg ;
  assign \piso.data_r [1472] = \piso.data_r_1472_sv2v_reg ;
  assign \piso.data_r [1471] = \piso.data_r_1471_sv2v_reg ;
  assign \piso.data_r [1470] = \piso.data_r_1470_sv2v_reg ;
  assign \piso.data_r [1469] = \piso.data_r_1469_sv2v_reg ;
  assign \piso.data_r [1468] = \piso.data_r_1468_sv2v_reg ;
  assign \piso.data_r [1467] = \piso.data_r_1467_sv2v_reg ;
  assign \piso.data_r [1466] = \piso.data_r_1466_sv2v_reg ;
  assign \piso.data_r [1465] = \piso.data_r_1465_sv2v_reg ;
  assign \piso.data_r [1464] = \piso.data_r_1464_sv2v_reg ;
  assign \piso.data_r [1463] = \piso.data_r_1463_sv2v_reg ;
  assign \piso.data_r [1462] = \piso.data_r_1462_sv2v_reg ;
  assign \piso.data_r [1461] = \piso.data_r_1461_sv2v_reg ;
  assign \piso.data_r [1460] = \piso.data_r_1460_sv2v_reg ;
  assign \piso.data_r [1459] = \piso.data_r_1459_sv2v_reg ;
  assign \piso.data_r [1458] = \piso.data_r_1458_sv2v_reg ;
  assign \piso.data_r [1457] = \piso.data_r_1457_sv2v_reg ;
  assign \piso.data_r [1456] = \piso.data_r_1456_sv2v_reg ;
  assign \piso.data_r [1455] = \piso.data_r_1455_sv2v_reg ;
  assign \piso.data_r [1454] = \piso.data_r_1454_sv2v_reg ;
  assign \piso.data_r [1453] = \piso.data_r_1453_sv2v_reg ;
  assign \piso.data_r [1452] = \piso.data_r_1452_sv2v_reg ;
  assign \piso.data_r [1451] = \piso.data_r_1451_sv2v_reg ;
  assign \piso.data_r [1450] = \piso.data_r_1450_sv2v_reg ;
  assign \piso.data_r [1449] = \piso.data_r_1449_sv2v_reg ;
  assign \piso.data_r [1448] = \piso.data_r_1448_sv2v_reg ;
  assign \piso.data_r [1447] = \piso.data_r_1447_sv2v_reg ;
  assign \piso.data_r [1446] = \piso.data_r_1446_sv2v_reg ;
  assign \piso.data_r [1445] = \piso.data_r_1445_sv2v_reg ;
  assign \piso.data_r [1444] = \piso.data_r_1444_sv2v_reg ;
  assign \piso.data_r [1443] = \piso.data_r_1443_sv2v_reg ;
  assign \piso.data_r [1442] = \piso.data_r_1442_sv2v_reg ;
  assign \piso.data_r [1441] = \piso.data_r_1441_sv2v_reg ;
  assign \piso.data_r [1440] = \piso.data_r_1440_sv2v_reg ;
  assign \piso.data_r [1439] = \piso.data_r_1439_sv2v_reg ;
  assign \piso.data_r [1438] = \piso.data_r_1438_sv2v_reg ;
  assign \piso.data_r [1437] = \piso.data_r_1437_sv2v_reg ;
  assign \piso.data_r [1436] = \piso.data_r_1436_sv2v_reg ;
  assign \piso.data_r [1435] = \piso.data_r_1435_sv2v_reg ;
  assign \piso.data_r [1434] = \piso.data_r_1434_sv2v_reg ;
  assign \piso.data_r [1433] = \piso.data_r_1433_sv2v_reg ;
  assign \piso.data_r [1432] = \piso.data_r_1432_sv2v_reg ;
  assign \piso.data_r [1431] = \piso.data_r_1431_sv2v_reg ;
  assign \piso.data_r [1430] = \piso.data_r_1430_sv2v_reg ;
  assign \piso.data_r [1429] = \piso.data_r_1429_sv2v_reg ;
  assign \piso.data_r [1428] = \piso.data_r_1428_sv2v_reg ;
  assign \piso.data_r [1427] = \piso.data_r_1427_sv2v_reg ;
  assign \piso.data_r [1426] = \piso.data_r_1426_sv2v_reg ;
  assign \piso.data_r [1425] = \piso.data_r_1425_sv2v_reg ;
  assign \piso.data_r [1424] = \piso.data_r_1424_sv2v_reg ;
  assign \piso.data_r [1423] = \piso.data_r_1423_sv2v_reg ;
  assign \piso.data_r [1422] = \piso.data_r_1422_sv2v_reg ;
  assign \piso.data_r [1421] = \piso.data_r_1421_sv2v_reg ;
  assign \piso.data_r [1420] = \piso.data_r_1420_sv2v_reg ;
  assign \piso.data_r [1419] = \piso.data_r_1419_sv2v_reg ;
  assign \piso.data_r [1418] = \piso.data_r_1418_sv2v_reg ;
  assign \piso.data_r [1417] = \piso.data_r_1417_sv2v_reg ;
  assign \piso.data_r [1416] = \piso.data_r_1416_sv2v_reg ;
  assign \piso.data_r [1415] = \piso.data_r_1415_sv2v_reg ;
  assign \piso.data_r [1414] = \piso.data_r_1414_sv2v_reg ;
  assign \piso.data_r [1413] = \piso.data_r_1413_sv2v_reg ;
  assign \piso.data_r [1412] = \piso.data_r_1412_sv2v_reg ;
  assign \piso.data_r [1411] = \piso.data_r_1411_sv2v_reg ;
  assign \piso.data_r [1410] = \piso.data_r_1410_sv2v_reg ;
  assign \piso.data_r [1409] = \piso.data_r_1409_sv2v_reg ;
  assign \piso.data_r [1408] = \piso.data_r_1408_sv2v_reg ;
  assign \piso.data_r [1407] = \piso.data_r_1407_sv2v_reg ;
  assign \piso.data_r [1406] = \piso.data_r_1406_sv2v_reg ;
  assign \piso.data_r [1405] = \piso.data_r_1405_sv2v_reg ;
  assign \piso.data_r [1404] = \piso.data_r_1404_sv2v_reg ;
  assign \piso.data_r [1403] = \piso.data_r_1403_sv2v_reg ;
  assign \piso.data_r [1402] = \piso.data_r_1402_sv2v_reg ;
  assign \piso.data_r [1401] = \piso.data_r_1401_sv2v_reg ;
  assign \piso.data_r [1400] = \piso.data_r_1400_sv2v_reg ;
  assign \piso.data_r [1399] = \piso.data_r_1399_sv2v_reg ;
  assign \piso.data_r [1398] = \piso.data_r_1398_sv2v_reg ;
  assign \piso.data_r [1397] = \piso.data_r_1397_sv2v_reg ;
  assign \piso.data_r [1396] = \piso.data_r_1396_sv2v_reg ;
  assign \piso.data_r [1395] = \piso.data_r_1395_sv2v_reg ;
  assign \piso.data_r [1394] = \piso.data_r_1394_sv2v_reg ;
  assign \piso.data_r [1393] = \piso.data_r_1393_sv2v_reg ;
  assign \piso.data_r [1392] = \piso.data_r_1392_sv2v_reg ;
  assign \piso.data_r [1391] = \piso.data_r_1391_sv2v_reg ;
  assign \piso.data_r [1390] = \piso.data_r_1390_sv2v_reg ;
  assign \piso.data_r [1389] = \piso.data_r_1389_sv2v_reg ;
  assign \piso.data_r [1388] = \piso.data_r_1388_sv2v_reg ;
  assign \piso.data_r [1387] = \piso.data_r_1387_sv2v_reg ;
  assign \piso.data_r [1386] = \piso.data_r_1386_sv2v_reg ;
  assign \piso.data_r [1385] = \piso.data_r_1385_sv2v_reg ;
  assign \piso.data_r [1384] = \piso.data_r_1384_sv2v_reg ;
  assign \piso.data_r [1383] = \piso.data_r_1383_sv2v_reg ;
  assign \piso.data_r [1382] = \piso.data_r_1382_sv2v_reg ;
  assign \piso.data_r [1381] = \piso.data_r_1381_sv2v_reg ;
  assign \piso.data_r [1380] = \piso.data_r_1380_sv2v_reg ;
  assign \piso.data_r [1379] = \piso.data_r_1379_sv2v_reg ;
  assign \piso.data_r [1378] = \piso.data_r_1378_sv2v_reg ;
  assign \piso.data_r [1377] = \piso.data_r_1377_sv2v_reg ;
  assign \piso.data_r [1376] = \piso.data_r_1376_sv2v_reg ;
  assign \piso.data_r [1375] = \piso.data_r_1375_sv2v_reg ;
  assign \piso.data_r [1374] = \piso.data_r_1374_sv2v_reg ;
  assign \piso.data_r [1373] = \piso.data_r_1373_sv2v_reg ;
  assign \piso.data_r [1372] = \piso.data_r_1372_sv2v_reg ;
  assign \piso.data_r [1371] = \piso.data_r_1371_sv2v_reg ;
  assign \piso.data_r [1370] = \piso.data_r_1370_sv2v_reg ;
  assign \piso.data_r [1369] = \piso.data_r_1369_sv2v_reg ;
  assign \piso.data_r [1368] = \piso.data_r_1368_sv2v_reg ;
  assign \piso.data_r [1367] = \piso.data_r_1367_sv2v_reg ;
  assign \piso.data_r [1366] = \piso.data_r_1366_sv2v_reg ;
  assign \piso.data_r [1365] = \piso.data_r_1365_sv2v_reg ;
  assign \piso.data_r [1364] = \piso.data_r_1364_sv2v_reg ;
  assign \piso.data_r [1363] = \piso.data_r_1363_sv2v_reg ;
  assign \piso.data_r [1362] = \piso.data_r_1362_sv2v_reg ;
  assign \piso.data_r [1361] = \piso.data_r_1361_sv2v_reg ;
  assign \piso.data_r [1360] = \piso.data_r_1360_sv2v_reg ;
  assign \piso.data_r [1359] = \piso.data_r_1359_sv2v_reg ;
  assign \piso.data_r [1358] = \piso.data_r_1358_sv2v_reg ;
  assign \piso.data_r [1357] = \piso.data_r_1357_sv2v_reg ;
  assign \piso.data_r [1356] = \piso.data_r_1356_sv2v_reg ;
  assign \piso.data_r [1355] = \piso.data_r_1355_sv2v_reg ;
  assign \piso.data_r [1354] = \piso.data_r_1354_sv2v_reg ;
  assign \piso.data_r [1353] = \piso.data_r_1353_sv2v_reg ;
  assign \piso.data_r [1352] = \piso.data_r_1352_sv2v_reg ;
  assign \piso.data_r [1351] = \piso.data_r_1351_sv2v_reg ;
  assign \piso.data_r [1350] = \piso.data_r_1350_sv2v_reg ;
  assign \piso.data_r [1349] = \piso.data_r_1349_sv2v_reg ;
  assign \piso.data_r [1348] = \piso.data_r_1348_sv2v_reg ;
  assign \piso.data_r [1347] = \piso.data_r_1347_sv2v_reg ;
  assign \piso.data_r [1346] = \piso.data_r_1346_sv2v_reg ;
  assign \piso.data_r [1345] = \piso.data_r_1345_sv2v_reg ;
  assign \piso.data_r [1344] = \piso.data_r_1344_sv2v_reg ;
  assign \piso.data_r [1343] = \piso.data_r_1343_sv2v_reg ;
  assign \piso.data_r [1342] = \piso.data_r_1342_sv2v_reg ;
  assign \piso.data_r [1341] = \piso.data_r_1341_sv2v_reg ;
  assign \piso.data_r [1340] = \piso.data_r_1340_sv2v_reg ;
  assign \piso.data_r [1339] = \piso.data_r_1339_sv2v_reg ;
  assign \piso.data_r [1338] = \piso.data_r_1338_sv2v_reg ;
  assign \piso.data_r [1337] = \piso.data_r_1337_sv2v_reg ;
  assign \piso.data_r [1336] = \piso.data_r_1336_sv2v_reg ;
  assign \piso.data_r [1335] = \piso.data_r_1335_sv2v_reg ;
  assign \piso.data_r [1334] = \piso.data_r_1334_sv2v_reg ;
  assign \piso.data_r [1333] = \piso.data_r_1333_sv2v_reg ;
  assign \piso.data_r [1332] = \piso.data_r_1332_sv2v_reg ;
  assign \piso.data_r [1331] = \piso.data_r_1331_sv2v_reg ;
  assign \piso.data_r [1330] = \piso.data_r_1330_sv2v_reg ;
  assign \piso.data_r [1329] = \piso.data_r_1329_sv2v_reg ;
  assign \piso.data_r [1328] = \piso.data_r_1328_sv2v_reg ;
  assign \piso.data_r [1327] = \piso.data_r_1327_sv2v_reg ;
  assign \piso.data_r [1326] = \piso.data_r_1326_sv2v_reg ;
  assign \piso.data_r [1325] = \piso.data_r_1325_sv2v_reg ;
  assign \piso.data_r [1324] = \piso.data_r_1324_sv2v_reg ;
  assign \piso.data_r [1323] = \piso.data_r_1323_sv2v_reg ;
  assign \piso.data_r [1322] = \piso.data_r_1322_sv2v_reg ;
  assign \piso.data_r [1321] = \piso.data_r_1321_sv2v_reg ;
  assign \piso.data_r [1320] = \piso.data_r_1320_sv2v_reg ;
  assign \piso.data_r [1319] = \piso.data_r_1319_sv2v_reg ;
  assign \piso.data_r [1318] = \piso.data_r_1318_sv2v_reg ;
  assign \piso.data_r [1317] = \piso.data_r_1317_sv2v_reg ;
  assign \piso.data_r [1316] = \piso.data_r_1316_sv2v_reg ;
  assign \piso.data_r [1315] = \piso.data_r_1315_sv2v_reg ;
  assign \piso.data_r [1314] = \piso.data_r_1314_sv2v_reg ;
  assign \piso.data_r [1313] = \piso.data_r_1313_sv2v_reg ;
  assign \piso.data_r [1312] = \piso.data_r_1312_sv2v_reg ;
  assign \piso.data_r [1311] = \piso.data_r_1311_sv2v_reg ;
  assign \piso.data_r [1310] = \piso.data_r_1310_sv2v_reg ;
  assign \piso.data_r [1309] = \piso.data_r_1309_sv2v_reg ;
  assign \piso.data_r [1308] = \piso.data_r_1308_sv2v_reg ;
  assign \piso.data_r [1307] = \piso.data_r_1307_sv2v_reg ;
  assign \piso.data_r [1306] = \piso.data_r_1306_sv2v_reg ;
  assign \piso.data_r [1305] = \piso.data_r_1305_sv2v_reg ;
  assign \piso.data_r [1304] = \piso.data_r_1304_sv2v_reg ;
  assign \piso.data_r [1303] = \piso.data_r_1303_sv2v_reg ;
  assign \piso.data_r [1302] = \piso.data_r_1302_sv2v_reg ;
  assign \piso.data_r [1301] = \piso.data_r_1301_sv2v_reg ;
  assign \piso.data_r [1300] = \piso.data_r_1300_sv2v_reg ;
  assign \piso.data_r [1299] = \piso.data_r_1299_sv2v_reg ;
  assign \piso.data_r [1298] = \piso.data_r_1298_sv2v_reg ;
  assign \piso.data_r [1297] = \piso.data_r_1297_sv2v_reg ;
  assign \piso.data_r [1296] = \piso.data_r_1296_sv2v_reg ;
  assign \piso.data_r [1295] = \piso.data_r_1295_sv2v_reg ;
  assign \piso.data_r [1294] = \piso.data_r_1294_sv2v_reg ;
  assign \piso.data_r [1293] = \piso.data_r_1293_sv2v_reg ;
  assign \piso.data_r [1292] = \piso.data_r_1292_sv2v_reg ;
  assign \piso.data_r [1291] = \piso.data_r_1291_sv2v_reg ;
  assign \piso.data_r [1290] = \piso.data_r_1290_sv2v_reg ;
  assign \piso.data_r [1289] = \piso.data_r_1289_sv2v_reg ;
  assign \piso.data_r [1288] = \piso.data_r_1288_sv2v_reg ;
  assign \piso.data_r [1287] = \piso.data_r_1287_sv2v_reg ;
  assign \piso.data_r [1286] = \piso.data_r_1286_sv2v_reg ;
  assign \piso.data_r [1285] = \piso.data_r_1285_sv2v_reg ;
  assign \piso.data_r [1284] = \piso.data_r_1284_sv2v_reg ;
  assign \piso.data_r [1283] = \piso.data_r_1283_sv2v_reg ;
  assign \piso.data_r [1282] = \piso.data_r_1282_sv2v_reg ;
  assign \piso.data_r [1281] = \piso.data_r_1281_sv2v_reg ;
  assign \piso.data_r [1280] = \piso.data_r_1280_sv2v_reg ;
  assign \piso.data_r [1279] = \piso.data_r_1279_sv2v_reg ;
  assign \piso.data_r [1278] = \piso.data_r_1278_sv2v_reg ;
  assign \piso.data_r [1277] = \piso.data_r_1277_sv2v_reg ;
  assign \piso.data_r [1276] = \piso.data_r_1276_sv2v_reg ;
  assign \piso.data_r [1275] = \piso.data_r_1275_sv2v_reg ;
  assign \piso.data_r [1274] = \piso.data_r_1274_sv2v_reg ;
  assign \piso.data_r [1273] = \piso.data_r_1273_sv2v_reg ;
  assign \piso.data_r [1272] = \piso.data_r_1272_sv2v_reg ;
  assign \piso.data_r [1271] = \piso.data_r_1271_sv2v_reg ;
  assign \piso.data_r [1270] = \piso.data_r_1270_sv2v_reg ;
  assign \piso.data_r [1269] = \piso.data_r_1269_sv2v_reg ;
  assign \piso.data_r [1268] = \piso.data_r_1268_sv2v_reg ;
  assign \piso.data_r [1267] = \piso.data_r_1267_sv2v_reg ;
  assign \piso.data_r [1266] = \piso.data_r_1266_sv2v_reg ;
  assign \piso.data_r [1265] = \piso.data_r_1265_sv2v_reg ;
  assign \piso.data_r [1264] = \piso.data_r_1264_sv2v_reg ;
  assign \piso.data_r [1263] = \piso.data_r_1263_sv2v_reg ;
  assign \piso.data_r [1262] = \piso.data_r_1262_sv2v_reg ;
  assign \piso.data_r [1261] = \piso.data_r_1261_sv2v_reg ;
  assign \piso.data_r [1260] = \piso.data_r_1260_sv2v_reg ;
  assign \piso.data_r [1259] = \piso.data_r_1259_sv2v_reg ;
  assign \piso.data_r [1258] = \piso.data_r_1258_sv2v_reg ;
  assign \piso.data_r [1257] = \piso.data_r_1257_sv2v_reg ;
  assign \piso.data_r [1256] = \piso.data_r_1256_sv2v_reg ;
  assign \piso.data_r [1255] = \piso.data_r_1255_sv2v_reg ;
  assign \piso.data_r [1254] = \piso.data_r_1254_sv2v_reg ;
  assign \piso.data_r [1253] = \piso.data_r_1253_sv2v_reg ;
  assign \piso.data_r [1252] = \piso.data_r_1252_sv2v_reg ;
  assign \piso.data_r [1251] = \piso.data_r_1251_sv2v_reg ;
  assign \piso.data_r [1250] = \piso.data_r_1250_sv2v_reg ;
  assign \piso.data_r [1249] = \piso.data_r_1249_sv2v_reg ;
  assign \piso.data_r [1248] = \piso.data_r_1248_sv2v_reg ;
  assign \piso.data_r [1247] = \piso.data_r_1247_sv2v_reg ;
  assign \piso.data_r [1246] = \piso.data_r_1246_sv2v_reg ;
  assign \piso.data_r [1245] = \piso.data_r_1245_sv2v_reg ;
  assign \piso.data_r [1244] = \piso.data_r_1244_sv2v_reg ;
  assign \piso.data_r [1243] = \piso.data_r_1243_sv2v_reg ;
  assign \piso.data_r [1242] = \piso.data_r_1242_sv2v_reg ;
  assign \piso.data_r [1241] = \piso.data_r_1241_sv2v_reg ;
  assign \piso.data_r [1240] = \piso.data_r_1240_sv2v_reg ;
  assign \piso.data_r [1239] = \piso.data_r_1239_sv2v_reg ;
  assign \piso.data_r [1238] = \piso.data_r_1238_sv2v_reg ;
  assign \piso.data_r [1237] = \piso.data_r_1237_sv2v_reg ;
  assign \piso.data_r [1236] = \piso.data_r_1236_sv2v_reg ;
  assign \piso.data_r [1235] = \piso.data_r_1235_sv2v_reg ;
  assign \piso.data_r [1234] = \piso.data_r_1234_sv2v_reg ;
  assign \piso.data_r [1233] = \piso.data_r_1233_sv2v_reg ;
  assign \piso.data_r [1232] = \piso.data_r_1232_sv2v_reg ;
  assign \piso.data_r [1231] = \piso.data_r_1231_sv2v_reg ;
  assign \piso.data_r [1230] = \piso.data_r_1230_sv2v_reg ;
  assign \piso.data_r [1229] = \piso.data_r_1229_sv2v_reg ;
  assign \piso.data_r [1228] = \piso.data_r_1228_sv2v_reg ;
  assign \piso.data_r [1227] = \piso.data_r_1227_sv2v_reg ;
  assign \piso.data_r [1226] = \piso.data_r_1226_sv2v_reg ;
  assign \piso.data_r [1225] = \piso.data_r_1225_sv2v_reg ;
  assign \piso.data_r [1224] = \piso.data_r_1224_sv2v_reg ;
  assign \piso.data_r [1223] = \piso.data_r_1223_sv2v_reg ;
  assign \piso.data_r [1222] = \piso.data_r_1222_sv2v_reg ;
  assign \piso.data_r [1221] = \piso.data_r_1221_sv2v_reg ;
  assign \piso.data_r [1220] = \piso.data_r_1220_sv2v_reg ;
  assign \piso.data_r [1219] = \piso.data_r_1219_sv2v_reg ;
  assign \piso.data_r [1218] = \piso.data_r_1218_sv2v_reg ;
  assign \piso.data_r [1217] = \piso.data_r_1217_sv2v_reg ;
  assign \piso.data_r [1216] = \piso.data_r_1216_sv2v_reg ;
  assign \piso.data_r [1215] = \piso.data_r_1215_sv2v_reg ;
  assign \piso.data_r [1214] = \piso.data_r_1214_sv2v_reg ;
  assign \piso.data_r [1213] = \piso.data_r_1213_sv2v_reg ;
  assign \piso.data_r [1212] = \piso.data_r_1212_sv2v_reg ;
  assign \piso.data_r [1211] = \piso.data_r_1211_sv2v_reg ;
  assign \piso.data_r [1210] = \piso.data_r_1210_sv2v_reg ;
  assign \piso.data_r [1209] = \piso.data_r_1209_sv2v_reg ;
  assign \piso.data_r [1208] = \piso.data_r_1208_sv2v_reg ;
  assign \piso.data_r [1207] = \piso.data_r_1207_sv2v_reg ;
  assign \piso.data_r [1206] = \piso.data_r_1206_sv2v_reg ;
  assign \piso.data_r [1205] = \piso.data_r_1205_sv2v_reg ;
  assign \piso.data_r [1204] = \piso.data_r_1204_sv2v_reg ;
  assign \piso.data_r [1203] = \piso.data_r_1203_sv2v_reg ;
  assign \piso.data_r [1202] = \piso.data_r_1202_sv2v_reg ;
  assign \piso.data_r [1201] = \piso.data_r_1201_sv2v_reg ;
  assign \piso.data_r [1200] = \piso.data_r_1200_sv2v_reg ;
  assign \piso.data_r [1199] = \piso.data_r_1199_sv2v_reg ;
  assign \piso.data_r [1198] = \piso.data_r_1198_sv2v_reg ;
  assign \piso.data_r [1197] = \piso.data_r_1197_sv2v_reg ;
  assign \piso.data_r [1196] = \piso.data_r_1196_sv2v_reg ;
  assign \piso.data_r [1195] = \piso.data_r_1195_sv2v_reg ;
  assign \piso.data_r [1194] = \piso.data_r_1194_sv2v_reg ;
  assign \piso.data_r [1193] = \piso.data_r_1193_sv2v_reg ;
  assign \piso.data_r [1192] = \piso.data_r_1192_sv2v_reg ;
  assign \piso.data_r [1191] = \piso.data_r_1191_sv2v_reg ;
  assign \piso.data_r [1190] = \piso.data_r_1190_sv2v_reg ;
  assign \piso.data_r [1189] = \piso.data_r_1189_sv2v_reg ;
  assign \piso.data_r [1188] = \piso.data_r_1188_sv2v_reg ;
  assign \piso.data_r [1187] = \piso.data_r_1187_sv2v_reg ;
  assign \piso.data_r [1186] = \piso.data_r_1186_sv2v_reg ;
  assign \piso.data_r [1185] = \piso.data_r_1185_sv2v_reg ;
  assign \piso.data_r [1184] = \piso.data_r_1184_sv2v_reg ;
  assign \piso.data_r [1183] = \piso.data_r_1183_sv2v_reg ;
  assign \piso.data_r [1182] = \piso.data_r_1182_sv2v_reg ;
  assign \piso.data_r [1181] = \piso.data_r_1181_sv2v_reg ;
  assign \piso.data_r [1180] = \piso.data_r_1180_sv2v_reg ;
  assign \piso.data_r [1179] = \piso.data_r_1179_sv2v_reg ;
  assign \piso.data_r [1178] = \piso.data_r_1178_sv2v_reg ;
  assign \piso.data_r [1177] = \piso.data_r_1177_sv2v_reg ;
  assign \piso.data_r [1176] = \piso.data_r_1176_sv2v_reg ;
  assign \piso.data_r [1175] = \piso.data_r_1175_sv2v_reg ;
  assign \piso.data_r [1174] = \piso.data_r_1174_sv2v_reg ;
  assign \piso.data_r [1173] = \piso.data_r_1173_sv2v_reg ;
  assign \piso.data_r [1172] = \piso.data_r_1172_sv2v_reg ;
  assign \piso.data_r [1171] = \piso.data_r_1171_sv2v_reg ;
  assign \piso.data_r [1170] = \piso.data_r_1170_sv2v_reg ;
  assign \piso.data_r [1169] = \piso.data_r_1169_sv2v_reg ;
  assign \piso.data_r [1168] = \piso.data_r_1168_sv2v_reg ;
  assign \piso.data_r [1167] = \piso.data_r_1167_sv2v_reg ;
  assign \piso.data_r [1166] = \piso.data_r_1166_sv2v_reg ;
  assign \piso.data_r [1165] = \piso.data_r_1165_sv2v_reg ;
  assign \piso.data_r [1164] = \piso.data_r_1164_sv2v_reg ;
  assign \piso.data_r [1163] = \piso.data_r_1163_sv2v_reg ;
  assign \piso.data_r [1162] = \piso.data_r_1162_sv2v_reg ;
  assign \piso.data_r [1161] = \piso.data_r_1161_sv2v_reg ;
  assign \piso.data_r [1160] = \piso.data_r_1160_sv2v_reg ;
  assign \piso.data_r [1159] = \piso.data_r_1159_sv2v_reg ;
  assign \piso.data_r [1158] = \piso.data_r_1158_sv2v_reg ;
  assign \piso.data_r [1157] = \piso.data_r_1157_sv2v_reg ;
  assign \piso.data_r [1156] = \piso.data_r_1156_sv2v_reg ;
  assign \piso.data_r [1155] = \piso.data_r_1155_sv2v_reg ;
  assign \piso.data_r [1154] = \piso.data_r_1154_sv2v_reg ;
  assign \piso.data_r [1153] = \piso.data_r_1153_sv2v_reg ;
  assign \piso.data_r [1152] = \piso.data_r_1152_sv2v_reg ;
  assign \piso.data_r [1151] = \piso.data_r_1151_sv2v_reg ;
  assign \piso.data_r [1150] = \piso.data_r_1150_sv2v_reg ;
  assign \piso.data_r [1149] = \piso.data_r_1149_sv2v_reg ;
  assign \piso.data_r [1148] = \piso.data_r_1148_sv2v_reg ;
  assign \piso.data_r [1147] = \piso.data_r_1147_sv2v_reg ;
  assign \piso.data_r [1146] = \piso.data_r_1146_sv2v_reg ;
  assign \piso.data_r [1145] = \piso.data_r_1145_sv2v_reg ;
  assign \piso.data_r [1144] = \piso.data_r_1144_sv2v_reg ;
  assign \piso.data_r [1143] = \piso.data_r_1143_sv2v_reg ;
  assign \piso.data_r [1142] = \piso.data_r_1142_sv2v_reg ;
  assign \piso.data_r [1141] = \piso.data_r_1141_sv2v_reg ;
  assign \piso.data_r [1140] = \piso.data_r_1140_sv2v_reg ;
  assign \piso.data_r [1139] = \piso.data_r_1139_sv2v_reg ;
  assign \piso.data_r [1138] = \piso.data_r_1138_sv2v_reg ;
  assign \piso.data_r [1137] = \piso.data_r_1137_sv2v_reg ;
  assign \piso.data_r [1136] = \piso.data_r_1136_sv2v_reg ;
  assign \piso.data_r [1135] = \piso.data_r_1135_sv2v_reg ;
  assign \piso.data_r [1134] = \piso.data_r_1134_sv2v_reg ;
  assign \piso.data_r [1133] = \piso.data_r_1133_sv2v_reg ;
  assign \piso.data_r [1132] = \piso.data_r_1132_sv2v_reg ;
  assign \piso.data_r [1131] = \piso.data_r_1131_sv2v_reg ;
  assign \piso.data_r [1130] = \piso.data_r_1130_sv2v_reg ;
  assign \piso.data_r [1129] = \piso.data_r_1129_sv2v_reg ;
  assign \piso.data_r [1128] = \piso.data_r_1128_sv2v_reg ;
  assign \piso.data_r [1127] = \piso.data_r_1127_sv2v_reg ;
  assign \piso.data_r [1126] = \piso.data_r_1126_sv2v_reg ;
  assign \piso.data_r [1125] = \piso.data_r_1125_sv2v_reg ;
  assign \piso.data_r [1124] = \piso.data_r_1124_sv2v_reg ;
  assign \piso.data_r [1123] = \piso.data_r_1123_sv2v_reg ;
  assign \piso.data_r [1122] = \piso.data_r_1122_sv2v_reg ;
  assign \piso.data_r [1121] = \piso.data_r_1121_sv2v_reg ;
  assign \piso.data_r [1120] = \piso.data_r_1120_sv2v_reg ;
  assign \piso.data_r [1119] = \piso.data_r_1119_sv2v_reg ;
  assign \piso.data_r [1118] = \piso.data_r_1118_sv2v_reg ;
  assign \piso.data_r [1117] = \piso.data_r_1117_sv2v_reg ;
  assign \piso.data_r [1116] = \piso.data_r_1116_sv2v_reg ;
  assign \piso.data_r [1115] = \piso.data_r_1115_sv2v_reg ;
  assign \piso.data_r [1114] = \piso.data_r_1114_sv2v_reg ;
  assign \piso.data_r [1113] = \piso.data_r_1113_sv2v_reg ;
  assign \piso.data_r [1112] = \piso.data_r_1112_sv2v_reg ;
  assign \piso.data_r [1111] = \piso.data_r_1111_sv2v_reg ;
  assign \piso.data_r [1110] = \piso.data_r_1110_sv2v_reg ;
  assign \piso.data_r [1109] = \piso.data_r_1109_sv2v_reg ;
  assign \piso.data_r [1108] = \piso.data_r_1108_sv2v_reg ;
  assign \piso.data_r [1107] = \piso.data_r_1107_sv2v_reg ;
  assign \piso.data_r [1106] = \piso.data_r_1106_sv2v_reg ;
  assign \piso.data_r [1105] = \piso.data_r_1105_sv2v_reg ;
  assign \piso.data_r [1104] = \piso.data_r_1104_sv2v_reg ;
  assign \piso.data_r [1103] = \piso.data_r_1103_sv2v_reg ;
  assign \piso.data_r [1102] = \piso.data_r_1102_sv2v_reg ;
  assign \piso.data_r [1101] = \piso.data_r_1101_sv2v_reg ;
  assign \piso.data_r [1100] = \piso.data_r_1100_sv2v_reg ;
  assign \piso.data_r [1099] = \piso.data_r_1099_sv2v_reg ;
  assign \piso.data_r [1098] = \piso.data_r_1098_sv2v_reg ;
  assign \piso.data_r [1097] = \piso.data_r_1097_sv2v_reg ;
  assign \piso.data_r [1096] = \piso.data_r_1096_sv2v_reg ;
  assign \piso.data_r [1095] = \piso.data_r_1095_sv2v_reg ;
  assign \piso.data_r [1094] = \piso.data_r_1094_sv2v_reg ;
  assign \piso.data_r [1093] = \piso.data_r_1093_sv2v_reg ;
  assign \piso.data_r [1092] = \piso.data_r_1092_sv2v_reg ;
  assign \piso.data_r [1091] = \piso.data_r_1091_sv2v_reg ;
  assign \piso.data_r [1090] = \piso.data_r_1090_sv2v_reg ;
  assign \piso.data_r [1089] = \piso.data_r_1089_sv2v_reg ;
  assign \piso.data_r [1088] = \piso.data_r_1088_sv2v_reg ;
  assign \piso.data_r [1087] = \piso.data_r_1087_sv2v_reg ;
  assign \piso.data_r [1086] = \piso.data_r_1086_sv2v_reg ;
  assign \piso.data_r [1085] = \piso.data_r_1085_sv2v_reg ;
  assign \piso.data_r [1084] = \piso.data_r_1084_sv2v_reg ;
  assign \piso.data_r [1083] = \piso.data_r_1083_sv2v_reg ;
  assign \piso.data_r [1082] = \piso.data_r_1082_sv2v_reg ;
  assign \piso.data_r [1081] = \piso.data_r_1081_sv2v_reg ;
  assign \piso.data_r [1080] = \piso.data_r_1080_sv2v_reg ;
  assign \piso.data_r [1079] = \piso.data_r_1079_sv2v_reg ;
  assign \piso.data_r [1078] = \piso.data_r_1078_sv2v_reg ;
  assign \piso.data_r [1077] = \piso.data_r_1077_sv2v_reg ;
  assign \piso.data_r [1076] = \piso.data_r_1076_sv2v_reg ;
  assign \piso.data_r [1075] = \piso.data_r_1075_sv2v_reg ;
  assign \piso.data_r [1074] = \piso.data_r_1074_sv2v_reg ;
  assign \piso.data_r [1073] = \piso.data_r_1073_sv2v_reg ;
  assign \piso.data_r [1072] = \piso.data_r_1072_sv2v_reg ;
  assign \piso.data_r [1071] = \piso.data_r_1071_sv2v_reg ;
  assign \piso.data_r [1070] = \piso.data_r_1070_sv2v_reg ;
  assign \piso.data_r [1069] = \piso.data_r_1069_sv2v_reg ;
  assign \piso.data_r [1068] = \piso.data_r_1068_sv2v_reg ;
  assign \piso.data_r [1067] = \piso.data_r_1067_sv2v_reg ;
  assign \piso.data_r [1066] = \piso.data_r_1066_sv2v_reg ;
  assign \piso.data_r [1065] = \piso.data_r_1065_sv2v_reg ;
  assign \piso.data_r [1064] = \piso.data_r_1064_sv2v_reg ;
  assign \piso.data_r [1063] = \piso.data_r_1063_sv2v_reg ;
  assign \piso.data_r [1062] = \piso.data_r_1062_sv2v_reg ;
  assign \piso.data_r [1061] = \piso.data_r_1061_sv2v_reg ;
  assign \piso.data_r [1060] = \piso.data_r_1060_sv2v_reg ;
  assign \piso.data_r [1059] = \piso.data_r_1059_sv2v_reg ;
  assign \piso.data_r [1058] = \piso.data_r_1058_sv2v_reg ;
  assign \piso.data_r [1057] = \piso.data_r_1057_sv2v_reg ;
  assign \piso.data_r [1056] = \piso.data_r_1056_sv2v_reg ;
  assign \piso.data_r [1055] = \piso.data_r_1055_sv2v_reg ;
  assign \piso.data_r [1054] = \piso.data_r_1054_sv2v_reg ;
  assign \piso.data_r [1053] = \piso.data_r_1053_sv2v_reg ;
  assign \piso.data_r [1052] = \piso.data_r_1052_sv2v_reg ;
  assign \piso.data_r [1051] = \piso.data_r_1051_sv2v_reg ;
  assign \piso.data_r [1050] = \piso.data_r_1050_sv2v_reg ;
  assign \piso.data_r [1049] = \piso.data_r_1049_sv2v_reg ;
  assign \piso.data_r [1048] = \piso.data_r_1048_sv2v_reg ;
  assign \piso.data_r [1047] = \piso.data_r_1047_sv2v_reg ;
  assign \piso.data_r [1046] = \piso.data_r_1046_sv2v_reg ;
  assign \piso.data_r [1045] = \piso.data_r_1045_sv2v_reg ;
  assign \piso.data_r [1044] = \piso.data_r_1044_sv2v_reg ;
  assign \piso.data_r [1043] = \piso.data_r_1043_sv2v_reg ;
  assign \piso.data_r [1042] = \piso.data_r_1042_sv2v_reg ;
  assign \piso.data_r [1041] = \piso.data_r_1041_sv2v_reg ;
  assign \piso.data_r [1040] = \piso.data_r_1040_sv2v_reg ;
  assign \piso.data_r [1039] = \piso.data_r_1039_sv2v_reg ;
  assign \piso.data_r [1038] = \piso.data_r_1038_sv2v_reg ;
  assign \piso.data_r [1037] = \piso.data_r_1037_sv2v_reg ;
  assign \piso.data_r [1036] = \piso.data_r_1036_sv2v_reg ;
  assign \piso.data_r [1035] = \piso.data_r_1035_sv2v_reg ;
  assign \piso.data_r [1034] = \piso.data_r_1034_sv2v_reg ;
  assign \piso.data_r [1033] = \piso.data_r_1033_sv2v_reg ;
  assign \piso.data_r [1032] = \piso.data_r_1032_sv2v_reg ;
  assign \piso.data_r [1031] = \piso.data_r_1031_sv2v_reg ;
  assign \piso.data_r [1030] = \piso.data_r_1030_sv2v_reg ;
  assign \piso.data_r [1029] = \piso.data_r_1029_sv2v_reg ;
  assign \piso.data_r [1028] = \piso.data_r_1028_sv2v_reg ;
  assign \piso.data_r [1027] = \piso.data_r_1027_sv2v_reg ;
  assign \piso.data_r [1026] = \piso.data_r_1026_sv2v_reg ;
  assign \piso.data_r [1025] = \piso.data_r_1025_sv2v_reg ;
  assign \piso.data_r [1024] = \piso.data_r_1024_sv2v_reg ;
  assign \piso.data_r [1023] = \piso.data_r_1023_sv2v_reg ;
  assign \piso.data_r [1022] = \piso.data_r_1022_sv2v_reg ;
  assign \piso.data_r [1021] = \piso.data_r_1021_sv2v_reg ;
  assign \piso.data_r [1020] = \piso.data_r_1020_sv2v_reg ;
  assign \piso.data_r [1019] = \piso.data_r_1019_sv2v_reg ;
  assign \piso.data_r [1018] = \piso.data_r_1018_sv2v_reg ;
  assign \piso.data_r [1017] = \piso.data_r_1017_sv2v_reg ;
  assign \piso.data_r [1016] = \piso.data_r_1016_sv2v_reg ;
  assign \piso.data_r [1015] = \piso.data_r_1015_sv2v_reg ;
  assign \piso.data_r [1014] = \piso.data_r_1014_sv2v_reg ;
  assign \piso.data_r [1013] = \piso.data_r_1013_sv2v_reg ;
  assign \piso.data_r [1012] = \piso.data_r_1012_sv2v_reg ;
  assign \piso.data_r [1011] = \piso.data_r_1011_sv2v_reg ;
  assign \piso.data_r [1010] = \piso.data_r_1010_sv2v_reg ;
  assign \piso.data_r [1009] = \piso.data_r_1009_sv2v_reg ;
  assign \piso.data_r [1008] = \piso.data_r_1008_sv2v_reg ;
  assign \piso.data_r [1007] = \piso.data_r_1007_sv2v_reg ;
  assign \piso.data_r [1006] = \piso.data_r_1006_sv2v_reg ;
  assign \piso.data_r [1005] = \piso.data_r_1005_sv2v_reg ;
  assign \piso.data_r [1004] = \piso.data_r_1004_sv2v_reg ;
  assign \piso.data_r [1003] = \piso.data_r_1003_sv2v_reg ;
  assign \piso.data_r [1002] = \piso.data_r_1002_sv2v_reg ;
  assign \piso.data_r [1001] = \piso.data_r_1001_sv2v_reg ;
  assign \piso.data_r [1000] = \piso.data_r_1000_sv2v_reg ;
  assign \piso.data_r [999] = \piso.data_r_999_sv2v_reg ;
  assign \piso.data_r [998] = \piso.data_r_998_sv2v_reg ;
  assign \piso.data_r [997] = \piso.data_r_997_sv2v_reg ;
  assign \piso.data_r [996] = \piso.data_r_996_sv2v_reg ;
  assign \piso.data_r [995] = \piso.data_r_995_sv2v_reg ;
  assign \piso.data_r [994] = \piso.data_r_994_sv2v_reg ;
  assign \piso.data_r [993] = \piso.data_r_993_sv2v_reg ;
  assign \piso.data_r [992] = \piso.data_r_992_sv2v_reg ;
  assign \piso.data_r [991] = \piso.data_r_991_sv2v_reg ;
  assign \piso.data_r [990] = \piso.data_r_990_sv2v_reg ;
  assign \piso.data_r [989] = \piso.data_r_989_sv2v_reg ;
  assign \piso.data_r [988] = \piso.data_r_988_sv2v_reg ;
  assign \piso.data_r [987] = \piso.data_r_987_sv2v_reg ;
  assign \piso.data_r [986] = \piso.data_r_986_sv2v_reg ;
  assign \piso.data_r [985] = \piso.data_r_985_sv2v_reg ;
  assign \piso.data_r [984] = \piso.data_r_984_sv2v_reg ;
  assign \piso.data_r [983] = \piso.data_r_983_sv2v_reg ;
  assign \piso.data_r [982] = \piso.data_r_982_sv2v_reg ;
  assign \piso.data_r [981] = \piso.data_r_981_sv2v_reg ;
  assign \piso.data_r [980] = \piso.data_r_980_sv2v_reg ;
  assign \piso.data_r [979] = \piso.data_r_979_sv2v_reg ;
  assign \piso.data_r [978] = \piso.data_r_978_sv2v_reg ;
  assign \piso.data_r [977] = \piso.data_r_977_sv2v_reg ;
  assign \piso.data_r [976] = \piso.data_r_976_sv2v_reg ;
  assign \piso.data_r [975] = \piso.data_r_975_sv2v_reg ;
  assign \piso.data_r [974] = \piso.data_r_974_sv2v_reg ;
  assign \piso.data_r [973] = \piso.data_r_973_sv2v_reg ;
  assign \piso.data_r [972] = \piso.data_r_972_sv2v_reg ;
  assign \piso.data_r [971] = \piso.data_r_971_sv2v_reg ;
  assign \piso.data_r [970] = \piso.data_r_970_sv2v_reg ;
  assign \piso.data_r [969] = \piso.data_r_969_sv2v_reg ;
  assign \piso.data_r [968] = \piso.data_r_968_sv2v_reg ;
  assign \piso.data_r [967] = \piso.data_r_967_sv2v_reg ;
  assign \piso.data_r [966] = \piso.data_r_966_sv2v_reg ;
  assign \piso.data_r [965] = \piso.data_r_965_sv2v_reg ;
  assign \piso.data_r [964] = \piso.data_r_964_sv2v_reg ;
  assign \piso.data_r [963] = \piso.data_r_963_sv2v_reg ;
  assign \piso.data_r [962] = \piso.data_r_962_sv2v_reg ;
  assign \piso.data_r [961] = \piso.data_r_961_sv2v_reg ;
  assign \piso.data_r [960] = \piso.data_r_960_sv2v_reg ;
  assign \piso.data_r [959] = \piso.data_r_959_sv2v_reg ;
  assign \piso.data_r [958] = \piso.data_r_958_sv2v_reg ;
  assign \piso.data_r [957] = \piso.data_r_957_sv2v_reg ;
  assign \piso.data_r [956] = \piso.data_r_956_sv2v_reg ;
  assign \piso.data_r [955] = \piso.data_r_955_sv2v_reg ;
  assign \piso.data_r [954] = \piso.data_r_954_sv2v_reg ;
  assign \piso.data_r [953] = \piso.data_r_953_sv2v_reg ;
  assign \piso.data_r [952] = \piso.data_r_952_sv2v_reg ;
  assign \piso.data_r [951] = \piso.data_r_951_sv2v_reg ;
  assign \piso.data_r [950] = \piso.data_r_950_sv2v_reg ;
  assign \piso.data_r [949] = \piso.data_r_949_sv2v_reg ;
  assign \piso.data_r [948] = \piso.data_r_948_sv2v_reg ;
  assign \piso.data_r [947] = \piso.data_r_947_sv2v_reg ;
  assign \piso.data_r [946] = \piso.data_r_946_sv2v_reg ;
  assign \piso.data_r [945] = \piso.data_r_945_sv2v_reg ;
  assign \piso.data_r [944] = \piso.data_r_944_sv2v_reg ;
  assign \piso.data_r [943] = \piso.data_r_943_sv2v_reg ;
  assign \piso.data_r [942] = \piso.data_r_942_sv2v_reg ;
  assign \piso.data_r [941] = \piso.data_r_941_sv2v_reg ;
  assign \piso.data_r [940] = \piso.data_r_940_sv2v_reg ;
  assign \piso.data_r [939] = \piso.data_r_939_sv2v_reg ;
  assign \piso.data_r [938] = \piso.data_r_938_sv2v_reg ;
  assign \piso.data_r [937] = \piso.data_r_937_sv2v_reg ;
  assign \piso.data_r [936] = \piso.data_r_936_sv2v_reg ;
  assign \piso.data_r [935] = \piso.data_r_935_sv2v_reg ;
  assign \piso.data_r [934] = \piso.data_r_934_sv2v_reg ;
  assign \piso.data_r [933] = \piso.data_r_933_sv2v_reg ;
  assign \piso.data_r [932] = \piso.data_r_932_sv2v_reg ;
  assign \piso.data_r [931] = \piso.data_r_931_sv2v_reg ;
  assign \piso.data_r [930] = \piso.data_r_930_sv2v_reg ;
  assign \piso.data_r [929] = \piso.data_r_929_sv2v_reg ;
  assign \piso.data_r [928] = \piso.data_r_928_sv2v_reg ;
  assign \piso.data_r [927] = \piso.data_r_927_sv2v_reg ;
  assign \piso.data_r [926] = \piso.data_r_926_sv2v_reg ;
  assign \piso.data_r [925] = \piso.data_r_925_sv2v_reg ;
  assign \piso.data_r [924] = \piso.data_r_924_sv2v_reg ;
  assign \piso.data_r [923] = \piso.data_r_923_sv2v_reg ;
  assign \piso.data_r [922] = \piso.data_r_922_sv2v_reg ;
  assign \piso.data_r [921] = \piso.data_r_921_sv2v_reg ;
  assign \piso.data_r [920] = \piso.data_r_920_sv2v_reg ;
  assign \piso.data_r [919] = \piso.data_r_919_sv2v_reg ;
  assign \piso.data_r [918] = \piso.data_r_918_sv2v_reg ;
  assign \piso.data_r [917] = \piso.data_r_917_sv2v_reg ;
  assign \piso.data_r [916] = \piso.data_r_916_sv2v_reg ;
  assign \piso.data_r [915] = \piso.data_r_915_sv2v_reg ;
  assign \piso.data_r [914] = \piso.data_r_914_sv2v_reg ;
  assign \piso.data_r [913] = \piso.data_r_913_sv2v_reg ;
  assign \piso.data_r [912] = \piso.data_r_912_sv2v_reg ;
  assign \piso.data_r [911] = \piso.data_r_911_sv2v_reg ;
  assign \piso.data_r [910] = \piso.data_r_910_sv2v_reg ;
  assign \piso.data_r [909] = \piso.data_r_909_sv2v_reg ;
  assign \piso.data_r [908] = \piso.data_r_908_sv2v_reg ;
  assign \piso.data_r [907] = \piso.data_r_907_sv2v_reg ;
  assign \piso.data_r [906] = \piso.data_r_906_sv2v_reg ;
  assign \piso.data_r [905] = \piso.data_r_905_sv2v_reg ;
  assign \piso.data_r [904] = \piso.data_r_904_sv2v_reg ;
  assign \piso.data_r [903] = \piso.data_r_903_sv2v_reg ;
  assign \piso.data_r [902] = \piso.data_r_902_sv2v_reg ;
  assign \piso.data_r [901] = \piso.data_r_901_sv2v_reg ;
  assign \piso.data_r [900] = \piso.data_r_900_sv2v_reg ;
  assign \piso.data_r [899] = \piso.data_r_899_sv2v_reg ;
  assign \piso.data_r [898] = \piso.data_r_898_sv2v_reg ;
  assign \piso.data_r [897] = \piso.data_r_897_sv2v_reg ;
  assign \piso.data_r [896] = \piso.data_r_896_sv2v_reg ;
  assign \piso.data_r [895] = \piso.data_r_895_sv2v_reg ;
  assign \piso.data_r [894] = \piso.data_r_894_sv2v_reg ;
  assign \piso.data_r [893] = \piso.data_r_893_sv2v_reg ;
  assign \piso.data_r [892] = \piso.data_r_892_sv2v_reg ;
  assign \piso.data_r [891] = \piso.data_r_891_sv2v_reg ;
  assign \piso.data_r [890] = \piso.data_r_890_sv2v_reg ;
  assign \piso.data_r [889] = \piso.data_r_889_sv2v_reg ;
  assign \piso.data_r [888] = \piso.data_r_888_sv2v_reg ;
  assign \piso.data_r [887] = \piso.data_r_887_sv2v_reg ;
  assign \piso.data_r [886] = \piso.data_r_886_sv2v_reg ;
  assign \piso.data_r [885] = \piso.data_r_885_sv2v_reg ;
  assign \piso.data_r [884] = \piso.data_r_884_sv2v_reg ;
  assign \piso.data_r [883] = \piso.data_r_883_sv2v_reg ;
  assign \piso.data_r [882] = \piso.data_r_882_sv2v_reg ;
  assign \piso.data_r [881] = \piso.data_r_881_sv2v_reg ;
  assign \piso.data_r [880] = \piso.data_r_880_sv2v_reg ;
  assign \piso.data_r [879] = \piso.data_r_879_sv2v_reg ;
  assign \piso.data_r [878] = \piso.data_r_878_sv2v_reg ;
  assign \piso.data_r [877] = \piso.data_r_877_sv2v_reg ;
  assign \piso.data_r [876] = \piso.data_r_876_sv2v_reg ;
  assign \piso.data_r [875] = \piso.data_r_875_sv2v_reg ;
  assign \piso.data_r [874] = \piso.data_r_874_sv2v_reg ;
  assign \piso.data_r [873] = \piso.data_r_873_sv2v_reg ;
  assign \piso.data_r [872] = \piso.data_r_872_sv2v_reg ;
  assign \piso.data_r [871] = \piso.data_r_871_sv2v_reg ;
  assign \piso.data_r [870] = \piso.data_r_870_sv2v_reg ;
  assign \piso.data_r [869] = \piso.data_r_869_sv2v_reg ;
  assign \piso.data_r [868] = \piso.data_r_868_sv2v_reg ;
  assign \piso.data_r [867] = \piso.data_r_867_sv2v_reg ;
  assign \piso.data_r [866] = \piso.data_r_866_sv2v_reg ;
  assign \piso.data_r [865] = \piso.data_r_865_sv2v_reg ;
  assign \piso.data_r [864] = \piso.data_r_864_sv2v_reg ;
  assign \piso.data_r [863] = \piso.data_r_863_sv2v_reg ;
  assign \piso.data_r [862] = \piso.data_r_862_sv2v_reg ;
  assign \piso.data_r [861] = \piso.data_r_861_sv2v_reg ;
  assign \piso.data_r [860] = \piso.data_r_860_sv2v_reg ;
  assign \piso.data_r [859] = \piso.data_r_859_sv2v_reg ;
  assign \piso.data_r [858] = \piso.data_r_858_sv2v_reg ;
  assign \piso.data_r [857] = \piso.data_r_857_sv2v_reg ;
  assign \piso.data_r [856] = \piso.data_r_856_sv2v_reg ;
  assign \piso.data_r [855] = \piso.data_r_855_sv2v_reg ;
  assign \piso.data_r [854] = \piso.data_r_854_sv2v_reg ;
  assign \piso.data_r [853] = \piso.data_r_853_sv2v_reg ;
  assign \piso.data_r [852] = \piso.data_r_852_sv2v_reg ;
  assign \piso.data_r [851] = \piso.data_r_851_sv2v_reg ;
  assign \piso.data_r [850] = \piso.data_r_850_sv2v_reg ;
  assign \piso.data_r [849] = \piso.data_r_849_sv2v_reg ;
  assign \piso.data_r [848] = \piso.data_r_848_sv2v_reg ;
  assign \piso.data_r [847] = \piso.data_r_847_sv2v_reg ;
  assign \piso.data_r [846] = \piso.data_r_846_sv2v_reg ;
  assign \piso.data_r [845] = \piso.data_r_845_sv2v_reg ;
  assign \piso.data_r [844] = \piso.data_r_844_sv2v_reg ;
  assign \piso.data_r [843] = \piso.data_r_843_sv2v_reg ;
  assign \piso.data_r [842] = \piso.data_r_842_sv2v_reg ;
  assign \piso.data_r [841] = \piso.data_r_841_sv2v_reg ;
  assign \piso.data_r [840] = \piso.data_r_840_sv2v_reg ;
  assign \piso.data_r [839] = \piso.data_r_839_sv2v_reg ;
  assign \piso.data_r [838] = \piso.data_r_838_sv2v_reg ;
  assign \piso.data_r [837] = \piso.data_r_837_sv2v_reg ;
  assign \piso.data_r [836] = \piso.data_r_836_sv2v_reg ;
  assign \piso.data_r [835] = \piso.data_r_835_sv2v_reg ;
  assign \piso.data_r [834] = \piso.data_r_834_sv2v_reg ;
  assign \piso.data_r [833] = \piso.data_r_833_sv2v_reg ;
  assign \piso.data_r [832] = \piso.data_r_832_sv2v_reg ;
  assign \piso.data_r [831] = \piso.data_r_831_sv2v_reg ;
  assign \piso.data_r [830] = \piso.data_r_830_sv2v_reg ;
  assign \piso.data_r [829] = \piso.data_r_829_sv2v_reg ;
  assign \piso.data_r [828] = \piso.data_r_828_sv2v_reg ;
  assign \piso.data_r [827] = \piso.data_r_827_sv2v_reg ;
  assign \piso.data_r [826] = \piso.data_r_826_sv2v_reg ;
  assign \piso.data_r [825] = \piso.data_r_825_sv2v_reg ;
  assign \piso.data_r [824] = \piso.data_r_824_sv2v_reg ;
  assign \piso.data_r [823] = \piso.data_r_823_sv2v_reg ;
  assign \piso.data_r [822] = \piso.data_r_822_sv2v_reg ;
  assign \piso.data_r [821] = \piso.data_r_821_sv2v_reg ;
  assign \piso.data_r [820] = \piso.data_r_820_sv2v_reg ;
  assign \piso.data_r [819] = \piso.data_r_819_sv2v_reg ;
  assign \piso.data_r [818] = \piso.data_r_818_sv2v_reg ;
  assign \piso.data_r [817] = \piso.data_r_817_sv2v_reg ;
  assign \piso.data_r [816] = \piso.data_r_816_sv2v_reg ;
  assign \piso.data_r [815] = \piso.data_r_815_sv2v_reg ;
  assign \piso.data_r [814] = \piso.data_r_814_sv2v_reg ;
  assign \piso.data_r [813] = \piso.data_r_813_sv2v_reg ;
  assign \piso.data_r [812] = \piso.data_r_812_sv2v_reg ;
  assign \piso.data_r [811] = \piso.data_r_811_sv2v_reg ;
  assign \piso.data_r [810] = \piso.data_r_810_sv2v_reg ;
  assign \piso.data_r [809] = \piso.data_r_809_sv2v_reg ;
  assign \piso.data_r [808] = \piso.data_r_808_sv2v_reg ;
  assign \piso.data_r [807] = \piso.data_r_807_sv2v_reg ;
  assign \piso.data_r [806] = \piso.data_r_806_sv2v_reg ;
  assign \piso.data_r [805] = \piso.data_r_805_sv2v_reg ;
  assign \piso.data_r [804] = \piso.data_r_804_sv2v_reg ;
  assign \piso.data_r [803] = \piso.data_r_803_sv2v_reg ;
  assign \piso.data_r [802] = \piso.data_r_802_sv2v_reg ;
  assign \piso.data_r [801] = \piso.data_r_801_sv2v_reg ;
  assign \piso.data_r [800] = \piso.data_r_800_sv2v_reg ;
  assign \piso.data_r [799] = \piso.data_r_799_sv2v_reg ;
  assign \piso.data_r [798] = \piso.data_r_798_sv2v_reg ;
  assign \piso.data_r [797] = \piso.data_r_797_sv2v_reg ;
  assign \piso.data_r [796] = \piso.data_r_796_sv2v_reg ;
  assign \piso.data_r [795] = \piso.data_r_795_sv2v_reg ;
  assign \piso.data_r [794] = \piso.data_r_794_sv2v_reg ;
  assign \piso.data_r [793] = \piso.data_r_793_sv2v_reg ;
  assign \piso.data_r [792] = \piso.data_r_792_sv2v_reg ;
  assign \piso.data_r [791] = \piso.data_r_791_sv2v_reg ;
  assign \piso.data_r [790] = \piso.data_r_790_sv2v_reg ;
  assign \piso.data_r [789] = \piso.data_r_789_sv2v_reg ;
  assign \piso.data_r [788] = \piso.data_r_788_sv2v_reg ;
  assign \piso.data_r [787] = \piso.data_r_787_sv2v_reg ;
  assign \piso.data_r [786] = \piso.data_r_786_sv2v_reg ;
  assign \piso.data_r [785] = \piso.data_r_785_sv2v_reg ;
  assign \piso.data_r [784] = \piso.data_r_784_sv2v_reg ;
  assign \piso.data_r [783] = \piso.data_r_783_sv2v_reg ;
  assign \piso.data_r [782] = \piso.data_r_782_sv2v_reg ;
  assign \piso.data_r [781] = \piso.data_r_781_sv2v_reg ;
  assign \piso.data_r [780] = \piso.data_r_780_sv2v_reg ;
  assign \piso.data_r [779] = \piso.data_r_779_sv2v_reg ;
  assign \piso.data_r [778] = \piso.data_r_778_sv2v_reg ;
  assign \piso.data_r [777] = \piso.data_r_777_sv2v_reg ;
  assign \piso.data_r [776] = \piso.data_r_776_sv2v_reg ;
  assign \piso.data_r [775] = \piso.data_r_775_sv2v_reg ;
  assign \piso.data_r [774] = \piso.data_r_774_sv2v_reg ;
  assign \piso.data_r [773] = \piso.data_r_773_sv2v_reg ;
  assign \piso.data_r [772] = \piso.data_r_772_sv2v_reg ;
  assign \piso.data_r [771] = \piso.data_r_771_sv2v_reg ;
  assign \piso.data_r [770] = \piso.data_r_770_sv2v_reg ;
  assign \piso.data_r [769] = \piso.data_r_769_sv2v_reg ;
  assign \piso.data_r [768] = \piso.data_r_768_sv2v_reg ;
  assign \piso.data_r [767] = \piso.data_r_767_sv2v_reg ;
  assign \piso.data_r [766] = \piso.data_r_766_sv2v_reg ;
  assign \piso.data_r [765] = \piso.data_r_765_sv2v_reg ;
  assign \piso.data_r [764] = \piso.data_r_764_sv2v_reg ;
  assign \piso.data_r [763] = \piso.data_r_763_sv2v_reg ;
  assign \piso.data_r [762] = \piso.data_r_762_sv2v_reg ;
  assign \piso.data_r [761] = \piso.data_r_761_sv2v_reg ;
  assign \piso.data_r [760] = \piso.data_r_760_sv2v_reg ;
  assign \piso.data_r [759] = \piso.data_r_759_sv2v_reg ;
  assign \piso.data_r [758] = \piso.data_r_758_sv2v_reg ;
  assign \piso.data_r [757] = \piso.data_r_757_sv2v_reg ;
  assign \piso.data_r [756] = \piso.data_r_756_sv2v_reg ;
  assign \piso.data_r [755] = \piso.data_r_755_sv2v_reg ;
  assign \piso.data_r [754] = \piso.data_r_754_sv2v_reg ;
  assign \piso.data_r [753] = \piso.data_r_753_sv2v_reg ;
  assign \piso.data_r [752] = \piso.data_r_752_sv2v_reg ;
  assign \piso.data_r [751] = \piso.data_r_751_sv2v_reg ;
  assign \piso.data_r [750] = \piso.data_r_750_sv2v_reg ;
  assign \piso.data_r [749] = \piso.data_r_749_sv2v_reg ;
  assign \piso.data_r [748] = \piso.data_r_748_sv2v_reg ;
  assign \piso.data_r [747] = \piso.data_r_747_sv2v_reg ;
  assign \piso.data_r [746] = \piso.data_r_746_sv2v_reg ;
  assign \piso.data_r [745] = \piso.data_r_745_sv2v_reg ;
  assign \piso.data_r [744] = \piso.data_r_744_sv2v_reg ;
  assign \piso.data_r [743] = \piso.data_r_743_sv2v_reg ;
  assign \piso.data_r [742] = \piso.data_r_742_sv2v_reg ;
  assign \piso.data_r [741] = \piso.data_r_741_sv2v_reg ;
  assign \piso.data_r [740] = \piso.data_r_740_sv2v_reg ;
  assign \piso.data_r [739] = \piso.data_r_739_sv2v_reg ;
  assign \piso.data_r [738] = \piso.data_r_738_sv2v_reg ;
  assign \piso.data_r [737] = \piso.data_r_737_sv2v_reg ;
  assign \piso.data_r [736] = \piso.data_r_736_sv2v_reg ;
  assign \piso.data_r [735] = \piso.data_r_735_sv2v_reg ;
  assign \piso.data_r [734] = \piso.data_r_734_sv2v_reg ;
  assign \piso.data_r [733] = \piso.data_r_733_sv2v_reg ;
  assign \piso.data_r [732] = \piso.data_r_732_sv2v_reg ;
  assign \piso.data_r [731] = \piso.data_r_731_sv2v_reg ;
  assign \piso.data_r [730] = \piso.data_r_730_sv2v_reg ;
  assign \piso.data_r [729] = \piso.data_r_729_sv2v_reg ;
  assign \piso.data_r [728] = \piso.data_r_728_sv2v_reg ;
  assign \piso.data_r [727] = \piso.data_r_727_sv2v_reg ;
  assign \piso.data_r [726] = \piso.data_r_726_sv2v_reg ;
  assign \piso.data_r [725] = \piso.data_r_725_sv2v_reg ;
  assign \piso.data_r [724] = \piso.data_r_724_sv2v_reg ;
  assign \piso.data_r [723] = \piso.data_r_723_sv2v_reg ;
  assign \piso.data_r [722] = \piso.data_r_722_sv2v_reg ;
  assign \piso.data_r [721] = \piso.data_r_721_sv2v_reg ;
  assign \piso.data_r [720] = \piso.data_r_720_sv2v_reg ;
  assign \piso.data_r [719] = \piso.data_r_719_sv2v_reg ;
  assign \piso.data_r [718] = \piso.data_r_718_sv2v_reg ;
  assign \piso.data_r [717] = \piso.data_r_717_sv2v_reg ;
  assign \piso.data_r [716] = \piso.data_r_716_sv2v_reg ;
  assign \piso.data_r [715] = \piso.data_r_715_sv2v_reg ;
  assign \piso.data_r [714] = \piso.data_r_714_sv2v_reg ;
  assign \piso.data_r [713] = \piso.data_r_713_sv2v_reg ;
  assign \piso.data_r [712] = \piso.data_r_712_sv2v_reg ;
  assign \piso.data_r [711] = \piso.data_r_711_sv2v_reg ;
  assign \piso.data_r [710] = \piso.data_r_710_sv2v_reg ;
  assign \piso.data_r [709] = \piso.data_r_709_sv2v_reg ;
  assign \piso.data_r [708] = \piso.data_r_708_sv2v_reg ;
  assign \piso.data_r [707] = \piso.data_r_707_sv2v_reg ;
  assign \piso.data_r [706] = \piso.data_r_706_sv2v_reg ;
  assign \piso.data_r [705] = \piso.data_r_705_sv2v_reg ;
  assign \piso.data_r [704] = \piso.data_r_704_sv2v_reg ;
  assign \piso.data_r [703] = \piso.data_r_703_sv2v_reg ;
  assign \piso.data_r [702] = \piso.data_r_702_sv2v_reg ;
  assign \piso.data_r [701] = \piso.data_r_701_sv2v_reg ;
  assign \piso.data_r [700] = \piso.data_r_700_sv2v_reg ;
  assign \piso.data_r [699] = \piso.data_r_699_sv2v_reg ;
  assign \piso.data_r [698] = \piso.data_r_698_sv2v_reg ;
  assign \piso.data_r [697] = \piso.data_r_697_sv2v_reg ;
  assign \piso.data_r [696] = \piso.data_r_696_sv2v_reg ;
  assign \piso.data_r [695] = \piso.data_r_695_sv2v_reg ;
  assign \piso.data_r [694] = \piso.data_r_694_sv2v_reg ;
  assign \piso.data_r [693] = \piso.data_r_693_sv2v_reg ;
  assign \piso.data_r [692] = \piso.data_r_692_sv2v_reg ;
  assign \piso.data_r [691] = \piso.data_r_691_sv2v_reg ;
  assign \piso.data_r [690] = \piso.data_r_690_sv2v_reg ;
  assign \piso.data_r [689] = \piso.data_r_689_sv2v_reg ;
  assign \piso.data_r [688] = \piso.data_r_688_sv2v_reg ;
  assign \piso.data_r [687] = \piso.data_r_687_sv2v_reg ;
  assign \piso.data_r [686] = \piso.data_r_686_sv2v_reg ;
  assign \piso.data_r [685] = \piso.data_r_685_sv2v_reg ;
  assign \piso.data_r [684] = \piso.data_r_684_sv2v_reg ;
  assign \piso.data_r [683] = \piso.data_r_683_sv2v_reg ;
  assign \piso.data_r [682] = \piso.data_r_682_sv2v_reg ;
  assign \piso.data_r [681] = \piso.data_r_681_sv2v_reg ;
  assign \piso.data_r [680] = \piso.data_r_680_sv2v_reg ;
  assign \piso.data_r [679] = \piso.data_r_679_sv2v_reg ;
  assign \piso.data_r [678] = \piso.data_r_678_sv2v_reg ;
  assign \piso.data_r [677] = \piso.data_r_677_sv2v_reg ;
  assign \piso.data_r [676] = \piso.data_r_676_sv2v_reg ;
  assign \piso.data_r [675] = \piso.data_r_675_sv2v_reg ;
  assign \piso.data_r [674] = \piso.data_r_674_sv2v_reg ;
  assign \piso.data_r [673] = \piso.data_r_673_sv2v_reg ;
  assign \piso.data_r [672] = \piso.data_r_672_sv2v_reg ;
  assign \piso.data_r [671] = \piso.data_r_671_sv2v_reg ;
  assign \piso.data_r [670] = \piso.data_r_670_sv2v_reg ;
  assign \piso.data_r [669] = \piso.data_r_669_sv2v_reg ;
  assign \piso.data_r [668] = \piso.data_r_668_sv2v_reg ;
  assign \piso.data_r [667] = \piso.data_r_667_sv2v_reg ;
  assign \piso.data_r [666] = \piso.data_r_666_sv2v_reg ;
  assign \piso.data_r [665] = \piso.data_r_665_sv2v_reg ;
  assign \piso.data_r [664] = \piso.data_r_664_sv2v_reg ;
  assign \piso.data_r [663] = \piso.data_r_663_sv2v_reg ;
  assign \piso.data_r [662] = \piso.data_r_662_sv2v_reg ;
  assign \piso.data_r [661] = \piso.data_r_661_sv2v_reg ;
  assign \piso.data_r [660] = \piso.data_r_660_sv2v_reg ;
  assign \piso.data_r [659] = \piso.data_r_659_sv2v_reg ;
  assign \piso.data_r [658] = \piso.data_r_658_sv2v_reg ;
  assign \piso.data_r [657] = \piso.data_r_657_sv2v_reg ;
  assign \piso.data_r [656] = \piso.data_r_656_sv2v_reg ;
  assign \piso.data_r [655] = \piso.data_r_655_sv2v_reg ;
  assign \piso.data_r [654] = \piso.data_r_654_sv2v_reg ;
  assign \piso.data_r [653] = \piso.data_r_653_sv2v_reg ;
  assign \piso.data_r [652] = \piso.data_r_652_sv2v_reg ;
  assign \piso.data_r [651] = \piso.data_r_651_sv2v_reg ;
  assign \piso.data_r [650] = \piso.data_r_650_sv2v_reg ;
  assign \piso.data_r [649] = \piso.data_r_649_sv2v_reg ;
  assign \piso.data_r [648] = \piso.data_r_648_sv2v_reg ;
  assign \piso.data_r [647] = \piso.data_r_647_sv2v_reg ;
  assign \piso.data_r [646] = \piso.data_r_646_sv2v_reg ;
  assign \piso.data_r [645] = \piso.data_r_645_sv2v_reg ;
  assign \piso.data_r [644] = \piso.data_r_644_sv2v_reg ;
  assign \piso.data_r [643] = \piso.data_r_643_sv2v_reg ;
  assign \piso.data_r [642] = \piso.data_r_642_sv2v_reg ;
  assign \piso.data_r [641] = \piso.data_r_641_sv2v_reg ;
  assign \piso.data_r [640] = \piso.data_r_640_sv2v_reg ;
  assign \piso.data_r [639] = \piso.data_r_639_sv2v_reg ;
  assign \piso.data_r [638] = \piso.data_r_638_sv2v_reg ;
  assign \piso.data_r [637] = \piso.data_r_637_sv2v_reg ;
  assign \piso.data_r [636] = \piso.data_r_636_sv2v_reg ;
  assign \piso.data_r [635] = \piso.data_r_635_sv2v_reg ;
  assign \piso.data_r [634] = \piso.data_r_634_sv2v_reg ;
  assign \piso.data_r [633] = \piso.data_r_633_sv2v_reg ;
  assign \piso.data_r [632] = \piso.data_r_632_sv2v_reg ;
  assign \piso.data_r [631] = \piso.data_r_631_sv2v_reg ;
  assign \piso.data_r [630] = \piso.data_r_630_sv2v_reg ;
  assign \piso.data_r [629] = \piso.data_r_629_sv2v_reg ;
  assign \piso.data_r [628] = \piso.data_r_628_sv2v_reg ;
  assign \piso.data_r [627] = \piso.data_r_627_sv2v_reg ;
  assign \piso.data_r [626] = \piso.data_r_626_sv2v_reg ;
  assign \piso.data_r [625] = \piso.data_r_625_sv2v_reg ;
  assign \piso.data_r [624] = \piso.data_r_624_sv2v_reg ;
  assign \piso.data_r [623] = \piso.data_r_623_sv2v_reg ;
  assign \piso.data_r [622] = \piso.data_r_622_sv2v_reg ;
  assign \piso.data_r [621] = \piso.data_r_621_sv2v_reg ;
  assign \piso.data_r [620] = \piso.data_r_620_sv2v_reg ;
  assign \piso.data_r [619] = \piso.data_r_619_sv2v_reg ;
  assign \piso.data_r [618] = \piso.data_r_618_sv2v_reg ;
  assign \piso.data_r [617] = \piso.data_r_617_sv2v_reg ;
  assign \piso.data_r [616] = \piso.data_r_616_sv2v_reg ;
  assign \piso.data_r [615] = \piso.data_r_615_sv2v_reg ;
  assign \piso.data_r [614] = \piso.data_r_614_sv2v_reg ;
  assign \piso.data_r [613] = \piso.data_r_613_sv2v_reg ;
  assign \piso.data_r [612] = \piso.data_r_612_sv2v_reg ;
  assign \piso.data_r [611] = \piso.data_r_611_sv2v_reg ;
  assign \piso.data_r [610] = \piso.data_r_610_sv2v_reg ;
  assign \piso.data_r [609] = \piso.data_r_609_sv2v_reg ;
  assign \piso.data_r [608] = \piso.data_r_608_sv2v_reg ;
  assign \piso.data_r [607] = \piso.data_r_607_sv2v_reg ;
  assign \piso.data_r [606] = \piso.data_r_606_sv2v_reg ;
  assign \piso.data_r [605] = \piso.data_r_605_sv2v_reg ;
  assign \piso.data_r [604] = \piso.data_r_604_sv2v_reg ;
  assign \piso.data_r [603] = \piso.data_r_603_sv2v_reg ;
  assign \piso.data_r [602] = \piso.data_r_602_sv2v_reg ;
  assign \piso.data_r [601] = \piso.data_r_601_sv2v_reg ;
  assign \piso.data_r [600] = \piso.data_r_600_sv2v_reg ;
  assign \piso.data_r [599] = \piso.data_r_599_sv2v_reg ;
  assign \piso.data_r [598] = \piso.data_r_598_sv2v_reg ;
  assign \piso.data_r [597] = \piso.data_r_597_sv2v_reg ;
  assign \piso.data_r [596] = \piso.data_r_596_sv2v_reg ;
  assign \piso.data_r [595] = \piso.data_r_595_sv2v_reg ;
  assign \piso.data_r [594] = \piso.data_r_594_sv2v_reg ;
  assign \piso.data_r [593] = \piso.data_r_593_sv2v_reg ;
  assign \piso.data_r [592] = \piso.data_r_592_sv2v_reg ;
  assign \piso.data_r [591] = \piso.data_r_591_sv2v_reg ;
  assign \piso.data_r [590] = \piso.data_r_590_sv2v_reg ;
  assign \piso.data_r [589] = \piso.data_r_589_sv2v_reg ;
  assign \piso.data_r [588] = \piso.data_r_588_sv2v_reg ;
  assign \piso.data_r [587] = \piso.data_r_587_sv2v_reg ;
  assign \piso.data_r [586] = \piso.data_r_586_sv2v_reg ;
  assign \piso.data_r [585] = \piso.data_r_585_sv2v_reg ;
  assign \piso.data_r [584] = \piso.data_r_584_sv2v_reg ;
  assign \piso.data_r [583] = \piso.data_r_583_sv2v_reg ;
  assign \piso.data_r [582] = \piso.data_r_582_sv2v_reg ;
  assign \piso.data_r [581] = \piso.data_r_581_sv2v_reg ;
  assign \piso.data_r [580] = \piso.data_r_580_sv2v_reg ;
  assign \piso.data_r [579] = \piso.data_r_579_sv2v_reg ;
  assign \piso.data_r [578] = \piso.data_r_578_sv2v_reg ;
  assign \piso.data_r [577] = \piso.data_r_577_sv2v_reg ;
  assign \piso.data_r [576] = \piso.data_r_576_sv2v_reg ;
  assign \piso.data_r [575] = \piso.data_r_575_sv2v_reg ;
  assign \piso.data_r [574] = \piso.data_r_574_sv2v_reg ;
  assign \piso.data_r [573] = \piso.data_r_573_sv2v_reg ;
  assign \piso.data_r [572] = \piso.data_r_572_sv2v_reg ;
  assign \piso.data_r [571] = \piso.data_r_571_sv2v_reg ;
  assign \piso.data_r [570] = \piso.data_r_570_sv2v_reg ;
  assign \piso.data_r [569] = \piso.data_r_569_sv2v_reg ;
  assign \piso.data_r [568] = \piso.data_r_568_sv2v_reg ;
  assign \piso.data_r [567] = \piso.data_r_567_sv2v_reg ;
  assign \piso.data_r [566] = \piso.data_r_566_sv2v_reg ;
  assign \piso.data_r [565] = \piso.data_r_565_sv2v_reg ;
  assign \piso.data_r [564] = \piso.data_r_564_sv2v_reg ;
  assign \piso.data_r [563] = \piso.data_r_563_sv2v_reg ;
  assign \piso.data_r [562] = \piso.data_r_562_sv2v_reg ;
  assign \piso.data_r [561] = \piso.data_r_561_sv2v_reg ;
  assign \piso.data_r [560] = \piso.data_r_560_sv2v_reg ;
  assign \piso.data_r [559] = \piso.data_r_559_sv2v_reg ;
  assign \piso.data_r [558] = \piso.data_r_558_sv2v_reg ;
  assign \piso.data_r [557] = \piso.data_r_557_sv2v_reg ;
  assign \piso.data_r [556] = \piso.data_r_556_sv2v_reg ;
  assign \piso.data_r [555] = \piso.data_r_555_sv2v_reg ;
  assign \piso.data_r [554] = \piso.data_r_554_sv2v_reg ;
  assign \piso.data_r [553] = \piso.data_r_553_sv2v_reg ;
  assign \piso.data_r [552] = \piso.data_r_552_sv2v_reg ;
  assign \piso.data_r [551] = \piso.data_r_551_sv2v_reg ;
  assign \piso.data_r [550] = \piso.data_r_550_sv2v_reg ;
  assign \piso.data_r [549] = \piso.data_r_549_sv2v_reg ;
  assign \piso.data_r [548] = \piso.data_r_548_sv2v_reg ;
  assign \piso.data_r [547] = \piso.data_r_547_sv2v_reg ;
  assign \piso.data_r [546] = \piso.data_r_546_sv2v_reg ;
  assign \piso.data_r [545] = \piso.data_r_545_sv2v_reg ;
  assign \piso.data_r [544] = \piso.data_r_544_sv2v_reg ;
  assign \piso.data_r [543] = \piso.data_r_543_sv2v_reg ;
  assign \piso.data_r [542] = \piso.data_r_542_sv2v_reg ;
  assign \piso.data_r [541] = \piso.data_r_541_sv2v_reg ;
  assign \piso.data_r [540] = \piso.data_r_540_sv2v_reg ;
  assign \piso.data_r [539] = \piso.data_r_539_sv2v_reg ;
  assign \piso.data_r [538] = \piso.data_r_538_sv2v_reg ;
  assign \piso.data_r [537] = \piso.data_r_537_sv2v_reg ;
  assign \piso.data_r [536] = \piso.data_r_536_sv2v_reg ;
  assign \piso.data_r [535] = \piso.data_r_535_sv2v_reg ;
  assign \piso.data_r [534] = \piso.data_r_534_sv2v_reg ;
  assign \piso.data_r [533] = \piso.data_r_533_sv2v_reg ;
  assign \piso.data_r [532] = \piso.data_r_532_sv2v_reg ;
  assign \piso.data_r [531] = \piso.data_r_531_sv2v_reg ;
  assign \piso.data_r [530] = \piso.data_r_530_sv2v_reg ;
  assign \piso.data_r [529] = \piso.data_r_529_sv2v_reg ;
  assign \piso.data_r [528] = \piso.data_r_528_sv2v_reg ;
  assign \piso.data_r [527] = \piso.data_r_527_sv2v_reg ;
  assign \piso.data_r [526] = \piso.data_r_526_sv2v_reg ;
  assign \piso.data_r [525] = \piso.data_r_525_sv2v_reg ;
  assign \piso.data_r [524] = \piso.data_r_524_sv2v_reg ;
  assign \piso.data_r [523] = \piso.data_r_523_sv2v_reg ;
  assign \piso.data_r [522] = \piso.data_r_522_sv2v_reg ;
  assign \piso.data_r [521] = \piso.data_r_521_sv2v_reg ;
  assign \piso.data_r [520] = \piso.data_r_520_sv2v_reg ;
  assign \piso.data_r [519] = \piso.data_r_519_sv2v_reg ;
  assign \piso.data_r [518] = \piso.data_r_518_sv2v_reg ;
  assign \piso.data_r [517] = \piso.data_r_517_sv2v_reg ;
  assign \piso.data_r [516] = \piso.data_r_516_sv2v_reg ;
  assign \piso.data_r [515] = \piso.data_r_515_sv2v_reg ;
  assign \piso.data_r [514] = \piso.data_r_514_sv2v_reg ;
  assign \piso.data_r [513] = \piso.data_r_513_sv2v_reg ;
  assign \piso.data_r [512] = \piso.data_r_512_sv2v_reg ;
  assign \piso.data_r [511] = \piso.data_r_511_sv2v_reg ;
  assign \piso.data_r [510] = \piso.data_r_510_sv2v_reg ;
  assign \piso.data_r [509] = \piso.data_r_509_sv2v_reg ;
  assign \piso.data_r [508] = \piso.data_r_508_sv2v_reg ;
  assign \piso.data_r [507] = \piso.data_r_507_sv2v_reg ;
  assign \piso.data_r [506] = \piso.data_r_506_sv2v_reg ;
  assign \piso.data_r [505] = \piso.data_r_505_sv2v_reg ;
  assign \piso.data_r [504] = \piso.data_r_504_sv2v_reg ;
  assign \piso.data_r [503] = \piso.data_r_503_sv2v_reg ;
  assign \piso.data_r [502] = \piso.data_r_502_sv2v_reg ;
  assign \piso.data_r [501] = \piso.data_r_501_sv2v_reg ;
  assign \piso.data_r [500] = \piso.data_r_500_sv2v_reg ;
  assign \piso.data_r [499] = \piso.data_r_499_sv2v_reg ;
  assign \piso.data_r [498] = \piso.data_r_498_sv2v_reg ;
  assign \piso.data_r [497] = \piso.data_r_497_sv2v_reg ;
  assign \piso.data_r [496] = \piso.data_r_496_sv2v_reg ;
  assign \piso.data_r [495] = \piso.data_r_495_sv2v_reg ;
  assign \piso.data_r [494] = \piso.data_r_494_sv2v_reg ;
  assign \piso.data_r [493] = \piso.data_r_493_sv2v_reg ;
  assign \piso.data_r [492] = \piso.data_r_492_sv2v_reg ;
  assign \piso.data_r [491] = \piso.data_r_491_sv2v_reg ;
  assign \piso.data_r [490] = \piso.data_r_490_sv2v_reg ;
  assign \piso.data_r [489] = \piso.data_r_489_sv2v_reg ;
  assign \piso.data_r [488] = \piso.data_r_488_sv2v_reg ;
  assign \piso.data_r [487] = \piso.data_r_487_sv2v_reg ;
  assign \piso.data_r [486] = \piso.data_r_486_sv2v_reg ;
  assign \piso.data_r [485] = \piso.data_r_485_sv2v_reg ;
  assign \piso.data_r [484] = \piso.data_r_484_sv2v_reg ;
  assign \piso.data_r [483] = \piso.data_r_483_sv2v_reg ;
  assign \piso.data_r [482] = \piso.data_r_482_sv2v_reg ;
  assign \piso.data_r [481] = \piso.data_r_481_sv2v_reg ;
  assign \piso.data_r [480] = \piso.data_r_480_sv2v_reg ;
  assign \piso.data_r [479] = \piso.data_r_479_sv2v_reg ;
  assign \piso.data_r [478] = \piso.data_r_478_sv2v_reg ;
  assign \piso.data_r [477] = \piso.data_r_477_sv2v_reg ;
  assign \piso.data_r [476] = \piso.data_r_476_sv2v_reg ;
  assign \piso.data_r [475] = \piso.data_r_475_sv2v_reg ;
  assign \piso.data_r [474] = \piso.data_r_474_sv2v_reg ;
  assign \piso.data_r [473] = \piso.data_r_473_sv2v_reg ;
  assign \piso.data_r [472] = \piso.data_r_472_sv2v_reg ;
  assign \piso.data_r [471] = \piso.data_r_471_sv2v_reg ;
  assign \piso.data_r [470] = \piso.data_r_470_sv2v_reg ;
  assign \piso.data_r [469] = \piso.data_r_469_sv2v_reg ;
  assign \piso.data_r [468] = \piso.data_r_468_sv2v_reg ;
  assign \piso.data_r [467] = \piso.data_r_467_sv2v_reg ;
  assign \piso.data_r [466] = \piso.data_r_466_sv2v_reg ;
  assign \piso.data_r [465] = \piso.data_r_465_sv2v_reg ;
  assign \piso.data_r [464] = \piso.data_r_464_sv2v_reg ;
  assign \piso.data_r [463] = \piso.data_r_463_sv2v_reg ;
  assign \piso.data_r [462] = \piso.data_r_462_sv2v_reg ;
  assign \piso.data_r [461] = \piso.data_r_461_sv2v_reg ;
  assign \piso.data_r [460] = \piso.data_r_460_sv2v_reg ;
  assign \piso.data_r [459] = \piso.data_r_459_sv2v_reg ;
  assign \piso.data_r [458] = \piso.data_r_458_sv2v_reg ;
  assign \piso.data_r [457] = \piso.data_r_457_sv2v_reg ;
  assign \piso.data_r [456] = \piso.data_r_456_sv2v_reg ;
  assign \piso.data_r [455] = \piso.data_r_455_sv2v_reg ;
  assign \piso.data_r [454] = \piso.data_r_454_sv2v_reg ;
  assign \piso.data_r [453] = \piso.data_r_453_sv2v_reg ;
  assign \piso.data_r [452] = \piso.data_r_452_sv2v_reg ;
  assign \piso.data_r [451] = \piso.data_r_451_sv2v_reg ;
  assign \piso.data_r [450] = \piso.data_r_450_sv2v_reg ;
  assign \piso.data_r [449] = \piso.data_r_449_sv2v_reg ;
  assign \piso.data_r [448] = \piso.data_r_448_sv2v_reg ;
  assign \piso.data_r [447] = \piso.data_r_447_sv2v_reg ;
  assign \piso.data_r [446] = \piso.data_r_446_sv2v_reg ;
  assign \piso.data_r [445] = \piso.data_r_445_sv2v_reg ;
  assign \piso.data_r [444] = \piso.data_r_444_sv2v_reg ;
  assign \piso.data_r [443] = \piso.data_r_443_sv2v_reg ;
  assign \piso.data_r [442] = \piso.data_r_442_sv2v_reg ;
  assign \piso.data_r [441] = \piso.data_r_441_sv2v_reg ;
  assign \piso.data_r [440] = \piso.data_r_440_sv2v_reg ;
  assign \piso.data_r [439] = \piso.data_r_439_sv2v_reg ;
  assign \piso.data_r [438] = \piso.data_r_438_sv2v_reg ;
  assign \piso.data_r [437] = \piso.data_r_437_sv2v_reg ;
  assign \piso.data_r [436] = \piso.data_r_436_sv2v_reg ;
  assign \piso.data_r [435] = \piso.data_r_435_sv2v_reg ;
  assign \piso.data_r [434] = \piso.data_r_434_sv2v_reg ;
  assign \piso.data_r [433] = \piso.data_r_433_sv2v_reg ;
  assign \piso.data_r [432] = \piso.data_r_432_sv2v_reg ;
  assign \piso.data_r [431] = \piso.data_r_431_sv2v_reg ;
  assign \piso.data_r [430] = \piso.data_r_430_sv2v_reg ;
  assign \piso.data_r [429] = \piso.data_r_429_sv2v_reg ;
  assign \piso.data_r [428] = \piso.data_r_428_sv2v_reg ;
  assign \piso.data_r [427] = \piso.data_r_427_sv2v_reg ;
  assign \piso.data_r [426] = \piso.data_r_426_sv2v_reg ;
  assign \piso.data_r [425] = \piso.data_r_425_sv2v_reg ;
  assign \piso.data_r [424] = \piso.data_r_424_sv2v_reg ;
  assign \piso.data_r [423] = \piso.data_r_423_sv2v_reg ;
  assign \piso.data_r [422] = \piso.data_r_422_sv2v_reg ;
  assign \piso.data_r [421] = \piso.data_r_421_sv2v_reg ;
  assign \piso.data_r [420] = \piso.data_r_420_sv2v_reg ;
  assign \piso.data_r [419] = \piso.data_r_419_sv2v_reg ;
  assign \piso.data_r [418] = \piso.data_r_418_sv2v_reg ;
  assign \piso.data_r [417] = \piso.data_r_417_sv2v_reg ;
  assign \piso.data_r [416] = \piso.data_r_416_sv2v_reg ;
  assign \piso.data_r [415] = \piso.data_r_415_sv2v_reg ;
  assign \piso.data_r [414] = \piso.data_r_414_sv2v_reg ;
  assign \piso.data_r [413] = \piso.data_r_413_sv2v_reg ;
  assign \piso.data_r [412] = \piso.data_r_412_sv2v_reg ;
  assign \piso.data_r [411] = \piso.data_r_411_sv2v_reg ;
  assign \piso.data_r [410] = \piso.data_r_410_sv2v_reg ;
  assign \piso.data_r [409] = \piso.data_r_409_sv2v_reg ;
  assign \piso.data_r [408] = \piso.data_r_408_sv2v_reg ;
  assign \piso.data_r [407] = \piso.data_r_407_sv2v_reg ;
  assign \piso.data_r [406] = \piso.data_r_406_sv2v_reg ;
  assign \piso.data_r [405] = \piso.data_r_405_sv2v_reg ;
  assign \piso.data_r [404] = \piso.data_r_404_sv2v_reg ;
  assign \piso.data_r [403] = \piso.data_r_403_sv2v_reg ;
  assign \piso.data_r [402] = \piso.data_r_402_sv2v_reg ;
  assign \piso.data_r [401] = \piso.data_r_401_sv2v_reg ;
  assign \piso.data_r [400] = \piso.data_r_400_sv2v_reg ;
  assign \piso.data_r [399] = \piso.data_r_399_sv2v_reg ;
  assign \piso.data_r [398] = \piso.data_r_398_sv2v_reg ;
  assign \piso.data_r [397] = \piso.data_r_397_sv2v_reg ;
  assign \piso.data_r [396] = \piso.data_r_396_sv2v_reg ;
  assign \piso.data_r [395] = \piso.data_r_395_sv2v_reg ;
  assign \piso.data_r [394] = \piso.data_r_394_sv2v_reg ;
  assign \piso.data_r [393] = \piso.data_r_393_sv2v_reg ;
  assign \piso.data_r [392] = \piso.data_r_392_sv2v_reg ;
  assign \piso.data_r [391] = \piso.data_r_391_sv2v_reg ;
  assign \piso.data_r [390] = \piso.data_r_390_sv2v_reg ;
  assign \piso.data_r [389] = \piso.data_r_389_sv2v_reg ;
  assign \piso.data_r [388] = \piso.data_r_388_sv2v_reg ;
  assign \piso.data_r [387] = \piso.data_r_387_sv2v_reg ;
  assign \piso.data_r [386] = \piso.data_r_386_sv2v_reg ;
  assign \piso.data_r [385] = \piso.data_r_385_sv2v_reg ;
  assign \piso.data_r [384] = \piso.data_r_384_sv2v_reg ;
  assign \piso.data_r [383] = \piso.data_r_383_sv2v_reg ;
  assign \piso.data_r [382] = \piso.data_r_382_sv2v_reg ;
  assign \piso.data_r [381] = \piso.data_r_381_sv2v_reg ;
  assign \piso.data_r [380] = \piso.data_r_380_sv2v_reg ;
  assign \piso.data_r [379] = \piso.data_r_379_sv2v_reg ;
  assign \piso.data_r [378] = \piso.data_r_378_sv2v_reg ;
  assign \piso.data_r [377] = \piso.data_r_377_sv2v_reg ;
  assign \piso.data_r [376] = \piso.data_r_376_sv2v_reg ;
  assign \piso.data_r [375] = \piso.data_r_375_sv2v_reg ;
  assign \piso.data_r [374] = \piso.data_r_374_sv2v_reg ;
  assign \piso.data_r [373] = \piso.data_r_373_sv2v_reg ;
  assign \piso.data_r [372] = \piso.data_r_372_sv2v_reg ;
  assign \piso.data_r [371] = \piso.data_r_371_sv2v_reg ;
  assign \piso.data_r [370] = \piso.data_r_370_sv2v_reg ;
  assign \piso.data_r [369] = \piso.data_r_369_sv2v_reg ;
  assign \piso.data_r [368] = \piso.data_r_368_sv2v_reg ;
  assign \piso.data_r [367] = \piso.data_r_367_sv2v_reg ;
  assign \piso.data_r [366] = \piso.data_r_366_sv2v_reg ;
  assign \piso.data_r [365] = \piso.data_r_365_sv2v_reg ;
  assign \piso.data_r [364] = \piso.data_r_364_sv2v_reg ;
  assign \piso.data_r [363] = \piso.data_r_363_sv2v_reg ;
  assign \piso.data_r [362] = \piso.data_r_362_sv2v_reg ;
  assign \piso.data_r [361] = \piso.data_r_361_sv2v_reg ;
  assign \piso.data_r [360] = \piso.data_r_360_sv2v_reg ;
  assign \piso.data_r [359] = \piso.data_r_359_sv2v_reg ;
  assign \piso.data_r [358] = \piso.data_r_358_sv2v_reg ;
  assign \piso.data_r [357] = \piso.data_r_357_sv2v_reg ;
  assign \piso.data_r [356] = \piso.data_r_356_sv2v_reg ;
  assign \piso.data_r [355] = \piso.data_r_355_sv2v_reg ;
  assign \piso.data_r [354] = \piso.data_r_354_sv2v_reg ;
  assign \piso.data_r [353] = \piso.data_r_353_sv2v_reg ;
  assign \piso.data_r [352] = \piso.data_r_352_sv2v_reg ;
  assign \piso.data_r [351] = \piso.data_r_351_sv2v_reg ;
  assign \piso.data_r [350] = \piso.data_r_350_sv2v_reg ;
  assign \piso.data_r [349] = \piso.data_r_349_sv2v_reg ;
  assign \piso.data_r [348] = \piso.data_r_348_sv2v_reg ;
  assign \piso.data_r [347] = \piso.data_r_347_sv2v_reg ;
  assign \piso.data_r [346] = \piso.data_r_346_sv2v_reg ;
  assign \piso.data_r [345] = \piso.data_r_345_sv2v_reg ;
  assign \piso.data_r [344] = \piso.data_r_344_sv2v_reg ;
  assign \piso.data_r [343] = \piso.data_r_343_sv2v_reg ;
  assign \piso.data_r [342] = \piso.data_r_342_sv2v_reg ;
  assign \piso.data_r [341] = \piso.data_r_341_sv2v_reg ;
  assign \piso.data_r [340] = \piso.data_r_340_sv2v_reg ;
  assign \piso.data_r [339] = \piso.data_r_339_sv2v_reg ;
  assign \piso.data_r [338] = \piso.data_r_338_sv2v_reg ;
  assign \piso.data_r [337] = \piso.data_r_337_sv2v_reg ;
  assign \piso.data_r [336] = \piso.data_r_336_sv2v_reg ;
  assign \piso.data_r [335] = \piso.data_r_335_sv2v_reg ;
  assign \piso.data_r [334] = \piso.data_r_334_sv2v_reg ;
  assign \piso.data_r [333] = \piso.data_r_333_sv2v_reg ;
  assign \piso.data_r [332] = \piso.data_r_332_sv2v_reg ;
  assign \piso.data_r [331] = \piso.data_r_331_sv2v_reg ;
  assign \piso.data_r [330] = \piso.data_r_330_sv2v_reg ;
  assign \piso.data_r [329] = \piso.data_r_329_sv2v_reg ;
  assign \piso.data_r [328] = \piso.data_r_328_sv2v_reg ;
  assign \piso.data_r [327] = \piso.data_r_327_sv2v_reg ;
  assign \piso.data_r [326] = \piso.data_r_326_sv2v_reg ;
  assign \piso.data_r [325] = \piso.data_r_325_sv2v_reg ;
  assign \piso.data_r [324] = \piso.data_r_324_sv2v_reg ;
  assign \piso.data_r [323] = \piso.data_r_323_sv2v_reg ;
  assign \piso.data_r [322] = \piso.data_r_322_sv2v_reg ;
  assign \piso.data_r [321] = \piso.data_r_321_sv2v_reg ;
  assign \piso.data_r [320] = \piso.data_r_320_sv2v_reg ;
  assign \piso.data_r [319] = \piso.data_r_319_sv2v_reg ;
  assign \piso.data_r [318] = \piso.data_r_318_sv2v_reg ;
  assign \piso.data_r [317] = \piso.data_r_317_sv2v_reg ;
  assign \piso.data_r [316] = \piso.data_r_316_sv2v_reg ;
  assign \piso.data_r [315] = \piso.data_r_315_sv2v_reg ;
  assign \piso.data_r [314] = \piso.data_r_314_sv2v_reg ;
  assign \piso.data_r [313] = \piso.data_r_313_sv2v_reg ;
  assign \piso.data_r [312] = \piso.data_r_312_sv2v_reg ;
  assign \piso.data_r [311] = \piso.data_r_311_sv2v_reg ;
  assign \piso.data_r [310] = \piso.data_r_310_sv2v_reg ;
  assign \piso.data_r [309] = \piso.data_r_309_sv2v_reg ;
  assign \piso.data_r [308] = \piso.data_r_308_sv2v_reg ;
  assign \piso.data_r [307] = \piso.data_r_307_sv2v_reg ;
  assign \piso.data_r [306] = \piso.data_r_306_sv2v_reg ;
  assign \piso.data_r [305] = \piso.data_r_305_sv2v_reg ;
  assign \piso.data_r [304] = \piso.data_r_304_sv2v_reg ;
  assign \piso.data_r [303] = \piso.data_r_303_sv2v_reg ;
  assign \piso.data_r [302] = \piso.data_r_302_sv2v_reg ;
  assign \piso.data_r [301] = \piso.data_r_301_sv2v_reg ;
  assign \piso.data_r [300] = \piso.data_r_300_sv2v_reg ;
  assign \piso.data_r [299] = \piso.data_r_299_sv2v_reg ;
  assign \piso.data_r [298] = \piso.data_r_298_sv2v_reg ;
  assign \piso.data_r [297] = \piso.data_r_297_sv2v_reg ;
  assign \piso.data_r [296] = \piso.data_r_296_sv2v_reg ;
  assign \piso.data_r [295] = \piso.data_r_295_sv2v_reg ;
  assign \piso.data_r [294] = \piso.data_r_294_sv2v_reg ;
  assign \piso.data_r [293] = \piso.data_r_293_sv2v_reg ;
  assign \piso.data_r [292] = \piso.data_r_292_sv2v_reg ;
  assign \piso.data_r [291] = \piso.data_r_291_sv2v_reg ;
  assign \piso.data_r [290] = \piso.data_r_290_sv2v_reg ;
  assign \piso.data_r [289] = \piso.data_r_289_sv2v_reg ;
  assign \piso.data_r [288] = \piso.data_r_288_sv2v_reg ;
  assign \piso.data_r [287] = \piso.data_r_287_sv2v_reg ;
  assign \piso.data_r [286] = \piso.data_r_286_sv2v_reg ;
  assign \piso.data_r [285] = \piso.data_r_285_sv2v_reg ;
  assign \piso.data_r [284] = \piso.data_r_284_sv2v_reg ;
  assign \piso.data_r [283] = \piso.data_r_283_sv2v_reg ;
  assign \piso.data_r [282] = \piso.data_r_282_sv2v_reg ;
  assign \piso.data_r [281] = \piso.data_r_281_sv2v_reg ;
  assign \piso.data_r [280] = \piso.data_r_280_sv2v_reg ;
  assign \piso.data_r [279] = \piso.data_r_279_sv2v_reg ;
  assign \piso.data_r [278] = \piso.data_r_278_sv2v_reg ;
  assign \piso.data_r [277] = \piso.data_r_277_sv2v_reg ;
  assign \piso.data_r [276] = \piso.data_r_276_sv2v_reg ;
  assign \piso.data_r [275] = \piso.data_r_275_sv2v_reg ;
  assign \piso.data_r [274] = \piso.data_r_274_sv2v_reg ;
  assign \piso.data_r [273] = \piso.data_r_273_sv2v_reg ;
  assign \piso.data_r [272] = \piso.data_r_272_sv2v_reg ;
  assign \piso.data_r [271] = \piso.data_r_271_sv2v_reg ;
  assign \piso.data_r [270] = \piso.data_r_270_sv2v_reg ;
  assign \piso.data_r [269] = \piso.data_r_269_sv2v_reg ;
  assign \piso.data_r [268] = \piso.data_r_268_sv2v_reg ;
  assign \piso.data_r [267] = \piso.data_r_267_sv2v_reg ;
  assign \piso.data_r [266] = \piso.data_r_266_sv2v_reg ;
  assign \piso.data_r [265] = \piso.data_r_265_sv2v_reg ;
  assign \piso.data_r [264] = \piso.data_r_264_sv2v_reg ;
  assign \piso.data_r [263] = \piso.data_r_263_sv2v_reg ;
  assign \piso.data_r [262] = \piso.data_r_262_sv2v_reg ;
  assign \piso.data_r [261] = \piso.data_r_261_sv2v_reg ;
  assign \piso.data_r [260] = \piso.data_r_260_sv2v_reg ;
  assign \piso.data_r [259] = \piso.data_r_259_sv2v_reg ;
  assign \piso.data_r [258] = \piso.data_r_258_sv2v_reg ;
  assign \piso.data_r [257] = \piso.data_r_257_sv2v_reg ;
  assign \piso.data_r [256] = \piso.data_r_256_sv2v_reg ;
  assign \piso.data_r [255] = \piso.data_r_255_sv2v_reg ;
  assign \piso.data_r [254] = \piso.data_r_254_sv2v_reg ;
  assign \piso.data_r [253] = \piso.data_r_253_sv2v_reg ;
  assign \piso.data_r [252] = \piso.data_r_252_sv2v_reg ;
  assign \piso.data_r [251] = \piso.data_r_251_sv2v_reg ;
  assign \piso.data_r [250] = \piso.data_r_250_sv2v_reg ;
  assign \piso.data_r [249] = \piso.data_r_249_sv2v_reg ;
  assign \piso.data_r [248] = \piso.data_r_248_sv2v_reg ;
  assign \piso.data_r [247] = \piso.data_r_247_sv2v_reg ;
  assign \piso.data_r [246] = \piso.data_r_246_sv2v_reg ;
  assign \piso.data_r [245] = \piso.data_r_245_sv2v_reg ;
  assign \piso.data_r [244] = \piso.data_r_244_sv2v_reg ;
  assign \piso.data_r [243] = \piso.data_r_243_sv2v_reg ;
  assign \piso.data_r [242] = \piso.data_r_242_sv2v_reg ;
  assign \piso.data_r [241] = \piso.data_r_241_sv2v_reg ;
  assign \piso.data_r [240] = \piso.data_r_240_sv2v_reg ;
  assign \piso.data_r [239] = \piso.data_r_239_sv2v_reg ;
  assign \piso.data_r [238] = \piso.data_r_238_sv2v_reg ;
  assign \piso.data_r [237] = \piso.data_r_237_sv2v_reg ;
  assign \piso.data_r [236] = \piso.data_r_236_sv2v_reg ;
  assign \piso.data_r [235] = \piso.data_r_235_sv2v_reg ;
  assign \piso.data_r [234] = \piso.data_r_234_sv2v_reg ;
  assign \piso.data_r [233] = \piso.data_r_233_sv2v_reg ;
  assign \piso.data_r [232] = \piso.data_r_232_sv2v_reg ;
  assign \piso.data_r [231] = \piso.data_r_231_sv2v_reg ;
  assign \piso.data_r [230] = \piso.data_r_230_sv2v_reg ;
  assign \piso.data_r [229] = \piso.data_r_229_sv2v_reg ;
  assign \piso.data_r [228] = \piso.data_r_228_sv2v_reg ;
  assign \piso.data_r [227] = \piso.data_r_227_sv2v_reg ;
  assign \piso.data_r [226] = \piso.data_r_226_sv2v_reg ;
  assign \piso.data_r [225] = \piso.data_r_225_sv2v_reg ;
  assign \piso.data_r [224] = \piso.data_r_224_sv2v_reg ;
  assign \piso.data_r [223] = \piso.data_r_223_sv2v_reg ;
  assign \piso.data_r [222] = \piso.data_r_222_sv2v_reg ;
  assign \piso.data_r [221] = \piso.data_r_221_sv2v_reg ;
  assign \piso.data_r [220] = \piso.data_r_220_sv2v_reg ;
  assign \piso.data_r [219] = \piso.data_r_219_sv2v_reg ;
  assign \piso.data_r [218] = \piso.data_r_218_sv2v_reg ;
  assign \piso.data_r [217] = \piso.data_r_217_sv2v_reg ;
  assign \piso.data_r [216] = \piso.data_r_216_sv2v_reg ;
  assign \piso.data_r [215] = \piso.data_r_215_sv2v_reg ;
  assign \piso.data_r [214] = \piso.data_r_214_sv2v_reg ;
  assign \piso.data_r [213] = \piso.data_r_213_sv2v_reg ;
  assign \piso.data_r [212] = \piso.data_r_212_sv2v_reg ;
  assign \piso.data_r [211] = \piso.data_r_211_sv2v_reg ;
  assign \piso.data_r [210] = \piso.data_r_210_sv2v_reg ;
  assign \piso.data_r [209] = \piso.data_r_209_sv2v_reg ;
  assign \piso.data_r [208] = \piso.data_r_208_sv2v_reg ;
  assign \piso.data_r [207] = \piso.data_r_207_sv2v_reg ;
  assign \piso.data_r [206] = \piso.data_r_206_sv2v_reg ;
  assign \piso.data_r [205] = \piso.data_r_205_sv2v_reg ;
  assign \piso.data_r [204] = \piso.data_r_204_sv2v_reg ;
  assign \piso.data_r [203] = \piso.data_r_203_sv2v_reg ;
  assign \piso.data_r [202] = \piso.data_r_202_sv2v_reg ;
  assign \piso.data_r [201] = \piso.data_r_201_sv2v_reg ;
  assign \piso.data_r [200] = \piso.data_r_200_sv2v_reg ;
  assign \piso.data_r [199] = \piso.data_r_199_sv2v_reg ;
  assign \piso.data_r [198] = \piso.data_r_198_sv2v_reg ;
  assign \piso.data_r [197] = \piso.data_r_197_sv2v_reg ;
  assign \piso.data_r [196] = \piso.data_r_196_sv2v_reg ;
  assign \piso.data_r [195] = \piso.data_r_195_sv2v_reg ;
  assign \piso.data_r [194] = \piso.data_r_194_sv2v_reg ;
  assign \piso.data_r [193] = \piso.data_r_193_sv2v_reg ;
  assign \piso.data_r [192] = \piso.data_r_192_sv2v_reg ;
  assign \piso.data_r [191] = \piso.data_r_191_sv2v_reg ;
  assign \piso.data_r [190] = \piso.data_r_190_sv2v_reg ;
  assign \piso.data_r [189] = \piso.data_r_189_sv2v_reg ;
  assign \piso.data_r [188] = \piso.data_r_188_sv2v_reg ;
  assign \piso.data_r [187] = \piso.data_r_187_sv2v_reg ;
  assign \piso.data_r [186] = \piso.data_r_186_sv2v_reg ;
  assign \piso.data_r [185] = \piso.data_r_185_sv2v_reg ;
  assign \piso.data_r [184] = \piso.data_r_184_sv2v_reg ;
  assign \piso.data_r [183] = \piso.data_r_183_sv2v_reg ;
  assign \piso.data_r [182] = \piso.data_r_182_sv2v_reg ;
  assign \piso.data_r [181] = \piso.data_r_181_sv2v_reg ;
  assign \piso.data_r [180] = \piso.data_r_180_sv2v_reg ;
  assign \piso.data_r [179] = \piso.data_r_179_sv2v_reg ;
  assign \piso.data_r [178] = \piso.data_r_178_sv2v_reg ;
  assign \piso.data_r [177] = \piso.data_r_177_sv2v_reg ;
  assign \piso.data_r [176] = \piso.data_r_176_sv2v_reg ;
  assign \piso.data_r [175] = \piso.data_r_175_sv2v_reg ;
  assign \piso.data_r [174] = \piso.data_r_174_sv2v_reg ;
  assign \piso.data_r [173] = \piso.data_r_173_sv2v_reg ;
  assign \piso.data_r [172] = \piso.data_r_172_sv2v_reg ;
  assign \piso.data_r [171] = \piso.data_r_171_sv2v_reg ;
  assign \piso.data_r [170] = \piso.data_r_170_sv2v_reg ;
  assign \piso.data_r [169] = \piso.data_r_169_sv2v_reg ;
  assign \piso.data_r [168] = \piso.data_r_168_sv2v_reg ;
  assign \piso.data_r [167] = \piso.data_r_167_sv2v_reg ;
  assign \piso.data_r [166] = \piso.data_r_166_sv2v_reg ;
  assign \piso.data_r [165] = \piso.data_r_165_sv2v_reg ;
  assign \piso.data_r [164] = \piso.data_r_164_sv2v_reg ;
  assign \piso.data_r [163] = \piso.data_r_163_sv2v_reg ;
  assign \piso.data_r [162] = \piso.data_r_162_sv2v_reg ;
  assign \piso.data_r [161] = \piso.data_r_161_sv2v_reg ;
  assign \piso.data_r [160] = \piso.data_r_160_sv2v_reg ;
  assign \piso.data_r [159] = \piso.data_r_159_sv2v_reg ;
  assign \piso.data_r [158] = \piso.data_r_158_sv2v_reg ;
  assign \piso.data_r [157] = \piso.data_r_157_sv2v_reg ;
  assign \piso.data_r [156] = \piso.data_r_156_sv2v_reg ;
  assign \piso.data_r [155] = \piso.data_r_155_sv2v_reg ;
  assign \piso.data_r [154] = \piso.data_r_154_sv2v_reg ;
  assign \piso.data_r [153] = \piso.data_r_153_sv2v_reg ;
  assign \piso.data_r [152] = \piso.data_r_152_sv2v_reg ;
  assign \piso.data_r [151] = \piso.data_r_151_sv2v_reg ;
  assign \piso.data_r [150] = \piso.data_r_150_sv2v_reg ;
  assign \piso.data_r [149] = \piso.data_r_149_sv2v_reg ;
  assign \piso.data_r [148] = \piso.data_r_148_sv2v_reg ;
  assign \piso.data_r [147] = \piso.data_r_147_sv2v_reg ;
  assign \piso.data_r [146] = \piso.data_r_146_sv2v_reg ;
  assign \piso.data_r [145] = \piso.data_r_145_sv2v_reg ;
  assign \piso.data_r [144] = \piso.data_r_144_sv2v_reg ;
  assign \piso.data_r [143] = \piso.data_r_143_sv2v_reg ;
  assign \piso.data_r [142] = \piso.data_r_142_sv2v_reg ;
  assign \piso.data_r [141] = \piso.data_r_141_sv2v_reg ;
  assign \piso.data_r [140] = \piso.data_r_140_sv2v_reg ;
  assign \piso.data_r [139] = \piso.data_r_139_sv2v_reg ;
  assign \piso.data_r [138] = \piso.data_r_138_sv2v_reg ;
  assign \piso.data_r [137] = \piso.data_r_137_sv2v_reg ;
  assign \piso.data_r [136] = \piso.data_r_136_sv2v_reg ;
  assign \piso.data_r [135] = \piso.data_r_135_sv2v_reg ;
  assign \piso.data_r [134] = \piso.data_r_134_sv2v_reg ;
  assign \piso.data_r [133] = \piso.data_r_133_sv2v_reg ;
  assign \piso.data_r [132] = \piso.data_r_132_sv2v_reg ;
  assign \piso.data_r [131] = \piso.data_r_131_sv2v_reg ;
  assign \piso.data_r [130] = \piso.data_r_130_sv2v_reg ;
  assign \piso.data_r [129] = \piso.data_r_129_sv2v_reg ;
  assign \piso.data_r [128] = \piso.data_r_128_sv2v_reg ;
  assign \piso.data_r [127] = \piso.data_r_127_sv2v_reg ;
  assign \piso.data_r [126] = \piso.data_r_126_sv2v_reg ;
  assign \piso.data_r [125] = \piso.data_r_125_sv2v_reg ;
  assign \piso.data_r [124] = \piso.data_r_124_sv2v_reg ;
  assign \piso.data_r [123] = \piso.data_r_123_sv2v_reg ;
  assign \piso.data_r [122] = \piso.data_r_122_sv2v_reg ;
  assign \piso.data_r [121] = \piso.data_r_121_sv2v_reg ;
  assign \piso.data_r [120] = \piso.data_r_120_sv2v_reg ;
  assign \piso.data_r [119] = \piso.data_r_119_sv2v_reg ;
  assign \piso.data_r [118] = \piso.data_r_118_sv2v_reg ;
  assign \piso.data_r [117] = \piso.data_r_117_sv2v_reg ;
  assign \piso.data_r [116] = \piso.data_r_116_sv2v_reg ;
  assign \piso.data_r [115] = \piso.data_r_115_sv2v_reg ;
  assign \piso.data_r [114] = \piso.data_r_114_sv2v_reg ;
  assign \piso.data_r [113] = \piso.data_r_113_sv2v_reg ;
  assign \piso.data_r [112] = \piso.data_r_112_sv2v_reg ;
  assign \piso.data_r [111] = \piso.data_r_111_sv2v_reg ;
  assign \piso.data_r [110] = \piso.data_r_110_sv2v_reg ;
  assign \piso.data_r [109] = \piso.data_r_109_sv2v_reg ;
  assign \piso.data_r [108] = \piso.data_r_108_sv2v_reg ;
  assign \piso.data_r [107] = \piso.data_r_107_sv2v_reg ;
  assign \piso.data_r [106] = \piso.data_r_106_sv2v_reg ;
  assign \piso.data_r [105] = \piso.data_r_105_sv2v_reg ;
  assign \piso.data_r [104] = \piso.data_r_104_sv2v_reg ;
  assign \piso.data_r [103] = \piso.data_r_103_sv2v_reg ;
  assign \piso.data_r [102] = \piso.data_r_102_sv2v_reg ;
  assign \piso.data_r [101] = \piso.data_r_101_sv2v_reg ;
  assign \piso.data_r [100] = \piso.data_r_100_sv2v_reg ;
  assign \piso.data_r [99] = \piso.data_r_99_sv2v_reg ;
  assign \piso.data_r [98] = \piso.data_r_98_sv2v_reg ;
  assign \piso.data_r [97] = \piso.data_r_97_sv2v_reg ;
  assign \piso.data_r [96] = \piso.data_r_96_sv2v_reg ;
  assign \piso.data_r [95] = \piso.data_r_95_sv2v_reg ;
  assign \piso.data_r [94] = \piso.data_r_94_sv2v_reg ;
  assign \piso.data_r [93] = \piso.data_r_93_sv2v_reg ;
  assign \piso.data_r [92] = \piso.data_r_92_sv2v_reg ;
  assign \piso.data_r [91] = \piso.data_r_91_sv2v_reg ;
  assign \piso.data_r [90] = \piso.data_r_90_sv2v_reg ;
  assign \piso.data_r [89] = \piso.data_r_89_sv2v_reg ;
  assign \piso.data_r [88] = \piso.data_r_88_sv2v_reg ;
  assign \piso.data_r [87] = \piso.data_r_87_sv2v_reg ;
  assign \piso.data_r [86] = \piso.data_r_86_sv2v_reg ;
  assign \piso.data_r [85] = \piso.data_r_85_sv2v_reg ;
  assign \piso.data_r [84] = \piso.data_r_84_sv2v_reg ;
  assign \piso.data_r [83] = \piso.data_r_83_sv2v_reg ;
  assign \piso.data_r [82] = \piso.data_r_82_sv2v_reg ;
  assign \piso.data_r [81] = \piso.data_r_81_sv2v_reg ;
  assign \piso.data_r [80] = \piso.data_r_80_sv2v_reg ;
  assign \piso.data_r [79] = \piso.data_r_79_sv2v_reg ;
  assign \piso.data_r [78] = \piso.data_r_78_sv2v_reg ;
  assign \piso.data_r [77] = \piso.data_r_77_sv2v_reg ;
  assign \piso.data_r [76] = \piso.data_r_76_sv2v_reg ;
  assign \piso.data_r [75] = \piso.data_r_75_sv2v_reg ;
  assign \piso.data_r [74] = \piso.data_r_74_sv2v_reg ;
  assign \piso.data_r [73] = \piso.data_r_73_sv2v_reg ;
  assign \piso.data_r [72] = \piso.data_r_72_sv2v_reg ;
  assign \piso.data_r [71] = \piso.data_r_71_sv2v_reg ;
  assign \piso.data_r [70] = \piso.data_r_70_sv2v_reg ;
  assign \piso.data_r [69] = \piso.data_r_69_sv2v_reg ;
  assign \piso.data_r [68] = \piso.data_r_68_sv2v_reg ;
  assign \piso.data_r [67] = \piso.data_r_67_sv2v_reg ;
  assign \piso.data_r [66] = \piso.data_r_66_sv2v_reg ;
  assign \piso.data_r [65] = \piso.data_r_65_sv2v_reg ;
  assign \piso.data_r [64] = \piso.data_r_64_sv2v_reg ;
  assign \piso.data_r [63] = \piso.data_r_63_sv2v_reg ;
  assign \piso.data_r [62] = \piso.data_r_62_sv2v_reg ;
  assign \piso.data_r [61] = \piso.data_r_61_sv2v_reg ;
  assign \piso.data_r [60] = \piso.data_r_60_sv2v_reg ;
  assign \piso.data_r [59] = \piso.data_r_59_sv2v_reg ;
  assign \piso.data_r [58] = \piso.data_r_58_sv2v_reg ;
  assign \piso.data_r [57] = \piso.data_r_57_sv2v_reg ;
  assign \piso.data_r [56] = \piso.data_r_56_sv2v_reg ;
  assign \piso.data_r [55] = \piso.data_r_55_sv2v_reg ;
  assign \piso.data_r [54] = \piso.data_r_54_sv2v_reg ;
  assign \piso.data_r [53] = \piso.data_r_53_sv2v_reg ;
  assign \piso.data_r [52] = \piso.data_r_52_sv2v_reg ;
  assign \piso.data_r [51] = \piso.data_r_51_sv2v_reg ;
  assign \piso.data_r [50] = \piso.data_r_50_sv2v_reg ;
  assign \piso.data_r [49] = \piso.data_r_49_sv2v_reg ;
  assign \piso.data_r [48] = \piso.data_r_48_sv2v_reg ;
  assign \piso.data_r [47] = \piso.data_r_47_sv2v_reg ;
  assign \piso.data_r [46] = \piso.data_r_46_sv2v_reg ;
  assign \piso.data_r [45] = \piso.data_r_45_sv2v_reg ;
  assign \piso.data_r [44] = \piso.data_r_44_sv2v_reg ;
  assign \piso.data_r [43] = \piso.data_r_43_sv2v_reg ;
  assign \piso.data_r [42] = \piso.data_r_42_sv2v_reg ;
  assign \piso.data_r [41] = \piso.data_r_41_sv2v_reg ;
  assign \piso.data_r [40] = \piso.data_r_40_sv2v_reg ;
  assign \piso.data_r [39] = \piso.data_r_39_sv2v_reg ;
  assign \piso.data_r [38] = \piso.data_r_38_sv2v_reg ;
  assign \piso.data_r [37] = \piso.data_r_37_sv2v_reg ;
  assign \piso.data_r [36] = \piso.data_r_36_sv2v_reg ;
  assign \piso.data_r [35] = \piso.data_r_35_sv2v_reg ;
  assign \piso.data_r [34] = \piso.data_r_34_sv2v_reg ;
  assign \piso.data_r [33] = \piso.data_r_33_sv2v_reg ;
  assign \piso.data_r [32] = \piso.data_r_32_sv2v_reg ;
  assign \piso.data_r [31] = \piso.data_r_31_sv2v_reg ;
  assign \piso.data_r [30] = \piso.data_r_30_sv2v_reg ;
  assign \piso.data_r [29] = \piso.data_r_29_sv2v_reg ;
  assign \piso.data_r [28] = \piso.data_r_28_sv2v_reg ;
  assign \piso.data_r [27] = \piso.data_r_27_sv2v_reg ;
  assign \piso.data_r [26] = \piso.data_r_26_sv2v_reg ;
  assign \piso.data_r [25] = \piso.data_r_25_sv2v_reg ;
  assign \piso.data_r [24] = \piso.data_r_24_sv2v_reg ;
  assign \piso.data_r [23] = \piso.data_r_23_sv2v_reg ;
  assign \piso.data_r [22] = \piso.data_r_22_sv2v_reg ;
  assign \piso.data_r [21] = \piso.data_r_21_sv2v_reg ;
  assign \piso.data_r [20] = \piso.data_r_20_sv2v_reg ;
  assign \piso.data_r [19] = \piso.data_r_19_sv2v_reg ;
  assign \piso.data_r [18] = \piso.data_r_18_sv2v_reg ;
  assign \piso.data_r [17] = \piso.data_r_17_sv2v_reg ;
  assign \piso.data_r [16] = \piso.data_r_16_sv2v_reg ;
  assign \piso.data_r [15] = \piso.data_r_15_sv2v_reg ;
  assign \piso.data_r [14] = \piso.data_r_14_sv2v_reg ;
  assign \piso.data_r [13] = \piso.data_r_13_sv2v_reg ;
  assign \piso.data_r [12] = \piso.data_r_12_sv2v_reg ;
  assign \piso.data_r [11] = \piso.data_r_11_sv2v_reg ;
  assign \piso.data_r [10] = \piso.data_r_10_sv2v_reg ;
  assign \piso.data_r [9] = \piso.data_r_9_sv2v_reg ;
  assign \piso.data_r [8] = \piso.data_r_8_sv2v_reg ;
  assign \piso.data_r [7] = \piso.data_r_7_sv2v_reg ;
  assign \piso.data_r [6] = \piso.data_r_6_sv2v_reg ;
  assign \piso.data_r [5] = \piso.data_r_5_sv2v_reg ;
  assign \piso.data_r [4] = \piso.data_r_4_sv2v_reg ;
  assign \piso.data_r [3] = \piso.data_r_3_sv2v_reg ;
  assign \piso.data_r [2] = \piso.data_r_2_sv2v_reg ;
  assign \piso.data_r [1] = \piso.data_r_1_sv2v_reg ;
  assign \piso.data_r [0] = \piso.data_r_0_sv2v_reg ;
  assign \piso.shift_ctr_r [5] = \piso.shift_ctr_r_5_sv2v_reg ;
  assign \piso.shift_ctr_r [4] = \piso.shift_ctr_r_4_sv2v_reg ;
  assign \piso.shift_ctr_r [3] = \piso.shift_ctr_r_3_sv2v_reg ;
  assign \piso.shift_ctr_r [2] = \piso.shift_ctr_r_2_sv2v_reg ;
  assign \piso.shift_ctr_r [1] = \piso.shift_ctr_r_1_sv2v_reg ;
  assign \piso.shift_ctr_r [0] = \piso.shift_ctr_r_0_sv2v_reg ;

  bsg_array_reverse_width_p32_els_p64
  \piso.hi2lo.bar 
  (
    .i(data_i),
    .o(\piso.data_li )
  );

  assign data_o[31] = (N89)? \piso.data_r [31] : 
                      (N91)? \piso.data_r [63] : 
                      (N93)? \piso.data_r [95] : 
                      (N95)? \piso.data_r [127] : 
                      (N97)? \piso.data_r [159] : 
                      (N99)? \piso.data_r [191] : 
                      (N101)? \piso.data_r [223] : 
                      (N103)? \piso.data_r [255] : 
                      (N105)? \piso.data_r [287] : 
                      (N107)? \piso.data_r [319] : 
                      (N109)? \piso.data_r [351] : 
                      (N111)? \piso.data_r [383] : 
                      (N113)? \piso.data_r [415] : 
                      (N115)? \piso.data_r [447] : 
                      (N117)? \piso.data_r [479] : 
                      (N119)? \piso.data_r [511] : 
                      (N121)? \piso.data_r [543] : 
                      (N123)? \piso.data_r [575] : 
                      (N125)? \piso.data_r [607] : 
                      (N127)? \piso.data_r [639] : 
                      (N129)? \piso.data_r [671] : 
                      (N131)? \piso.data_r [703] : 
                      (N133)? \piso.data_r [735] : 
                      (N135)? \piso.data_r [767] : 
                      (N137)? \piso.data_r [799] : 
                      (N139)? \piso.data_r [831] : 
                      (N141)? \piso.data_r [863] : 
                      (N143)? \piso.data_r [895] : 
                      (N145)? \piso.data_r [927] : 
                      (N147)? \piso.data_r [959] : 
                      (N149)? \piso.data_r [991] : 
                      (N151)? \piso.data_r [1023] : 
                      (N90)? \piso.data_r [1055] : 
                      (N92)? \piso.data_r [1087] : 
                      (N94)? \piso.data_r [1119] : 
                      (N96)? \piso.data_r [1151] : 
                      (N98)? \piso.data_r [1183] : 
                      (N100)? \piso.data_r [1215] : 
                      (N102)? \piso.data_r [1247] : 
                      (N104)? \piso.data_r [1279] : 
                      (N106)? \piso.data_r [1311] : 
                      (N108)? \piso.data_r [1343] : 
                      (N110)? \piso.data_r [1375] : 
                      (N112)? \piso.data_r [1407] : 
                      (N114)? \piso.data_r [1439] : 
                      (N116)? \piso.data_r [1471] : 
                      (N118)? \piso.data_r [1503] : 
                      (N120)? \piso.data_r [1535] : 
                      (N122)? \piso.data_r [1567] : 
                      (N124)? \piso.data_r [1599] : 
                      (N126)? \piso.data_r [1631] : 
                      (N128)? \piso.data_r [1663] : 
                      (N130)? \piso.data_r [1695] : 
                      (N132)? \piso.data_r [1727] : 
                      (N134)? \piso.data_r [1759] : 
                      (N136)? \piso.data_r [1791] : 
                      (N138)? \piso.data_r [1823] : 
                      (N140)? \piso.data_r [1855] : 
                      (N142)? \piso.data_r [1887] : 
                      (N144)? \piso.data_r [1919] : 
                      (N146)? \piso.data_r [1951] : 
                      (N148)? \piso.data_r [1983] : 
                      (N150)? \piso.data_r [2015] : 
                      (N152)? \piso.data_r [2047] : 1'b0;
  assign data_o[30] = (N89)? \piso.data_r [30] : 
                      (N91)? \piso.data_r [62] : 
                      (N93)? \piso.data_r [94] : 
                      (N95)? \piso.data_r [126] : 
                      (N97)? \piso.data_r [158] : 
                      (N99)? \piso.data_r [190] : 
                      (N101)? \piso.data_r [222] : 
                      (N103)? \piso.data_r [254] : 
                      (N105)? \piso.data_r [286] : 
                      (N107)? \piso.data_r [318] : 
                      (N109)? \piso.data_r [350] : 
                      (N111)? \piso.data_r [382] : 
                      (N113)? \piso.data_r [414] : 
                      (N115)? \piso.data_r [446] : 
                      (N117)? \piso.data_r [478] : 
                      (N119)? \piso.data_r [510] : 
                      (N121)? \piso.data_r [542] : 
                      (N123)? \piso.data_r [574] : 
                      (N125)? \piso.data_r [606] : 
                      (N127)? \piso.data_r [638] : 
                      (N129)? \piso.data_r [670] : 
                      (N131)? \piso.data_r [702] : 
                      (N133)? \piso.data_r [734] : 
                      (N135)? \piso.data_r [766] : 
                      (N137)? \piso.data_r [798] : 
                      (N139)? \piso.data_r [830] : 
                      (N141)? \piso.data_r [862] : 
                      (N143)? \piso.data_r [894] : 
                      (N145)? \piso.data_r [926] : 
                      (N147)? \piso.data_r [958] : 
                      (N149)? \piso.data_r [990] : 
                      (N151)? \piso.data_r [1022] : 
                      (N90)? \piso.data_r [1054] : 
                      (N92)? \piso.data_r [1086] : 
                      (N94)? \piso.data_r [1118] : 
                      (N96)? \piso.data_r [1150] : 
                      (N98)? \piso.data_r [1182] : 
                      (N100)? \piso.data_r [1214] : 
                      (N102)? \piso.data_r [1246] : 
                      (N104)? \piso.data_r [1278] : 
                      (N106)? \piso.data_r [1310] : 
                      (N108)? \piso.data_r [1342] : 
                      (N110)? \piso.data_r [1374] : 
                      (N112)? \piso.data_r [1406] : 
                      (N114)? \piso.data_r [1438] : 
                      (N116)? \piso.data_r [1470] : 
                      (N118)? \piso.data_r [1502] : 
                      (N120)? \piso.data_r [1534] : 
                      (N122)? \piso.data_r [1566] : 
                      (N124)? \piso.data_r [1598] : 
                      (N126)? \piso.data_r [1630] : 
                      (N128)? \piso.data_r [1662] : 
                      (N130)? \piso.data_r [1694] : 
                      (N132)? \piso.data_r [1726] : 
                      (N134)? \piso.data_r [1758] : 
                      (N136)? \piso.data_r [1790] : 
                      (N138)? \piso.data_r [1822] : 
                      (N140)? \piso.data_r [1854] : 
                      (N142)? \piso.data_r [1886] : 
                      (N144)? \piso.data_r [1918] : 
                      (N146)? \piso.data_r [1950] : 
                      (N148)? \piso.data_r [1982] : 
                      (N150)? \piso.data_r [2014] : 
                      (N152)? \piso.data_r [2046] : 1'b0;
  assign data_o[29] = (N89)? \piso.data_r [29] : 
                      (N91)? \piso.data_r [61] : 
                      (N93)? \piso.data_r [93] : 
                      (N95)? \piso.data_r [125] : 
                      (N97)? \piso.data_r [157] : 
                      (N99)? \piso.data_r [189] : 
                      (N101)? \piso.data_r [221] : 
                      (N103)? \piso.data_r [253] : 
                      (N105)? \piso.data_r [285] : 
                      (N107)? \piso.data_r [317] : 
                      (N109)? \piso.data_r [349] : 
                      (N111)? \piso.data_r [381] : 
                      (N113)? \piso.data_r [413] : 
                      (N115)? \piso.data_r [445] : 
                      (N117)? \piso.data_r [477] : 
                      (N119)? \piso.data_r [509] : 
                      (N121)? \piso.data_r [541] : 
                      (N123)? \piso.data_r [573] : 
                      (N125)? \piso.data_r [605] : 
                      (N127)? \piso.data_r [637] : 
                      (N129)? \piso.data_r [669] : 
                      (N131)? \piso.data_r [701] : 
                      (N133)? \piso.data_r [733] : 
                      (N135)? \piso.data_r [765] : 
                      (N137)? \piso.data_r [797] : 
                      (N139)? \piso.data_r [829] : 
                      (N141)? \piso.data_r [861] : 
                      (N143)? \piso.data_r [893] : 
                      (N145)? \piso.data_r [925] : 
                      (N147)? \piso.data_r [957] : 
                      (N149)? \piso.data_r [989] : 
                      (N151)? \piso.data_r [1021] : 
                      (N90)? \piso.data_r [1053] : 
                      (N92)? \piso.data_r [1085] : 
                      (N94)? \piso.data_r [1117] : 
                      (N96)? \piso.data_r [1149] : 
                      (N98)? \piso.data_r [1181] : 
                      (N100)? \piso.data_r [1213] : 
                      (N102)? \piso.data_r [1245] : 
                      (N104)? \piso.data_r [1277] : 
                      (N106)? \piso.data_r [1309] : 
                      (N108)? \piso.data_r [1341] : 
                      (N110)? \piso.data_r [1373] : 
                      (N112)? \piso.data_r [1405] : 
                      (N114)? \piso.data_r [1437] : 
                      (N116)? \piso.data_r [1469] : 
                      (N118)? \piso.data_r [1501] : 
                      (N120)? \piso.data_r [1533] : 
                      (N122)? \piso.data_r [1565] : 
                      (N124)? \piso.data_r [1597] : 
                      (N126)? \piso.data_r [1629] : 
                      (N128)? \piso.data_r [1661] : 
                      (N130)? \piso.data_r [1693] : 
                      (N132)? \piso.data_r [1725] : 
                      (N134)? \piso.data_r [1757] : 
                      (N136)? \piso.data_r [1789] : 
                      (N138)? \piso.data_r [1821] : 
                      (N140)? \piso.data_r [1853] : 
                      (N142)? \piso.data_r [1885] : 
                      (N144)? \piso.data_r [1917] : 
                      (N146)? \piso.data_r [1949] : 
                      (N148)? \piso.data_r [1981] : 
                      (N150)? \piso.data_r [2013] : 
                      (N152)? \piso.data_r [2045] : 1'b0;
  assign data_o[28] = (N89)? \piso.data_r [28] : 
                      (N91)? \piso.data_r [60] : 
                      (N93)? \piso.data_r [92] : 
                      (N95)? \piso.data_r [124] : 
                      (N97)? \piso.data_r [156] : 
                      (N99)? \piso.data_r [188] : 
                      (N101)? \piso.data_r [220] : 
                      (N103)? \piso.data_r [252] : 
                      (N105)? \piso.data_r [284] : 
                      (N107)? \piso.data_r [316] : 
                      (N109)? \piso.data_r [348] : 
                      (N111)? \piso.data_r [380] : 
                      (N113)? \piso.data_r [412] : 
                      (N115)? \piso.data_r [444] : 
                      (N117)? \piso.data_r [476] : 
                      (N119)? \piso.data_r [508] : 
                      (N121)? \piso.data_r [540] : 
                      (N123)? \piso.data_r [572] : 
                      (N125)? \piso.data_r [604] : 
                      (N127)? \piso.data_r [636] : 
                      (N129)? \piso.data_r [668] : 
                      (N131)? \piso.data_r [700] : 
                      (N133)? \piso.data_r [732] : 
                      (N135)? \piso.data_r [764] : 
                      (N137)? \piso.data_r [796] : 
                      (N139)? \piso.data_r [828] : 
                      (N141)? \piso.data_r [860] : 
                      (N143)? \piso.data_r [892] : 
                      (N145)? \piso.data_r [924] : 
                      (N147)? \piso.data_r [956] : 
                      (N149)? \piso.data_r [988] : 
                      (N151)? \piso.data_r [1020] : 
                      (N90)? \piso.data_r [1052] : 
                      (N92)? \piso.data_r [1084] : 
                      (N94)? \piso.data_r [1116] : 
                      (N96)? \piso.data_r [1148] : 
                      (N98)? \piso.data_r [1180] : 
                      (N100)? \piso.data_r [1212] : 
                      (N102)? \piso.data_r [1244] : 
                      (N104)? \piso.data_r [1276] : 
                      (N106)? \piso.data_r [1308] : 
                      (N108)? \piso.data_r [1340] : 
                      (N110)? \piso.data_r [1372] : 
                      (N112)? \piso.data_r [1404] : 
                      (N114)? \piso.data_r [1436] : 
                      (N116)? \piso.data_r [1468] : 
                      (N118)? \piso.data_r [1500] : 
                      (N120)? \piso.data_r [1532] : 
                      (N122)? \piso.data_r [1564] : 
                      (N124)? \piso.data_r [1596] : 
                      (N126)? \piso.data_r [1628] : 
                      (N128)? \piso.data_r [1660] : 
                      (N130)? \piso.data_r [1692] : 
                      (N132)? \piso.data_r [1724] : 
                      (N134)? \piso.data_r [1756] : 
                      (N136)? \piso.data_r [1788] : 
                      (N138)? \piso.data_r [1820] : 
                      (N140)? \piso.data_r [1852] : 
                      (N142)? \piso.data_r [1884] : 
                      (N144)? \piso.data_r [1916] : 
                      (N146)? \piso.data_r [1948] : 
                      (N148)? \piso.data_r [1980] : 
                      (N150)? \piso.data_r [2012] : 
                      (N152)? \piso.data_r [2044] : 1'b0;
  assign data_o[27] = (N89)? \piso.data_r [27] : 
                      (N91)? \piso.data_r [59] : 
                      (N93)? \piso.data_r [91] : 
                      (N95)? \piso.data_r [123] : 
                      (N97)? \piso.data_r [155] : 
                      (N99)? \piso.data_r [187] : 
                      (N101)? \piso.data_r [219] : 
                      (N103)? \piso.data_r [251] : 
                      (N105)? \piso.data_r [283] : 
                      (N107)? \piso.data_r [315] : 
                      (N109)? \piso.data_r [347] : 
                      (N111)? \piso.data_r [379] : 
                      (N113)? \piso.data_r [411] : 
                      (N115)? \piso.data_r [443] : 
                      (N117)? \piso.data_r [475] : 
                      (N119)? \piso.data_r [507] : 
                      (N121)? \piso.data_r [539] : 
                      (N123)? \piso.data_r [571] : 
                      (N125)? \piso.data_r [603] : 
                      (N127)? \piso.data_r [635] : 
                      (N129)? \piso.data_r [667] : 
                      (N131)? \piso.data_r [699] : 
                      (N133)? \piso.data_r [731] : 
                      (N135)? \piso.data_r [763] : 
                      (N137)? \piso.data_r [795] : 
                      (N139)? \piso.data_r [827] : 
                      (N141)? \piso.data_r [859] : 
                      (N143)? \piso.data_r [891] : 
                      (N145)? \piso.data_r [923] : 
                      (N147)? \piso.data_r [955] : 
                      (N149)? \piso.data_r [987] : 
                      (N151)? \piso.data_r [1019] : 
                      (N90)? \piso.data_r [1051] : 
                      (N92)? \piso.data_r [1083] : 
                      (N94)? \piso.data_r [1115] : 
                      (N96)? \piso.data_r [1147] : 
                      (N98)? \piso.data_r [1179] : 
                      (N100)? \piso.data_r [1211] : 
                      (N102)? \piso.data_r [1243] : 
                      (N104)? \piso.data_r [1275] : 
                      (N106)? \piso.data_r [1307] : 
                      (N108)? \piso.data_r [1339] : 
                      (N110)? \piso.data_r [1371] : 
                      (N112)? \piso.data_r [1403] : 
                      (N114)? \piso.data_r [1435] : 
                      (N116)? \piso.data_r [1467] : 
                      (N118)? \piso.data_r [1499] : 
                      (N120)? \piso.data_r [1531] : 
                      (N122)? \piso.data_r [1563] : 
                      (N124)? \piso.data_r [1595] : 
                      (N126)? \piso.data_r [1627] : 
                      (N128)? \piso.data_r [1659] : 
                      (N130)? \piso.data_r [1691] : 
                      (N132)? \piso.data_r [1723] : 
                      (N134)? \piso.data_r [1755] : 
                      (N136)? \piso.data_r [1787] : 
                      (N138)? \piso.data_r [1819] : 
                      (N140)? \piso.data_r [1851] : 
                      (N142)? \piso.data_r [1883] : 
                      (N144)? \piso.data_r [1915] : 
                      (N146)? \piso.data_r [1947] : 
                      (N148)? \piso.data_r [1979] : 
                      (N150)? \piso.data_r [2011] : 
                      (N152)? \piso.data_r [2043] : 1'b0;
  assign data_o[26] = (N89)? \piso.data_r [26] : 
                      (N91)? \piso.data_r [58] : 
                      (N93)? \piso.data_r [90] : 
                      (N95)? \piso.data_r [122] : 
                      (N97)? \piso.data_r [154] : 
                      (N99)? \piso.data_r [186] : 
                      (N101)? \piso.data_r [218] : 
                      (N103)? \piso.data_r [250] : 
                      (N105)? \piso.data_r [282] : 
                      (N107)? \piso.data_r [314] : 
                      (N109)? \piso.data_r [346] : 
                      (N111)? \piso.data_r [378] : 
                      (N113)? \piso.data_r [410] : 
                      (N115)? \piso.data_r [442] : 
                      (N117)? \piso.data_r [474] : 
                      (N119)? \piso.data_r [506] : 
                      (N121)? \piso.data_r [538] : 
                      (N123)? \piso.data_r [570] : 
                      (N125)? \piso.data_r [602] : 
                      (N127)? \piso.data_r [634] : 
                      (N129)? \piso.data_r [666] : 
                      (N131)? \piso.data_r [698] : 
                      (N133)? \piso.data_r [730] : 
                      (N135)? \piso.data_r [762] : 
                      (N137)? \piso.data_r [794] : 
                      (N139)? \piso.data_r [826] : 
                      (N141)? \piso.data_r [858] : 
                      (N143)? \piso.data_r [890] : 
                      (N145)? \piso.data_r [922] : 
                      (N147)? \piso.data_r [954] : 
                      (N149)? \piso.data_r [986] : 
                      (N151)? \piso.data_r [1018] : 
                      (N90)? \piso.data_r [1050] : 
                      (N92)? \piso.data_r [1082] : 
                      (N94)? \piso.data_r [1114] : 
                      (N96)? \piso.data_r [1146] : 
                      (N98)? \piso.data_r [1178] : 
                      (N100)? \piso.data_r [1210] : 
                      (N102)? \piso.data_r [1242] : 
                      (N104)? \piso.data_r [1274] : 
                      (N106)? \piso.data_r [1306] : 
                      (N108)? \piso.data_r [1338] : 
                      (N110)? \piso.data_r [1370] : 
                      (N112)? \piso.data_r [1402] : 
                      (N114)? \piso.data_r [1434] : 
                      (N116)? \piso.data_r [1466] : 
                      (N118)? \piso.data_r [1498] : 
                      (N120)? \piso.data_r [1530] : 
                      (N122)? \piso.data_r [1562] : 
                      (N124)? \piso.data_r [1594] : 
                      (N126)? \piso.data_r [1626] : 
                      (N128)? \piso.data_r [1658] : 
                      (N130)? \piso.data_r [1690] : 
                      (N132)? \piso.data_r [1722] : 
                      (N134)? \piso.data_r [1754] : 
                      (N136)? \piso.data_r [1786] : 
                      (N138)? \piso.data_r [1818] : 
                      (N140)? \piso.data_r [1850] : 
                      (N142)? \piso.data_r [1882] : 
                      (N144)? \piso.data_r [1914] : 
                      (N146)? \piso.data_r [1946] : 
                      (N148)? \piso.data_r [1978] : 
                      (N150)? \piso.data_r [2010] : 
                      (N152)? \piso.data_r [2042] : 1'b0;
  assign data_o[25] = (N89)? \piso.data_r [25] : 
                      (N91)? \piso.data_r [57] : 
                      (N93)? \piso.data_r [89] : 
                      (N95)? \piso.data_r [121] : 
                      (N97)? \piso.data_r [153] : 
                      (N99)? \piso.data_r [185] : 
                      (N101)? \piso.data_r [217] : 
                      (N103)? \piso.data_r [249] : 
                      (N105)? \piso.data_r [281] : 
                      (N107)? \piso.data_r [313] : 
                      (N109)? \piso.data_r [345] : 
                      (N111)? \piso.data_r [377] : 
                      (N113)? \piso.data_r [409] : 
                      (N115)? \piso.data_r [441] : 
                      (N117)? \piso.data_r [473] : 
                      (N119)? \piso.data_r [505] : 
                      (N121)? \piso.data_r [537] : 
                      (N123)? \piso.data_r [569] : 
                      (N125)? \piso.data_r [601] : 
                      (N127)? \piso.data_r [633] : 
                      (N129)? \piso.data_r [665] : 
                      (N131)? \piso.data_r [697] : 
                      (N133)? \piso.data_r [729] : 
                      (N135)? \piso.data_r [761] : 
                      (N137)? \piso.data_r [793] : 
                      (N139)? \piso.data_r [825] : 
                      (N141)? \piso.data_r [857] : 
                      (N143)? \piso.data_r [889] : 
                      (N145)? \piso.data_r [921] : 
                      (N147)? \piso.data_r [953] : 
                      (N149)? \piso.data_r [985] : 
                      (N151)? \piso.data_r [1017] : 
                      (N90)? \piso.data_r [1049] : 
                      (N92)? \piso.data_r [1081] : 
                      (N94)? \piso.data_r [1113] : 
                      (N96)? \piso.data_r [1145] : 
                      (N98)? \piso.data_r [1177] : 
                      (N100)? \piso.data_r [1209] : 
                      (N102)? \piso.data_r [1241] : 
                      (N104)? \piso.data_r [1273] : 
                      (N106)? \piso.data_r [1305] : 
                      (N108)? \piso.data_r [1337] : 
                      (N110)? \piso.data_r [1369] : 
                      (N112)? \piso.data_r [1401] : 
                      (N114)? \piso.data_r [1433] : 
                      (N116)? \piso.data_r [1465] : 
                      (N118)? \piso.data_r [1497] : 
                      (N120)? \piso.data_r [1529] : 
                      (N122)? \piso.data_r [1561] : 
                      (N124)? \piso.data_r [1593] : 
                      (N126)? \piso.data_r [1625] : 
                      (N128)? \piso.data_r [1657] : 
                      (N130)? \piso.data_r [1689] : 
                      (N132)? \piso.data_r [1721] : 
                      (N134)? \piso.data_r [1753] : 
                      (N136)? \piso.data_r [1785] : 
                      (N138)? \piso.data_r [1817] : 
                      (N140)? \piso.data_r [1849] : 
                      (N142)? \piso.data_r [1881] : 
                      (N144)? \piso.data_r [1913] : 
                      (N146)? \piso.data_r [1945] : 
                      (N148)? \piso.data_r [1977] : 
                      (N150)? \piso.data_r [2009] : 
                      (N152)? \piso.data_r [2041] : 1'b0;
  assign data_o[24] = (N89)? \piso.data_r [24] : 
                      (N91)? \piso.data_r [56] : 
                      (N93)? \piso.data_r [88] : 
                      (N95)? \piso.data_r [120] : 
                      (N97)? \piso.data_r [152] : 
                      (N99)? \piso.data_r [184] : 
                      (N101)? \piso.data_r [216] : 
                      (N103)? \piso.data_r [248] : 
                      (N105)? \piso.data_r [280] : 
                      (N107)? \piso.data_r [312] : 
                      (N109)? \piso.data_r [344] : 
                      (N111)? \piso.data_r [376] : 
                      (N113)? \piso.data_r [408] : 
                      (N115)? \piso.data_r [440] : 
                      (N117)? \piso.data_r [472] : 
                      (N119)? \piso.data_r [504] : 
                      (N121)? \piso.data_r [536] : 
                      (N123)? \piso.data_r [568] : 
                      (N125)? \piso.data_r [600] : 
                      (N127)? \piso.data_r [632] : 
                      (N129)? \piso.data_r [664] : 
                      (N131)? \piso.data_r [696] : 
                      (N133)? \piso.data_r [728] : 
                      (N135)? \piso.data_r [760] : 
                      (N137)? \piso.data_r [792] : 
                      (N139)? \piso.data_r [824] : 
                      (N141)? \piso.data_r [856] : 
                      (N143)? \piso.data_r [888] : 
                      (N145)? \piso.data_r [920] : 
                      (N147)? \piso.data_r [952] : 
                      (N149)? \piso.data_r [984] : 
                      (N151)? \piso.data_r [1016] : 
                      (N90)? \piso.data_r [1048] : 
                      (N92)? \piso.data_r [1080] : 
                      (N94)? \piso.data_r [1112] : 
                      (N96)? \piso.data_r [1144] : 
                      (N98)? \piso.data_r [1176] : 
                      (N100)? \piso.data_r [1208] : 
                      (N102)? \piso.data_r [1240] : 
                      (N104)? \piso.data_r [1272] : 
                      (N106)? \piso.data_r [1304] : 
                      (N108)? \piso.data_r [1336] : 
                      (N110)? \piso.data_r [1368] : 
                      (N112)? \piso.data_r [1400] : 
                      (N114)? \piso.data_r [1432] : 
                      (N116)? \piso.data_r [1464] : 
                      (N118)? \piso.data_r [1496] : 
                      (N120)? \piso.data_r [1528] : 
                      (N122)? \piso.data_r [1560] : 
                      (N124)? \piso.data_r [1592] : 
                      (N126)? \piso.data_r [1624] : 
                      (N128)? \piso.data_r [1656] : 
                      (N130)? \piso.data_r [1688] : 
                      (N132)? \piso.data_r [1720] : 
                      (N134)? \piso.data_r [1752] : 
                      (N136)? \piso.data_r [1784] : 
                      (N138)? \piso.data_r [1816] : 
                      (N140)? \piso.data_r [1848] : 
                      (N142)? \piso.data_r [1880] : 
                      (N144)? \piso.data_r [1912] : 
                      (N146)? \piso.data_r [1944] : 
                      (N148)? \piso.data_r [1976] : 
                      (N150)? \piso.data_r [2008] : 
                      (N152)? \piso.data_r [2040] : 1'b0;
  assign data_o[23] = (N89)? \piso.data_r [23] : 
                      (N91)? \piso.data_r [55] : 
                      (N93)? \piso.data_r [87] : 
                      (N95)? \piso.data_r [119] : 
                      (N97)? \piso.data_r [151] : 
                      (N99)? \piso.data_r [183] : 
                      (N101)? \piso.data_r [215] : 
                      (N103)? \piso.data_r [247] : 
                      (N105)? \piso.data_r [279] : 
                      (N107)? \piso.data_r [311] : 
                      (N109)? \piso.data_r [343] : 
                      (N111)? \piso.data_r [375] : 
                      (N113)? \piso.data_r [407] : 
                      (N115)? \piso.data_r [439] : 
                      (N117)? \piso.data_r [471] : 
                      (N119)? \piso.data_r [503] : 
                      (N121)? \piso.data_r [535] : 
                      (N123)? \piso.data_r [567] : 
                      (N125)? \piso.data_r [599] : 
                      (N127)? \piso.data_r [631] : 
                      (N129)? \piso.data_r [663] : 
                      (N131)? \piso.data_r [695] : 
                      (N133)? \piso.data_r [727] : 
                      (N135)? \piso.data_r [759] : 
                      (N137)? \piso.data_r [791] : 
                      (N139)? \piso.data_r [823] : 
                      (N141)? \piso.data_r [855] : 
                      (N143)? \piso.data_r [887] : 
                      (N145)? \piso.data_r [919] : 
                      (N147)? \piso.data_r [951] : 
                      (N149)? \piso.data_r [983] : 
                      (N151)? \piso.data_r [1015] : 
                      (N90)? \piso.data_r [1047] : 
                      (N92)? \piso.data_r [1079] : 
                      (N94)? \piso.data_r [1111] : 
                      (N96)? \piso.data_r [1143] : 
                      (N98)? \piso.data_r [1175] : 
                      (N100)? \piso.data_r [1207] : 
                      (N102)? \piso.data_r [1239] : 
                      (N104)? \piso.data_r [1271] : 
                      (N106)? \piso.data_r [1303] : 
                      (N108)? \piso.data_r [1335] : 
                      (N110)? \piso.data_r [1367] : 
                      (N112)? \piso.data_r [1399] : 
                      (N114)? \piso.data_r [1431] : 
                      (N116)? \piso.data_r [1463] : 
                      (N118)? \piso.data_r [1495] : 
                      (N120)? \piso.data_r [1527] : 
                      (N122)? \piso.data_r [1559] : 
                      (N124)? \piso.data_r [1591] : 
                      (N126)? \piso.data_r [1623] : 
                      (N128)? \piso.data_r [1655] : 
                      (N130)? \piso.data_r [1687] : 
                      (N132)? \piso.data_r [1719] : 
                      (N134)? \piso.data_r [1751] : 
                      (N136)? \piso.data_r [1783] : 
                      (N138)? \piso.data_r [1815] : 
                      (N140)? \piso.data_r [1847] : 
                      (N142)? \piso.data_r [1879] : 
                      (N144)? \piso.data_r [1911] : 
                      (N146)? \piso.data_r [1943] : 
                      (N148)? \piso.data_r [1975] : 
                      (N150)? \piso.data_r [2007] : 
                      (N152)? \piso.data_r [2039] : 1'b0;
  assign data_o[22] = (N89)? \piso.data_r [22] : 
                      (N91)? \piso.data_r [54] : 
                      (N93)? \piso.data_r [86] : 
                      (N95)? \piso.data_r [118] : 
                      (N97)? \piso.data_r [150] : 
                      (N99)? \piso.data_r [182] : 
                      (N101)? \piso.data_r [214] : 
                      (N103)? \piso.data_r [246] : 
                      (N105)? \piso.data_r [278] : 
                      (N107)? \piso.data_r [310] : 
                      (N109)? \piso.data_r [342] : 
                      (N111)? \piso.data_r [374] : 
                      (N113)? \piso.data_r [406] : 
                      (N115)? \piso.data_r [438] : 
                      (N117)? \piso.data_r [470] : 
                      (N119)? \piso.data_r [502] : 
                      (N121)? \piso.data_r [534] : 
                      (N123)? \piso.data_r [566] : 
                      (N125)? \piso.data_r [598] : 
                      (N127)? \piso.data_r [630] : 
                      (N129)? \piso.data_r [662] : 
                      (N131)? \piso.data_r [694] : 
                      (N133)? \piso.data_r [726] : 
                      (N135)? \piso.data_r [758] : 
                      (N137)? \piso.data_r [790] : 
                      (N139)? \piso.data_r [822] : 
                      (N141)? \piso.data_r [854] : 
                      (N143)? \piso.data_r [886] : 
                      (N145)? \piso.data_r [918] : 
                      (N147)? \piso.data_r [950] : 
                      (N149)? \piso.data_r [982] : 
                      (N151)? \piso.data_r [1014] : 
                      (N90)? \piso.data_r [1046] : 
                      (N92)? \piso.data_r [1078] : 
                      (N94)? \piso.data_r [1110] : 
                      (N96)? \piso.data_r [1142] : 
                      (N98)? \piso.data_r [1174] : 
                      (N100)? \piso.data_r [1206] : 
                      (N102)? \piso.data_r [1238] : 
                      (N104)? \piso.data_r [1270] : 
                      (N106)? \piso.data_r [1302] : 
                      (N108)? \piso.data_r [1334] : 
                      (N110)? \piso.data_r [1366] : 
                      (N112)? \piso.data_r [1398] : 
                      (N114)? \piso.data_r [1430] : 
                      (N116)? \piso.data_r [1462] : 
                      (N118)? \piso.data_r [1494] : 
                      (N120)? \piso.data_r [1526] : 
                      (N122)? \piso.data_r [1558] : 
                      (N124)? \piso.data_r [1590] : 
                      (N126)? \piso.data_r [1622] : 
                      (N128)? \piso.data_r [1654] : 
                      (N130)? \piso.data_r [1686] : 
                      (N132)? \piso.data_r [1718] : 
                      (N134)? \piso.data_r [1750] : 
                      (N136)? \piso.data_r [1782] : 
                      (N138)? \piso.data_r [1814] : 
                      (N140)? \piso.data_r [1846] : 
                      (N142)? \piso.data_r [1878] : 
                      (N144)? \piso.data_r [1910] : 
                      (N146)? \piso.data_r [1942] : 
                      (N148)? \piso.data_r [1974] : 
                      (N150)? \piso.data_r [2006] : 
                      (N152)? \piso.data_r [2038] : 1'b0;
  assign data_o[21] = (N89)? \piso.data_r [21] : 
                      (N91)? \piso.data_r [53] : 
                      (N93)? \piso.data_r [85] : 
                      (N95)? \piso.data_r [117] : 
                      (N97)? \piso.data_r [149] : 
                      (N99)? \piso.data_r [181] : 
                      (N101)? \piso.data_r [213] : 
                      (N103)? \piso.data_r [245] : 
                      (N105)? \piso.data_r [277] : 
                      (N107)? \piso.data_r [309] : 
                      (N109)? \piso.data_r [341] : 
                      (N111)? \piso.data_r [373] : 
                      (N113)? \piso.data_r [405] : 
                      (N115)? \piso.data_r [437] : 
                      (N117)? \piso.data_r [469] : 
                      (N119)? \piso.data_r [501] : 
                      (N121)? \piso.data_r [533] : 
                      (N123)? \piso.data_r [565] : 
                      (N125)? \piso.data_r [597] : 
                      (N127)? \piso.data_r [629] : 
                      (N129)? \piso.data_r [661] : 
                      (N131)? \piso.data_r [693] : 
                      (N133)? \piso.data_r [725] : 
                      (N135)? \piso.data_r [757] : 
                      (N137)? \piso.data_r [789] : 
                      (N139)? \piso.data_r [821] : 
                      (N141)? \piso.data_r [853] : 
                      (N143)? \piso.data_r [885] : 
                      (N145)? \piso.data_r [917] : 
                      (N147)? \piso.data_r [949] : 
                      (N149)? \piso.data_r [981] : 
                      (N151)? \piso.data_r [1013] : 
                      (N90)? \piso.data_r [1045] : 
                      (N92)? \piso.data_r [1077] : 
                      (N94)? \piso.data_r [1109] : 
                      (N96)? \piso.data_r [1141] : 
                      (N98)? \piso.data_r [1173] : 
                      (N100)? \piso.data_r [1205] : 
                      (N102)? \piso.data_r [1237] : 
                      (N104)? \piso.data_r [1269] : 
                      (N106)? \piso.data_r [1301] : 
                      (N108)? \piso.data_r [1333] : 
                      (N110)? \piso.data_r [1365] : 
                      (N112)? \piso.data_r [1397] : 
                      (N114)? \piso.data_r [1429] : 
                      (N116)? \piso.data_r [1461] : 
                      (N118)? \piso.data_r [1493] : 
                      (N120)? \piso.data_r [1525] : 
                      (N122)? \piso.data_r [1557] : 
                      (N124)? \piso.data_r [1589] : 
                      (N126)? \piso.data_r [1621] : 
                      (N128)? \piso.data_r [1653] : 
                      (N130)? \piso.data_r [1685] : 
                      (N132)? \piso.data_r [1717] : 
                      (N134)? \piso.data_r [1749] : 
                      (N136)? \piso.data_r [1781] : 
                      (N138)? \piso.data_r [1813] : 
                      (N140)? \piso.data_r [1845] : 
                      (N142)? \piso.data_r [1877] : 
                      (N144)? \piso.data_r [1909] : 
                      (N146)? \piso.data_r [1941] : 
                      (N148)? \piso.data_r [1973] : 
                      (N150)? \piso.data_r [2005] : 
                      (N152)? \piso.data_r [2037] : 1'b0;
  assign data_o[20] = (N89)? \piso.data_r [20] : 
                      (N91)? \piso.data_r [52] : 
                      (N93)? \piso.data_r [84] : 
                      (N95)? \piso.data_r [116] : 
                      (N97)? \piso.data_r [148] : 
                      (N99)? \piso.data_r [180] : 
                      (N101)? \piso.data_r [212] : 
                      (N103)? \piso.data_r [244] : 
                      (N105)? \piso.data_r [276] : 
                      (N107)? \piso.data_r [308] : 
                      (N109)? \piso.data_r [340] : 
                      (N111)? \piso.data_r [372] : 
                      (N113)? \piso.data_r [404] : 
                      (N115)? \piso.data_r [436] : 
                      (N117)? \piso.data_r [468] : 
                      (N119)? \piso.data_r [500] : 
                      (N121)? \piso.data_r [532] : 
                      (N123)? \piso.data_r [564] : 
                      (N125)? \piso.data_r [596] : 
                      (N127)? \piso.data_r [628] : 
                      (N129)? \piso.data_r [660] : 
                      (N131)? \piso.data_r [692] : 
                      (N133)? \piso.data_r [724] : 
                      (N135)? \piso.data_r [756] : 
                      (N137)? \piso.data_r [788] : 
                      (N139)? \piso.data_r [820] : 
                      (N141)? \piso.data_r [852] : 
                      (N143)? \piso.data_r [884] : 
                      (N145)? \piso.data_r [916] : 
                      (N147)? \piso.data_r [948] : 
                      (N149)? \piso.data_r [980] : 
                      (N151)? \piso.data_r [1012] : 
                      (N90)? \piso.data_r [1044] : 
                      (N92)? \piso.data_r [1076] : 
                      (N94)? \piso.data_r [1108] : 
                      (N96)? \piso.data_r [1140] : 
                      (N98)? \piso.data_r [1172] : 
                      (N100)? \piso.data_r [1204] : 
                      (N102)? \piso.data_r [1236] : 
                      (N104)? \piso.data_r [1268] : 
                      (N106)? \piso.data_r [1300] : 
                      (N108)? \piso.data_r [1332] : 
                      (N110)? \piso.data_r [1364] : 
                      (N112)? \piso.data_r [1396] : 
                      (N114)? \piso.data_r [1428] : 
                      (N116)? \piso.data_r [1460] : 
                      (N118)? \piso.data_r [1492] : 
                      (N120)? \piso.data_r [1524] : 
                      (N122)? \piso.data_r [1556] : 
                      (N124)? \piso.data_r [1588] : 
                      (N126)? \piso.data_r [1620] : 
                      (N128)? \piso.data_r [1652] : 
                      (N130)? \piso.data_r [1684] : 
                      (N132)? \piso.data_r [1716] : 
                      (N134)? \piso.data_r [1748] : 
                      (N136)? \piso.data_r [1780] : 
                      (N138)? \piso.data_r [1812] : 
                      (N140)? \piso.data_r [1844] : 
                      (N142)? \piso.data_r [1876] : 
                      (N144)? \piso.data_r [1908] : 
                      (N146)? \piso.data_r [1940] : 
                      (N148)? \piso.data_r [1972] : 
                      (N150)? \piso.data_r [2004] : 
                      (N152)? \piso.data_r [2036] : 1'b0;
  assign data_o[19] = (N89)? \piso.data_r [19] : 
                      (N91)? \piso.data_r [51] : 
                      (N93)? \piso.data_r [83] : 
                      (N95)? \piso.data_r [115] : 
                      (N97)? \piso.data_r [147] : 
                      (N99)? \piso.data_r [179] : 
                      (N101)? \piso.data_r [211] : 
                      (N103)? \piso.data_r [243] : 
                      (N105)? \piso.data_r [275] : 
                      (N107)? \piso.data_r [307] : 
                      (N109)? \piso.data_r [339] : 
                      (N111)? \piso.data_r [371] : 
                      (N113)? \piso.data_r [403] : 
                      (N115)? \piso.data_r [435] : 
                      (N117)? \piso.data_r [467] : 
                      (N119)? \piso.data_r [499] : 
                      (N121)? \piso.data_r [531] : 
                      (N123)? \piso.data_r [563] : 
                      (N125)? \piso.data_r [595] : 
                      (N127)? \piso.data_r [627] : 
                      (N129)? \piso.data_r [659] : 
                      (N131)? \piso.data_r [691] : 
                      (N133)? \piso.data_r [723] : 
                      (N135)? \piso.data_r [755] : 
                      (N137)? \piso.data_r [787] : 
                      (N139)? \piso.data_r [819] : 
                      (N141)? \piso.data_r [851] : 
                      (N143)? \piso.data_r [883] : 
                      (N145)? \piso.data_r [915] : 
                      (N147)? \piso.data_r [947] : 
                      (N149)? \piso.data_r [979] : 
                      (N151)? \piso.data_r [1011] : 
                      (N90)? \piso.data_r [1043] : 
                      (N92)? \piso.data_r [1075] : 
                      (N94)? \piso.data_r [1107] : 
                      (N96)? \piso.data_r [1139] : 
                      (N98)? \piso.data_r [1171] : 
                      (N100)? \piso.data_r [1203] : 
                      (N102)? \piso.data_r [1235] : 
                      (N104)? \piso.data_r [1267] : 
                      (N106)? \piso.data_r [1299] : 
                      (N108)? \piso.data_r [1331] : 
                      (N110)? \piso.data_r [1363] : 
                      (N112)? \piso.data_r [1395] : 
                      (N114)? \piso.data_r [1427] : 
                      (N116)? \piso.data_r [1459] : 
                      (N118)? \piso.data_r [1491] : 
                      (N120)? \piso.data_r [1523] : 
                      (N122)? \piso.data_r [1555] : 
                      (N124)? \piso.data_r [1587] : 
                      (N126)? \piso.data_r [1619] : 
                      (N128)? \piso.data_r [1651] : 
                      (N130)? \piso.data_r [1683] : 
                      (N132)? \piso.data_r [1715] : 
                      (N134)? \piso.data_r [1747] : 
                      (N136)? \piso.data_r [1779] : 
                      (N138)? \piso.data_r [1811] : 
                      (N140)? \piso.data_r [1843] : 
                      (N142)? \piso.data_r [1875] : 
                      (N144)? \piso.data_r [1907] : 
                      (N146)? \piso.data_r [1939] : 
                      (N148)? \piso.data_r [1971] : 
                      (N150)? \piso.data_r [2003] : 
                      (N152)? \piso.data_r [2035] : 1'b0;
  assign data_o[18] = (N89)? \piso.data_r [18] : 
                      (N91)? \piso.data_r [50] : 
                      (N93)? \piso.data_r [82] : 
                      (N95)? \piso.data_r [114] : 
                      (N97)? \piso.data_r [146] : 
                      (N99)? \piso.data_r [178] : 
                      (N101)? \piso.data_r [210] : 
                      (N103)? \piso.data_r [242] : 
                      (N105)? \piso.data_r [274] : 
                      (N107)? \piso.data_r [306] : 
                      (N109)? \piso.data_r [338] : 
                      (N111)? \piso.data_r [370] : 
                      (N113)? \piso.data_r [402] : 
                      (N115)? \piso.data_r [434] : 
                      (N117)? \piso.data_r [466] : 
                      (N119)? \piso.data_r [498] : 
                      (N121)? \piso.data_r [530] : 
                      (N123)? \piso.data_r [562] : 
                      (N125)? \piso.data_r [594] : 
                      (N127)? \piso.data_r [626] : 
                      (N129)? \piso.data_r [658] : 
                      (N131)? \piso.data_r [690] : 
                      (N133)? \piso.data_r [722] : 
                      (N135)? \piso.data_r [754] : 
                      (N137)? \piso.data_r [786] : 
                      (N139)? \piso.data_r [818] : 
                      (N141)? \piso.data_r [850] : 
                      (N143)? \piso.data_r [882] : 
                      (N145)? \piso.data_r [914] : 
                      (N147)? \piso.data_r [946] : 
                      (N149)? \piso.data_r [978] : 
                      (N151)? \piso.data_r [1010] : 
                      (N90)? \piso.data_r [1042] : 
                      (N92)? \piso.data_r [1074] : 
                      (N94)? \piso.data_r [1106] : 
                      (N96)? \piso.data_r [1138] : 
                      (N98)? \piso.data_r [1170] : 
                      (N100)? \piso.data_r [1202] : 
                      (N102)? \piso.data_r [1234] : 
                      (N104)? \piso.data_r [1266] : 
                      (N106)? \piso.data_r [1298] : 
                      (N108)? \piso.data_r [1330] : 
                      (N110)? \piso.data_r [1362] : 
                      (N112)? \piso.data_r [1394] : 
                      (N114)? \piso.data_r [1426] : 
                      (N116)? \piso.data_r [1458] : 
                      (N118)? \piso.data_r [1490] : 
                      (N120)? \piso.data_r [1522] : 
                      (N122)? \piso.data_r [1554] : 
                      (N124)? \piso.data_r [1586] : 
                      (N126)? \piso.data_r [1618] : 
                      (N128)? \piso.data_r [1650] : 
                      (N130)? \piso.data_r [1682] : 
                      (N132)? \piso.data_r [1714] : 
                      (N134)? \piso.data_r [1746] : 
                      (N136)? \piso.data_r [1778] : 
                      (N138)? \piso.data_r [1810] : 
                      (N140)? \piso.data_r [1842] : 
                      (N142)? \piso.data_r [1874] : 
                      (N144)? \piso.data_r [1906] : 
                      (N146)? \piso.data_r [1938] : 
                      (N148)? \piso.data_r [1970] : 
                      (N150)? \piso.data_r [2002] : 
                      (N152)? \piso.data_r [2034] : 1'b0;
  assign data_o[17] = (N89)? \piso.data_r [17] : 
                      (N91)? \piso.data_r [49] : 
                      (N93)? \piso.data_r [81] : 
                      (N95)? \piso.data_r [113] : 
                      (N97)? \piso.data_r [145] : 
                      (N99)? \piso.data_r [177] : 
                      (N101)? \piso.data_r [209] : 
                      (N103)? \piso.data_r [241] : 
                      (N105)? \piso.data_r [273] : 
                      (N107)? \piso.data_r [305] : 
                      (N109)? \piso.data_r [337] : 
                      (N111)? \piso.data_r [369] : 
                      (N113)? \piso.data_r [401] : 
                      (N115)? \piso.data_r [433] : 
                      (N117)? \piso.data_r [465] : 
                      (N119)? \piso.data_r [497] : 
                      (N121)? \piso.data_r [529] : 
                      (N123)? \piso.data_r [561] : 
                      (N125)? \piso.data_r [593] : 
                      (N127)? \piso.data_r [625] : 
                      (N129)? \piso.data_r [657] : 
                      (N131)? \piso.data_r [689] : 
                      (N133)? \piso.data_r [721] : 
                      (N135)? \piso.data_r [753] : 
                      (N137)? \piso.data_r [785] : 
                      (N139)? \piso.data_r [817] : 
                      (N141)? \piso.data_r [849] : 
                      (N143)? \piso.data_r [881] : 
                      (N145)? \piso.data_r [913] : 
                      (N147)? \piso.data_r [945] : 
                      (N149)? \piso.data_r [977] : 
                      (N151)? \piso.data_r [1009] : 
                      (N90)? \piso.data_r [1041] : 
                      (N92)? \piso.data_r [1073] : 
                      (N94)? \piso.data_r [1105] : 
                      (N96)? \piso.data_r [1137] : 
                      (N98)? \piso.data_r [1169] : 
                      (N100)? \piso.data_r [1201] : 
                      (N102)? \piso.data_r [1233] : 
                      (N104)? \piso.data_r [1265] : 
                      (N106)? \piso.data_r [1297] : 
                      (N108)? \piso.data_r [1329] : 
                      (N110)? \piso.data_r [1361] : 
                      (N112)? \piso.data_r [1393] : 
                      (N114)? \piso.data_r [1425] : 
                      (N116)? \piso.data_r [1457] : 
                      (N118)? \piso.data_r [1489] : 
                      (N120)? \piso.data_r [1521] : 
                      (N122)? \piso.data_r [1553] : 
                      (N124)? \piso.data_r [1585] : 
                      (N126)? \piso.data_r [1617] : 
                      (N128)? \piso.data_r [1649] : 
                      (N130)? \piso.data_r [1681] : 
                      (N132)? \piso.data_r [1713] : 
                      (N134)? \piso.data_r [1745] : 
                      (N136)? \piso.data_r [1777] : 
                      (N138)? \piso.data_r [1809] : 
                      (N140)? \piso.data_r [1841] : 
                      (N142)? \piso.data_r [1873] : 
                      (N144)? \piso.data_r [1905] : 
                      (N146)? \piso.data_r [1937] : 
                      (N148)? \piso.data_r [1969] : 
                      (N150)? \piso.data_r [2001] : 
                      (N152)? \piso.data_r [2033] : 1'b0;
  assign data_o[16] = (N89)? \piso.data_r [16] : 
                      (N91)? \piso.data_r [48] : 
                      (N93)? \piso.data_r [80] : 
                      (N95)? \piso.data_r [112] : 
                      (N97)? \piso.data_r [144] : 
                      (N99)? \piso.data_r [176] : 
                      (N101)? \piso.data_r [208] : 
                      (N103)? \piso.data_r [240] : 
                      (N105)? \piso.data_r [272] : 
                      (N107)? \piso.data_r [304] : 
                      (N109)? \piso.data_r [336] : 
                      (N111)? \piso.data_r [368] : 
                      (N113)? \piso.data_r [400] : 
                      (N115)? \piso.data_r [432] : 
                      (N117)? \piso.data_r [464] : 
                      (N119)? \piso.data_r [496] : 
                      (N121)? \piso.data_r [528] : 
                      (N123)? \piso.data_r [560] : 
                      (N125)? \piso.data_r [592] : 
                      (N127)? \piso.data_r [624] : 
                      (N129)? \piso.data_r [656] : 
                      (N131)? \piso.data_r [688] : 
                      (N133)? \piso.data_r [720] : 
                      (N135)? \piso.data_r [752] : 
                      (N137)? \piso.data_r [784] : 
                      (N139)? \piso.data_r [816] : 
                      (N141)? \piso.data_r [848] : 
                      (N143)? \piso.data_r [880] : 
                      (N145)? \piso.data_r [912] : 
                      (N147)? \piso.data_r [944] : 
                      (N149)? \piso.data_r [976] : 
                      (N151)? \piso.data_r [1008] : 
                      (N90)? \piso.data_r [1040] : 
                      (N92)? \piso.data_r [1072] : 
                      (N94)? \piso.data_r [1104] : 
                      (N96)? \piso.data_r [1136] : 
                      (N98)? \piso.data_r [1168] : 
                      (N100)? \piso.data_r [1200] : 
                      (N102)? \piso.data_r [1232] : 
                      (N104)? \piso.data_r [1264] : 
                      (N106)? \piso.data_r [1296] : 
                      (N108)? \piso.data_r [1328] : 
                      (N110)? \piso.data_r [1360] : 
                      (N112)? \piso.data_r [1392] : 
                      (N114)? \piso.data_r [1424] : 
                      (N116)? \piso.data_r [1456] : 
                      (N118)? \piso.data_r [1488] : 
                      (N120)? \piso.data_r [1520] : 
                      (N122)? \piso.data_r [1552] : 
                      (N124)? \piso.data_r [1584] : 
                      (N126)? \piso.data_r [1616] : 
                      (N128)? \piso.data_r [1648] : 
                      (N130)? \piso.data_r [1680] : 
                      (N132)? \piso.data_r [1712] : 
                      (N134)? \piso.data_r [1744] : 
                      (N136)? \piso.data_r [1776] : 
                      (N138)? \piso.data_r [1808] : 
                      (N140)? \piso.data_r [1840] : 
                      (N142)? \piso.data_r [1872] : 
                      (N144)? \piso.data_r [1904] : 
                      (N146)? \piso.data_r [1936] : 
                      (N148)? \piso.data_r [1968] : 
                      (N150)? \piso.data_r [2000] : 
                      (N152)? \piso.data_r [2032] : 1'b0;
  assign data_o[15] = (N89)? \piso.data_r [15] : 
                      (N91)? \piso.data_r [47] : 
                      (N93)? \piso.data_r [79] : 
                      (N95)? \piso.data_r [111] : 
                      (N97)? \piso.data_r [143] : 
                      (N99)? \piso.data_r [175] : 
                      (N101)? \piso.data_r [207] : 
                      (N103)? \piso.data_r [239] : 
                      (N105)? \piso.data_r [271] : 
                      (N107)? \piso.data_r [303] : 
                      (N109)? \piso.data_r [335] : 
                      (N111)? \piso.data_r [367] : 
                      (N113)? \piso.data_r [399] : 
                      (N115)? \piso.data_r [431] : 
                      (N117)? \piso.data_r [463] : 
                      (N119)? \piso.data_r [495] : 
                      (N121)? \piso.data_r [527] : 
                      (N123)? \piso.data_r [559] : 
                      (N125)? \piso.data_r [591] : 
                      (N127)? \piso.data_r [623] : 
                      (N129)? \piso.data_r [655] : 
                      (N131)? \piso.data_r [687] : 
                      (N133)? \piso.data_r [719] : 
                      (N135)? \piso.data_r [751] : 
                      (N137)? \piso.data_r [783] : 
                      (N139)? \piso.data_r [815] : 
                      (N141)? \piso.data_r [847] : 
                      (N143)? \piso.data_r [879] : 
                      (N145)? \piso.data_r [911] : 
                      (N147)? \piso.data_r [943] : 
                      (N149)? \piso.data_r [975] : 
                      (N151)? \piso.data_r [1007] : 
                      (N90)? \piso.data_r [1039] : 
                      (N92)? \piso.data_r [1071] : 
                      (N94)? \piso.data_r [1103] : 
                      (N96)? \piso.data_r [1135] : 
                      (N98)? \piso.data_r [1167] : 
                      (N100)? \piso.data_r [1199] : 
                      (N102)? \piso.data_r [1231] : 
                      (N104)? \piso.data_r [1263] : 
                      (N106)? \piso.data_r [1295] : 
                      (N108)? \piso.data_r [1327] : 
                      (N110)? \piso.data_r [1359] : 
                      (N112)? \piso.data_r [1391] : 
                      (N114)? \piso.data_r [1423] : 
                      (N116)? \piso.data_r [1455] : 
                      (N118)? \piso.data_r [1487] : 
                      (N120)? \piso.data_r [1519] : 
                      (N122)? \piso.data_r [1551] : 
                      (N124)? \piso.data_r [1583] : 
                      (N126)? \piso.data_r [1615] : 
                      (N128)? \piso.data_r [1647] : 
                      (N130)? \piso.data_r [1679] : 
                      (N132)? \piso.data_r [1711] : 
                      (N134)? \piso.data_r [1743] : 
                      (N136)? \piso.data_r [1775] : 
                      (N138)? \piso.data_r [1807] : 
                      (N140)? \piso.data_r [1839] : 
                      (N142)? \piso.data_r [1871] : 
                      (N144)? \piso.data_r [1903] : 
                      (N146)? \piso.data_r [1935] : 
                      (N148)? \piso.data_r [1967] : 
                      (N150)? \piso.data_r [1999] : 
                      (N152)? \piso.data_r [2031] : 1'b0;
  assign data_o[14] = (N89)? \piso.data_r [14] : 
                      (N91)? \piso.data_r [46] : 
                      (N93)? \piso.data_r [78] : 
                      (N95)? \piso.data_r [110] : 
                      (N97)? \piso.data_r [142] : 
                      (N99)? \piso.data_r [174] : 
                      (N101)? \piso.data_r [206] : 
                      (N103)? \piso.data_r [238] : 
                      (N105)? \piso.data_r [270] : 
                      (N107)? \piso.data_r [302] : 
                      (N109)? \piso.data_r [334] : 
                      (N111)? \piso.data_r [366] : 
                      (N113)? \piso.data_r [398] : 
                      (N115)? \piso.data_r [430] : 
                      (N117)? \piso.data_r [462] : 
                      (N119)? \piso.data_r [494] : 
                      (N121)? \piso.data_r [526] : 
                      (N123)? \piso.data_r [558] : 
                      (N125)? \piso.data_r [590] : 
                      (N127)? \piso.data_r [622] : 
                      (N129)? \piso.data_r [654] : 
                      (N131)? \piso.data_r [686] : 
                      (N133)? \piso.data_r [718] : 
                      (N135)? \piso.data_r [750] : 
                      (N137)? \piso.data_r [782] : 
                      (N139)? \piso.data_r [814] : 
                      (N141)? \piso.data_r [846] : 
                      (N143)? \piso.data_r [878] : 
                      (N145)? \piso.data_r [910] : 
                      (N147)? \piso.data_r [942] : 
                      (N149)? \piso.data_r [974] : 
                      (N151)? \piso.data_r [1006] : 
                      (N90)? \piso.data_r [1038] : 
                      (N92)? \piso.data_r [1070] : 
                      (N94)? \piso.data_r [1102] : 
                      (N96)? \piso.data_r [1134] : 
                      (N98)? \piso.data_r [1166] : 
                      (N100)? \piso.data_r [1198] : 
                      (N102)? \piso.data_r [1230] : 
                      (N104)? \piso.data_r [1262] : 
                      (N106)? \piso.data_r [1294] : 
                      (N108)? \piso.data_r [1326] : 
                      (N110)? \piso.data_r [1358] : 
                      (N112)? \piso.data_r [1390] : 
                      (N114)? \piso.data_r [1422] : 
                      (N116)? \piso.data_r [1454] : 
                      (N118)? \piso.data_r [1486] : 
                      (N120)? \piso.data_r [1518] : 
                      (N122)? \piso.data_r [1550] : 
                      (N124)? \piso.data_r [1582] : 
                      (N126)? \piso.data_r [1614] : 
                      (N128)? \piso.data_r [1646] : 
                      (N130)? \piso.data_r [1678] : 
                      (N132)? \piso.data_r [1710] : 
                      (N134)? \piso.data_r [1742] : 
                      (N136)? \piso.data_r [1774] : 
                      (N138)? \piso.data_r [1806] : 
                      (N140)? \piso.data_r [1838] : 
                      (N142)? \piso.data_r [1870] : 
                      (N144)? \piso.data_r [1902] : 
                      (N146)? \piso.data_r [1934] : 
                      (N148)? \piso.data_r [1966] : 
                      (N150)? \piso.data_r [1998] : 
                      (N152)? \piso.data_r [2030] : 1'b0;
  assign data_o[13] = (N89)? \piso.data_r [13] : 
                      (N91)? \piso.data_r [45] : 
                      (N93)? \piso.data_r [77] : 
                      (N95)? \piso.data_r [109] : 
                      (N97)? \piso.data_r [141] : 
                      (N99)? \piso.data_r [173] : 
                      (N101)? \piso.data_r [205] : 
                      (N103)? \piso.data_r [237] : 
                      (N105)? \piso.data_r [269] : 
                      (N107)? \piso.data_r [301] : 
                      (N109)? \piso.data_r [333] : 
                      (N111)? \piso.data_r [365] : 
                      (N113)? \piso.data_r [397] : 
                      (N115)? \piso.data_r [429] : 
                      (N117)? \piso.data_r [461] : 
                      (N119)? \piso.data_r [493] : 
                      (N121)? \piso.data_r [525] : 
                      (N123)? \piso.data_r [557] : 
                      (N125)? \piso.data_r [589] : 
                      (N127)? \piso.data_r [621] : 
                      (N129)? \piso.data_r [653] : 
                      (N131)? \piso.data_r [685] : 
                      (N133)? \piso.data_r [717] : 
                      (N135)? \piso.data_r [749] : 
                      (N137)? \piso.data_r [781] : 
                      (N139)? \piso.data_r [813] : 
                      (N141)? \piso.data_r [845] : 
                      (N143)? \piso.data_r [877] : 
                      (N145)? \piso.data_r [909] : 
                      (N147)? \piso.data_r [941] : 
                      (N149)? \piso.data_r [973] : 
                      (N151)? \piso.data_r [1005] : 
                      (N90)? \piso.data_r [1037] : 
                      (N92)? \piso.data_r [1069] : 
                      (N94)? \piso.data_r [1101] : 
                      (N96)? \piso.data_r [1133] : 
                      (N98)? \piso.data_r [1165] : 
                      (N100)? \piso.data_r [1197] : 
                      (N102)? \piso.data_r [1229] : 
                      (N104)? \piso.data_r [1261] : 
                      (N106)? \piso.data_r [1293] : 
                      (N108)? \piso.data_r [1325] : 
                      (N110)? \piso.data_r [1357] : 
                      (N112)? \piso.data_r [1389] : 
                      (N114)? \piso.data_r [1421] : 
                      (N116)? \piso.data_r [1453] : 
                      (N118)? \piso.data_r [1485] : 
                      (N120)? \piso.data_r [1517] : 
                      (N122)? \piso.data_r [1549] : 
                      (N124)? \piso.data_r [1581] : 
                      (N126)? \piso.data_r [1613] : 
                      (N128)? \piso.data_r [1645] : 
                      (N130)? \piso.data_r [1677] : 
                      (N132)? \piso.data_r [1709] : 
                      (N134)? \piso.data_r [1741] : 
                      (N136)? \piso.data_r [1773] : 
                      (N138)? \piso.data_r [1805] : 
                      (N140)? \piso.data_r [1837] : 
                      (N142)? \piso.data_r [1869] : 
                      (N144)? \piso.data_r [1901] : 
                      (N146)? \piso.data_r [1933] : 
                      (N148)? \piso.data_r [1965] : 
                      (N150)? \piso.data_r [1997] : 
                      (N152)? \piso.data_r [2029] : 1'b0;
  assign data_o[12] = (N89)? \piso.data_r [12] : 
                      (N91)? \piso.data_r [44] : 
                      (N93)? \piso.data_r [76] : 
                      (N95)? \piso.data_r [108] : 
                      (N97)? \piso.data_r [140] : 
                      (N99)? \piso.data_r [172] : 
                      (N101)? \piso.data_r [204] : 
                      (N103)? \piso.data_r [236] : 
                      (N105)? \piso.data_r [268] : 
                      (N107)? \piso.data_r [300] : 
                      (N109)? \piso.data_r [332] : 
                      (N111)? \piso.data_r [364] : 
                      (N113)? \piso.data_r [396] : 
                      (N115)? \piso.data_r [428] : 
                      (N117)? \piso.data_r [460] : 
                      (N119)? \piso.data_r [492] : 
                      (N121)? \piso.data_r [524] : 
                      (N123)? \piso.data_r [556] : 
                      (N125)? \piso.data_r [588] : 
                      (N127)? \piso.data_r [620] : 
                      (N129)? \piso.data_r [652] : 
                      (N131)? \piso.data_r [684] : 
                      (N133)? \piso.data_r [716] : 
                      (N135)? \piso.data_r [748] : 
                      (N137)? \piso.data_r [780] : 
                      (N139)? \piso.data_r [812] : 
                      (N141)? \piso.data_r [844] : 
                      (N143)? \piso.data_r [876] : 
                      (N145)? \piso.data_r [908] : 
                      (N147)? \piso.data_r [940] : 
                      (N149)? \piso.data_r [972] : 
                      (N151)? \piso.data_r [1004] : 
                      (N90)? \piso.data_r [1036] : 
                      (N92)? \piso.data_r [1068] : 
                      (N94)? \piso.data_r [1100] : 
                      (N96)? \piso.data_r [1132] : 
                      (N98)? \piso.data_r [1164] : 
                      (N100)? \piso.data_r [1196] : 
                      (N102)? \piso.data_r [1228] : 
                      (N104)? \piso.data_r [1260] : 
                      (N106)? \piso.data_r [1292] : 
                      (N108)? \piso.data_r [1324] : 
                      (N110)? \piso.data_r [1356] : 
                      (N112)? \piso.data_r [1388] : 
                      (N114)? \piso.data_r [1420] : 
                      (N116)? \piso.data_r [1452] : 
                      (N118)? \piso.data_r [1484] : 
                      (N120)? \piso.data_r [1516] : 
                      (N122)? \piso.data_r [1548] : 
                      (N124)? \piso.data_r [1580] : 
                      (N126)? \piso.data_r [1612] : 
                      (N128)? \piso.data_r [1644] : 
                      (N130)? \piso.data_r [1676] : 
                      (N132)? \piso.data_r [1708] : 
                      (N134)? \piso.data_r [1740] : 
                      (N136)? \piso.data_r [1772] : 
                      (N138)? \piso.data_r [1804] : 
                      (N140)? \piso.data_r [1836] : 
                      (N142)? \piso.data_r [1868] : 
                      (N144)? \piso.data_r [1900] : 
                      (N146)? \piso.data_r [1932] : 
                      (N148)? \piso.data_r [1964] : 
                      (N150)? \piso.data_r [1996] : 
                      (N152)? \piso.data_r [2028] : 1'b0;
  assign data_o[11] = (N89)? \piso.data_r [11] : 
                      (N91)? \piso.data_r [43] : 
                      (N93)? \piso.data_r [75] : 
                      (N95)? \piso.data_r [107] : 
                      (N97)? \piso.data_r [139] : 
                      (N99)? \piso.data_r [171] : 
                      (N101)? \piso.data_r [203] : 
                      (N103)? \piso.data_r [235] : 
                      (N105)? \piso.data_r [267] : 
                      (N107)? \piso.data_r [299] : 
                      (N109)? \piso.data_r [331] : 
                      (N111)? \piso.data_r [363] : 
                      (N113)? \piso.data_r [395] : 
                      (N115)? \piso.data_r [427] : 
                      (N117)? \piso.data_r [459] : 
                      (N119)? \piso.data_r [491] : 
                      (N121)? \piso.data_r [523] : 
                      (N123)? \piso.data_r [555] : 
                      (N125)? \piso.data_r [587] : 
                      (N127)? \piso.data_r [619] : 
                      (N129)? \piso.data_r [651] : 
                      (N131)? \piso.data_r [683] : 
                      (N133)? \piso.data_r [715] : 
                      (N135)? \piso.data_r [747] : 
                      (N137)? \piso.data_r [779] : 
                      (N139)? \piso.data_r [811] : 
                      (N141)? \piso.data_r [843] : 
                      (N143)? \piso.data_r [875] : 
                      (N145)? \piso.data_r [907] : 
                      (N147)? \piso.data_r [939] : 
                      (N149)? \piso.data_r [971] : 
                      (N151)? \piso.data_r [1003] : 
                      (N90)? \piso.data_r [1035] : 
                      (N92)? \piso.data_r [1067] : 
                      (N94)? \piso.data_r [1099] : 
                      (N96)? \piso.data_r [1131] : 
                      (N98)? \piso.data_r [1163] : 
                      (N100)? \piso.data_r [1195] : 
                      (N102)? \piso.data_r [1227] : 
                      (N104)? \piso.data_r [1259] : 
                      (N106)? \piso.data_r [1291] : 
                      (N108)? \piso.data_r [1323] : 
                      (N110)? \piso.data_r [1355] : 
                      (N112)? \piso.data_r [1387] : 
                      (N114)? \piso.data_r [1419] : 
                      (N116)? \piso.data_r [1451] : 
                      (N118)? \piso.data_r [1483] : 
                      (N120)? \piso.data_r [1515] : 
                      (N122)? \piso.data_r [1547] : 
                      (N124)? \piso.data_r [1579] : 
                      (N126)? \piso.data_r [1611] : 
                      (N128)? \piso.data_r [1643] : 
                      (N130)? \piso.data_r [1675] : 
                      (N132)? \piso.data_r [1707] : 
                      (N134)? \piso.data_r [1739] : 
                      (N136)? \piso.data_r [1771] : 
                      (N138)? \piso.data_r [1803] : 
                      (N140)? \piso.data_r [1835] : 
                      (N142)? \piso.data_r [1867] : 
                      (N144)? \piso.data_r [1899] : 
                      (N146)? \piso.data_r [1931] : 
                      (N148)? \piso.data_r [1963] : 
                      (N150)? \piso.data_r [1995] : 
                      (N152)? \piso.data_r [2027] : 1'b0;
  assign data_o[10] = (N89)? \piso.data_r [10] : 
                      (N91)? \piso.data_r [42] : 
                      (N93)? \piso.data_r [74] : 
                      (N95)? \piso.data_r [106] : 
                      (N97)? \piso.data_r [138] : 
                      (N99)? \piso.data_r [170] : 
                      (N101)? \piso.data_r [202] : 
                      (N103)? \piso.data_r [234] : 
                      (N105)? \piso.data_r [266] : 
                      (N107)? \piso.data_r [298] : 
                      (N109)? \piso.data_r [330] : 
                      (N111)? \piso.data_r [362] : 
                      (N113)? \piso.data_r [394] : 
                      (N115)? \piso.data_r [426] : 
                      (N117)? \piso.data_r [458] : 
                      (N119)? \piso.data_r [490] : 
                      (N121)? \piso.data_r [522] : 
                      (N123)? \piso.data_r [554] : 
                      (N125)? \piso.data_r [586] : 
                      (N127)? \piso.data_r [618] : 
                      (N129)? \piso.data_r [650] : 
                      (N131)? \piso.data_r [682] : 
                      (N133)? \piso.data_r [714] : 
                      (N135)? \piso.data_r [746] : 
                      (N137)? \piso.data_r [778] : 
                      (N139)? \piso.data_r [810] : 
                      (N141)? \piso.data_r [842] : 
                      (N143)? \piso.data_r [874] : 
                      (N145)? \piso.data_r [906] : 
                      (N147)? \piso.data_r [938] : 
                      (N149)? \piso.data_r [970] : 
                      (N151)? \piso.data_r [1002] : 
                      (N90)? \piso.data_r [1034] : 
                      (N92)? \piso.data_r [1066] : 
                      (N94)? \piso.data_r [1098] : 
                      (N96)? \piso.data_r [1130] : 
                      (N98)? \piso.data_r [1162] : 
                      (N100)? \piso.data_r [1194] : 
                      (N102)? \piso.data_r [1226] : 
                      (N104)? \piso.data_r [1258] : 
                      (N106)? \piso.data_r [1290] : 
                      (N108)? \piso.data_r [1322] : 
                      (N110)? \piso.data_r [1354] : 
                      (N112)? \piso.data_r [1386] : 
                      (N114)? \piso.data_r [1418] : 
                      (N116)? \piso.data_r [1450] : 
                      (N118)? \piso.data_r [1482] : 
                      (N120)? \piso.data_r [1514] : 
                      (N122)? \piso.data_r [1546] : 
                      (N124)? \piso.data_r [1578] : 
                      (N126)? \piso.data_r [1610] : 
                      (N128)? \piso.data_r [1642] : 
                      (N130)? \piso.data_r [1674] : 
                      (N132)? \piso.data_r [1706] : 
                      (N134)? \piso.data_r [1738] : 
                      (N136)? \piso.data_r [1770] : 
                      (N138)? \piso.data_r [1802] : 
                      (N140)? \piso.data_r [1834] : 
                      (N142)? \piso.data_r [1866] : 
                      (N144)? \piso.data_r [1898] : 
                      (N146)? \piso.data_r [1930] : 
                      (N148)? \piso.data_r [1962] : 
                      (N150)? \piso.data_r [1994] : 
                      (N152)? \piso.data_r [2026] : 1'b0;
  assign data_o[9] = (N89)? \piso.data_r [9] : 
                     (N91)? \piso.data_r [41] : 
                     (N93)? \piso.data_r [73] : 
                     (N95)? \piso.data_r [105] : 
                     (N97)? \piso.data_r [137] : 
                     (N99)? \piso.data_r [169] : 
                     (N101)? \piso.data_r [201] : 
                     (N103)? \piso.data_r [233] : 
                     (N105)? \piso.data_r [265] : 
                     (N107)? \piso.data_r [297] : 
                     (N109)? \piso.data_r [329] : 
                     (N111)? \piso.data_r [361] : 
                     (N113)? \piso.data_r [393] : 
                     (N115)? \piso.data_r [425] : 
                     (N117)? \piso.data_r [457] : 
                     (N119)? \piso.data_r [489] : 
                     (N121)? \piso.data_r [521] : 
                     (N123)? \piso.data_r [553] : 
                     (N125)? \piso.data_r [585] : 
                     (N127)? \piso.data_r [617] : 
                     (N129)? \piso.data_r [649] : 
                     (N131)? \piso.data_r [681] : 
                     (N133)? \piso.data_r [713] : 
                     (N135)? \piso.data_r [745] : 
                     (N137)? \piso.data_r [777] : 
                     (N139)? \piso.data_r [809] : 
                     (N141)? \piso.data_r [841] : 
                     (N143)? \piso.data_r [873] : 
                     (N145)? \piso.data_r [905] : 
                     (N147)? \piso.data_r [937] : 
                     (N149)? \piso.data_r [969] : 
                     (N151)? \piso.data_r [1001] : 
                     (N90)? \piso.data_r [1033] : 
                     (N92)? \piso.data_r [1065] : 
                     (N94)? \piso.data_r [1097] : 
                     (N96)? \piso.data_r [1129] : 
                     (N98)? \piso.data_r [1161] : 
                     (N100)? \piso.data_r [1193] : 
                     (N102)? \piso.data_r [1225] : 
                     (N104)? \piso.data_r [1257] : 
                     (N106)? \piso.data_r [1289] : 
                     (N108)? \piso.data_r [1321] : 
                     (N110)? \piso.data_r [1353] : 
                     (N112)? \piso.data_r [1385] : 
                     (N114)? \piso.data_r [1417] : 
                     (N116)? \piso.data_r [1449] : 
                     (N118)? \piso.data_r [1481] : 
                     (N120)? \piso.data_r [1513] : 
                     (N122)? \piso.data_r [1545] : 
                     (N124)? \piso.data_r [1577] : 
                     (N126)? \piso.data_r [1609] : 
                     (N128)? \piso.data_r [1641] : 
                     (N130)? \piso.data_r [1673] : 
                     (N132)? \piso.data_r [1705] : 
                     (N134)? \piso.data_r [1737] : 
                     (N136)? \piso.data_r [1769] : 
                     (N138)? \piso.data_r [1801] : 
                     (N140)? \piso.data_r [1833] : 
                     (N142)? \piso.data_r [1865] : 
                     (N144)? \piso.data_r [1897] : 
                     (N146)? \piso.data_r [1929] : 
                     (N148)? \piso.data_r [1961] : 
                     (N150)? \piso.data_r [1993] : 
                     (N152)? \piso.data_r [2025] : 1'b0;
  assign data_o[8] = (N89)? \piso.data_r [8] : 
                     (N91)? \piso.data_r [40] : 
                     (N93)? \piso.data_r [72] : 
                     (N95)? \piso.data_r [104] : 
                     (N97)? \piso.data_r [136] : 
                     (N99)? \piso.data_r [168] : 
                     (N101)? \piso.data_r [200] : 
                     (N103)? \piso.data_r [232] : 
                     (N105)? \piso.data_r [264] : 
                     (N107)? \piso.data_r [296] : 
                     (N109)? \piso.data_r [328] : 
                     (N111)? \piso.data_r [360] : 
                     (N113)? \piso.data_r [392] : 
                     (N115)? \piso.data_r [424] : 
                     (N117)? \piso.data_r [456] : 
                     (N119)? \piso.data_r [488] : 
                     (N121)? \piso.data_r [520] : 
                     (N123)? \piso.data_r [552] : 
                     (N125)? \piso.data_r [584] : 
                     (N127)? \piso.data_r [616] : 
                     (N129)? \piso.data_r [648] : 
                     (N131)? \piso.data_r [680] : 
                     (N133)? \piso.data_r [712] : 
                     (N135)? \piso.data_r [744] : 
                     (N137)? \piso.data_r [776] : 
                     (N139)? \piso.data_r [808] : 
                     (N141)? \piso.data_r [840] : 
                     (N143)? \piso.data_r [872] : 
                     (N145)? \piso.data_r [904] : 
                     (N147)? \piso.data_r [936] : 
                     (N149)? \piso.data_r [968] : 
                     (N151)? \piso.data_r [1000] : 
                     (N90)? \piso.data_r [1032] : 
                     (N92)? \piso.data_r [1064] : 
                     (N94)? \piso.data_r [1096] : 
                     (N96)? \piso.data_r [1128] : 
                     (N98)? \piso.data_r [1160] : 
                     (N100)? \piso.data_r [1192] : 
                     (N102)? \piso.data_r [1224] : 
                     (N104)? \piso.data_r [1256] : 
                     (N106)? \piso.data_r [1288] : 
                     (N108)? \piso.data_r [1320] : 
                     (N110)? \piso.data_r [1352] : 
                     (N112)? \piso.data_r [1384] : 
                     (N114)? \piso.data_r [1416] : 
                     (N116)? \piso.data_r [1448] : 
                     (N118)? \piso.data_r [1480] : 
                     (N120)? \piso.data_r [1512] : 
                     (N122)? \piso.data_r [1544] : 
                     (N124)? \piso.data_r [1576] : 
                     (N126)? \piso.data_r [1608] : 
                     (N128)? \piso.data_r [1640] : 
                     (N130)? \piso.data_r [1672] : 
                     (N132)? \piso.data_r [1704] : 
                     (N134)? \piso.data_r [1736] : 
                     (N136)? \piso.data_r [1768] : 
                     (N138)? \piso.data_r [1800] : 
                     (N140)? \piso.data_r [1832] : 
                     (N142)? \piso.data_r [1864] : 
                     (N144)? \piso.data_r [1896] : 
                     (N146)? \piso.data_r [1928] : 
                     (N148)? \piso.data_r [1960] : 
                     (N150)? \piso.data_r [1992] : 
                     (N152)? \piso.data_r [2024] : 1'b0;
  assign data_o[7] = (N89)? \piso.data_r [7] : 
                     (N91)? \piso.data_r [39] : 
                     (N93)? \piso.data_r [71] : 
                     (N95)? \piso.data_r [103] : 
                     (N97)? \piso.data_r [135] : 
                     (N99)? \piso.data_r [167] : 
                     (N101)? \piso.data_r [199] : 
                     (N103)? \piso.data_r [231] : 
                     (N105)? \piso.data_r [263] : 
                     (N107)? \piso.data_r [295] : 
                     (N109)? \piso.data_r [327] : 
                     (N111)? \piso.data_r [359] : 
                     (N113)? \piso.data_r [391] : 
                     (N115)? \piso.data_r [423] : 
                     (N117)? \piso.data_r [455] : 
                     (N119)? \piso.data_r [487] : 
                     (N121)? \piso.data_r [519] : 
                     (N123)? \piso.data_r [551] : 
                     (N125)? \piso.data_r [583] : 
                     (N127)? \piso.data_r [615] : 
                     (N129)? \piso.data_r [647] : 
                     (N131)? \piso.data_r [679] : 
                     (N133)? \piso.data_r [711] : 
                     (N135)? \piso.data_r [743] : 
                     (N137)? \piso.data_r [775] : 
                     (N139)? \piso.data_r [807] : 
                     (N141)? \piso.data_r [839] : 
                     (N143)? \piso.data_r [871] : 
                     (N145)? \piso.data_r [903] : 
                     (N147)? \piso.data_r [935] : 
                     (N149)? \piso.data_r [967] : 
                     (N151)? \piso.data_r [999] : 
                     (N90)? \piso.data_r [1031] : 
                     (N92)? \piso.data_r [1063] : 
                     (N94)? \piso.data_r [1095] : 
                     (N96)? \piso.data_r [1127] : 
                     (N98)? \piso.data_r [1159] : 
                     (N100)? \piso.data_r [1191] : 
                     (N102)? \piso.data_r [1223] : 
                     (N104)? \piso.data_r [1255] : 
                     (N106)? \piso.data_r [1287] : 
                     (N108)? \piso.data_r [1319] : 
                     (N110)? \piso.data_r [1351] : 
                     (N112)? \piso.data_r [1383] : 
                     (N114)? \piso.data_r [1415] : 
                     (N116)? \piso.data_r [1447] : 
                     (N118)? \piso.data_r [1479] : 
                     (N120)? \piso.data_r [1511] : 
                     (N122)? \piso.data_r [1543] : 
                     (N124)? \piso.data_r [1575] : 
                     (N126)? \piso.data_r [1607] : 
                     (N128)? \piso.data_r [1639] : 
                     (N130)? \piso.data_r [1671] : 
                     (N132)? \piso.data_r [1703] : 
                     (N134)? \piso.data_r [1735] : 
                     (N136)? \piso.data_r [1767] : 
                     (N138)? \piso.data_r [1799] : 
                     (N140)? \piso.data_r [1831] : 
                     (N142)? \piso.data_r [1863] : 
                     (N144)? \piso.data_r [1895] : 
                     (N146)? \piso.data_r [1927] : 
                     (N148)? \piso.data_r [1959] : 
                     (N150)? \piso.data_r [1991] : 
                     (N152)? \piso.data_r [2023] : 1'b0;
  assign data_o[6] = (N89)? \piso.data_r [6] : 
                     (N91)? \piso.data_r [38] : 
                     (N93)? \piso.data_r [70] : 
                     (N95)? \piso.data_r [102] : 
                     (N97)? \piso.data_r [134] : 
                     (N99)? \piso.data_r [166] : 
                     (N101)? \piso.data_r [198] : 
                     (N103)? \piso.data_r [230] : 
                     (N105)? \piso.data_r [262] : 
                     (N107)? \piso.data_r [294] : 
                     (N109)? \piso.data_r [326] : 
                     (N111)? \piso.data_r [358] : 
                     (N113)? \piso.data_r [390] : 
                     (N115)? \piso.data_r [422] : 
                     (N117)? \piso.data_r [454] : 
                     (N119)? \piso.data_r [486] : 
                     (N121)? \piso.data_r [518] : 
                     (N123)? \piso.data_r [550] : 
                     (N125)? \piso.data_r [582] : 
                     (N127)? \piso.data_r [614] : 
                     (N129)? \piso.data_r [646] : 
                     (N131)? \piso.data_r [678] : 
                     (N133)? \piso.data_r [710] : 
                     (N135)? \piso.data_r [742] : 
                     (N137)? \piso.data_r [774] : 
                     (N139)? \piso.data_r [806] : 
                     (N141)? \piso.data_r [838] : 
                     (N143)? \piso.data_r [870] : 
                     (N145)? \piso.data_r [902] : 
                     (N147)? \piso.data_r [934] : 
                     (N149)? \piso.data_r [966] : 
                     (N151)? \piso.data_r [998] : 
                     (N90)? \piso.data_r [1030] : 
                     (N92)? \piso.data_r [1062] : 
                     (N94)? \piso.data_r [1094] : 
                     (N96)? \piso.data_r [1126] : 
                     (N98)? \piso.data_r [1158] : 
                     (N100)? \piso.data_r [1190] : 
                     (N102)? \piso.data_r [1222] : 
                     (N104)? \piso.data_r [1254] : 
                     (N106)? \piso.data_r [1286] : 
                     (N108)? \piso.data_r [1318] : 
                     (N110)? \piso.data_r [1350] : 
                     (N112)? \piso.data_r [1382] : 
                     (N114)? \piso.data_r [1414] : 
                     (N116)? \piso.data_r [1446] : 
                     (N118)? \piso.data_r [1478] : 
                     (N120)? \piso.data_r [1510] : 
                     (N122)? \piso.data_r [1542] : 
                     (N124)? \piso.data_r [1574] : 
                     (N126)? \piso.data_r [1606] : 
                     (N128)? \piso.data_r [1638] : 
                     (N130)? \piso.data_r [1670] : 
                     (N132)? \piso.data_r [1702] : 
                     (N134)? \piso.data_r [1734] : 
                     (N136)? \piso.data_r [1766] : 
                     (N138)? \piso.data_r [1798] : 
                     (N140)? \piso.data_r [1830] : 
                     (N142)? \piso.data_r [1862] : 
                     (N144)? \piso.data_r [1894] : 
                     (N146)? \piso.data_r [1926] : 
                     (N148)? \piso.data_r [1958] : 
                     (N150)? \piso.data_r [1990] : 
                     (N152)? \piso.data_r [2022] : 1'b0;
  assign data_o[5] = (N89)? \piso.data_r [5] : 
                     (N91)? \piso.data_r [37] : 
                     (N93)? \piso.data_r [69] : 
                     (N95)? \piso.data_r [101] : 
                     (N97)? \piso.data_r [133] : 
                     (N99)? \piso.data_r [165] : 
                     (N101)? \piso.data_r [197] : 
                     (N103)? \piso.data_r [229] : 
                     (N105)? \piso.data_r [261] : 
                     (N107)? \piso.data_r [293] : 
                     (N109)? \piso.data_r [325] : 
                     (N111)? \piso.data_r [357] : 
                     (N113)? \piso.data_r [389] : 
                     (N115)? \piso.data_r [421] : 
                     (N117)? \piso.data_r [453] : 
                     (N119)? \piso.data_r [485] : 
                     (N121)? \piso.data_r [517] : 
                     (N123)? \piso.data_r [549] : 
                     (N125)? \piso.data_r [581] : 
                     (N127)? \piso.data_r [613] : 
                     (N129)? \piso.data_r [645] : 
                     (N131)? \piso.data_r [677] : 
                     (N133)? \piso.data_r [709] : 
                     (N135)? \piso.data_r [741] : 
                     (N137)? \piso.data_r [773] : 
                     (N139)? \piso.data_r [805] : 
                     (N141)? \piso.data_r [837] : 
                     (N143)? \piso.data_r [869] : 
                     (N145)? \piso.data_r [901] : 
                     (N147)? \piso.data_r [933] : 
                     (N149)? \piso.data_r [965] : 
                     (N151)? \piso.data_r [997] : 
                     (N90)? \piso.data_r [1029] : 
                     (N92)? \piso.data_r [1061] : 
                     (N94)? \piso.data_r [1093] : 
                     (N96)? \piso.data_r [1125] : 
                     (N98)? \piso.data_r [1157] : 
                     (N100)? \piso.data_r [1189] : 
                     (N102)? \piso.data_r [1221] : 
                     (N104)? \piso.data_r [1253] : 
                     (N106)? \piso.data_r [1285] : 
                     (N108)? \piso.data_r [1317] : 
                     (N110)? \piso.data_r [1349] : 
                     (N112)? \piso.data_r [1381] : 
                     (N114)? \piso.data_r [1413] : 
                     (N116)? \piso.data_r [1445] : 
                     (N118)? \piso.data_r [1477] : 
                     (N120)? \piso.data_r [1509] : 
                     (N122)? \piso.data_r [1541] : 
                     (N124)? \piso.data_r [1573] : 
                     (N126)? \piso.data_r [1605] : 
                     (N128)? \piso.data_r [1637] : 
                     (N130)? \piso.data_r [1669] : 
                     (N132)? \piso.data_r [1701] : 
                     (N134)? \piso.data_r [1733] : 
                     (N136)? \piso.data_r [1765] : 
                     (N138)? \piso.data_r [1797] : 
                     (N140)? \piso.data_r [1829] : 
                     (N142)? \piso.data_r [1861] : 
                     (N144)? \piso.data_r [1893] : 
                     (N146)? \piso.data_r [1925] : 
                     (N148)? \piso.data_r [1957] : 
                     (N150)? \piso.data_r [1989] : 
                     (N152)? \piso.data_r [2021] : 1'b0;
  assign data_o[4] = (N89)? \piso.data_r [4] : 
                     (N91)? \piso.data_r [36] : 
                     (N93)? \piso.data_r [68] : 
                     (N95)? \piso.data_r [100] : 
                     (N97)? \piso.data_r [132] : 
                     (N99)? \piso.data_r [164] : 
                     (N101)? \piso.data_r [196] : 
                     (N103)? \piso.data_r [228] : 
                     (N105)? \piso.data_r [260] : 
                     (N107)? \piso.data_r [292] : 
                     (N109)? \piso.data_r [324] : 
                     (N111)? \piso.data_r [356] : 
                     (N113)? \piso.data_r [388] : 
                     (N115)? \piso.data_r [420] : 
                     (N117)? \piso.data_r [452] : 
                     (N119)? \piso.data_r [484] : 
                     (N121)? \piso.data_r [516] : 
                     (N123)? \piso.data_r [548] : 
                     (N125)? \piso.data_r [580] : 
                     (N127)? \piso.data_r [612] : 
                     (N129)? \piso.data_r [644] : 
                     (N131)? \piso.data_r [676] : 
                     (N133)? \piso.data_r [708] : 
                     (N135)? \piso.data_r [740] : 
                     (N137)? \piso.data_r [772] : 
                     (N139)? \piso.data_r [804] : 
                     (N141)? \piso.data_r [836] : 
                     (N143)? \piso.data_r [868] : 
                     (N145)? \piso.data_r [900] : 
                     (N147)? \piso.data_r [932] : 
                     (N149)? \piso.data_r [964] : 
                     (N151)? \piso.data_r [996] : 
                     (N90)? \piso.data_r [1028] : 
                     (N92)? \piso.data_r [1060] : 
                     (N94)? \piso.data_r [1092] : 
                     (N96)? \piso.data_r [1124] : 
                     (N98)? \piso.data_r [1156] : 
                     (N100)? \piso.data_r [1188] : 
                     (N102)? \piso.data_r [1220] : 
                     (N104)? \piso.data_r [1252] : 
                     (N106)? \piso.data_r [1284] : 
                     (N108)? \piso.data_r [1316] : 
                     (N110)? \piso.data_r [1348] : 
                     (N112)? \piso.data_r [1380] : 
                     (N114)? \piso.data_r [1412] : 
                     (N116)? \piso.data_r [1444] : 
                     (N118)? \piso.data_r [1476] : 
                     (N120)? \piso.data_r [1508] : 
                     (N122)? \piso.data_r [1540] : 
                     (N124)? \piso.data_r [1572] : 
                     (N126)? \piso.data_r [1604] : 
                     (N128)? \piso.data_r [1636] : 
                     (N130)? \piso.data_r [1668] : 
                     (N132)? \piso.data_r [1700] : 
                     (N134)? \piso.data_r [1732] : 
                     (N136)? \piso.data_r [1764] : 
                     (N138)? \piso.data_r [1796] : 
                     (N140)? \piso.data_r [1828] : 
                     (N142)? \piso.data_r [1860] : 
                     (N144)? \piso.data_r [1892] : 
                     (N146)? \piso.data_r [1924] : 
                     (N148)? \piso.data_r [1956] : 
                     (N150)? \piso.data_r [1988] : 
                     (N152)? \piso.data_r [2020] : 1'b0;
  assign data_o[3] = (N89)? \piso.data_r [3] : 
                     (N91)? \piso.data_r [35] : 
                     (N93)? \piso.data_r [67] : 
                     (N95)? \piso.data_r [99] : 
                     (N97)? \piso.data_r [131] : 
                     (N99)? \piso.data_r [163] : 
                     (N101)? \piso.data_r [195] : 
                     (N103)? \piso.data_r [227] : 
                     (N105)? \piso.data_r [259] : 
                     (N107)? \piso.data_r [291] : 
                     (N109)? \piso.data_r [323] : 
                     (N111)? \piso.data_r [355] : 
                     (N113)? \piso.data_r [387] : 
                     (N115)? \piso.data_r [419] : 
                     (N117)? \piso.data_r [451] : 
                     (N119)? \piso.data_r [483] : 
                     (N121)? \piso.data_r [515] : 
                     (N123)? \piso.data_r [547] : 
                     (N125)? \piso.data_r [579] : 
                     (N127)? \piso.data_r [611] : 
                     (N129)? \piso.data_r [643] : 
                     (N131)? \piso.data_r [675] : 
                     (N133)? \piso.data_r [707] : 
                     (N135)? \piso.data_r [739] : 
                     (N137)? \piso.data_r [771] : 
                     (N139)? \piso.data_r [803] : 
                     (N141)? \piso.data_r [835] : 
                     (N143)? \piso.data_r [867] : 
                     (N145)? \piso.data_r [899] : 
                     (N147)? \piso.data_r [931] : 
                     (N149)? \piso.data_r [963] : 
                     (N151)? \piso.data_r [995] : 
                     (N90)? \piso.data_r [1027] : 
                     (N92)? \piso.data_r [1059] : 
                     (N94)? \piso.data_r [1091] : 
                     (N96)? \piso.data_r [1123] : 
                     (N98)? \piso.data_r [1155] : 
                     (N100)? \piso.data_r [1187] : 
                     (N102)? \piso.data_r [1219] : 
                     (N104)? \piso.data_r [1251] : 
                     (N106)? \piso.data_r [1283] : 
                     (N108)? \piso.data_r [1315] : 
                     (N110)? \piso.data_r [1347] : 
                     (N112)? \piso.data_r [1379] : 
                     (N114)? \piso.data_r [1411] : 
                     (N116)? \piso.data_r [1443] : 
                     (N118)? \piso.data_r [1475] : 
                     (N120)? \piso.data_r [1507] : 
                     (N122)? \piso.data_r [1539] : 
                     (N124)? \piso.data_r [1571] : 
                     (N126)? \piso.data_r [1603] : 
                     (N128)? \piso.data_r [1635] : 
                     (N130)? \piso.data_r [1667] : 
                     (N132)? \piso.data_r [1699] : 
                     (N134)? \piso.data_r [1731] : 
                     (N136)? \piso.data_r [1763] : 
                     (N138)? \piso.data_r [1795] : 
                     (N140)? \piso.data_r [1827] : 
                     (N142)? \piso.data_r [1859] : 
                     (N144)? \piso.data_r [1891] : 
                     (N146)? \piso.data_r [1923] : 
                     (N148)? \piso.data_r [1955] : 
                     (N150)? \piso.data_r [1987] : 
                     (N152)? \piso.data_r [2019] : 1'b0;
  assign data_o[2] = (N89)? \piso.data_r [2] : 
                     (N91)? \piso.data_r [34] : 
                     (N93)? \piso.data_r [66] : 
                     (N95)? \piso.data_r [98] : 
                     (N97)? \piso.data_r [130] : 
                     (N99)? \piso.data_r [162] : 
                     (N101)? \piso.data_r [194] : 
                     (N103)? \piso.data_r [226] : 
                     (N105)? \piso.data_r [258] : 
                     (N107)? \piso.data_r [290] : 
                     (N109)? \piso.data_r [322] : 
                     (N111)? \piso.data_r [354] : 
                     (N113)? \piso.data_r [386] : 
                     (N115)? \piso.data_r [418] : 
                     (N117)? \piso.data_r [450] : 
                     (N119)? \piso.data_r [482] : 
                     (N121)? \piso.data_r [514] : 
                     (N123)? \piso.data_r [546] : 
                     (N125)? \piso.data_r [578] : 
                     (N127)? \piso.data_r [610] : 
                     (N129)? \piso.data_r [642] : 
                     (N131)? \piso.data_r [674] : 
                     (N133)? \piso.data_r [706] : 
                     (N135)? \piso.data_r [738] : 
                     (N137)? \piso.data_r [770] : 
                     (N139)? \piso.data_r [802] : 
                     (N141)? \piso.data_r [834] : 
                     (N143)? \piso.data_r [866] : 
                     (N145)? \piso.data_r [898] : 
                     (N147)? \piso.data_r [930] : 
                     (N149)? \piso.data_r [962] : 
                     (N151)? \piso.data_r [994] : 
                     (N90)? \piso.data_r [1026] : 
                     (N92)? \piso.data_r [1058] : 
                     (N94)? \piso.data_r [1090] : 
                     (N96)? \piso.data_r [1122] : 
                     (N98)? \piso.data_r [1154] : 
                     (N100)? \piso.data_r [1186] : 
                     (N102)? \piso.data_r [1218] : 
                     (N104)? \piso.data_r [1250] : 
                     (N106)? \piso.data_r [1282] : 
                     (N108)? \piso.data_r [1314] : 
                     (N110)? \piso.data_r [1346] : 
                     (N112)? \piso.data_r [1378] : 
                     (N114)? \piso.data_r [1410] : 
                     (N116)? \piso.data_r [1442] : 
                     (N118)? \piso.data_r [1474] : 
                     (N120)? \piso.data_r [1506] : 
                     (N122)? \piso.data_r [1538] : 
                     (N124)? \piso.data_r [1570] : 
                     (N126)? \piso.data_r [1602] : 
                     (N128)? \piso.data_r [1634] : 
                     (N130)? \piso.data_r [1666] : 
                     (N132)? \piso.data_r [1698] : 
                     (N134)? \piso.data_r [1730] : 
                     (N136)? \piso.data_r [1762] : 
                     (N138)? \piso.data_r [1794] : 
                     (N140)? \piso.data_r [1826] : 
                     (N142)? \piso.data_r [1858] : 
                     (N144)? \piso.data_r [1890] : 
                     (N146)? \piso.data_r [1922] : 
                     (N148)? \piso.data_r [1954] : 
                     (N150)? \piso.data_r [1986] : 
                     (N152)? \piso.data_r [2018] : 1'b0;
  assign data_o[1] = (N89)? \piso.data_r [1] : 
                     (N91)? \piso.data_r [33] : 
                     (N93)? \piso.data_r [65] : 
                     (N95)? \piso.data_r [97] : 
                     (N97)? \piso.data_r [129] : 
                     (N99)? \piso.data_r [161] : 
                     (N101)? \piso.data_r [193] : 
                     (N103)? \piso.data_r [225] : 
                     (N105)? \piso.data_r [257] : 
                     (N107)? \piso.data_r [289] : 
                     (N109)? \piso.data_r [321] : 
                     (N111)? \piso.data_r [353] : 
                     (N113)? \piso.data_r [385] : 
                     (N115)? \piso.data_r [417] : 
                     (N117)? \piso.data_r [449] : 
                     (N119)? \piso.data_r [481] : 
                     (N121)? \piso.data_r [513] : 
                     (N123)? \piso.data_r [545] : 
                     (N125)? \piso.data_r [577] : 
                     (N127)? \piso.data_r [609] : 
                     (N129)? \piso.data_r [641] : 
                     (N131)? \piso.data_r [673] : 
                     (N133)? \piso.data_r [705] : 
                     (N135)? \piso.data_r [737] : 
                     (N137)? \piso.data_r [769] : 
                     (N139)? \piso.data_r [801] : 
                     (N141)? \piso.data_r [833] : 
                     (N143)? \piso.data_r [865] : 
                     (N145)? \piso.data_r [897] : 
                     (N147)? \piso.data_r [929] : 
                     (N149)? \piso.data_r [961] : 
                     (N151)? \piso.data_r [993] : 
                     (N90)? \piso.data_r [1025] : 
                     (N92)? \piso.data_r [1057] : 
                     (N94)? \piso.data_r [1089] : 
                     (N96)? \piso.data_r [1121] : 
                     (N98)? \piso.data_r [1153] : 
                     (N100)? \piso.data_r [1185] : 
                     (N102)? \piso.data_r [1217] : 
                     (N104)? \piso.data_r [1249] : 
                     (N106)? \piso.data_r [1281] : 
                     (N108)? \piso.data_r [1313] : 
                     (N110)? \piso.data_r [1345] : 
                     (N112)? \piso.data_r [1377] : 
                     (N114)? \piso.data_r [1409] : 
                     (N116)? \piso.data_r [1441] : 
                     (N118)? \piso.data_r [1473] : 
                     (N120)? \piso.data_r [1505] : 
                     (N122)? \piso.data_r [1537] : 
                     (N124)? \piso.data_r [1569] : 
                     (N126)? \piso.data_r [1601] : 
                     (N128)? \piso.data_r [1633] : 
                     (N130)? \piso.data_r [1665] : 
                     (N132)? \piso.data_r [1697] : 
                     (N134)? \piso.data_r [1729] : 
                     (N136)? \piso.data_r [1761] : 
                     (N138)? \piso.data_r [1793] : 
                     (N140)? \piso.data_r [1825] : 
                     (N142)? \piso.data_r [1857] : 
                     (N144)? \piso.data_r [1889] : 
                     (N146)? \piso.data_r [1921] : 
                     (N148)? \piso.data_r [1953] : 
                     (N150)? \piso.data_r [1985] : 
                     (N152)? \piso.data_r [2017] : 1'b0;
  assign data_o[0] = (N89)? \piso.data_r [0] : 
                     (N91)? \piso.data_r [32] : 
                     (N93)? \piso.data_r [64] : 
                     (N95)? \piso.data_r [96] : 
                     (N97)? \piso.data_r [128] : 
                     (N99)? \piso.data_r [160] : 
                     (N101)? \piso.data_r [192] : 
                     (N103)? \piso.data_r [224] : 
                     (N105)? \piso.data_r [256] : 
                     (N107)? \piso.data_r [288] : 
                     (N109)? \piso.data_r [320] : 
                     (N111)? \piso.data_r [352] : 
                     (N113)? \piso.data_r [384] : 
                     (N115)? \piso.data_r [416] : 
                     (N117)? \piso.data_r [448] : 
                     (N119)? \piso.data_r [480] : 
                     (N121)? \piso.data_r [512] : 
                     (N123)? \piso.data_r [544] : 
                     (N125)? \piso.data_r [576] : 
                     (N127)? \piso.data_r [608] : 
                     (N129)? \piso.data_r [640] : 
                     (N131)? \piso.data_r [672] : 
                     (N133)? \piso.data_r [704] : 
                     (N135)? \piso.data_r [736] : 
                     (N137)? \piso.data_r [768] : 
                     (N139)? \piso.data_r [800] : 
                     (N141)? \piso.data_r [832] : 
                     (N143)? \piso.data_r [864] : 
                     (N145)? \piso.data_r [896] : 
                     (N147)? \piso.data_r [928] : 
                     (N149)? \piso.data_r [960] : 
                     (N151)? \piso.data_r [992] : 
                     (N90)? \piso.data_r [1024] : 
                     (N92)? \piso.data_r [1056] : 
                     (N94)? \piso.data_r [1088] : 
                     (N96)? \piso.data_r [1120] : 
                     (N98)? \piso.data_r [1152] : 
                     (N100)? \piso.data_r [1184] : 
                     (N102)? \piso.data_r [1216] : 
                     (N104)? \piso.data_r [1248] : 
                     (N106)? \piso.data_r [1280] : 
                     (N108)? \piso.data_r [1312] : 
                     (N110)? \piso.data_r [1344] : 
                     (N112)? \piso.data_r [1376] : 
                     (N114)? \piso.data_r [1408] : 
                     (N116)? \piso.data_r [1440] : 
                     (N118)? \piso.data_r [1472] : 
                     (N120)? \piso.data_r [1504] : 
                     (N122)? \piso.data_r [1536] : 
                     (N124)? \piso.data_r [1568] : 
                     (N126)? \piso.data_r [1600] : 
                     (N128)? \piso.data_r [1632] : 
                     (N130)? \piso.data_r [1664] : 
                     (N132)? \piso.data_r [1696] : 
                     (N134)? \piso.data_r [1728] : 
                     (N136)? \piso.data_r [1760] : 
                     (N138)? \piso.data_r [1792] : 
                     (N140)? \piso.data_r [1824] : 
                     (N142)? \piso.data_r [1856] : 
                     (N144)? \piso.data_r [1888] : 
                     (N146)? \piso.data_r [1920] : 
                     (N148)? \piso.data_r [1952] : 
                     (N150)? \piso.data_r [1984] : 
                     (N152)? \piso.data_r [2016] : 1'b0;
  assign N155 = ~valid_o;
  assign N156 = \piso.shift_ctr_r [4] & \piso.shift_ctr_r [5];
  assign N157 = \piso.shift_ctr_r [3] & N156;
  assign N158 = \piso.shift_ctr_r [2] & N157;
  assign N159 = \piso.shift_ctr_r [1] & N158;
  assign N160 = \piso.shift_ctr_r [0] & N159;
  assign { N22, N21, N20, N19, N18, N17 } = \piso.shift_ctr_r  + 1'b1;
  assign \piso.state_n [0] = (N0)? 1'b1 : 
                             (N5)? 1'b0 : 1'b0;
  assign N0 = N2;
  assign { N14, N13, N12, N11, N10, N9 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                           (N8)? { N22, N21, N20, N19, N18, N17 } : 1'b0;
  assign N1 = N7;
  assign \piso.done_tx_n  = N161 & yumi_i;
  assign N161 = valid_o & N160;
  assign ready_o = N155 | \piso.done_tx_n ;
  assign N2 = ready_o & valid_i;
  assign N3 = \piso.done_tx_n  | N2;
  assign N4 = ~N2;
  assign N5 = \piso.done_tx_n  & N4;
  assign N6 = ready_o & valid_i;
  assign N7 = ready_o & valid_i;
  assign N8 = ~N7;
  assign N15 = N162 & N163;
  assign N162 = valid_o & yumi_i;
  assign N163 = ~\piso.done_tx_n ;
  assign N16 = ~N15;
  assign N23 = ~\piso.shift_ctr_r [0];
  assign N24 = ~\piso.shift_ctr_r [1];
  assign N25 = N23 & N24;
  assign N26 = N23 & \piso.shift_ctr_r [1];
  assign N27 = \piso.shift_ctr_r [0] & N24;
  assign N28 = \piso.shift_ctr_r [0] & \piso.shift_ctr_r [1];
  assign N29 = ~\piso.shift_ctr_r [2];
  assign N30 = N25 & N29;
  assign N31 = N25 & \piso.shift_ctr_r [2];
  assign N32 = N27 & N29;
  assign N33 = N27 & \piso.shift_ctr_r [2];
  assign N34 = N26 & N29;
  assign N35 = N26 & \piso.shift_ctr_r [2];
  assign N36 = N28 & N29;
  assign N37 = N28 & \piso.shift_ctr_r [2];
  assign N38 = ~\piso.shift_ctr_r [3];
  assign N39 = N30 & N38;
  assign N40 = N30 & \piso.shift_ctr_r [3];
  assign N41 = N32 & N38;
  assign N42 = N32 & \piso.shift_ctr_r [3];
  assign N43 = N34 & N38;
  assign N44 = N34 & \piso.shift_ctr_r [3];
  assign N45 = N36 & N38;
  assign N46 = N36 & \piso.shift_ctr_r [3];
  assign N47 = N31 & N38;
  assign N48 = N31 & \piso.shift_ctr_r [3];
  assign N49 = N33 & N38;
  assign N50 = N33 & \piso.shift_ctr_r [3];
  assign N51 = N35 & N38;
  assign N52 = N35 & \piso.shift_ctr_r [3];
  assign N53 = N37 & N38;
  assign N54 = N37 & \piso.shift_ctr_r [3];
  assign N55 = ~\piso.shift_ctr_r [4];
  assign N56 = N39 & N55;
  assign N57 = N39 & \piso.shift_ctr_r [4];
  assign N58 = N41 & N55;
  assign N59 = N41 & \piso.shift_ctr_r [4];
  assign N60 = N43 & N55;
  assign N61 = N43 & \piso.shift_ctr_r [4];
  assign N62 = N45 & N55;
  assign N63 = N45 & \piso.shift_ctr_r [4];
  assign N64 = N47 & N55;
  assign N65 = N47 & \piso.shift_ctr_r [4];
  assign N66 = N49 & N55;
  assign N67 = N49 & \piso.shift_ctr_r [4];
  assign N68 = N51 & N55;
  assign N69 = N51 & \piso.shift_ctr_r [4];
  assign N70 = N53 & N55;
  assign N71 = N53 & \piso.shift_ctr_r [4];
  assign N72 = N40 & N55;
  assign N73 = N40 & \piso.shift_ctr_r [4];
  assign N74 = N42 & N55;
  assign N75 = N42 & \piso.shift_ctr_r [4];
  assign N76 = N44 & N55;
  assign N77 = N44 & \piso.shift_ctr_r [4];
  assign N78 = N46 & N55;
  assign N79 = N46 & \piso.shift_ctr_r [4];
  assign N80 = N48 & N55;
  assign N81 = N48 & \piso.shift_ctr_r [4];
  assign N82 = N50 & N55;
  assign N83 = N50 & \piso.shift_ctr_r [4];
  assign N84 = N52 & N55;
  assign N85 = N52 & \piso.shift_ctr_r [4];
  assign N86 = N54 & N55;
  assign N87 = N54 & \piso.shift_ctr_r [4];
  assign N88 = ~\piso.shift_ctr_r [5];
  assign N89 = N56 & N88;
  assign N90 = N56 & \piso.shift_ctr_r [5];
  assign N91 = N58 & N88;
  assign N92 = N58 & \piso.shift_ctr_r [5];
  assign N93 = N60 & N88;
  assign N94 = N60 & \piso.shift_ctr_r [5];
  assign N95 = N62 & N88;
  assign N96 = N62 & \piso.shift_ctr_r [5];
  assign N97 = N64 & N88;
  assign N98 = N64 & \piso.shift_ctr_r [5];
  assign N99 = N66 & N88;
  assign N100 = N66 & \piso.shift_ctr_r [5];
  assign N101 = N68 & N88;
  assign N102 = N68 & \piso.shift_ctr_r [5];
  assign N103 = N70 & N88;
  assign N104 = N70 & \piso.shift_ctr_r [5];
  assign N105 = N72 & N88;
  assign N106 = N72 & \piso.shift_ctr_r [5];
  assign N107 = N74 & N88;
  assign N108 = N74 & \piso.shift_ctr_r [5];
  assign N109 = N76 & N88;
  assign N110 = N76 & \piso.shift_ctr_r [5];
  assign N111 = N78 & N88;
  assign N112 = N78 & \piso.shift_ctr_r [5];
  assign N113 = N80 & N88;
  assign N114 = N80 & \piso.shift_ctr_r [5];
  assign N115 = N82 & N88;
  assign N116 = N82 & \piso.shift_ctr_r [5];
  assign N117 = N84 & N88;
  assign N118 = N84 & \piso.shift_ctr_r [5];
  assign N119 = N86 & N88;
  assign N120 = N86 & \piso.shift_ctr_r [5];
  assign N121 = N57 & N88;
  assign N122 = N57 & \piso.shift_ctr_r [5];
  assign N123 = N59 & N88;
  assign N124 = N59 & \piso.shift_ctr_r [5];
  assign N125 = N61 & N88;
  assign N126 = N61 & \piso.shift_ctr_r [5];
  assign N127 = N63 & N88;
  assign N128 = N63 & \piso.shift_ctr_r [5];
  assign N129 = N65 & N88;
  assign N130 = N65 & \piso.shift_ctr_r [5];
  assign N131 = N67 & N88;
  assign N132 = N67 & \piso.shift_ctr_r [5];
  assign N133 = N69 & N88;
  assign N134 = N69 & \piso.shift_ctr_r [5];
  assign N135 = N71 & N88;
  assign N136 = N71 & \piso.shift_ctr_r [5];
  assign N137 = N73 & N88;
  assign N138 = N73 & \piso.shift_ctr_r [5];
  assign N139 = N75 & N88;
  assign N140 = N75 & \piso.shift_ctr_r [5];
  assign N141 = N77 & N88;
  assign N142 = N77 & \piso.shift_ctr_r [5];
  assign N143 = N79 & N88;
  assign N144 = N79 & \piso.shift_ctr_r [5];
  assign N145 = N81 & N88;
  assign N146 = N81 & \piso.shift_ctr_r [5];
  assign N147 = N83 & N88;
  assign N148 = N83 & \piso.shift_ctr_r [5];
  assign N149 = N85 & N88;
  assign N150 = N85 & \piso.shift_ctr_r [5];
  assign N151 = N87 & N88;
  assign N152 = N87 & \piso.shift_ctr_r [5];
  assign N153 = N16 & N8;
  assign N154 = ~N153;

  always @(posedge clk_i) begin
    if(reset_i) begin
      valid_o_sv2v_reg <= 1'b0;
    end else if(N3) begin
      valid_o_sv2v_reg <= \piso.state_n [0];
    end 
    if(reset_i) begin
      \piso.data_r_2047_sv2v_reg  <= 1'b0;
      \piso.data_r_2046_sv2v_reg  <= 1'b0;
      \piso.data_r_2045_sv2v_reg  <= 1'b0;
      \piso.data_r_2044_sv2v_reg  <= 1'b0;
      \piso.data_r_2043_sv2v_reg  <= 1'b0;
      \piso.data_r_2042_sv2v_reg  <= 1'b0;
      \piso.data_r_2041_sv2v_reg  <= 1'b0;
      \piso.data_r_2040_sv2v_reg  <= 1'b0;
      \piso.data_r_2039_sv2v_reg  <= 1'b0;
      \piso.data_r_2038_sv2v_reg  <= 1'b0;
      \piso.data_r_2037_sv2v_reg  <= 1'b0;
      \piso.data_r_2036_sv2v_reg  <= 1'b0;
      \piso.data_r_2035_sv2v_reg  <= 1'b0;
      \piso.data_r_2034_sv2v_reg  <= 1'b0;
      \piso.data_r_2033_sv2v_reg  <= 1'b0;
      \piso.data_r_2032_sv2v_reg  <= 1'b0;
      \piso.data_r_2031_sv2v_reg  <= 1'b0;
      \piso.data_r_2030_sv2v_reg  <= 1'b0;
      \piso.data_r_2029_sv2v_reg  <= 1'b0;
      \piso.data_r_2028_sv2v_reg  <= 1'b0;
      \piso.data_r_2027_sv2v_reg  <= 1'b0;
      \piso.data_r_2026_sv2v_reg  <= 1'b0;
      \piso.data_r_2025_sv2v_reg  <= 1'b0;
      \piso.data_r_2024_sv2v_reg  <= 1'b0;
      \piso.data_r_2023_sv2v_reg  <= 1'b0;
      \piso.data_r_2022_sv2v_reg  <= 1'b0;
      \piso.data_r_2021_sv2v_reg  <= 1'b0;
      \piso.data_r_2020_sv2v_reg  <= 1'b0;
      \piso.data_r_2019_sv2v_reg  <= 1'b0;
      \piso.data_r_2018_sv2v_reg  <= 1'b0;
      \piso.data_r_2017_sv2v_reg  <= 1'b0;
      \piso.data_r_2016_sv2v_reg  <= 1'b0;
      \piso.data_r_2015_sv2v_reg  <= 1'b0;
      \piso.data_r_2014_sv2v_reg  <= 1'b0;
      \piso.data_r_2013_sv2v_reg  <= 1'b0;
      \piso.data_r_2012_sv2v_reg  <= 1'b0;
      \piso.data_r_2011_sv2v_reg  <= 1'b0;
      \piso.data_r_2010_sv2v_reg  <= 1'b0;
      \piso.data_r_2009_sv2v_reg  <= 1'b0;
      \piso.data_r_2008_sv2v_reg  <= 1'b0;
      \piso.data_r_2007_sv2v_reg  <= 1'b0;
      \piso.data_r_2006_sv2v_reg  <= 1'b0;
      \piso.data_r_2005_sv2v_reg  <= 1'b0;
      \piso.data_r_2004_sv2v_reg  <= 1'b0;
      \piso.data_r_2003_sv2v_reg  <= 1'b0;
      \piso.data_r_2002_sv2v_reg  <= 1'b0;
      \piso.data_r_2001_sv2v_reg  <= 1'b0;
      \piso.data_r_2000_sv2v_reg  <= 1'b0;
      \piso.data_r_1999_sv2v_reg  <= 1'b0;
      \piso.data_r_1998_sv2v_reg  <= 1'b0;
      \piso.data_r_1997_sv2v_reg  <= 1'b0;
      \piso.data_r_1996_sv2v_reg  <= 1'b0;
      \piso.data_r_1995_sv2v_reg  <= 1'b0;
      \piso.data_r_1994_sv2v_reg  <= 1'b0;
      \piso.data_r_1993_sv2v_reg  <= 1'b0;
      \piso.data_r_1992_sv2v_reg  <= 1'b0;
      \piso.data_r_1991_sv2v_reg  <= 1'b0;
      \piso.data_r_1990_sv2v_reg  <= 1'b0;
      \piso.data_r_1989_sv2v_reg  <= 1'b0;
      \piso.data_r_1988_sv2v_reg  <= 1'b0;
      \piso.data_r_1987_sv2v_reg  <= 1'b0;
      \piso.data_r_1986_sv2v_reg  <= 1'b0;
      \piso.data_r_1985_sv2v_reg  <= 1'b0;
      \piso.data_r_1984_sv2v_reg  <= 1'b0;
      \piso.data_r_1983_sv2v_reg  <= 1'b0;
      \piso.data_r_1982_sv2v_reg  <= 1'b0;
      \piso.data_r_1981_sv2v_reg  <= 1'b0;
      \piso.data_r_1980_sv2v_reg  <= 1'b0;
      \piso.data_r_1979_sv2v_reg  <= 1'b0;
      \piso.data_r_1978_sv2v_reg  <= 1'b0;
      \piso.data_r_1977_sv2v_reg  <= 1'b0;
      \piso.data_r_1976_sv2v_reg  <= 1'b0;
      \piso.data_r_1975_sv2v_reg  <= 1'b0;
      \piso.data_r_1974_sv2v_reg  <= 1'b0;
      \piso.data_r_1973_sv2v_reg  <= 1'b0;
      \piso.data_r_1972_sv2v_reg  <= 1'b0;
      \piso.data_r_1971_sv2v_reg  <= 1'b0;
      \piso.data_r_1970_sv2v_reg  <= 1'b0;
      \piso.data_r_1969_sv2v_reg  <= 1'b0;
      \piso.data_r_1968_sv2v_reg  <= 1'b0;
      \piso.data_r_1967_sv2v_reg  <= 1'b0;
      \piso.data_r_1966_sv2v_reg  <= 1'b0;
      \piso.data_r_1965_sv2v_reg  <= 1'b0;
      \piso.data_r_1964_sv2v_reg  <= 1'b0;
      \piso.data_r_1963_sv2v_reg  <= 1'b0;
      \piso.data_r_1962_sv2v_reg  <= 1'b0;
      \piso.data_r_1961_sv2v_reg  <= 1'b0;
      \piso.data_r_1960_sv2v_reg  <= 1'b0;
      \piso.data_r_1959_sv2v_reg  <= 1'b0;
      \piso.data_r_1958_sv2v_reg  <= 1'b0;
      \piso.data_r_1957_sv2v_reg  <= 1'b0;
      \piso.data_r_1956_sv2v_reg  <= 1'b0;
      \piso.data_r_1955_sv2v_reg  <= 1'b0;
      \piso.data_r_1954_sv2v_reg  <= 1'b0;
      \piso.data_r_1953_sv2v_reg  <= 1'b0;
      \piso.data_r_1952_sv2v_reg  <= 1'b0;
      \piso.data_r_1951_sv2v_reg  <= 1'b0;
      \piso.data_r_1950_sv2v_reg  <= 1'b0;
      \piso.data_r_1949_sv2v_reg  <= 1'b0;
      \piso.data_r_1948_sv2v_reg  <= 1'b0;
      \piso.data_r_1947_sv2v_reg  <= 1'b0;
      \piso.data_r_1946_sv2v_reg  <= 1'b0;
      \piso.data_r_1945_sv2v_reg  <= 1'b0;
      \piso.data_r_1944_sv2v_reg  <= 1'b0;
      \piso.data_r_1943_sv2v_reg  <= 1'b0;
      \piso.data_r_1942_sv2v_reg  <= 1'b0;
      \piso.data_r_1941_sv2v_reg  <= 1'b0;
      \piso.data_r_1940_sv2v_reg  <= 1'b0;
      \piso.data_r_1939_sv2v_reg  <= 1'b0;
      \piso.data_r_1938_sv2v_reg  <= 1'b0;
      \piso.data_r_1937_sv2v_reg  <= 1'b0;
      \piso.data_r_1936_sv2v_reg  <= 1'b0;
      \piso.data_r_1935_sv2v_reg  <= 1'b0;
      \piso.data_r_1934_sv2v_reg  <= 1'b0;
      \piso.data_r_1933_sv2v_reg  <= 1'b0;
      \piso.data_r_1932_sv2v_reg  <= 1'b0;
      \piso.data_r_1931_sv2v_reg  <= 1'b0;
      \piso.data_r_1930_sv2v_reg  <= 1'b0;
      \piso.data_r_1929_sv2v_reg  <= 1'b0;
      \piso.data_r_1928_sv2v_reg  <= 1'b0;
      \piso.data_r_1927_sv2v_reg  <= 1'b0;
      \piso.data_r_1926_sv2v_reg  <= 1'b0;
      \piso.data_r_1925_sv2v_reg  <= 1'b0;
      \piso.data_r_1924_sv2v_reg  <= 1'b0;
      \piso.data_r_1923_sv2v_reg  <= 1'b0;
      \piso.data_r_1922_sv2v_reg  <= 1'b0;
      \piso.data_r_1921_sv2v_reg  <= 1'b0;
      \piso.data_r_1920_sv2v_reg  <= 1'b0;
      \piso.data_r_1919_sv2v_reg  <= 1'b0;
      \piso.data_r_1918_sv2v_reg  <= 1'b0;
      \piso.data_r_1917_sv2v_reg  <= 1'b0;
      \piso.data_r_1916_sv2v_reg  <= 1'b0;
      \piso.data_r_1915_sv2v_reg  <= 1'b0;
      \piso.data_r_1914_sv2v_reg  <= 1'b0;
      \piso.data_r_1913_sv2v_reg  <= 1'b0;
      \piso.data_r_1912_sv2v_reg  <= 1'b0;
      \piso.data_r_1911_sv2v_reg  <= 1'b0;
      \piso.data_r_1910_sv2v_reg  <= 1'b0;
      \piso.data_r_1909_sv2v_reg  <= 1'b0;
      \piso.data_r_1908_sv2v_reg  <= 1'b0;
      \piso.data_r_1907_sv2v_reg  <= 1'b0;
      \piso.data_r_1906_sv2v_reg  <= 1'b0;
      \piso.data_r_1905_sv2v_reg  <= 1'b0;
      \piso.data_r_1904_sv2v_reg  <= 1'b0;
      \piso.data_r_1903_sv2v_reg  <= 1'b0;
      \piso.data_r_1902_sv2v_reg  <= 1'b0;
      \piso.data_r_1901_sv2v_reg  <= 1'b0;
      \piso.data_r_1900_sv2v_reg  <= 1'b0;
      \piso.data_r_1899_sv2v_reg  <= 1'b0;
      \piso.data_r_1898_sv2v_reg  <= 1'b0;
      \piso.data_r_1897_sv2v_reg  <= 1'b0;
      \piso.data_r_1896_sv2v_reg  <= 1'b0;
      \piso.data_r_1895_sv2v_reg  <= 1'b0;
      \piso.data_r_1894_sv2v_reg  <= 1'b0;
      \piso.data_r_1893_sv2v_reg  <= 1'b0;
      \piso.data_r_1892_sv2v_reg  <= 1'b0;
      \piso.data_r_1891_sv2v_reg  <= 1'b0;
      \piso.data_r_1890_sv2v_reg  <= 1'b0;
      \piso.data_r_1889_sv2v_reg  <= 1'b0;
      \piso.data_r_1888_sv2v_reg  <= 1'b0;
      \piso.data_r_1887_sv2v_reg  <= 1'b0;
      \piso.data_r_1886_sv2v_reg  <= 1'b0;
      \piso.data_r_1885_sv2v_reg  <= 1'b0;
      \piso.data_r_1884_sv2v_reg  <= 1'b0;
      \piso.data_r_1883_sv2v_reg  <= 1'b0;
      \piso.data_r_1882_sv2v_reg  <= 1'b0;
      \piso.data_r_1881_sv2v_reg  <= 1'b0;
      \piso.data_r_1880_sv2v_reg  <= 1'b0;
      \piso.data_r_1879_sv2v_reg  <= 1'b0;
      \piso.data_r_1878_sv2v_reg  <= 1'b0;
      \piso.data_r_1877_sv2v_reg  <= 1'b0;
      \piso.data_r_1876_sv2v_reg  <= 1'b0;
      \piso.data_r_1875_sv2v_reg  <= 1'b0;
      \piso.data_r_1874_sv2v_reg  <= 1'b0;
      \piso.data_r_1873_sv2v_reg  <= 1'b0;
      \piso.data_r_1872_sv2v_reg  <= 1'b0;
      \piso.data_r_1871_sv2v_reg  <= 1'b0;
      \piso.data_r_1870_sv2v_reg  <= 1'b0;
      \piso.data_r_1869_sv2v_reg  <= 1'b0;
      \piso.data_r_1868_sv2v_reg  <= 1'b0;
      \piso.data_r_1867_sv2v_reg  <= 1'b0;
      \piso.data_r_1866_sv2v_reg  <= 1'b0;
      \piso.data_r_1865_sv2v_reg  <= 1'b0;
      \piso.data_r_1864_sv2v_reg  <= 1'b0;
      \piso.data_r_1863_sv2v_reg  <= 1'b0;
      \piso.data_r_1862_sv2v_reg  <= 1'b0;
      \piso.data_r_1861_sv2v_reg  <= 1'b0;
      \piso.data_r_1860_sv2v_reg  <= 1'b0;
      \piso.data_r_1859_sv2v_reg  <= 1'b0;
      \piso.data_r_1858_sv2v_reg  <= 1'b0;
      \piso.data_r_1857_sv2v_reg  <= 1'b0;
      \piso.data_r_1856_sv2v_reg  <= 1'b0;
      \piso.data_r_1855_sv2v_reg  <= 1'b0;
      \piso.data_r_1854_sv2v_reg  <= 1'b0;
      \piso.data_r_1853_sv2v_reg  <= 1'b0;
      \piso.data_r_1852_sv2v_reg  <= 1'b0;
      \piso.data_r_1851_sv2v_reg  <= 1'b0;
      \piso.data_r_1850_sv2v_reg  <= 1'b0;
      \piso.data_r_1849_sv2v_reg  <= 1'b0;
      \piso.data_r_1848_sv2v_reg  <= 1'b0;
      \piso.data_r_1847_sv2v_reg  <= 1'b0;
      \piso.data_r_1846_sv2v_reg  <= 1'b0;
      \piso.data_r_1845_sv2v_reg  <= 1'b0;
      \piso.data_r_1844_sv2v_reg  <= 1'b0;
      \piso.data_r_1843_sv2v_reg  <= 1'b0;
      \piso.data_r_1842_sv2v_reg  <= 1'b0;
      \piso.data_r_1841_sv2v_reg  <= 1'b0;
      \piso.data_r_1840_sv2v_reg  <= 1'b0;
      \piso.data_r_1839_sv2v_reg  <= 1'b0;
      \piso.data_r_1838_sv2v_reg  <= 1'b0;
      \piso.data_r_1837_sv2v_reg  <= 1'b0;
      \piso.data_r_1836_sv2v_reg  <= 1'b0;
      \piso.data_r_1835_sv2v_reg  <= 1'b0;
      \piso.data_r_1834_sv2v_reg  <= 1'b0;
      \piso.data_r_1833_sv2v_reg  <= 1'b0;
      \piso.data_r_1832_sv2v_reg  <= 1'b0;
      \piso.data_r_1831_sv2v_reg  <= 1'b0;
      \piso.data_r_1830_sv2v_reg  <= 1'b0;
      \piso.data_r_1829_sv2v_reg  <= 1'b0;
      \piso.data_r_1828_sv2v_reg  <= 1'b0;
      \piso.data_r_1827_sv2v_reg  <= 1'b0;
      \piso.data_r_1826_sv2v_reg  <= 1'b0;
      \piso.data_r_1825_sv2v_reg  <= 1'b0;
      \piso.data_r_1824_sv2v_reg  <= 1'b0;
      \piso.data_r_1823_sv2v_reg  <= 1'b0;
      \piso.data_r_1822_sv2v_reg  <= 1'b0;
      \piso.data_r_1821_sv2v_reg  <= 1'b0;
      \piso.data_r_1820_sv2v_reg  <= 1'b0;
      \piso.data_r_1819_sv2v_reg  <= 1'b0;
      \piso.data_r_1818_sv2v_reg  <= 1'b0;
      \piso.data_r_1817_sv2v_reg  <= 1'b0;
      \piso.data_r_1816_sv2v_reg  <= 1'b0;
      \piso.data_r_1815_sv2v_reg  <= 1'b0;
      \piso.data_r_1814_sv2v_reg  <= 1'b0;
      \piso.data_r_1813_sv2v_reg  <= 1'b0;
      \piso.data_r_1812_sv2v_reg  <= 1'b0;
      \piso.data_r_1811_sv2v_reg  <= 1'b0;
      \piso.data_r_1810_sv2v_reg  <= 1'b0;
      \piso.data_r_1809_sv2v_reg  <= 1'b0;
      \piso.data_r_1808_sv2v_reg  <= 1'b0;
      \piso.data_r_1807_sv2v_reg  <= 1'b0;
      \piso.data_r_1806_sv2v_reg  <= 1'b0;
      \piso.data_r_1805_sv2v_reg  <= 1'b0;
      \piso.data_r_1804_sv2v_reg  <= 1'b0;
      \piso.data_r_1803_sv2v_reg  <= 1'b0;
      \piso.data_r_1802_sv2v_reg  <= 1'b0;
      \piso.data_r_1801_sv2v_reg  <= 1'b0;
      \piso.data_r_1800_sv2v_reg  <= 1'b0;
      \piso.data_r_1799_sv2v_reg  <= 1'b0;
      \piso.data_r_1798_sv2v_reg  <= 1'b0;
      \piso.data_r_1797_sv2v_reg  <= 1'b0;
      \piso.data_r_1796_sv2v_reg  <= 1'b0;
      \piso.data_r_1795_sv2v_reg  <= 1'b0;
      \piso.data_r_1794_sv2v_reg  <= 1'b0;
      \piso.data_r_1793_sv2v_reg  <= 1'b0;
      \piso.data_r_1792_sv2v_reg  <= 1'b0;
      \piso.data_r_1791_sv2v_reg  <= 1'b0;
      \piso.data_r_1790_sv2v_reg  <= 1'b0;
      \piso.data_r_1789_sv2v_reg  <= 1'b0;
      \piso.data_r_1788_sv2v_reg  <= 1'b0;
      \piso.data_r_1787_sv2v_reg  <= 1'b0;
      \piso.data_r_1786_sv2v_reg  <= 1'b0;
      \piso.data_r_1785_sv2v_reg  <= 1'b0;
      \piso.data_r_1784_sv2v_reg  <= 1'b0;
      \piso.data_r_1783_sv2v_reg  <= 1'b0;
      \piso.data_r_1782_sv2v_reg  <= 1'b0;
      \piso.data_r_1781_sv2v_reg  <= 1'b0;
      \piso.data_r_1780_sv2v_reg  <= 1'b0;
      \piso.data_r_1779_sv2v_reg  <= 1'b0;
      \piso.data_r_1778_sv2v_reg  <= 1'b0;
      \piso.data_r_1777_sv2v_reg  <= 1'b0;
      \piso.data_r_1776_sv2v_reg  <= 1'b0;
      \piso.data_r_1775_sv2v_reg  <= 1'b0;
      \piso.data_r_1774_sv2v_reg  <= 1'b0;
      \piso.data_r_1773_sv2v_reg  <= 1'b0;
      \piso.data_r_1772_sv2v_reg  <= 1'b0;
      \piso.data_r_1771_sv2v_reg  <= 1'b0;
      \piso.data_r_1770_sv2v_reg  <= 1'b0;
      \piso.data_r_1769_sv2v_reg  <= 1'b0;
      \piso.data_r_1768_sv2v_reg  <= 1'b0;
      \piso.data_r_1767_sv2v_reg  <= 1'b0;
      \piso.data_r_1766_sv2v_reg  <= 1'b0;
      \piso.data_r_1765_sv2v_reg  <= 1'b0;
      \piso.data_r_1764_sv2v_reg  <= 1'b0;
      \piso.data_r_1763_sv2v_reg  <= 1'b0;
      \piso.data_r_1762_sv2v_reg  <= 1'b0;
      \piso.data_r_1761_sv2v_reg  <= 1'b0;
      \piso.data_r_1760_sv2v_reg  <= 1'b0;
      \piso.data_r_1759_sv2v_reg  <= 1'b0;
      \piso.data_r_1758_sv2v_reg  <= 1'b0;
      \piso.data_r_1757_sv2v_reg  <= 1'b0;
      \piso.data_r_1756_sv2v_reg  <= 1'b0;
      \piso.data_r_1755_sv2v_reg  <= 1'b0;
      \piso.data_r_1754_sv2v_reg  <= 1'b0;
      \piso.data_r_1753_sv2v_reg  <= 1'b0;
      \piso.data_r_1752_sv2v_reg  <= 1'b0;
      \piso.data_r_1751_sv2v_reg  <= 1'b0;
      \piso.data_r_1750_sv2v_reg  <= 1'b0;
      \piso.data_r_1749_sv2v_reg  <= 1'b0;
      \piso.data_r_1748_sv2v_reg  <= 1'b0;
      \piso.data_r_1747_sv2v_reg  <= 1'b0;
      \piso.data_r_1746_sv2v_reg  <= 1'b0;
      \piso.data_r_1745_sv2v_reg  <= 1'b0;
      \piso.data_r_1744_sv2v_reg  <= 1'b0;
      \piso.data_r_1743_sv2v_reg  <= 1'b0;
      \piso.data_r_1742_sv2v_reg  <= 1'b0;
      \piso.data_r_1741_sv2v_reg  <= 1'b0;
      \piso.data_r_1740_sv2v_reg  <= 1'b0;
      \piso.data_r_1739_sv2v_reg  <= 1'b0;
      \piso.data_r_1738_sv2v_reg  <= 1'b0;
      \piso.data_r_1737_sv2v_reg  <= 1'b0;
      \piso.data_r_1736_sv2v_reg  <= 1'b0;
      \piso.data_r_1735_sv2v_reg  <= 1'b0;
      \piso.data_r_1734_sv2v_reg  <= 1'b0;
      \piso.data_r_1733_sv2v_reg  <= 1'b0;
      \piso.data_r_1732_sv2v_reg  <= 1'b0;
      \piso.data_r_1731_sv2v_reg  <= 1'b0;
      \piso.data_r_1730_sv2v_reg  <= 1'b0;
      \piso.data_r_1729_sv2v_reg  <= 1'b0;
      \piso.data_r_1728_sv2v_reg  <= 1'b0;
      \piso.data_r_1727_sv2v_reg  <= 1'b0;
      \piso.data_r_1726_sv2v_reg  <= 1'b0;
      \piso.data_r_1725_sv2v_reg  <= 1'b0;
      \piso.data_r_1724_sv2v_reg  <= 1'b0;
      \piso.data_r_1723_sv2v_reg  <= 1'b0;
      \piso.data_r_1722_sv2v_reg  <= 1'b0;
      \piso.data_r_1721_sv2v_reg  <= 1'b0;
      \piso.data_r_1720_sv2v_reg  <= 1'b0;
      \piso.data_r_1719_sv2v_reg  <= 1'b0;
      \piso.data_r_1718_sv2v_reg  <= 1'b0;
      \piso.data_r_1717_sv2v_reg  <= 1'b0;
      \piso.data_r_1716_sv2v_reg  <= 1'b0;
      \piso.data_r_1715_sv2v_reg  <= 1'b0;
      \piso.data_r_1714_sv2v_reg  <= 1'b0;
      \piso.data_r_1713_sv2v_reg  <= 1'b0;
      \piso.data_r_1712_sv2v_reg  <= 1'b0;
      \piso.data_r_1711_sv2v_reg  <= 1'b0;
      \piso.data_r_1710_sv2v_reg  <= 1'b0;
      \piso.data_r_1709_sv2v_reg  <= 1'b0;
      \piso.data_r_1708_sv2v_reg  <= 1'b0;
      \piso.data_r_1707_sv2v_reg  <= 1'b0;
      \piso.data_r_1706_sv2v_reg  <= 1'b0;
      \piso.data_r_1705_sv2v_reg  <= 1'b0;
      \piso.data_r_1704_sv2v_reg  <= 1'b0;
      \piso.data_r_1703_sv2v_reg  <= 1'b0;
      \piso.data_r_1702_sv2v_reg  <= 1'b0;
      \piso.data_r_1701_sv2v_reg  <= 1'b0;
      \piso.data_r_1700_sv2v_reg  <= 1'b0;
      \piso.data_r_1699_sv2v_reg  <= 1'b0;
      \piso.data_r_1698_sv2v_reg  <= 1'b0;
      \piso.data_r_1697_sv2v_reg  <= 1'b0;
      \piso.data_r_1696_sv2v_reg  <= 1'b0;
      \piso.data_r_1695_sv2v_reg  <= 1'b0;
      \piso.data_r_1694_sv2v_reg  <= 1'b0;
      \piso.data_r_1693_sv2v_reg  <= 1'b0;
      \piso.data_r_1692_sv2v_reg  <= 1'b0;
      \piso.data_r_1691_sv2v_reg  <= 1'b0;
      \piso.data_r_1690_sv2v_reg  <= 1'b0;
      \piso.data_r_1689_sv2v_reg  <= 1'b0;
      \piso.data_r_1688_sv2v_reg  <= 1'b0;
      \piso.data_r_1687_sv2v_reg  <= 1'b0;
      \piso.data_r_1686_sv2v_reg  <= 1'b0;
      \piso.data_r_1685_sv2v_reg  <= 1'b0;
      \piso.data_r_1684_sv2v_reg  <= 1'b0;
      \piso.data_r_1683_sv2v_reg  <= 1'b0;
      \piso.data_r_1682_sv2v_reg  <= 1'b0;
      \piso.data_r_1681_sv2v_reg  <= 1'b0;
      \piso.data_r_1680_sv2v_reg  <= 1'b0;
      \piso.data_r_1679_sv2v_reg  <= 1'b0;
      \piso.data_r_1678_sv2v_reg  <= 1'b0;
      \piso.data_r_1677_sv2v_reg  <= 1'b0;
      \piso.data_r_1676_sv2v_reg  <= 1'b0;
      \piso.data_r_1675_sv2v_reg  <= 1'b0;
      \piso.data_r_1674_sv2v_reg  <= 1'b0;
      \piso.data_r_1673_sv2v_reg  <= 1'b0;
      \piso.data_r_1672_sv2v_reg  <= 1'b0;
      \piso.data_r_1671_sv2v_reg  <= 1'b0;
      \piso.data_r_1670_sv2v_reg  <= 1'b0;
      \piso.data_r_1669_sv2v_reg  <= 1'b0;
      \piso.data_r_1668_sv2v_reg  <= 1'b0;
      \piso.data_r_1667_sv2v_reg  <= 1'b0;
      \piso.data_r_1666_sv2v_reg  <= 1'b0;
      \piso.data_r_1665_sv2v_reg  <= 1'b0;
      \piso.data_r_1664_sv2v_reg  <= 1'b0;
      \piso.data_r_1663_sv2v_reg  <= 1'b0;
      \piso.data_r_1662_sv2v_reg  <= 1'b0;
      \piso.data_r_1661_sv2v_reg  <= 1'b0;
      \piso.data_r_1660_sv2v_reg  <= 1'b0;
      \piso.data_r_1659_sv2v_reg  <= 1'b0;
      \piso.data_r_1658_sv2v_reg  <= 1'b0;
      \piso.data_r_1657_sv2v_reg  <= 1'b0;
      \piso.data_r_1656_sv2v_reg  <= 1'b0;
      \piso.data_r_1655_sv2v_reg  <= 1'b0;
      \piso.data_r_1654_sv2v_reg  <= 1'b0;
      \piso.data_r_1653_sv2v_reg  <= 1'b0;
      \piso.data_r_1652_sv2v_reg  <= 1'b0;
      \piso.data_r_1651_sv2v_reg  <= 1'b0;
      \piso.data_r_1650_sv2v_reg  <= 1'b0;
      \piso.data_r_1649_sv2v_reg  <= 1'b0;
      \piso.data_r_1648_sv2v_reg  <= 1'b0;
      \piso.data_r_1647_sv2v_reg  <= 1'b0;
      \piso.data_r_1646_sv2v_reg  <= 1'b0;
      \piso.data_r_1645_sv2v_reg  <= 1'b0;
      \piso.data_r_1644_sv2v_reg  <= 1'b0;
      \piso.data_r_1643_sv2v_reg  <= 1'b0;
      \piso.data_r_1642_sv2v_reg  <= 1'b0;
      \piso.data_r_1641_sv2v_reg  <= 1'b0;
      \piso.data_r_1640_sv2v_reg  <= 1'b0;
      \piso.data_r_1639_sv2v_reg  <= 1'b0;
      \piso.data_r_1638_sv2v_reg  <= 1'b0;
      \piso.data_r_1637_sv2v_reg  <= 1'b0;
      \piso.data_r_1636_sv2v_reg  <= 1'b0;
      \piso.data_r_1635_sv2v_reg  <= 1'b0;
      \piso.data_r_1634_sv2v_reg  <= 1'b0;
      \piso.data_r_1633_sv2v_reg  <= 1'b0;
      \piso.data_r_1632_sv2v_reg  <= 1'b0;
      \piso.data_r_1631_sv2v_reg  <= 1'b0;
      \piso.data_r_1630_sv2v_reg  <= 1'b0;
      \piso.data_r_1629_sv2v_reg  <= 1'b0;
      \piso.data_r_1628_sv2v_reg  <= 1'b0;
      \piso.data_r_1627_sv2v_reg  <= 1'b0;
      \piso.data_r_1626_sv2v_reg  <= 1'b0;
      \piso.data_r_1625_sv2v_reg  <= 1'b0;
      \piso.data_r_1624_sv2v_reg  <= 1'b0;
      \piso.data_r_1623_sv2v_reg  <= 1'b0;
      \piso.data_r_1622_sv2v_reg  <= 1'b0;
      \piso.data_r_1621_sv2v_reg  <= 1'b0;
      \piso.data_r_1620_sv2v_reg  <= 1'b0;
      \piso.data_r_1619_sv2v_reg  <= 1'b0;
      \piso.data_r_1618_sv2v_reg  <= 1'b0;
      \piso.data_r_1617_sv2v_reg  <= 1'b0;
      \piso.data_r_1616_sv2v_reg  <= 1'b0;
      \piso.data_r_1615_sv2v_reg  <= 1'b0;
      \piso.data_r_1614_sv2v_reg  <= 1'b0;
      \piso.data_r_1613_sv2v_reg  <= 1'b0;
      \piso.data_r_1612_sv2v_reg  <= 1'b0;
      \piso.data_r_1611_sv2v_reg  <= 1'b0;
      \piso.data_r_1610_sv2v_reg  <= 1'b0;
      \piso.data_r_1609_sv2v_reg  <= 1'b0;
      \piso.data_r_1608_sv2v_reg  <= 1'b0;
      \piso.data_r_1607_sv2v_reg  <= 1'b0;
      \piso.data_r_1606_sv2v_reg  <= 1'b0;
      \piso.data_r_1605_sv2v_reg  <= 1'b0;
      \piso.data_r_1604_sv2v_reg  <= 1'b0;
      \piso.data_r_1603_sv2v_reg  <= 1'b0;
      \piso.data_r_1602_sv2v_reg  <= 1'b0;
      \piso.data_r_1601_sv2v_reg  <= 1'b0;
      \piso.data_r_1600_sv2v_reg  <= 1'b0;
      \piso.data_r_1599_sv2v_reg  <= 1'b0;
      \piso.data_r_1598_sv2v_reg  <= 1'b0;
      \piso.data_r_1597_sv2v_reg  <= 1'b0;
      \piso.data_r_1596_sv2v_reg  <= 1'b0;
      \piso.data_r_1595_sv2v_reg  <= 1'b0;
      \piso.data_r_1594_sv2v_reg  <= 1'b0;
      \piso.data_r_1593_sv2v_reg  <= 1'b0;
      \piso.data_r_1592_sv2v_reg  <= 1'b0;
      \piso.data_r_1591_sv2v_reg  <= 1'b0;
      \piso.data_r_1590_sv2v_reg  <= 1'b0;
      \piso.data_r_1589_sv2v_reg  <= 1'b0;
      \piso.data_r_1588_sv2v_reg  <= 1'b0;
      \piso.data_r_1587_sv2v_reg  <= 1'b0;
      \piso.data_r_1586_sv2v_reg  <= 1'b0;
      \piso.data_r_1585_sv2v_reg  <= 1'b0;
      \piso.data_r_1584_sv2v_reg  <= 1'b0;
      \piso.data_r_1583_sv2v_reg  <= 1'b0;
      \piso.data_r_1582_sv2v_reg  <= 1'b0;
      \piso.data_r_1581_sv2v_reg  <= 1'b0;
      \piso.data_r_1580_sv2v_reg  <= 1'b0;
      \piso.data_r_1579_sv2v_reg  <= 1'b0;
      \piso.data_r_1578_sv2v_reg  <= 1'b0;
      \piso.data_r_1577_sv2v_reg  <= 1'b0;
      \piso.data_r_1576_sv2v_reg  <= 1'b0;
      \piso.data_r_1575_sv2v_reg  <= 1'b0;
      \piso.data_r_1574_sv2v_reg  <= 1'b0;
      \piso.data_r_1573_sv2v_reg  <= 1'b0;
      \piso.data_r_1572_sv2v_reg  <= 1'b0;
      \piso.data_r_1571_sv2v_reg  <= 1'b0;
      \piso.data_r_1570_sv2v_reg  <= 1'b0;
      \piso.data_r_1569_sv2v_reg  <= 1'b0;
      \piso.data_r_1568_sv2v_reg  <= 1'b0;
      \piso.data_r_1567_sv2v_reg  <= 1'b0;
      \piso.data_r_1566_sv2v_reg  <= 1'b0;
      \piso.data_r_1565_sv2v_reg  <= 1'b0;
      \piso.data_r_1564_sv2v_reg  <= 1'b0;
      \piso.data_r_1563_sv2v_reg  <= 1'b0;
      \piso.data_r_1562_sv2v_reg  <= 1'b0;
      \piso.data_r_1561_sv2v_reg  <= 1'b0;
      \piso.data_r_1560_sv2v_reg  <= 1'b0;
      \piso.data_r_1559_sv2v_reg  <= 1'b0;
      \piso.data_r_1558_sv2v_reg  <= 1'b0;
      \piso.data_r_1557_sv2v_reg  <= 1'b0;
      \piso.data_r_1556_sv2v_reg  <= 1'b0;
      \piso.data_r_1555_sv2v_reg  <= 1'b0;
      \piso.data_r_1554_sv2v_reg  <= 1'b0;
      \piso.data_r_1553_sv2v_reg  <= 1'b0;
      \piso.data_r_1552_sv2v_reg  <= 1'b0;
      \piso.data_r_1551_sv2v_reg  <= 1'b0;
      \piso.data_r_1550_sv2v_reg  <= 1'b0;
      \piso.data_r_1549_sv2v_reg  <= 1'b0;
      \piso.data_r_1548_sv2v_reg  <= 1'b0;
      \piso.data_r_1547_sv2v_reg  <= 1'b0;
      \piso.data_r_1546_sv2v_reg  <= 1'b0;
      \piso.data_r_1545_sv2v_reg  <= 1'b0;
      \piso.data_r_1544_sv2v_reg  <= 1'b0;
      \piso.data_r_1543_sv2v_reg  <= 1'b0;
      \piso.data_r_1542_sv2v_reg  <= 1'b0;
      \piso.data_r_1541_sv2v_reg  <= 1'b0;
      \piso.data_r_1540_sv2v_reg  <= 1'b0;
      \piso.data_r_1539_sv2v_reg  <= 1'b0;
      \piso.data_r_1538_sv2v_reg  <= 1'b0;
      \piso.data_r_1537_sv2v_reg  <= 1'b0;
      \piso.data_r_1536_sv2v_reg  <= 1'b0;
      \piso.data_r_1535_sv2v_reg  <= 1'b0;
      \piso.data_r_1534_sv2v_reg  <= 1'b0;
      \piso.data_r_1533_sv2v_reg  <= 1'b0;
      \piso.data_r_1532_sv2v_reg  <= 1'b0;
      \piso.data_r_1531_sv2v_reg  <= 1'b0;
      \piso.data_r_1530_sv2v_reg  <= 1'b0;
      \piso.data_r_1529_sv2v_reg  <= 1'b0;
      \piso.data_r_1528_sv2v_reg  <= 1'b0;
      \piso.data_r_1527_sv2v_reg  <= 1'b0;
      \piso.data_r_1526_sv2v_reg  <= 1'b0;
      \piso.data_r_1525_sv2v_reg  <= 1'b0;
      \piso.data_r_1524_sv2v_reg  <= 1'b0;
      \piso.data_r_1523_sv2v_reg  <= 1'b0;
      \piso.data_r_1522_sv2v_reg  <= 1'b0;
      \piso.data_r_1521_sv2v_reg  <= 1'b0;
      \piso.data_r_1520_sv2v_reg  <= 1'b0;
      \piso.data_r_1519_sv2v_reg  <= 1'b0;
      \piso.data_r_1518_sv2v_reg  <= 1'b0;
      \piso.data_r_1517_sv2v_reg  <= 1'b0;
      \piso.data_r_1516_sv2v_reg  <= 1'b0;
      \piso.data_r_1515_sv2v_reg  <= 1'b0;
      \piso.data_r_1514_sv2v_reg  <= 1'b0;
      \piso.data_r_1513_sv2v_reg  <= 1'b0;
      \piso.data_r_1512_sv2v_reg  <= 1'b0;
      \piso.data_r_1511_sv2v_reg  <= 1'b0;
      \piso.data_r_1510_sv2v_reg  <= 1'b0;
      \piso.data_r_1509_sv2v_reg  <= 1'b0;
      \piso.data_r_1508_sv2v_reg  <= 1'b0;
      \piso.data_r_1507_sv2v_reg  <= 1'b0;
      \piso.data_r_1506_sv2v_reg  <= 1'b0;
      \piso.data_r_1505_sv2v_reg  <= 1'b0;
      \piso.data_r_1504_sv2v_reg  <= 1'b0;
      \piso.data_r_1503_sv2v_reg  <= 1'b0;
      \piso.data_r_1502_sv2v_reg  <= 1'b0;
      \piso.data_r_1501_sv2v_reg  <= 1'b0;
      \piso.data_r_1500_sv2v_reg  <= 1'b0;
      \piso.data_r_1499_sv2v_reg  <= 1'b0;
      \piso.data_r_1498_sv2v_reg  <= 1'b0;
      \piso.data_r_1497_sv2v_reg  <= 1'b0;
      \piso.data_r_1496_sv2v_reg  <= 1'b0;
      \piso.data_r_1495_sv2v_reg  <= 1'b0;
      \piso.data_r_1494_sv2v_reg  <= 1'b0;
      \piso.data_r_1493_sv2v_reg  <= 1'b0;
      \piso.data_r_1492_sv2v_reg  <= 1'b0;
      \piso.data_r_1491_sv2v_reg  <= 1'b0;
      \piso.data_r_1490_sv2v_reg  <= 1'b0;
      \piso.data_r_1489_sv2v_reg  <= 1'b0;
      \piso.data_r_1488_sv2v_reg  <= 1'b0;
      \piso.data_r_1487_sv2v_reg  <= 1'b0;
      \piso.data_r_1486_sv2v_reg  <= 1'b0;
      \piso.data_r_1485_sv2v_reg  <= 1'b0;
      \piso.data_r_1484_sv2v_reg  <= 1'b0;
      \piso.data_r_1483_sv2v_reg  <= 1'b0;
      \piso.data_r_1482_sv2v_reg  <= 1'b0;
      \piso.data_r_1481_sv2v_reg  <= 1'b0;
      \piso.data_r_1480_sv2v_reg  <= 1'b0;
      \piso.data_r_1479_sv2v_reg  <= 1'b0;
      \piso.data_r_1478_sv2v_reg  <= 1'b0;
      \piso.data_r_1477_sv2v_reg  <= 1'b0;
      \piso.data_r_1476_sv2v_reg  <= 1'b0;
      \piso.data_r_1475_sv2v_reg  <= 1'b0;
      \piso.data_r_1474_sv2v_reg  <= 1'b0;
      \piso.data_r_1473_sv2v_reg  <= 1'b0;
      \piso.data_r_1472_sv2v_reg  <= 1'b0;
      \piso.data_r_1471_sv2v_reg  <= 1'b0;
      \piso.data_r_1470_sv2v_reg  <= 1'b0;
      \piso.data_r_1469_sv2v_reg  <= 1'b0;
      \piso.data_r_1468_sv2v_reg  <= 1'b0;
      \piso.data_r_1467_sv2v_reg  <= 1'b0;
      \piso.data_r_1466_sv2v_reg  <= 1'b0;
      \piso.data_r_1465_sv2v_reg  <= 1'b0;
      \piso.data_r_1464_sv2v_reg  <= 1'b0;
      \piso.data_r_1463_sv2v_reg  <= 1'b0;
      \piso.data_r_1462_sv2v_reg  <= 1'b0;
      \piso.data_r_1461_sv2v_reg  <= 1'b0;
      \piso.data_r_1460_sv2v_reg  <= 1'b0;
      \piso.data_r_1459_sv2v_reg  <= 1'b0;
      \piso.data_r_1458_sv2v_reg  <= 1'b0;
      \piso.data_r_1457_sv2v_reg  <= 1'b0;
      \piso.data_r_1456_sv2v_reg  <= 1'b0;
      \piso.data_r_1455_sv2v_reg  <= 1'b0;
      \piso.data_r_1454_sv2v_reg  <= 1'b0;
      \piso.data_r_1453_sv2v_reg  <= 1'b0;
      \piso.data_r_1452_sv2v_reg  <= 1'b0;
      \piso.data_r_1451_sv2v_reg  <= 1'b0;
      \piso.data_r_1450_sv2v_reg  <= 1'b0;
      \piso.data_r_1449_sv2v_reg  <= 1'b0;
      \piso.data_r_1448_sv2v_reg  <= 1'b0;
      \piso.data_r_1447_sv2v_reg  <= 1'b0;
      \piso.data_r_1446_sv2v_reg  <= 1'b0;
      \piso.data_r_1445_sv2v_reg  <= 1'b0;
      \piso.data_r_1444_sv2v_reg  <= 1'b0;
      \piso.data_r_1443_sv2v_reg  <= 1'b0;
      \piso.data_r_1442_sv2v_reg  <= 1'b0;
      \piso.data_r_1441_sv2v_reg  <= 1'b0;
      \piso.data_r_1440_sv2v_reg  <= 1'b0;
      \piso.data_r_1439_sv2v_reg  <= 1'b0;
      \piso.data_r_1438_sv2v_reg  <= 1'b0;
      \piso.data_r_1437_sv2v_reg  <= 1'b0;
      \piso.data_r_1436_sv2v_reg  <= 1'b0;
      \piso.data_r_1435_sv2v_reg  <= 1'b0;
      \piso.data_r_1434_sv2v_reg  <= 1'b0;
      \piso.data_r_1433_sv2v_reg  <= 1'b0;
      \piso.data_r_1432_sv2v_reg  <= 1'b0;
      \piso.data_r_1431_sv2v_reg  <= 1'b0;
      \piso.data_r_1430_sv2v_reg  <= 1'b0;
      \piso.data_r_1429_sv2v_reg  <= 1'b0;
      \piso.data_r_1428_sv2v_reg  <= 1'b0;
      \piso.data_r_1427_sv2v_reg  <= 1'b0;
      \piso.data_r_1426_sv2v_reg  <= 1'b0;
      \piso.data_r_1425_sv2v_reg  <= 1'b0;
      \piso.data_r_1424_sv2v_reg  <= 1'b0;
      \piso.data_r_1423_sv2v_reg  <= 1'b0;
      \piso.data_r_1422_sv2v_reg  <= 1'b0;
      \piso.data_r_1421_sv2v_reg  <= 1'b0;
      \piso.data_r_1420_sv2v_reg  <= 1'b0;
      \piso.data_r_1419_sv2v_reg  <= 1'b0;
      \piso.data_r_1418_sv2v_reg  <= 1'b0;
      \piso.data_r_1417_sv2v_reg  <= 1'b0;
      \piso.data_r_1416_sv2v_reg  <= 1'b0;
      \piso.data_r_1415_sv2v_reg  <= 1'b0;
      \piso.data_r_1414_sv2v_reg  <= 1'b0;
      \piso.data_r_1413_sv2v_reg  <= 1'b0;
      \piso.data_r_1412_sv2v_reg  <= 1'b0;
      \piso.data_r_1411_sv2v_reg  <= 1'b0;
      \piso.data_r_1410_sv2v_reg  <= 1'b0;
      \piso.data_r_1409_sv2v_reg  <= 1'b0;
      \piso.data_r_1408_sv2v_reg  <= 1'b0;
      \piso.data_r_1407_sv2v_reg  <= 1'b0;
      \piso.data_r_1406_sv2v_reg  <= 1'b0;
      \piso.data_r_1405_sv2v_reg  <= 1'b0;
      \piso.data_r_1404_sv2v_reg  <= 1'b0;
      \piso.data_r_1403_sv2v_reg  <= 1'b0;
      \piso.data_r_1402_sv2v_reg  <= 1'b0;
      \piso.data_r_1401_sv2v_reg  <= 1'b0;
      \piso.data_r_1400_sv2v_reg  <= 1'b0;
      \piso.data_r_1399_sv2v_reg  <= 1'b0;
      \piso.data_r_1398_sv2v_reg  <= 1'b0;
      \piso.data_r_1397_sv2v_reg  <= 1'b0;
      \piso.data_r_1396_sv2v_reg  <= 1'b0;
      \piso.data_r_1395_sv2v_reg  <= 1'b0;
      \piso.data_r_1394_sv2v_reg  <= 1'b0;
      \piso.data_r_1393_sv2v_reg  <= 1'b0;
      \piso.data_r_1392_sv2v_reg  <= 1'b0;
      \piso.data_r_1391_sv2v_reg  <= 1'b0;
      \piso.data_r_1390_sv2v_reg  <= 1'b0;
      \piso.data_r_1389_sv2v_reg  <= 1'b0;
      \piso.data_r_1388_sv2v_reg  <= 1'b0;
      \piso.data_r_1387_sv2v_reg  <= 1'b0;
      \piso.data_r_1386_sv2v_reg  <= 1'b0;
      \piso.data_r_1385_sv2v_reg  <= 1'b0;
      \piso.data_r_1384_sv2v_reg  <= 1'b0;
      \piso.data_r_1383_sv2v_reg  <= 1'b0;
      \piso.data_r_1382_sv2v_reg  <= 1'b0;
      \piso.data_r_1381_sv2v_reg  <= 1'b0;
      \piso.data_r_1380_sv2v_reg  <= 1'b0;
      \piso.data_r_1379_sv2v_reg  <= 1'b0;
      \piso.data_r_1378_sv2v_reg  <= 1'b0;
      \piso.data_r_1377_sv2v_reg  <= 1'b0;
      \piso.data_r_1376_sv2v_reg  <= 1'b0;
      \piso.data_r_1375_sv2v_reg  <= 1'b0;
      \piso.data_r_1374_sv2v_reg  <= 1'b0;
      \piso.data_r_1373_sv2v_reg  <= 1'b0;
      \piso.data_r_1372_sv2v_reg  <= 1'b0;
      \piso.data_r_1371_sv2v_reg  <= 1'b0;
      \piso.data_r_1370_sv2v_reg  <= 1'b0;
      \piso.data_r_1369_sv2v_reg  <= 1'b0;
      \piso.data_r_1368_sv2v_reg  <= 1'b0;
      \piso.data_r_1367_sv2v_reg  <= 1'b0;
      \piso.data_r_1366_sv2v_reg  <= 1'b0;
      \piso.data_r_1365_sv2v_reg  <= 1'b0;
      \piso.data_r_1364_sv2v_reg  <= 1'b0;
      \piso.data_r_1363_sv2v_reg  <= 1'b0;
      \piso.data_r_1362_sv2v_reg  <= 1'b0;
      \piso.data_r_1361_sv2v_reg  <= 1'b0;
      \piso.data_r_1360_sv2v_reg  <= 1'b0;
      \piso.data_r_1359_sv2v_reg  <= 1'b0;
      \piso.data_r_1358_sv2v_reg  <= 1'b0;
      \piso.data_r_1357_sv2v_reg  <= 1'b0;
      \piso.data_r_1356_sv2v_reg  <= 1'b0;
      \piso.data_r_1355_sv2v_reg  <= 1'b0;
      \piso.data_r_1354_sv2v_reg  <= 1'b0;
      \piso.data_r_1353_sv2v_reg  <= 1'b0;
      \piso.data_r_1352_sv2v_reg  <= 1'b0;
      \piso.data_r_1351_sv2v_reg  <= 1'b0;
      \piso.data_r_1350_sv2v_reg  <= 1'b0;
      \piso.data_r_1349_sv2v_reg  <= 1'b0;
      \piso.data_r_1348_sv2v_reg  <= 1'b0;
      \piso.data_r_1347_sv2v_reg  <= 1'b0;
      \piso.data_r_1346_sv2v_reg  <= 1'b0;
      \piso.data_r_1345_sv2v_reg  <= 1'b0;
      \piso.data_r_1344_sv2v_reg  <= 1'b0;
      \piso.data_r_1343_sv2v_reg  <= 1'b0;
      \piso.data_r_1342_sv2v_reg  <= 1'b0;
      \piso.data_r_1341_sv2v_reg  <= 1'b0;
      \piso.data_r_1340_sv2v_reg  <= 1'b0;
      \piso.data_r_1339_sv2v_reg  <= 1'b0;
      \piso.data_r_1338_sv2v_reg  <= 1'b0;
      \piso.data_r_1337_sv2v_reg  <= 1'b0;
      \piso.data_r_1336_sv2v_reg  <= 1'b0;
      \piso.data_r_1335_sv2v_reg  <= 1'b0;
      \piso.data_r_1334_sv2v_reg  <= 1'b0;
      \piso.data_r_1333_sv2v_reg  <= 1'b0;
      \piso.data_r_1332_sv2v_reg  <= 1'b0;
      \piso.data_r_1331_sv2v_reg  <= 1'b0;
      \piso.data_r_1330_sv2v_reg  <= 1'b0;
      \piso.data_r_1329_sv2v_reg  <= 1'b0;
      \piso.data_r_1328_sv2v_reg  <= 1'b0;
      \piso.data_r_1327_sv2v_reg  <= 1'b0;
      \piso.data_r_1326_sv2v_reg  <= 1'b0;
      \piso.data_r_1325_sv2v_reg  <= 1'b0;
      \piso.data_r_1324_sv2v_reg  <= 1'b0;
      \piso.data_r_1323_sv2v_reg  <= 1'b0;
      \piso.data_r_1322_sv2v_reg  <= 1'b0;
      \piso.data_r_1321_sv2v_reg  <= 1'b0;
      \piso.data_r_1320_sv2v_reg  <= 1'b0;
      \piso.data_r_1319_sv2v_reg  <= 1'b0;
      \piso.data_r_1318_sv2v_reg  <= 1'b0;
      \piso.data_r_1317_sv2v_reg  <= 1'b0;
      \piso.data_r_1316_sv2v_reg  <= 1'b0;
      \piso.data_r_1315_sv2v_reg  <= 1'b0;
      \piso.data_r_1314_sv2v_reg  <= 1'b0;
      \piso.data_r_1313_sv2v_reg  <= 1'b0;
      \piso.data_r_1312_sv2v_reg  <= 1'b0;
      \piso.data_r_1311_sv2v_reg  <= 1'b0;
      \piso.data_r_1310_sv2v_reg  <= 1'b0;
      \piso.data_r_1309_sv2v_reg  <= 1'b0;
      \piso.data_r_1308_sv2v_reg  <= 1'b0;
      \piso.data_r_1307_sv2v_reg  <= 1'b0;
      \piso.data_r_1306_sv2v_reg  <= 1'b0;
      \piso.data_r_1305_sv2v_reg  <= 1'b0;
      \piso.data_r_1304_sv2v_reg  <= 1'b0;
      \piso.data_r_1303_sv2v_reg  <= 1'b0;
      \piso.data_r_1302_sv2v_reg  <= 1'b0;
      \piso.data_r_1301_sv2v_reg  <= 1'b0;
      \piso.data_r_1300_sv2v_reg  <= 1'b0;
      \piso.data_r_1299_sv2v_reg  <= 1'b0;
      \piso.data_r_1298_sv2v_reg  <= 1'b0;
      \piso.data_r_1297_sv2v_reg  <= 1'b0;
      \piso.data_r_1296_sv2v_reg  <= 1'b0;
      \piso.data_r_1295_sv2v_reg  <= 1'b0;
      \piso.data_r_1294_sv2v_reg  <= 1'b0;
      \piso.data_r_1293_sv2v_reg  <= 1'b0;
      \piso.data_r_1292_sv2v_reg  <= 1'b0;
      \piso.data_r_1291_sv2v_reg  <= 1'b0;
      \piso.data_r_1290_sv2v_reg  <= 1'b0;
      \piso.data_r_1289_sv2v_reg  <= 1'b0;
      \piso.data_r_1288_sv2v_reg  <= 1'b0;
      \piso.data_r_1287_sv2v_reg  <= 1'b0;
      \piso.data_r_1286_sv2v_reg  <= 1'b0;
      \piso.data_r_1285_sv2v_reg  <= 1'b0;
      \piso.data_r_1284_sv2v_reg  <= 1'b0;
      \piso.data_r_1283_sv2v_reg  <= 1'b0;
      \piso.data_r_1282_sv2v_reg  <= 1'b0;
      \piso.data_r_1281_sv2v_reg  <= 1'b0;
      \piso.data_r_1280_sv2v_reg  <= 1'b0;
      \piso.data_r_1279_sv2v_reg  <= 1'b0;
      \piso.data_r_1278_sv2v_reg  <= 1'b0;
      \piso.data_r_1277_sv2v_reg  <= 1'b0;
      \piso.data_r_1276_sv2v_reg  <= 1'b0;
      \piso.data_r_1275_sv2v_reg  <= 1'b0;
      \piso.data_r_1274_sv2v_reg  <= 1'b0;
      \piso.data_r_1273_sv2v_reg  <= 1'b0;
      \piso.data_r_1272_sv2v_reg  <= 1'b0;
      \piso.data_r_1271_sv2v_reg  <= 1'b0;
      \piso.data_r_1270_sv2v_reg  <= 1'b0;
      \piso.data_r_1269_sv2v_reg  <= 1'b0;
      \piso.data_r_1268_sv2v_reg  <= 1'b0;
      \piso.data_r_1267_sv2v_reg  <= 1'b0;
      \piso.data_r_1266_sv2v_reg  <= 1'b0;
      \piso.data_r_1265_sv2v_reg  <= 1'b0;
      \piso.data_r_1264_sv2v_reg  <= 1'b0;
      \piso.data_r_1263_sv2v_reg  <= 1'b0;
      \piso.data_r_1262_sv2v_reg  <= 1'b0;
      \piso.data_r_1261_sv2v_reg  <= 1'b0;
      \piso.data_r_1260_sv2v_reg  <= 1'b0;
      \piso.data_r_1259_sv2v_reg  <= 1'b0;
      \piso.data_r_1258_sv2v_reg  <= 1'b0;
      \piso.data_r_1257_sv2v_reg  <= 1'b0;
      \piso.data_r_1256_sv2v_reg  <= 1'b0;
      \piso.data_r_1255_sv2v_reg  <= 1'b0;
      \piso.data_r_1254_sv2v_reg  <= 1'b0;
      \piso.data_r_1253_sv2v_reg  <= 1'b0;
      \piso.data_r_1252_sv2v_reg  <= 1'b0;
      \piso.data_r_1251_sv2v_reg  <= 1'b0;
      \piso.data_r_1250_sv2v_reg  <= 1'b0;
      \piso.data_r_1249_sv2v_reg  <= 1'b0;
      \piso.data_r_1248_sv2v_reg  <= 1'b0;
      \piso.data_r_1247_sv2v_reg  <= 1'b0;
      \piso.data_r_1246_sv2v_reg  <= 1'b0;
      \piso.data_r_1245_sv2v_reg  <= 1'b0;
      \piso.data_r_1244_sv2v_reg  <= 1'b0;
      \piso.data_r_1243_sv2v_reg  <= 1'b0;
      \piso.data_r_1242_sv2v_reg  <= 1'b0;
      \piso.data_r_1241_sv2v_reg  <= 1'b0;
      \piso.data_r_1240_sv2v_reg  <= 1'b0;
      \piso.data_r_1239_sv2v_reg  <= 1'b0;
      \piso.data_r_1238_sv2v_reg  <= 1'b0;
      \piso.data_r_1237_sv2v_reg  <= 1'b0;
      \piso.data_r_1236_sv2v_reg  <= 1'b0;
      \piso.data_r_1235_sv2v_reg  <= 1'b0;
      \piso.data_r_1234_sv2v_reg  <= 1'b0;
      \piso.data_r_1233_sv2v_reg  <= 1'b0;
      \piso.data_r_1232_sv2v_reg  <= 1'b0;
      \piso.data_r_1231_sv2v_reg  <= 1'b0;
      \piso.data_r_1230_sv2v_reg  <= 1'b0;
      \piso.data_r_1229_sv2v_reg  <= 1'b0;
      \piso.data_r_1228_sv2v_reg  <= 1'b0;
      \piso.data_r_1227_sv2v_reg  <= 1'b0;
      \piso.data_r_1226_sv2v_reg  <= 1'b0;
      \piso.data_r_1225_sv2v_reg  <= 1'b0;
      \piso.data_r_1224_sv2v_reg  <= 1'b0;
      \piso.data_r_1223_sv2v_reg  <= 1'b0;
      \piso.data_r_1222_sv2v_reg  <= 1'b0;
      \piso.data_r_1221_sv2v_reg  <= 1'b0;
      \piso.data_r_1220_sv2v_reg  <= 1'b0;
      \piso.data_r_1219_sv2v_reg  <= 1'b0;
      \piso.data_r_1218_sv2v_reg  <= 1'b0;
      \piso.data_r_1217_sv2v_reg  <= 1'b0;
      \piso.data_r_1216_sv2v_reg  <= 1'b0;
      \piso.data_r_1215_sv2v_reg  <= 1'b0;
      \piso.data_r_1214_sv2v_reg  <= 1'b0;
      \piso.data_r_1213_sv2v_reg  <= 1'b0;
      \piso.data_r_1212_sv2v_reg  <= 1'b0;
      \piso.data_r_1211_sv2v_reg  <= 1'b0;
      \piso.data_r_1210_sv2v_reg  <= 1'b0;
      \piso.data_r_1209_sv2v_reg  <= 1'b0;
      \piso.data_r_1208_sv2v_reg  <= 1'b0;
      \piso.data_r_1207_sv2v_reg  <= 1'b0;
      \piso.data_r_1206_sv2v_reg  <= 1'b0;
      \piso.data_r_1205_sv2v_reg  <= 1'b0;
      \piso.data_r_1204_sv2v_reg  <= 1'b0;
      \piso.data_r_1203_sv2v_reg  <= 1'b0;
      \piso.data_r_1202_sv2v_reg  <= 1'b0;
      \piso.data_r_1201_sv2v_reg  <= 1'b0;
      \piso.data_r_1200_sv2v_reg  <= 1'b0;
      \piso.data_r_1199_sv2v_reg  <= 1'b0;
      \piso.data_r_1198_sv2v_reg  <= 1'b0;
      \piso.data_r_1197_sv2v_reg  <= 1'b0;
      \piso.data_r_1196_sv2v_reg  <= 1'b0;
      \piso.data_r_1195_sv2v_reg  <= 1'b0;
      \piso.data_r_1194_sv2v_reg  <= 1'b0;
      \piso.data_r_1193_sv2v_reg  <= 1'b0;
      \piso.data_r_1192_sv2v_reg  <= 1'b0;
      \piso.data_r_1191_sv2v_reg  <= 1'b0;
      \piso.data_r_1190_sv2v_reg  <= 1'b0;
      \piso.data_r_1189_sv2v_reg  <= 1'b0;
      \piso.data_r_1188_sv2v_reg  <= 1'b0;
      \piso.data_r_1187_sv2v_reg  <= 1'b0;
      \piso.data_r_1186_sv2v_reg  <= 1'b0;
      \piso.data_r_1185_sv2v_reg  <= 1'b0;
      \piso.data_r_1184_sv2v_reg  <= 1'b0;
      \piso.data_r_1183_sv2v_reg  <= 1'b0;
      \piso.data_r_1182_sv2v_reg  <= 1'b0;
      \piso.data_r_1181_sv2v_reg  <= 1'b0;
      \piso.data_r_1180_sv2v_reg  <= 1'b0;
      \piso.data_r_1179_sv2v_reg  <= 1'b0;
      \piso.data_r_1178_sv2v_reg  <= 1'b0;
      \piso.data_r_1177_sv2v_reg  <= 1'b0;
      \piso.data_r_1176_sv2v_reg  <= 1'b0;
      \piso.data_r_1175_sv2v_reg  <= 1'b0;
      \piso.data_r_1174_sv2v_reg  <= 1'b0;
      \piso.data_r_1173_sv2v_reg  <= 1'b0;
      \piso.data_r_1172_sv2v_reg  <= 1'b0;
      \piso.data_r_1171_sv2v_reg  <= 1'b0;
      \piso.data_r_1170_sv2v_reg  <= 1'b0;
      \piso.data_r_1169_sv2v_reg  <= 1'b0;
      \piso.data_r_1168_sv2v_reg  <= 1'b0;
      \piso.data_r_1167_sv2v_reg  <= 1'b0;
      \piso.data_r_1166_sv2v_reg  <= 1'b0;
      \piso.data_r_1165_sv2v_reg  <= 1'b0;
      \piso.data_r_1164_sv2v_reg  <= 1'b0;
      \piso.data_r_1163_sv2v_reg  <= 1'b0;
      \piso.data_r_1162_sv2v_reg  <= 1'b0;
      \piso.data_r_1161_sv2v_reg  <= 1'b0;
      \piso.data_r_1160_sv2v_reg  <= 1'b0;
      \piso.data_r_1159_sv2v_reg  <= 1'b0;
      \piso.data_r_1158_sv2v_reg  <= 1'b0;
      \piso.data_r_1157_sv2v_reg  <= 1'b0;
      \piso.data_r_1156_sv2v_reg  <= 1'b0;
      \piso.data_r_1155_sv2v_reg  <= 1'b0;
      \piso.data_r_1154_sv2v_reg  <= 1'b0;
      \piso.data_r_1153_sv2v_reg  <= 1'b0;
      \piso.data_r_1152_sv2v_reg  <= 1'b0;
      \piso.data_r_1151_sv2v_reg  <= 1'b0;
      \piso.data_r_1150_sv2v_reg  <= 1'b0;
      \piso.data_r_1149_sv2v_reg  <= 1'b0;
      \piso.data_r_1148_sv2v_reg  <= 1'b0;
      \piso.data_r_1147_sv2v_reg  <= 1'b0;
      \piso.data_r_1146_sv2v_reg  <= 1'b0;
      \piso.data_r_1145_sv2v_reg  <= 1'b0;
      \piso.data_r_1144_sv2v_reg  <= 1'b0;
      \piso.data_r_1143_sv2v_reg  <= 1'b0;
      \piso.data_r_1142_sv2v_reg  <= 1'b0;
      \piso.data_r_1141_sv2v_reg  <= 1'b0;
      \piso.data_r_1140_sv2v_reg  <= 1'b0;
      \piso.data_r_1139_sv2v_reg  <= 1'b0;
      \piso.data_r_1138_sv2v_reg  <= 1'b0;
      \piso.data_r_1137_sv2v_reg  <= 1'b0;
      \piso.data_r_1136_sv2v_reg  <= 1'b0;
      \piso.data_r_1135_sv2v_reg  <= 1'b0;
      \piso.data_r_1134_sv2v_reg  <= 1'b0;
      \piso.data_r_1133_sv2v_reg  <= 1'b0;
      \piso.data_r_1132_sv2v_reg  <= 1'b0;
      \piso.data_r_1131_sv2v_reg  <= 1'b0;
      \piso.data_r_1130_sv2v_reg  <= 1'b0;
      \piso.data_r_1129_sv2v_reg  <= 1'b0;
      \piso.data_r_1128_sv2v_reg  <= 1'b0;
      \piso.data_r_1127_sv2v_reg  <= 1'b0;
      \piso.data_r_1126_sv2v_reg  <= 1'b0;
      \piso.data_r_1125_sv2v_reg  <= 1'b0;
      \piso.data_r_1124_sv2v_reg  <= 1'b0;
      \piso.data_r_1123_sv2v_reg  <= 1'b0;
      \piso.data_r_1122_sv2v_reg  <= 1'b0;
      \piso.data_r_1121_sv2v_reg  <= 1'b0;
      \piso.data_r_1120_sv2v_reg  <= 1'b0;
      \piso.data_r_1119_sv2v_reg  <= 1'b0;
      \piso.data_r_1118_sv2v_reg  <= 1'b0;
      \piso.data_r_1117_sv2v_reg  <= 1'b0;
      \piso.data_r_1116_sv2v_reg  <= 1'b0;
      \piso.data_r_1115_sv2v_reg  <= 1'b0;
      \piso.data_r_1114_sv2v_reg  <= 1'b0;
      \piso.data_r_1113_sv2v_reg  <= 1'b0;
      \piso.data_r_1112_sv2v_reg  <= 1'b0;
      \piso.data_r_1111_sv2v_reg  <= 1'b0;
      \piso.data_r_1110_sv2v_reg  <= 1'b0;
      \piso.data_r_1109_sv2v_reg  <= 1'b0;
      \piso.data_r_1108_sv2v_reg  <= 1'b0;
      \piso.data_r_1107_sv2v_reg  <= 1'b0;
      \piso.data_r_1106_sv2v_reg  <= 1'b0;
      \piso.data_r_1105_sv2v_reg  <= 1'b0;
      \piso.data_r_1104_sv2v_reg  <= 1'b0;
      \piso.data_r_1103_sv2v_reg  <= 1'b0;
      \piso.data_r_1102_sv2v_reg  <= 1'b0;
      \piso.data_r_1101_sv2v_reg  <= 1'b0;
      \piso.data_r_1100_sv2v_reg  <= 1'b0;
      \piso.data_r_1099_sv2v_reg  <= 1'b0;
      \piso.data_r_1098_sv2v_reg  <= 1'b0;
      \piso.data_r_1097_sv2v_reg  <= 1'b0;
      \piso.data_r_1096_sv2v_reg  <= 1'b0;
      \piso.data_r_1095_sv2v_reg  <= 1'b0;
      \piso.data_r_1094_sv2v_reg  <= 1'b0;
      \piso.data_r_1093_sv2v_reg  <= 1'b0;
      \piso.data_r_1092_sv2v_reg  <= 1'b0;
      \piso.data_r_1091_sv2v_reg  <= 1'b0;
      \piso.data_r_1090_sv2v_reg  <= 1'b0;
      \piso.data_r_1089_sv2v_reg  <= 1'b0;
      \piso.data_r_1088_sv2v_reg  <= 1'b0;
      \piso.data_r_1087_sv2v_reg  <= 1'b0;
      \piso.data_r_1086_sv2v_reg  <= 1'b0;
      \piso.data_r_1085_sv2v_reg  <= 1'b0;
      \piso.data_r_1084_sv2v_reg  <= 1'b0;
      \piso.data_r_1083_sv2v_reg  <= 1'b0;
      \piso.data_r_1082_sv2v_reg  <= 1'b0;
      \piso.data_r_1081_sv2v_reg  <= 1'b0;
      \piso.data_r_1080_sv2v_reg  <= 1'b0;
      \piso.data_r_1079_sv2v_reg  <= 1'b0;
      \piso.data_r_1078_sv2v_reg  <= 1'b0;
      \piso.data_r_1077_sv2v_reg  <= 1'b0;
      \piso.data_r_1076_sv2v_reg  <= 1'b0;
      \piso.data_r_1075_sv2v_reg  <= 1'b0;
      \piso.data_r_1074_sv2v_reg  <= 1'b0;
      \piso.data_r_1073_sv2v_reg  <= 1'b0;
      \piso.data_r_1072_sv2v_reg  <= 1'b0;
      \piso.data_r_1071_sv2v_reg  <= 1'b0;
      \piso.data_r_1070_sv2v_reg  <= 1'b0;
      \piso.data_r_1069_sv2v_reg  <= 1'b0;
      \piso.data_r_1068_sv2v_reg  <= 1'b0;
      \piso.data_r_1067_sv2v_reg  <= 1'b0;
      \piso.data_r_1066_sv2v_reg  <= 1'b0;
      \piso.data_r_1065_sv2v_reg  <= 1'b0;
      \piso.data_r_1064_sv2v_reg  <= 1'b0;
      \piso.data_r_1063_sv2v_reg  <= 1'b0;
      \piso.data_r_1062_sv2v_reg  <= 1'b0;
      \piso.data_r_1061_sv2v_reg  <= 1'b0;
      \piso.data_r_1060_sv2v_reg  <= 1'b0;
      \piso.data_r_1059_sv2v_reg  <= 1'b0;
      \piso.data_r_1058_sv2v_reg  <= 1'b0;
      \piso.data_r_1057_sv2v_reg  <= 1'b0;
      \piso.data_r_1056_sv2v_reg  <= 1'b0;
      \piso.data_r_1055_sv2v_reg  <= 1'b0;
      \piso.data_r_1054_sv2v_reg  <= 1'b0;
      \piso.data_r_1053_sv2v_reg  <= 1'b0;
      \piso.data_r_1052_sv2v_reg  <= 1'b0;
      \piso.data_r_1051_sv2v_reg  <= 1'b0;
      \piso.data_r_1050_sv2v_reg  <= 1'b0;
      \piso.data_r_1049_sv2v_reg  <= 1'b0;
      \piso.data_r_1048_sv2v_reg  <= 1'b0;
      \piso.data_r_1047_sv2v_reg  <= 1'b0;
      \piso.data_r_1046_sv2v_reg  <= 1'b0;
      \piso.data_r_1045_sv2v_reg  <= 1'b0;
      \piso.data_r_1044_sv2v_reg  <= 1'b0;
      \piso.data_r_1043_sv2v_reg  <= 1'b0;
      \piso.data_r_1042_sv2v_reg  <= 1'b0;
      \piso.data_r_1041_sv2v_reg  <= 1'b0;
      \piso.data_r_1040_sv2v_reg  <= 1'b0;
      \piso.data_r_1039_sv2v_reg  <= 1'b0;
      \piso.data_r_1038_sv2v_reg  <= 1'b0;
      \piso.data_r_1037_sv2v_reg  <= 1'b0;
      \piso.data_r_1036_sv2v_reg  <= 1'b0;
      \piso.data_r_1035_sv2v_reg  <= 1'b0;
      \piso.data_r_1034_sv2v_reg  <= 1'b0;
      \piso.data_r_1033_sv2v_reg  <= 1'b0;
      \piso.data_r_1032_sv2v_reg  <= 1'b0;
      \piso.data_r_1031_sv2v_reg  <= 1'b0;
      \piso.data_r_1030_sv2v_reg  <= 1'b0;
      \piso.data_r_1029_sv2v_reg  <= 1'b0;
      \piso.data_r_1028_sv2v_reg  <= 1'b0;
      \piso.data_r_1027_sv2v_reg  <= 1'b0;
      \piso.data_r_1026_sv2v_reg  <= 1'b0;
      \piso.data_r_1025_sv2v_reg  <= 1'b0;
      \piso.data_r_1024_sv2v_reg  <= 1'b0;
      \piso.data_r_1023_sv2v_reg  <= 1'b0;
      \piso.data_r_1022_sv2v_reg  <= 1'b0;
      \piso.data_r_1021_sv2v_reg  <= 1'b0;
      \piso.data_r_1020_sv2v_reg  <= 1'b0;
      \piso.data_r_1019_sv2v_reg  <= 1'b0;
      \piso.data_r_1018_sv2v_reg  <= 1'b0;
      \piso.data_r_1017_sv2v_reg  <= 1'b0;
      \piso.data_r_1016_sv2v_reg  <= 1'b0;
      \piso.data_r_1015_sv2v_reg  <= 1'b0;
      \piso.data_r_1014_sv2v_reg  <= 1'b0;
      \piso.data_r_1013_sv2v_reg  <= 1'b0;
      \piso.data_r_1012_sv2v_reg  <= 1'b0;
      \piso.data_r_1011_sv2v_reg  <= 1'b0;
      \piso.data_r_1010_sv2v_reg  <= 1'b0;
      \piso.data_r_1009_sv2v_reg  <= 1'b0;
      \piso.data_r_1008_sv2v_reg  <= 1'b0;
      \piso.data_r_1007_sv2v_reg  <= 1'b0;
      \piso.data_r_1006_sv2v_reg  <= 1'b0;
      \piso.data_r_1005_sv2v_reg  <= 1'b0;
      \piso.data_r_1004_sv2v_reg  <= 1'b0;
      \piso.data_r_1003_sv2v_reg  <= 1'b0;
      \piso.data_r_1002_sv2v_reg  <= 1'b0;
      \piso.data_r_1001_sv2v_reg  <= 1'b0;
      \piso.data_r_1000_sv2v_reg  <= 1'b0;
      \piso.data_r_999_sv2v_reg  <= 1'b0;
      \piso.data_r_998_sv2v_reg  <= 1'b0;
      \piso.data_r_997_sv2v_reg  <= 1'b0;
      \piso.data_r_996_sv2v_reg  <= 1'b0;
      \piso.data_r_995_sv2v_reg  <= 1'b0;
      \piso.data_r_994_sv2v_reg  <= 1'b0;
      \piso.data_r_993_sv2v_reg  <= 1'b0;
      \piso.data_r_992_sv2v_reg  <= 1'b0;
      \piso.data_r_991_sv2v_reg  <= 1'b0;
      \piso.data_r_990_sv2v_reg  <= 1'b0;
      \piso.data_r_989_sv2v_reg  <= 1'b0;
      \piso.data_r_988_sv2v_reg  <= 1'b0;
      \piso.data_r_987_sv2v_reg  <= 1'b0;
      \piso.data_r_986_sv2v_reg  <= 1'b0;
      \piso.data_r_985_sv2v_reg  <= 1'b0;
      \piso.data_r_984_sv2v_reg  <= 1'b0;
      \piso.data_r_983_sv2v_reg  <= 1'b0;
      \piso.data_r_982_sv2v_reg  <= 1'b0;
      \piso.data_r_981_sv2v_reg  <= 1'b0;
      \piso.data_r_980_sv2v_reg  <= 1'b0;
      \piso.data_r_979_sv2v_reg  <= 1'b0;
      \piso.data_r_978_sv2v_reg  <= 1'b0;
      \piso.data_r_977_sv2v_reg  <= 1'b0;
      \piso.data_r_976_sv2v_reg  <= 1'b0;
      \piso.data_r_975_sv2v_reg  <= 1'b0;
      \piso.data_r_974_sv2v_reg  <= 1'b0;
      \piso.data_r_973_sv2v_reg  <= 1'b0;
      \piso.data_r_972_sv2v_reg  <= 1'b0;
      \piso.data_r_971_sv2v_reg  <= 1'b0;
      \piso.data_r_970_sv2v_reg  <= 1'b0;
      \piso.data_r_969_sv2v_reg  <= 1'b0;
      \piso.data_r_968_sv2v_reg  <= 1'b0;
      \piso.data_r_967_sv2v_reg  <= 1'b0;
      \piso.data_r_966_sv2v_reg  <= 1'b0;
      \piso.data_r_965_sv2v_reg  <= 1'b0;
      \piso.data_r_964_sv2v_reg  <= 1'b0;
      \piso.data_r_963_sv2v_reg  <= 1'b0;
      \piso.data_r_962_sv2v_reg  <= 1'b0;
      \piso.data_r_961_sv2v_reg  <= 1'b0;
      \piso.data_r_960_sv2v_reg  <= 1'b0;
      \piso.data_r_959_sv2v_reg  <= 1'b0;
      \piso.data_r_958_sv2v_reg  <= 1'b0;
      \piso.data_r_957_sv2v_reg  <= 1'b0;
      \piso.data_r_956_sv2v_reg  <= 1'b0;
      \piso.data_r_955_sv2v_reg  <= 1'b0;
      \piso.data_r_954_sv2v_reg  <= 1'b0;
      \piso.data_r_953_sv2v_reg  <= 1'b0;
      \piso.data_r_952_sv2v_reg  <= 1'b0;
      \piso.data_r_951_sv2v_reg  <= 1'b0;
      \piso.data_r_950_sv2v_reg  <= 1'b0;
      \piso.data_r_949_sv2v_reg  <= 1'b0;
      \piso.data_r_948_sv2v_reg  <= 1'b0;
      \piso.data_r_947_sv2v_reg  <= 1'b0;
      \piso.data_r_946_sv2v_reg  <= 1'b0;
      \piso.data_r_945_sv2v_reg  <= 1'b0;
      \piso.data_r_944_sv2v_reg  <= 1'b0;
      \piso.data_r_943_sv2v_reg  <= 1'b0;
      \piso.data_r_942_sv2v_reg  <= 1'b0;
      \piso.data_r_941_sv2v_reg  <= 1'b0;
      \piso.data_r_940_sv2v_reg  <= 1'b0;
      \piso.data_r_939_sv2v_reg  <= 1'b0;
      \piso.data_r_938_sv2v_reg  <= 1'b0;
      \piso.data_r_937_sv2v_reg  <= 1'b0;
      \piso.data_r_936_sv2v_reg  <= 1'b0;
      \piso.data_r_935_sv2v_reg  <= 1'b0;
      \piso.data_r_934_sv2v_reg  <= 1'b0;
      \piso.data_r_933_sv2v_reg  <= 1'b0;
      \piso.data_r_932_sv2v_reg  <= 1'b0;
      \piso.data_r_931_sv2v_reg  <= 1'b0;
      \piso.data_r_930_sv2v_reg  <= 1'b0;
      \piso.data_r_929_sv2v_reg  <= 1'b0;
      \piso.data_r_928_sv2v_reg  <= 1'b0;
      \piso.data_r_927_sv2v_reg  <= 1'b0;
      \piso.data_r_926_sv2v_reg  <= 1'b0;
      \piso.data_r_925_sv2v_reg  <= 1'b0;
      \piso.data_r_924_sv2v_reg  <= 1'b0;
      \piso.data_r_923_sv2v_reg  <= 1'b0;
      \piso.data_r_922_sv2v_reg  <= 1'b0;
      \piso.data_r_921_sv2v_reg  <= 1'b0;
      \piso.data_r_920_sv2v_reg  <= 1'b0;
      \piso.data_r_919_sv2v_reg  <= 1'b0;
      \piso.data_r_918_sv2v_reg  <= 1'b0;
      \piso.data_r_917_sv2v_reg  <= 1'b0;
      \piso.data_r_916_sv2v_reg  <= 1'b0;
      \piso.data_r_915_sv2v_reg  <= 1'b0;
      \piso.data_r_914_sv2v_reg  <= 1'b0;
      \piso.data_r_913_sv2v_reg  <= 1'b0;
      \piso.data_r_912_sv2v_reg  <= 1'b0;
      \piso.data_r_911_sv2v_reg  <= 1'b0;
      \piso.data_r_910_sv2v_reg  <= 1'b0;
      \piso.data_r_909_sv2v_reg  <= 1'b0;
      \piso.data_r_908_sv2v_reg  <= 1'b0;
      \piso.data_r_907_sv2v_reg  <= 1'b0;
      \piso.data_r_906_sv2v_reg  <= 1'b0;
      \piso.data_r_905_sv2v_reg  <= 1'b0;
      \piso.data_r_904_sv2v_reg  <= 1'b0;
      \piso.data_r_903_sv2v_reg  <= 1'b0;
      \piso.data_r_902_sv2v_reg  <= 1'b0;
      \piso.data_r_901_sv2v_reg  <= 1'b0;
      \piso.data_r_900_sv2v_reg  <= 1'b0;
      \piso.data_r_899_sv2v_reg  <= 1'b0;
      \piso.data_r_898_sv2v_reg  <= 1'b0;
      \piso.data_r_897_sv2v_reg  <= 1'b0;
      \piso.data_r_896_sv2v_reg  <= 1'b0;
      \piso.data_r_895_sv2v_reg  <= 1'b0;
      \piso.data_r_894_sv2v_reg  <= 1'b0;
      \piso.data_r_893_sv2v_reg  <= 1'b0;
      \piso.data_r_892_sv2v_reg  <= 1'b0;
      \piso.data_r_891_sv2v_reg  <= 1'b0;
      \piso.data_r_890_sv2v_reg  <= 1'b0;
      \piso.data_r_889_sv2v_reg  <= 1'b0;
      \piso.data_r_888_sv2v_reg  <= 1'b0;
      \piso.data_r_887_sv2v_reg  <= 1'b0;
      \piso.data_r_886_sv2v_reg  <= 1'b0;
      \piso.data_r_885_sv2v_reg  <= 1'b0;
      \piso.data_r_884_sv2v_reg  <= 1'b0;
      \piso.data_r_883_sv2v_reg  <= 1'b0;
      \piso.data_r_882_sv2v_reg  <= 1'b0;
      \piso.data_r_881_sv2v_reg  <= 1'b0;
      \piso.data_r_880_sv2v_reg  <= 1'b0;
      \piso.data_r_879_sv2v_reg  <= 1'b0;
      \piso.data_r_878_sv2v_reg  <= 1'b0;
      \piso.data_r_877_sv2v_reg  <= 1'b0;
      \piso.data_r_876_sv2v_reg  <= 1'b0;
      \piso.data_r_875_sv2v_reg  <= 1'b0;
      \piso.data_r_874_sv2v_reg  <= 1'b0;
      \piso.data_r_873_sv2v_reg  <= 1'b0;
      \piso.data_r_872_sv2v_reg  <= 1'b0;
      \piso.data_r_871_sv2v_reg  <= 1'b0;
      \piso.data_r_870_sv2v_reg  <= 1'b0;
      \piso.data_r_869_sv2v_reg  <= 1'b0;
      \piso.data_r_868_sv2v_reg  <= 1'b0;
      \piso.data_r_867_sv2v_reg  <= 1'b0;
      \piso.data_r_866_sv2v_reg  <= 1'b0;
      \piso.data_r_865_sv2v_reg  <= 1'b0;
      \piso.data_r_864_sv2v_reg  <= 1'b0;
      \piso.data_r_863_sv2v_reg  <= 1'b0;
      \piso.data_r_862_sv2v_reg  <= 1'b0;
      \piso.data_r_861_sv2v_reg  <= 1'b0;
      \piso.data_r_860_sv2v_reg  <= 1'b0;
      \piso.data_r_859_sv2v_reg  <= 1'b0;
      \piso.data_r_858_sv2v_reg  <= 1'b0;
      \piso.data_r_857_sv2v_reg  <= 1'b0;
      \piso.data_r_856_sv2v_reg  <= 1'b0;
      \piso.data_r_855_sv2v_reg  <= 1'b0;
      \piso.data_r_854_sv2v_reg  <= 1'b0;
      \piso.data_r_853_sv2v_reg  <= 1'b0;
      \piso.data_r_852_sv2v_reg  <= 1'b0;
      \piso.data_r_851_sv2v_reg  <= 1'b0;
      \piso.data_r_850_sv2v_reg  <= 1'b0;
      \piso.data_r_849_sv2v_reg  <= 1'b0;
      \piso.data_r_848_sv2v_reg  <= 1'b0;
      \piso.data_r_847_sv2v_reg  <= 1'b0;
      \piso.data_r_846_sv2v_reg  <= 1'b0;
      \piso.data_r_845_sv2v_reg  <= 1'b0;
      \piso.data_r_844_sv2v_reg  <= 1'b0;
      \piso.data_r_843_sv2v_reg  <= 1'b0;
      \piso.data_r_842_sv2v_reg  <= 1'b0;
      \piso.data_r_841_sv2v_reg  <= 1'b0;
      \piso.data_r_840_sv2v_reg  <= 1'b0;
      \piso.data_r_839_sv2v_reg  <= 1'b0;
      \piso.data_r_838_sv2v_reg  <= 1'b0;
      \piso.data_r_837_sv2v_reg  <= 1'b0;
      \piso.data_r_836_sv2v_reg  <= 1'b0;
      \piso.data_r_835_sv2v_reg  <= 1'b0;
      \piso.data_r_834_sv2v_reg  <= 1'b0;
      \piso.data_r_833_sv2v_reg  <= 1'b0;
      \piso.data_r_832_sv2v_reg  <= 1'b0;
      \piso.data_r_831_sv2v_reg  <= 1'b0;
      \piso.data_r_830_sv2v_reg  <= 1'b0;
      \piso.data_r_829_sv2v_reg  <= 1'b0;
      \piso.data_r_828_sv2v_reg  <= 1'b0;
      \piso.data_r_827_sv2v_reg  <= 1'b0;
      \piso.data_r_826_sv2v_reg  <= 1'b0;
      \piso.data_r_825_sv2v_reg  <= 1'b0;
      \piso.data_r_824_sv2v_reg  <= 1'b0;
      \piso.data_r_823_sv2v_reg  <= 1'b0;
      \piso.data_r_822_sv2v_reg  <= 1'b0;
      \piso.data_r_821_sv2v_reg  <= 1'b0;
      \piso.data_r_820_sv2v_reg  <= 1'b0;
      \piso.data_r_819_sv2v_reg  <= 1'b0;
      \piso.data_r_818_sv2v_reg  <= 1'b0;
      \piso.data_r_817_sv2v_reg  <= 1'b0;
      \piso.data_r_816_sv2v_reg  <= 1'b0;
      \piso.data_r_815_sv2v_reg  <= 1'b0;
      \piso.data_r_814_sv2v_reg  <= 1'b0;
      \piso.data_r_813_sv2v_reg  <= 1'b0;
      \piso.data_r_812_sv2v_reg  <= 1'b0;
      \piso.data_r_811_sv2v_reg  <= 1'b0;
      \piso.data_r_810_sv2v_reg  <= 1'b0;
      \piso.data_r_809_sv2v_reg  <= 1'b0;
      \piso.data_r_808_sv2v_reg  <= 1'b0;
      \piso.data_r_807_sv2v_reg  <= 1'b0;
      \piso.data_r_806_sv2v_reg  <= 1'b0;
      \piso.data_r_805_sv2v_reg  <= 1'b0;
      \piso.data_r_804_sv2v_reg  <= 1'b0;
      \piso.data_r_803_sv2v_reg  <= 1'b0;
      \piso.data_r_802_sv2v_reg  <= 1'b0;
      \piso.data_r_801_sv2v_reg  <= 1'b0;
      \piso.data_r_800_sv2v_reg  <= 1'b0;
      \piso.data_r_799_sv2v_reg  <= 1'b0;
      \piso.data_r_798_sv2v_reg  <= 1'b0;
      \piso.data_r_797_sv2v_reg  <= 1'b0;
      \piso.data_r_796_sv2v_reg  <= 1'b0;
      \piso.data_r_795_sv2v_reg  <= 1'b0;
      \piso.data_r_794_sv2v_reg  <= 1'b0;
      \piso.data_r_793_sv2v_reg  <= 1'b0;
      \piso.data_r_792_sv2v_reg  <= 1'b0;
      \piso.data_r_791_sv2v_reg  <= 1'b0;
      \piso.data_r_790_sv2v_reg  <= 1'b0;
      \piso.data_r_789_sv2v_reg  <= 1'b0;
      \piso.data_r_788_sv2v_reg  <= 1'b0;
      \piso.data_r_787_sv2v_reg  <= 1'b0;
      \piso.data_r_786_sv2v_reg  <= 1'b0;
      \piso.data_r_785_sv2v_reg  <= 1'b0;
      \piso.data_r_784_sv2v_reg  <= 1'b0;
      \piso.data_r_783_sv2v_reg  <= 1'b0;
      \piso.data_r_782_sv2v_reg  <= 1'b0;
      \piso.data_r_781_sv2v_reg  <= 1'b0;
      \piso.data_r_780_sv2v_reg  <= 1'b0;
      \piso.data_r_779_sv2v_reg  <= 1'b0;
      \piso.data_r_778_sv2v_reg  <= 1'b0;
      \piso.data_r_777_sv2v_reg  <= 1'b0;
      \piso.data_r_776_sv2v_reg  <= 1'b0;
      \piso.data_r_775_sv2v_reg  <= 1'b0;
      \piso.data_r_774_sv2v_reg  <= 1'b0;
      \piso.data_r_773_sv2v_reg  <= 1'b0;
      \piso.data_r_772_sv2v_reg  <= 1'b0;
      \piso.data_r_771_sv2v_reg  <= 1'b0;
      \piso.data_r_770_sv2v_reg  <= 1'b0;
      \piso.data_r_769_sv2v_reg  <= 1'b0;
      \piso.data_r_768_sv2v_reg  <= 1'b0;
      \piso.data_r_767_sv2v_reg  <= 1'b0;
      \piso.data_r_766_sv2v_reg  <= 1'b0;
      \piso.data_r_765_sv2v_reg  <= 1'b0;
      \piso.data_r_764_sv2v_reg  <= 1'b0;
      \piso.data_r_763_sv2v_reg  <= 1'b0;
      \piso.data_r_762_sv2v_reg  <= 1'b0;
      \piso.data_r_761_sv2v_reg  <= 1'b0;
      \piso.data_r_760_sv2v_reg  <= 1'b0;
      \piso.data_r_759_sv2v_reg  <= 1'b0;
      \piso.data_r_758_sv2v_reg  <= 1'b0;
      \piso.data_r_757_sv2v_reg  <= 1'b0;
      \piso.data_r_756_sv2v_reg  <= 1'b0;
      \piso.data_r_755_sv2v_reg  <= 1'b0;
      \piso.data_r_754_sv2v_reg  <= 1'b0;
      \piso.data_r_753_sv2v_reg  <= 1'b0;
      \piso.data_r_752_sv2v_reg  <= 1'b0;
      \piso.data_r_751_sv2v_reg  <= 1'b0;
      \piso.data_r_750_sv2v_reg  <= 1'b0;
      \piso.data_r_749_sv2v_reg  <= 1'b0;
      \piso.data_r_748_sv2v_reg  <= 1'b0;
      \piso.data_r_747_sv2v_reg  <= 1'b0;
      \piso.data_r_746_sv2v_reg  <= 1'b0;
      \piso.data_r_745_sv2v_reg  <= 1'b0;
      \piso.data_r_744_sv2v_reg  <= 1'b0;
      \piso.data_r_743_sv2v_reg  <= 1'b0;
      \piso.data_r_742_sv2v_reg  <= 1'b0;
      \piso.data_r_741_sv2v_reg  <= 1'b0;
      \piso.data_r_740_sv2v_reg  <= 1'b0;
      \piso.data_r_739_sv2v_reg  <= 1'b0;
      \piso.data_r_738_sv2v_reg  <= 1'b0;
      \piso.data_r_737_sv2v_reg  <= 1'b0;
      \piso.data_r_736_sv2v_reg  <= 1'b0;
      \piso.data_r_735_sv2v_reg  <= 1'b0;
      \piso.data_r_734_sv2v_reg  <= 1'b0;
      \piso.data_r_733_sv2v_reg  <= 1'b0;
      \piso.data_r_732_sv2v_reg  <= 1'b0;
      \piso.data_r_731_sv2v_reg  <= 1'b0;
      \piso.data_r_730_sv2v_reg  <= 1'b0;
      \piso.data_r_729_sv2v_reg  <= 1'b0;
      \piso.data_r_728_sv2v_reg  <= 1'b0;
      \piso.data_r_727_sv2v_reg  <= 1'b0;
      \piso.data_r_726_sv2v_reg  <= 1'b0;
      \piso.data_r_725_sv2v_reg  <= 1'b0;
      \piso.data_r_724_sv2v_reg  <= 1'b0;
      \piso.data_r_723_sv2v_reg  <= 1'b0;
      \piso.data_r_722_sv2v_reg  <= 1'b0;
      \piso.data_r_721_sv2v_reg  <= 1'b0;
      \piso.data_r_720_sv2v_reg  <= 1'b0;
      \piso.data_r_719_sv2v_reg  <= 1'b0;
      \piso.data_r_718_sv2v_reg  <= 1'b0;
      \piso.data_r_717_sv2v_reg  <= 1'b0;
      \piso.data_r_716_sv2v_reg  <= 1'b0;
      \piso.data_r_715_sv2v_reg  <= 1'b0;
      \piso.data_r_714_sv2v_reg  <= 1'b0;
      \piso.data_r_713_sv2v_reg  <= 1'b0;
      \piso.data_r_712_sv2v_reg  <= 1'b0;
      \piso.data_r_711_sv2v_reg  <= 1'b0;
      \piso.data_r_710_sv2v_reg  <= 1'b0;
      \piso.data_r_709_sv2v_reg  <= 1'b0;
      \piso.data_r_708_sv2v_reg  <= 1'b0;
      \piso.data_r_707_sv2v_reg  <= 1'b0;
      \piso.data_r_706_sv2v_reg  <= 1'b0;
      \piso.data_r_705_sv2v_reg  <= 1'b0;
      \piso.data_r_704_sv2v_reg  <= 1'b0;
      \piso.data_r_703_sv2v_reg  <= 1'b0;
      \piso.data_r_702_sv2v_reg  <= 1'b0;
      \piso.data_r_701_sv2v_reg  <= 1'b0;
      \piso.data_r_700_sv2v_reg  <= 1'b0;
      \piso.data_r_699_sv2v_reg  <= 1'b0;
      \piso.data_r_698_sv2v_reg  <= 1'b0;
      \piso.data_r_697_sv2v_reg  <= 1'b0;
      \piso.data_r_696_sv2v_reg  <= 1'b0;
      \piso.data_r_695_sv2v_reg  <= 1'b0;
      \piso.data_r_694_sv2v_reg  <= 1'b0;
      \piso.data_r_693_sv2v_reg  <= 1'b0;
      \piso.data_r_692_sv2v_reg  <= 1'b0;
      \piso.data_r_691_sv2v_reg  <= 1'b0;
      \piso.data_r_690_sv2v_reg  <= 1'b0;
      \piso.data_r_689_sv2v_reg  <= 1'b0;
      \piso.data_r_688_sv2v_reg  <= 1'b0;
      \piso.data_r_687_sv2v_reg  <= 1'b0;
      \piso.data_r_686_sv2v_reg  <= 1'b0;
      \piso.data_r_685_sv2v_reg  <= 1'b0;
      \piso.data_r_684_sv2v_reg  <= 1'b0;
      \piso.data_r_683_sv2v_reg  <= 1'b0;
      \piso.data_r_682_sv2v_reg  <= 1'b0;
      \piso.data_r_681_sv2v_reg  <= 1'b0;
      \piso.data_r_680_sv2v_reg  <= 1'b0;
      \piso.data_r_679_sv2v_reg  <= 1'b0;
      \piso.data_r_678_sv2v_reg  <= 1'b0;
      \piso.data_r_677_sv2v_reg  <= 1'b0;
      \piso.data_r_676_sv2v_reg  <= 1'b0;
      \piso.data_r_675_sv2v_reg  <= 1'b0;
      \piso.data_r_674_sv2v_reg  <= 1'b0;
      \piso.data_r_673_sv2v_reg  <= 1'b0;
      \piso.data_r_672_sv2v_reg  <= 1'b0;
      \piso.data_r_671_sv2v_reg  <= 1'b0;
      \piso.data_r_670_sv2v_reg  <= 1'b0;
      \piso.data_r_669_sv2v_reg  <= 1'b0;
      \piso.data_r_668_sv2v_reg  <= 1'b0;
      \piso.data_r_667_sv2v_reg  <= 1'b0;
      \piso.data_r_666_sv2v_reg  <= 1'b0;
      \piso.data_r_665_sv2v_reg  <= 1'b0;
      \piso.data_r_664_sv2v_reg  <= 1'b0;
      \piso.data_r_663_sv2v_reg  <= 1'b0;
      \piso.data_r_662_sv2v_reg  <= 1'b0;
      \piso.data_r_661_sv2v_reg  <= 1'b0;
      \piso.data_r_660_sv2v_reg  <= 1'b0;
      \piso.data_r_659_sv2v_reg  <= 1'b0;
      \piso.data_r_658_sv2v_reg  <= 1'b0;
      \piso.data_r_657_sv2v_reg  <= 1'b0;
      \piso.data_r_656_sv2v_reg  <= 1'b0;
      \piso.data_r_655_sv2v_reg  <= 1'b0;
      \piso.data_r_654_sv2v_reg  <= 1'b0;
      \piso.data_r_653_sv2v_reg  <= 1'b0;
      \piso.data_r_652_sv2v_reg  <= 1'b0;
      \piso.data_r_651_sv2v_reg  <= 1'b0;
      \piso.data_r_650_sv2v_reg  <= 1'b0;
      \piso.data_r_649_sv2v_reg  <= 1'b0;
      \piso.data_r_648_sv2v_reg  <= 1'b0;
      \piso.data_r_647_sv2v_reg  <= 1'b0;
      \piso.data_r_646_sv2v_reg  <= 1'b0;
      \piso.data_r_645_sv2v_reg  <= 1'b0;
      \piso.data_r_644_sv2v_reg  <= 1'b0;
      \piso.data_r_643_sv2v_reg  <= 1'b0;
      \piso.data_r_642_sv2v_reg  <= 1'b0;
      \piso.data_r_641_sv2v_reg  <= 1'b0;
      \piso.data_r_640_sv2v_reg  <= 1'b0;
      \piso.data_r_639_sv2v_reg  <= 1'b0;
      \piso.data_r_638_sv2v_reg  <= 1'b0;
      \piso.data_r_637_sv2v_reg  <= 1'b0;
      \piso.data_r_636_sv2v_reg  <= 1'b0;
      \piso.data_r_635_sv2v_reg  <= 1'b0;
      \piso.data_r_634_sv2v_reg  <= 1'b0;
      \piso.data_r_633_sv2v_reg  <= 1'b0;
      \piso.data_r_632_sv2v_reg  <= 1'b0;
      \piso.data_r_631_sv2v_reg  <= 1'b0;
      \piso.data_r_630_sv2v_reg  <= 1'b0;
      \piso.data_r_629_sv2v_reg  <= 1'b0;
      \piso.data_r_628_sv2v_reg  <= 1'b0;
      \piso.data_r_627_sv2v_reg  <= 1'b0;
      \piso.data_r_626_sv2v_reg  <= 1'b0;
      \piso.data_r_625_sv2v_reg  <= 1'b0;
      \piso.data_r_624_sv2v_reg  <= 1'b0;
      \piso.data_r_623_sv2v_reg  <= 1'b0;
      \piso.data_r_622_sv2v_reg  <= 1'b0;
      \piso.data_r_621_sv2v_reg  <= 1'b0;
      \piso.data_r_620_sv2v_reg  <= 1'b0;
      \piso.data_r_619_sv2v_reg  <= 1'b0;
      \piso.data_r_618_sv2v_reg  <= 1'b0;
      \piso.data_r_617_sv2v_reg  <= 1'b0;
      \piso.data_r_616_sv2v_reg  <= 1'b0;
      \piso.data_r_615_sv2v_reg  <= 1'b0;
      \piso.data_r_614_sv2v_reg  <= 1'b0;
      \piso.data_r_613_sv2v_reg  <= 1'b0;
      \piso.data_r_612_sv2v_reg  <= 1'b0;
      \piso.data_r_611_sv2v_reg  <= 1'b0;
      \piso.data_r_610_sv2v_reg  <= 1'b0;
      \piso.data_r_609_sv2v_reg  <= 1'b0;
      \piso.data_r_608_sv2v_reg  <= 1'b0;
      \piso.data_r_607_sv2v_reg  <= 1'b0;
      \piso.data_r_606_sv2v_reg  <= 1'b0;
      \piso.data_r_605_sv2v_reg  <= 1'b0;
      \piso.data_r_604_sv2v_reg  <= 1'b0;
      \piso.data_r_603_sv2v_reg  <= 1'b0;
      \piso.data_r_602_sv2v_reg  <= 1'b0;
      \piso.data_r_601_sv2v_reg  <= 1'b0;
      \piso.data_r_600_sv2v_reg  <= 1'b0;
      \piso.data_r_599_sv2v_reg  <= 1'b0;
      \piso.data_r_598_sv2v_reg  <= 1'b0;
      \piso.data_r_597_sv2v_reg  <= 1'b0;
      \piso.data_r_596_sv2v_reg  <= 1'b0;
      \piso.data_r_595_sv2v_reg  <= 1'b0;
      \piso.data_r_594_sv2v_reg  <= 1'b0;
      \piso.data_r_593_sv2v_reg  <= 1'b0;
      \piso.data_r_592_sv2v_reg  <= 1'b0;
      \piso.data_r_591_sv2v_reg  <= 1'b0;
      \piso.data_r_590_sv2v_reg  <= 1'b0;
      \piso.data_r_589_sv2v_reg  <= 1'b0;
      \piso.data_r_588_sv2v_reg  <= 1'b0;
      \piso.data_r_587_sv2v_reg  <= 1'b0;
      \piso.data_r_586_sv2v_reg  <= 1'b0;
      \piso.data_r_585_sv2v_reg  <= 1'b0;
      \piso.data_r_584_sv2v_reg  <= 1'b0;
      \piso.data_r_583_sv2v_reg  <= 1'b0;
      \piso.data_r_582_sv2v_reg  <= 1'b0;
      \piso.data_r_581_sv2v_reg  <= 1'b0;
      \piso.data_r_580_sv2v_reg  <= 1'b0;
      \piso.data_r_579_sv2v_reg  <= 1'b0;
      \piso.data_r_578_sv2v_reg  <= 1'b0;
      \piso.data_r_577_sv2v_reg  <= 1'b0;
      \piso.data_r_576_sv2v_reg  <= 1'b0;
      \piso.data_r_575_sv2v_reg  <= 1'b0;
      \piso.data_r_574_sv2v_reg  <= 1'b0;
      \piso.data_r_573_sv2v_reg  <= 1'b0;
      \piso.data_r_572_sv2v_reg  <= 1'b0;
      \piso.data_r_571_sv2v_reg  <= 1'b0;
      \piso.data_r_570_sv2v_reg  <= 1'b0;
      \piso.data_r_569_sv2v_reg  <= 1'b0;
      \piso.data_r_568_sv2v_reg  <= 1'b0;
      \piso.data_r_567_sv2v_reg  <= 1'b0;
      \piso.data_r_566_sv2v_reg  <= 1'b0;
      \piso.data_r_565_sv2v_reg  <= 1'b0;
      \piso.data_r_564_sv2v_reg  <= 1'b0;
      \piso.data_r_563_sv2v_reg  <= 1'b0;
      \piso.data_r_562_sv2v_reg  <= 1'b0;
      \piso.data_r_561_sv2v_reg  <= 1'b0;
      \piso.data_r_560_sv2v_reg  <= 1'b0;
      \piso.data_r_559_sv2v_reg  <= 1'b0;
      \piso.data_r_558_sv2v_reg  <= 1'b0;
      \piso.data_r_557_sv2v_reg  <= 1'b0;
      \piso.data_r_556_sv2v_reg  <= 1'b0;
      \piso.data_r_555_sv2v_reg  <= 1'b0;
      \piso.data_r_554_sv2v_reg  <= 1'b0;
      \piso.data_r_553_sv2v_reg  <= 1'b0;
      \piso.data_r_552_sv2v_reg  <= 1'b0;
      \piso.data_r_551_sv2v_reg  <= 1'b0;
      \piso.data_r_550_sv2v_reg  <= 1'b0;
      \piso.data_r_549_sv2v_reg  <= 1'b0;
      \piso.data_r_548_sv2v_reg  <= 1'b0;
      \piso.data_r_547_sv2v_reg  <= 1'b0;
      \piso.data_r_546_sv2v_reg  <= 1'b0;
      \piso.data_r_545_sv2v_reg  <= 1'b0;
      \piso.data_r_544_sv2v_reg  <= 1'b0;
      \piso.data_r_543_sv2v_reg  <= 1'b0;
      \piso.data_r_542_sv2v_reg  <= 1'b0;
      \piso.data_r_541_sv2v_reg  <= 1'b0;
      \piso.data_r_540_sv2v_reg  <= 1'b0;
      \piso.data_r_539_sv2v_reg  <= 1'b0;
      \piso.data_r_538_sv2v_reg  <= 1'b0;
      \piso.data_r_537_sv2v_reg  <= 1'b0;
      \piso.data_r_536_sv2v_reg  <= 1'b0;
      \piso.data_r_535_sv2v_reg  <= 1'b0;
      \piso.data_r_534_sv2v_reg  <= 1'b0;
      \piso.data_r_533_sv2v_reg  <= 1'b0;
      \piso.data_r_532_sv2v_reg  <= 1'b0;
      \piso.data_r_531_sv2v_reg  <= 1'b0;
      \piso.data_r_530_sv2v_reg  <= 1'b0;
      \piso.data_r_529_sv2v_reg  <= 1'b0;
      \piso.data_r_528_sv2v_reg  <= 1'b0;
      \piso.data_r_527_sv2v_reg  <= 1'b0;
      \piso.data_r_526_sv2v_reg  <= 1'b0;
      \piso.data_r_525_sv2v_reg  <= 1'b0;
      \piso.data_r_524_sv2v_reg  <= 1'b0;
      \piso.data_r_523_sv2v_reg  <= 1'b0;
      \piso.data_r_522_sv2v_reg  <= 1'b0;
      \piso.data_r_521_sv2v_reg  <= 1'b0;
      \piso.data_r_520_sv2v_reg  <= 1'b0;
      \piso.data_r_519_sv2v_reg  <= 1'b0;
      \piso.data_r_518_sv2v_reg  <= 1'b0;
      \piso.data_r_517_sv2v_reg  <= 1'b0;
      \piso.data_r_516_sv2v_reg  <= 1'b0;
      \piso.data_r_515_sv2v_reg  <= 1'b0;
      \piso.data_r_514_sv2v_reg  <= 1'b0;
      \piso.data_r_513_sv2v_reg  <= 1'b0;
      \piso.data_r_512_sv2v_reg  <= 1'b0;
      \piso.data_r_511_sv2v_reg  <= 1'b0;
      \piso.data_r_510_sv2v_reg  <= 1'b0;
      \piso.data_r_509_sv2v_reg  <= 1'b0;
      \piso.data_r_508_sv2v_reg  <= 1'b0;
      \piso.data_r_507_sv2v_reg  <= 1'b0;
      \piso.data_r_506_sv2v_reg  <= 1'b0;
      \piso.data_r_505_sv2v_reg  <= 1'b0;
      \piso.data_r_504_sv2v_reg  <= 1'b0;
      \piso.data_r_503_sv2v_reg  <= 1'b0;
      \piso.data_r_502_sv2v_reg  <= 1'b0;
      \piso.data_r_501_sv2v_reg  <= 1'b0;
      \piso.data_r_500_sv2v_reg  <= 1'b0;
      \piso.data_r_499_sv2v_reg  <= 1'b0;
      \piso.data_r_498_sv2v_reg  <= 1'b0;
      \piso.data_r_497_sv2v_reg  <= 1'b0;
      \piso.data_r_496_sv2v_reg  <= 1'b0;
      \piso.data_r_495_sv2v_reg  <= 1'b0;
      \piso.data_r_494_sv2v_reg  <= 1'b0;
      \piso.data_r_493_sv2v_reg  <= 1'b0;
      \piso.data_r_492_sv2v_reg  <= 1'b0;
      \piso.data_r_491_sv2v_reg  <= 1'b0;
      \piso.data_r_490_sv2v_reg  <= 1'b0;
      \piso.data_r_489_sv2v_reg  <= 1'b0;
      \piso.data_r_488_sv2v_reg  <= 1'b0;
      \piso.data_r_487_sv2v_reg  <= 1'b0;
      \piso.data_r_486_sv2v_reg  <= 1'b0;
      \piso.data_r_485_sv2v_reg  <= 1'b0;
      \piso.data_r_484_sv2v_reg  <= 1'b0;
      \piso.data_r_483_sv2v_reg  <= 1'b0;
      \piso.data_r_482_sv2v_reg  <= 1'b0;
      \piso.data_r_481_sv2v_reg  <= 1'b0;
      \piso.data_r_480_sv2v_reg  <= 1'b0;
      \piso.data_r_479_sv2v_reg  <= 1'b0;
      \piso.data_r_478_sv2v_reg  <= 1'b0;
      \piso.data_r_477_sv2v_reg  <= 1'b0;
      \piso.data_r_476_sv2v_reg  <= 1'b0;
      \piso.data_r_475_sv2v_reg  <= 1'b0;
      \piso.data_r_474_sv2v_reg  <= 1'b0;
      \piso.data_r_473_sv2v_reg  <= 1'b0;
      \piso.data_r_472_sv2v_reg  <= 1'b0;
      \piso.data_r_471_sv2v_reg  <= 1'b0;
      \piso.data_r_470_sv2v_reg  <= 1'b0;
      \piso.data_r_469_sv2v_reg  <= 1'b0;
      \piso.data_r_468_sv2v_reg  <= 1'b0;
      \piso.data_r_467_sv2v_reg  <= 1'b0;
      \piso.data_r_466_sv2v_reg  <= 1'b0;
      \piso.data_r_465_sv2v_reg  <= 1'b0;
      \piso.data_r_464_sv2v_reg  <= 1'b0;
      \piso.data_r_463_sv2v_reg  <= 1'b0;
      \piso.data_r_462_sv2v_reg  <= 1'b0;
      \piso.data_r_461_sv2v_reg  <= 1'b0;
      \piso.data_r_460_sv2v_reg  <= 1'b0;
      \piso.data_r_459_sv2v_reg  <= 1'b0;
      \piso.data_r_458_sv2v_reg  <= 1'b0;
      \piso.data_r_457_sv2v_reg  <= 1'b0;
      \piso.data_r_456_sv2v_reg  <= 1'b0;
      \piso.data_r_455_sv2v_reg  <= 1'b0;
      \piso.data_r_454_sv2v_reg  <= 1'b0;
      \piso.data_r_453_sv2v_reg  <= 1'b0;
      \piso.data_r_452_sv2v_reg  <= 1'b0;
      \piso.data_r_451_sv2v_reg  <= 1'b0;
      \piso.data_r_450_sv2v_reg  <= 1'b0;
      \piso.data_r_449_sv2v_reg  <= 1'b0;
      \piso.data_r_448_sv2v_reg  <= 1'b0;
      \piso.data_r_447_sv2v_reg  <= 1'b0;
      \piso.data_r_446_sv2v_reg  <= 1'b0;
      \piso.data_r_445_sv2v_reg  <= 1'b0;
      \piso.data_r_444_sv2v_reg  <= 1'b0;
      \piso.data_r_443_sv2v_reg  <= 1'b0;
      \piso.data_r_442_sv2v_reg  <= 1'b0;
      \piso.data_r_441_sv2v_reg  <= 1'b0;
      \piso.data_r_440_sv2v_reg  <= 1'b0;
      \piso.data_r_439_sv2v_reg  <= 1'b0;
      \piso.data_r_438_sv2v_reg  <= 1'b0;
      \piso.data_r_437_sv2v_reg  <= 1'b0;
      \piso.data_r_436_sv2v_reg  <= 1'b0;
      \piso.data_r_435_sv2v_reg  <= 1'b0;
      \piso.data_r_434_sv2v_reg  <= 1'b0;
      \piso.data_r_433_sv2v_reg  <= 1'b0;
      \piso.data_r_432_sv2v_reg  <= 1'b0;
      \piso.data_r_431_sv2v_reg  <= 1'b0;
      \piso.data_r_430_sv2v_reg  <= 1'b0;
      \piso.data_r_429_sv2v_reg  <= 1'b0;
      \piso.data_r_428_sv2v_reg  <= 1'b0;
      \piso.data_r_427_sv2v_reg  <= 1'b0;
      \piso.data_r_426_sv2v_reg  <= 1'b0;
      \piso.data_r_425_sv2v_reg  <= 1'b0;
      \piso.data_r_424_sv2v_reg  <= 1'b0;
      \piso.data_r_423_sv2v_reg  <= 1'b0;
      \piso.data_r_422_sv2v_reg  <= 1'b0;
      \piso.data_r_421_sv2v_reg  <= 1'b0;
      \piso.data_r_420_sv2v_reg  <= 1'b0;
      \piso.data_r_419_sv2v_reg  <= 1'b0;
      \piso.data_r_418_sv2v_reg  <= 1'b0;
      \piso.data_r_417_sv2v_reg  <= 1'b0;
      \piso.data_r_416_sv2v_reg  <= 1'b0;
      \piso.data_r_415_sv2v_reg  <= 1'b0;
      \piso.data_r_414_sv2v_reg  <= 1'b0;
      \piso.data_r_413_sv2v_reg  <= 1'b0;
      \piso.data_r_412_sv2v_reg  <= 1'b0;
      \piso.data_r_411_sv2v_reg  <= 1'b0;
      \piso.data_r_410_sv2v_reg  <= 1'b0;
      \piso.data_r_409_sv2v_reg  <= 1'b0;
      \piso.data_r_408_sv2v_reg  <= 1'b0;
      \piso.data_r_407_sv2v_reg  <= 1'b0;
      \piso.data_r_406_sv2v_reg  <= 1'b0;
      \piso.data_r_405_sv2v_reg  <= 1'b0;
      \piso.data_r_404_sv2v_reg  <= 1'b0;
      \piso.data_r_403_sv2v_reg  <= 1'b0;
      \piso.data_r_402_sv2v_reg  <= 1'b0;
      \piso.data_r_401_sv2v_reg  <= 1'b0;
      \piso.data_r_400_sv2v_reg  <= 1'b0;
      \piso.data_r_399_sv2v_reg  <= 1'b0;
      \piso.data_r_398_sv2v_reg  <= 1'b0;
      \piso.data_r_397_sv2v_reg  <= 1'b0;
      \piso.data_r_396_sv2v_reg  <= 1'b0;
      \piso.data_r_395_sv2v_reg  <= 1'b0;
      \piso.data_r_394_sv2v_reg  <= 1'b0;
      \piso.data_r_393_sv2v_reg  <= 1'b0;
      \piso.data_r_392_sv2v_reg  <= 1'b0;
      \piso.data_r_391_sv2v_reg  <= 1'b0;
      \piso.data_r_390_sv2v_reg  <= 1'b0;
      \piso.data_r_389_sv2v_reg  <= 1'b0;
      \piso.data_r_388_sv2v_reg  <= 1'b0;
      \piso.data_r_387_sv2v_reg  <= 1'b0;
      \piso.data_r_386_sv2v_reg  <= 1'b0;
      \piso.data_r_385_sv2v_reg  <= 1'b0;
      \piso.data_r_384_sv2v_reg  <= 1'b0;
      \piso.data_r_383_sv2v_reg  <= 1'b0;
      \piso.data_r_382_sv2v_reg  <= 1'b0;
      \piso.data_r_381_sv2v_reg  <= 1'b0;
      \piso.data_r_380_sv2v_reg  <= 1'b0;
      \piso.data_r_379_sv2v_reg  <= 1'b0;
      \piso.data_r_378_sv2v_reg  <= 1'b0;
      \piso.data_r_377_sv2v_reg  <= 1'b0;
      \piso.data_r_376_sv2v_reg  <= 1'b0;
      \piso.data_r_375_sv2v_reg  <= 1'b0;
      \piso.data_r_374_sv2v_reg  <= 1'b0;
      \piso.data_r_373_sv2v_reg  <= 1'b0;
      \piso.data_r_372_sv2v_reg  <= 1'b0;
      \piso.data_r_371_sv2v_reg  <= 1'b0;
      \piso.data_r_370_sv2v_reg  <= 1'b0;
      \piso.data_r_369_sv2v_reg  <= 1'b0;
      \piso.data_r_368_sv2v_reg  <= 1'b0;
      \piso.data_r_367_sv2v_reg  <= 1'b0;
      \piso.data_r_366_sv2v_reg  <= 1'b0;
      \piso.data_r_365_sv2v_reg  <= 1'b0;
      \piso.data_r_364_sv2v_reg  <= 1'b0;
      \piso.data_r_363_sv2v_reg  <= 1'b0;
      \piso.data_r_362_sv2v_reg  <= 1'b0;
      \piso.data_r_361_sv2v_reg  <= 1'b0;
      \piso.data_r_360_sv2v_reg  <= 1'b0;
      \piso.data_r_359_sv2v_reg  <= 1'b0;
      \piso.data_r_358_sv2v_reg  <= 1'b0;
      \piso.data_r_357_sv2v_reg  <= 1'b0;
      \piso.data_r_356_sv2v_reg  <= 1'b0;
      \piso.data_r_355_sv2v_reg  <= 1'b0;
      \piso.data_r_354_sv2v_reg  <= 1'b0;
      \piso.data_r_353_sv2v_reg  <= 1'b0;
      \piso.data_r_352_sv2v_reg  <= 1'b0;
      \piso.data_r_351_sv2v_reg  <= 1'b0;
      \piso.data_r_350_sv2v_reg  <= 1'b0;
      \piso.data_r_349_sv2v_reg  <= 1'b0;
      \piso.data_r_348_sv2v_reg  <= 1'b0;
      \piso.data_r_347_sv2v_reg  <= 1'b0;
      \piso.data_r_346_sv2v_reg  <= 1'b0;
      \piso.data_r_345_sv2v_reg  <= 1'b0;
      \piso.data_r_344_sv2v_reg  <= 1'b0;
      \piso.data_r_343_sv2v_reg  <= 1'b0;
      \piso.data_r_342_sv2v_reg  <= 1'b0;
      \piso.data_r_341_sv2v_reg  <= 1'b0;
      \piso.data_r_340_sv2v_reg  <= 1'b0;
      \piso.data_r_339_sv2v_reg  <= 1'b0;
      \piso.data_r_338_sv2v_reg  <= 1'b0;
      \piso.data_r_337_sv2v_reg  <= 1'b0;
      \piso.data_r_336_sv2v_reg  <= 1'b0;
      \piso.data_r_335_sv2v_reg  <= 1'b0;
      \piso.data_r_334_sv2v_reg  <= 1'b0;
      \piso.data_r_333_sv2v_reg  <= 1'b0;
      \piso.data_r_332_sv2v_reg  <= 1'b0;
      \piso.data_r_331_sv2v_reg  <= 1'b0;
      \piso.data_r_330_sv2v_reg  <= 1'b0;
      \piso.data_r_329_sv2v_reg  <= 1'b0;
      \piso.data_r_328_sv2v_reg  <= 1'b0;
      \piso.data_r_327_sv2v_reg  <= 1'b0;
      \piso.data_r_326_sv2v_reg  <= 1'b0;
      \piso.data_r_325_sv2v_reg  <= 1'b0;
      \piso.data_r_324_sv2v_reg  <= 1'b0;
      \piso.data_r_323_sv2v_reg  <= 1'b0;
      \piso.data_r_322_sv2v_reg  <= 1'b0;
      \piso.data_r_321_sv2v_reg  <= 1'b0;
      \piso.data_r_320_sv2v_reg  <= 1'b0;
      \piso.data_r_319_sv2v_reg  <= 1'b0;
      \piso.data_r_318_sv2v_reg  <= 1'b0;
      \piso.data_r_317_sv2v_reg  <= 1'b0;
      \piso.data_r_316_sv2v_reg  <= 1'b0;
      \piso.data_r_315_sv2v_reg  <= 1'b0;
      \piso.data_r_314_sv2v_reg  <= 1'b0;
      \piso.data_r_313_sv2v_reg  <= 1'b0;
      \piso.data_r_312_sv2v_reg  <= 1'b0;
      \piso.data_r_311_sv2v_reg  <= 1'b0;
      \piso.data_r_310_sv2v_reg  <= 1'b0;
      \piso.data_r_309_sv2v_reg  <= 1'b0;
      \piso.data_r_308_sv2v_reg  <= 1'b0;
      \piso.data_r_307_sv2v_reg  <= 1'b0;
      \piso.data_r_306_sv2v_reg  <= 1'b0;
      \piso.data_r_305_sv2v_reg  <= 1'b0;
      \piso.data_r_304_sv2v_reg  <= 1'b0;
      \piso.data_r_303_sv2v_reg  <= 1'b0;
      \piso.data_r_302_sv2v_reg  <= 1'b0;
      \piso.data_r_301_sv2v_reg  <= 1'b0;
      \piso.data_r_300_sv2v_reg  <= 1'b0;
      \piso.data_r_299_sv2v_reg  <= 1'b0;
      \piso.data_r_298_sv2v_reg  <= 1'b0;
      \piso.data_r_297_sv2v_reg  <= 1'b0;
      \piso.data_r_296_sv2v_reg  <= 1'b0;
      \piso.data_r_295_sv2v_reg  <= 1'b0;
      \piso.data_r_294_sv2v_reg  <= 1'b0;
      \piso.data_r_293_sv2v_reg  <= 1'b0;
      \piso.data_r_292_sv2v_reg  <= 1'b0;
      \piso.data_r_291_sv2v_reg  <= 1'b0;
      \piso.data_r_290_sv2v_reg  <= 1'b0;
      \piso.data_r_289_sv2v_reg  <= 1'b0;
      \piso.data_r_288_sv2v_reg  <= 1'b0;
      \piso.data_r_287_sv2v_reg  <= 1'b0;
      \piso.data_r_286_sv2v_reg  <= 1'b0;
      \piso.data_r_285_sv2v_reg  <= 1'b0;
      \piso.data_r_284_sv2v_reg  <= 1'b0;
      \piso.data_r_283_sv2v_reg  <= 1'b0;
      \piso.data_r_282_sv2v_reg  <= 1'b0;
      \piso.data_r_281_sv2v_reg  <= 1'b0;
      \piso.data_r_280_sv2v_reg  <= 1'b0;
      \piso.data_r_279_sv2v_reg  <= 1'b0;
      \piso.data_r_278_sv2v_reg  <= 1'b0;
      \piso.data_r_277_sv2v_reg  <= 1'b0;
      \piso.data_r_276_sv2v_reg  <= 1'b0;
      \piso.data_r_275_sv2v_reg  <= 1'b0;
      \piso.data_r_274_sv2v_reg  <= 1'b0;
      \piso.data_r_273_sv2v_reg  <= 1'b0;
      \piso.data_r_272_sv2v_reg  <= 1'b0;
      \piso.data_r_271_sv2v_reg  <= 1'b0;
      \piso.data_r_270_sv2v_reg  <= 1'b0;
      \piso.data_r_269_sv2v_reg  <= 1'b0;
      \piso.data_r_268_sv2v_reg  <= 1'b0;
      \piso.data_r_267_sv2v_reg  <= 1'b0;
      \piso.data_r_266_sv2v_reg  <= 1'b0;
      \piso.data_r_265_sv2v_reg  <= 1'b0;
      \piso.data_r_264_sv2v_reg  <= 1'b0;
      \piso.data_r_263_sv2v_reg  <= 1'b0;
      \piso.data_r_262_sv2v_reg  <= 1'b0;
      \piso.data_r_261_sv2v_reg  <= 1'b0;
      \piso.data_r_260_sv2v_reg  <= 1'b0;
      \piso.data_r_259_sv2v_reg  <= 1'b0;
      \piso.data_r_258_sv2v_reg  <= 1'b0;
      \piso.data_r_257_sv2v_reg  <= 1'b0;
      \piso.data_r_256_sv2v_reg  <= 1'b0;
      \piso.data_r_255_sv2v_reg  <= 1'b0;
      \piso.data_r_254_sv2v_reg  <= 1'b0;
      \piso.data_r_253_sv2v_reg  <= 1'b0;
      \piso.data_r_252_sv2v_reg  <= 1'b0;
      \piso.data_r_251_sv2v_reg  <= 1'b0;
      \piso.data_r_250_sv2v_reg  <= 1'b0;
      \piso.data_r_249_sv2v_reg  <= 1'b0;
      \piso.data_r_248_sv2v_reg  <= 1'b0;
      \piso.data_r_247_sv2v_reg  <= 1'b0;
      \piso.data_r_246_sv2v_reg  <= 1'b0;
      \piso.data_r_245_sv2v_reg  <= 1'b0;
      \piso.data_r_244_sv2v_reg  <= 1'b0;
      \piso.data_r_243_sv2v_reg  <= 1'b0;
      \piso.data_r_242_sv2v_reg  <= 1'b0;
      \piso.data_r_241_sv2v_reg  <= 1'b0;
      \piso.data_r_240_sv2v_reg  <= 1'b0;
      \piso.data_r_239_sv2v_reg  <= 1'b0;
      \piso.data_r_238_sv2v_reg  <= 1'b0;
      \piso.data_r_237_sv2v_reg  <= 1'b0;
      \piso.data_r_236_sv2v_reg  <= 1'b0;
      \piso.data_r_235_sv2v_reg  <= 1'b0;
      \piso.data_r_234_sv2v_reg  <= 1'b0;
      \piso.data_r_233_sv2v_reg  <= 1'b0;
      \piso.data_r_232_sv2v_reg  <= 1'b0;
      \piso.data_r_231_sv2v_reg  <= 1'b0;
      \piso.data_r_230_sv2v_reg  <= 1'b0;
      \piso.data_r_229_sv2v_reg  <= 1'b0;
      \piso.data_r_228_sv2v_reg  <= 1'b0;
      \piso.data_r_227_sv2v_reg  <= 1'b0;
      \piso.data_r_226_sv2v_reg  <= 1'b0;
      \piso.data_r_225_sv2v_reg  <= 1'b0;
      \piso.data_r_224_sv2v_reg  <= 1'b0;
      \piso.data_r_223_sv2v_reg  <= 1'b0;
      \piso.data_r_222_sv2v_reg  <= 1'b0;
      \piso.data_r_221_sv2v_reg  <= 1'b0;
      \piso.data_r_220_sv2v_reg  <= 1'b0;
      \piso.data_r_219_sv2v_reg  <= 1'b0;
      \piso.data_r_218_sv2v_reg  <= 1'b0;
      \piso.data_r_217_sv2v_reg  <= 1'b0;
      \piso.data_r_216_sv2v_reg  <= 1'b0;
      \piso.data_r_215_sv2v_reg  <= 1'b0;
      \piso.data_r_214_sv2v_reg  <= 1'b0;
      \piso.data_r_213_sv2v_reg  <= 1'b0;
      \piso.data_r_212_sv2v_reg  <= 1'b0;
      \piso.data_r_211_sv2v_reg  <= 1'b0;
      \piso.data_r_210_sv2v_reg  <= 1'b0;
      \piso.data_r_209_sv2v_reg  <= 1'b0;
      \piso.data_r_208_sv2v_reg  <= 1'b0;
      \piso.data_r_207_sv2v_reg  <= 1'b0;
      \piso.data_r_206_sv2v_reg  <= 1'b0;
      \piso.data_r_205_sv2v_reg  <= 1'b0;
      \piso.data_r_204_sv2v_reg  <= 1'b0;
      \piso.data_r_203_sv2v_reg  <= 1'b0;
      \piso.data_r_202_sv2v_reg  <= 1'b0;
      \piso.data_r_201_sv2v_reg  <= 1'b0;
      \piso.data_r_200_sv2v_reg  <= 1'b0;
      \piso.data_r_199_sv2v_reg  <= 1'b0;
      \piso.data_r_198_sv2v_reg  <= 1'b0;
      \piso.data_r_197_sv2v_reg  <= 1'b0;
      \piso.data_r_196_sv2v_reg  <= 1'b0;
      \piso.data_r_195_sv2v_reg  <= 1'b0;
      \piso.data_r_194_sv2v_reg  <= 1'b0;
      \piso.data_r_193_sv2v_reg  <= 1'b0;
      \piso.data_r_192_sv2v_reg  <= 1'b0;
      \piso.data_r_191_sv2v_reg  <= 1'b0;
      \piso.data_r_190_sv2v_reg  <= 1'b0;
      \piso.data_r_189_sv2v_reg  <= 1'b0;
      \piso.data_r_188_sv2v_reg  <= 1'b0;
      \piso.data_r_187_sv2v_reg  <= 1'b0;
      \piso.data_r_186_sv2v_reg  <= 1'b0;
      \piso.data_r_185_sv2v_reg  <= 1'b0;
      \piso.data_r_184_sv2v_reg  <= 1'b0;
      \piso.data_r_183_sv2v_reg  <= 1'b0;
      \piso.data_r_182_sv2v_reg  <= 1'b0;
      \piso.data_r_181_sv2v_reg  <= 1'b0;
      \piso.data_r_180_sv2v_reg  <= 1'b0;
      \piso.data_r_179_sv2v_reg  <= 1'b0;
      \piso.data_r_178_sv2v_reg  <= 1'b0;
      \piso.data_r_177_sv2v_reg  <= 1'b0;
      \piso.data_r_176_sv2v_reg  <= 1'b0;
      \piso.data_r_175_sv2v_reg  <= 1'b0;
      \piso.data_r_174_sv2v_reg  <= 1'b0;
      \piso.data_r_173_sv2v_reg  <= 1'b0;
      \piso.data_r_172_sv2v_reg  <= 1'b0;
      \piso.data_r_171_sv2v_reg  <= 1'b0;
      \piso.data_r_170_sv2v_reg  <= 1'b0;
      \piso.data_r_169_sv2v_reg  <= 1'b0;
      \piso.data_r_168_sv2v_reg  <= 1'b0;
      \piso.data_r_167_sv2v_reg  <= 1'b0;
      \piso.data_r_166_sv2v_reg  <= 1'b0;
      \piso.data_r_165_sv2v_reg  <= 1'b0;
      \piso.data_r_164_sv2v_reg  <= 1'b0;
      \piso.data_r_163_sv2v_reg  <= 1'b0;
      \piso.data_r_162_sv2v_reg  <= 1'b0;
      \piso.data_r_161_sv2v_reg  <= 1'b0;
      \piso.data_r_160_sv2v_reg  <= 1'b0;
      \piso.data_r_159_sv2v_reg  <= 1'b0;
      \piso.data_r_158_sv2v_reg  <= 1'b0;
      \piso.data_r_157_sv2v_reg  <= 1'b0;
      \piso.data_r_156_sv2v_reg  <= 1'b0;
      \piso.data_r_155_sv2v_reg  <= 1'b0;
      \piso.data_r_154_sv2v_reg  <= 1'b0;
      \piso.data_r_153_sv2v_reg  <= 1'b0;
      \piso.data_r_152_sv2v_reg  <= 1'b0;
      \piso.data_r_151_sv2v_reg  <= 1'b0;
      \piso.data_r_150_sv2v_reg  <= 1'b0;
      \piso.data_r_149_sv2v_reg  <= 1'b0;
      \piso.data_r_148_sv2v_reg  <= 1'b0;
      \piso.data_r_147_sv2v_reg  <= 1'b0;
      \piso.data_r_146_sv2v_reg  <= 1'b0;
      \piso.data_r_145_sv2v_reg  <= 1'b0;
      \piso.data_r_144_sv2v_reg  <= 1'b0;
      \piso.data_r_143_sv2v_reg  <= 1'b0;
      \piso.data_r_142_sv2v_reg  <= 1'b0;
      \piso.data_r_141_sv2v_reg  <= 1'b0;
      \piso.data_r_140_sv2v_reg  <= 1'b0;
      \piso.data_r_139_sv2v_reg  <= 1'b0;
      \piso.data_r_138_sv2v_reg  <= 1'b0;
      \piso.data_r_137_sv2v_reg  <= 1'b0;
      \piso.data_r_136_sv2v_reg  <= 1'b0;
      \piso.data_r_135_sv2v_reg  <= 1'b0;
      \piso.data_r_134_sv2v_reg  <= 1'b0;
      \piso.data_r_133_sv2v_reg  <= 1'b0;
      \piso.data_r_132_sv2v_reg  <= 1'b0;
      \piso.data_r_131_sv2v_reg  <= 1'b0;
      \piso.data_r_130_sv2v_reg  <= 1'b0;
      \piso.data_r_129_sv2v_reg  <= 1'b0;
      \piso.data_r_128_sv2v_reg  <= 1'b0;
      \piso.data_r_127_sv2v_reg  <= 1'b0;
      \piso.data_r_126_sv2v_reg  <= 1'b0;
      \piso.data_r_125_sv2v_reg  <= 1'b0;
      \piso.data_r_124_sv2v_reg  <= 1'b0;
      \piso.data_r_123_sv2v_reg  <= 1'b0;
      \piso.data_r_122_sv2v_reg  <= 1'b0;
      \piso.data_r_121_sv2v_reg  <= 1'b0;
      \piso.data_r_120_sv2v_reg  <= 1'b0;
      \piso.data_r_119_sv2v_reg  <= 1'b0;
      \piso.data_r_118_sv2v_reg  <= 1'b0;
      \piso.data_r_117_sv2v_reg  <= 1'b0;
      \piso.data_r_116_sv2v_reg  <= 1'b0;
      \piso.data_r_115_sv2v_reg  <= 1'b0;
      \piso.data_r_114_sv2v_reg  <= 1'b0;
      \piso.data_r_113_sv2v_reg  <= 1'b0;
      \piso.data_r_112_sv2v_reg  <= 1'b0;
      \piso.data_r_111_sv2v_reg  <= 1'b0;
      \piso.data_r_110_sv2v_reg  <= 1'b0;
      \piso.data_r_109_sv2v_reg  <= 1'b0;
      \piso.data_r_108_sv2v_reg  <= 1'b0;
      \piso.data_r_107_sv2v_reg  <= 1'b0;
      \piso.data_r_106_sv2v_reg  <= 1'b0;
      \piso.data_r_105_sv2v_reg  <= 1'b0;
      \piso.data_r_104_sv2v_reg  <= 1'b0;
      \piso.data_r_103_sv2v_reg  <= 1'b0;
      \piso.data_r_102_sv2v_reg  <= 1'b0;
      \piso.data_r_101_sv2v_reg  <= 1'b0;
      \piso.data_r_100_sv2v_reg  <= 1'b0;
      \piso.data_r_99_sv2v_reg  <= 1'b0;
      \piso.data_r_98_sv2v_reg  <= 1'b0;
      \piso.data_r_97_sv2v_reg  <= 1'b0;
      \piso.data_r_96_sv2v_reg  <= 1'b0;
      \piso.data_r_95_sv2v_reg  <= 1'b0;
      \piso.data_r_94_sv2v_reg  <= 1'b0;
      \piso.data_r_93_sv2v_reg  <= 1'b0;
      \piso.data_r_92_sv2v_reg  <= 1'b0;
      \piso.data_r_91_sv2v_reg  <= 1'b0;
      \piso.data_r_90_sv2v_reg  <= 1'b0;
      \piso.data_r_89_sv2v_reg  <= 1'b0;
      \piso.data_r_88_sv2v_reg  <= 1'b0;
      \piso.data_r_87_sv2v_reg  <= 1'b0;
      \piso.data_r_86_sv2v_reg  <= 1'b0;
      \piso.data_r_85_sv2v_reg  <= 1'b0;
      \piso.data_r_84_sv2v_reg  <= 1'b0;
      \piso.data_r_83_sv2v_reg  <= 1'b0;
      \piso.data_r_82_sv2v_reg  <= 1'b0;
      \piso.data_r_81_sv2v_reg  <= 1'b0;
      \piso.data_r_80_sv2v_reg  <= 1'b0;
      \piso.data_r_79_sv2v_reg  <= 1'b0;
      \piso.data_r_78_sv2v_reg  <= 1'b0;
      \piso.data_r_77_sv2v_reg  <= 1'b0;
      \piso.data_r_76_sv2v_reg  <= 1'b0;
      \piso.data_r_75_sv2v_reg  <= 1'b0;
      \piso.data_r_74_sv2v_reg  <= 1'b0;
      \piso.data_r_73_sv2v_reg  <= 1'b0;
      \piso.data_r_72_sv2v_reg  <= 1'b0;
      \piso.data_r_71_sv2v_reg  <= 1'b0;
      \piso.data_r_70_sv2v_reg  <= 1'b0;
      \piso.data_r_69_sv2v_reg  <= 1'b0;
      \piso.data_r_68_sv2v_reg  <= 1'b0;
      \piso.data_r_67_sv2v_reg  <= 1'b0;
      \piso.data_r_66_sv2v_reg  <= 1'b0;
      \piso.data_r_65_sv2v_reg  <= 1'b0;
      \piso.data_r_64_sv2v_reg  <= 1'b0;
      \piso.data_r_63_sv2v_reg  <= 1'b0;
      \piso.data_r_62_sv2v_reg  <= 1'b0;
      \piso.data_r_61_sv2v_reg  <= 1'b0;
      \piso.data_r_60_sv2v_reg  <= 1'b0;
      \piso.data_r_59_sv2v_reg  <= 1'b0;
      \piso.data_r_58_sv2v_reg  <= 1'b0;
      \piso.data_r_57_sv2v_reg  <= 1'b0;
      \piso.data_r_56_sv2v_reg  <= 1'b0;
      \piso.data_r_55_sv2v_reg  <= 1'b0;
      \piso.data_r_54_sv2v_reg  <= 1'b0;
      \piso.data_r_53_sv2v_reg  <= 1'b0;
      \piso.data_r_52_sv2v_reg  <= 1'b0;
      \piso.data_r_51_sv2v_reg  <= 1'b0;
      \piso.data_r_50_sv2v_reg  <= 1'b0;
      \piso.data_r_49_sv2v_reg  <= 1'b0;
      \piso.data_r_48_sv2v_reg  <= 1'b0;
      \piso.data_r_47_sv2v_reg  <= 1'b0;
      \piso.data_r_46_sv2v_reg  <= 1'b0;
      \piso.data_r_45_sv2v_reg  <= 1'b0;
      \piso.data_r_44_sv2v_reg  <= 1'b0;
      \piso.data_r_43_sv2v_reg  <= 1'b0;
      \piso.data_r_42_sv2v_reg  <= 1'b0;
      \piso.data_r_41_sv2v_reg  <= 1'b0;
      \piso.data_r_40_sv2v_reg  <= 1'b0;
      \piso.data_r_39_sv2v_reg  <= 1'b0;
      \piso.data_r_38_sv2v_reg  <= 1'b0;
      \piso.data_r_37_sv2v_reg  <= 1'b0;
      \piso.data_r_36_sv2v_reg  <= 1'b0;
      \piso.data_r_35_sv2v_reg  <= 1'b0;
      \piso.data_r_34_sv2v_reg  <= 1'b0;
      \piso.data_r_33_sv2v_reg  <= 1'b0;
      \piso.data_r_32_sv2v_reg  <= 1'b0;
      \piso.data_r_31_sv2v_reg  <= 1'b0;
      \piso.data_r_30_sv2v_reg  <= 1'b0;
      \piso.data_r_29_sv2v_reg  <= 1'b0;
      \piso.data_r_28_sv2v_reg  <= 1'b0;
      \piso.data_r_27_sv2v_reg  <= 1'b0;
      \piso.data_r_26_sv2v_reg  <= 1'b0;
      \piso.data_r_25_sv2v_reg  <= 1'b0;
      \piso.data_r_24_sv2v_reg  <= 1'b0;
      \piso.data_r_23_sv2v_reg  <= 1'b0;
      \piso.data_r_22_sv2v_reg  <= 1'b0;
      \piso.data_r_21_sv2v_reg  <= 1'b0;
      \piso.data_r_20_sv2v_reg  <= 1'b0;
      \piso.data_r_19_sv2v_reg  <= 1'b0;
      \piso.data_r_18_sv2v_reg  <= 1'b0;
      \piso.data_r_17_sv2v_reg  <= 1'b0;
      \piso.data_r_16_sv2v_reg  <= 1'b0;
      \piso.data_r_15_sv2v_reg  <= 1'b0;
      \piso.data_r_14_sv2v_reg  <= 1'b0;
      \piso.data_r_13_sv2v_reg  <= 1'b0;
      \piso.data_r_12_sv2v_reg  <= 1'b0;
      \piso.data_r_11_sv2v_reg  <= 1'b0;
      \piso.data_r_10_sv2v_reg  <= 1'b0;
      \piso.data_r_9_sv2v_reg  <= 1'b0;
      \piso.data_r_8_sv2v_reg  <= 1'b0;
      \piso.data_r_7_sv2v_reg  <= 1'b0;
      \piso.data_r_6_sv2v_reg  <= 1'b0;
      \piso.data_r_5_sv2v_reg  <= 1'b0;
      \piso.data_r_4_sv2v_reg  <= 1'b0;
      \piso.data_r_3_sv2v_reg  <= 1'b0;
      \piso.data_r_2_sv2v_reg  <= 1'b0;
      \piso.data_r_1_sv2v_reg  <= 1'b0;
      \piso.data_r_0_sv2v_reg  <= 1'b0;
    end else if(N6) begin
      \piso.data_r_2047_sv2v_reg  <= \piso.data_li [2047];
      \piso.data_r_2046_sv2v_reg  <= \piso.data_li [2046];
      \piso.data_r_2045_sv2v_reg  <= \piso.data_li [2045];
      \piso.data_r_2044_sv2v_reg  <= \piso.data_li [2044];
      \piso.data_r_2043_sv2v_reg  <= \piso.data_li [2043];
      \piso.data_r_2042_sv2v_reg  <= \piso.data_li [2042];
      \piso.data_r_2041_sv2v_reg  <= \piso.data_li [2041];
      \piso.data_r_2040_sv2v_reg  <= \piso.data_li [2040];
      \piso.data_r_2039_sv2v_reg  <= \piso.data_li [2039];
      \piso.data_r_2038_sv2v_reg  <= \piso.data_li [2038];
      \piso.data_r_2037_sv2v_reg  <= \piso.data_li [2037];
      \piso.data_r_2036_sv2v_reg  <= \piso.data_li [2036];
      \piso.data_r_2035_sv2v_reg  <= \piso.data_li [2035];
      \piso.data_r_2034_sv2v_reg  <= \piso.data_li [2034];
      \piso.data_r_2033_sv2v_reg  <= \piso.data_li [2033];
      \piso.data_r_2032_sv2v_reg  <= \piso.data_li [2032];
      \piso.data_r_2031_sv2v_reg  <= \piso.data_li [2031];
      \piso.data_r_2030_sv2v_reg  <= \piso.data_li [2030];
      \piso.data_r_2029_sv2v_reg  <= \piso.data_li [2029];
      \piso.data_r_2028_sv2v_reg  <= \piso.data_li [2028];
      \piso.data_r_2027_sv2v_reg  <= \piso.data_li [2027];
      \piso.data_r_2026_sv2v_reg  <= \piso.data_li [2026];
      \piso.data_r_2025_sv2v_reg  <= \piso.data_li [2025];
      \piso.data_r_2024_sv2v_reg  <= \piso.data_li [2024];
      \piso.data_r_2023_sv2v_reg  <= \piso.data_li [2023];
      \piso.data_r_2022_sv2v_reg  <= \piso.data_li [2022];
      \piso.data_r_2021_sv2v_reg  <= \piso.data_li [2021];
      \piso.data_r_2020_sv2v_reg  <= \piso.data_li [2020];
      \piso.data_r_2019_sv2v_reg  <= \piso.data_li [2019];
      \piso.data_r_2018_sv2v_reg  <= \piso.data_li [2018];
      \piso.data_r_2017_sv2v_reg  <= \piso.data_li [2017];
      \piso.data_r_2016_sv2v_reg  <= \piso.data_li [2016];
      \piso.data_r_2015_sv2v_reg  <= \piso.data_li [2015];
      \piso.data_r_2014_sv2v_reg  <= \piso.data_li [2014];
      \piso.data_r_2013_sv2v_reg  <= \piso.data_li [2013];
      \piso.data_r_2012_sv2v_reg  <= \piso.data_li [2012];
      \piso.data_r_2011_sv2v_reg  <= \piso.data_li [2011];
      \piso.data_r_2010_sv2v_reg  <= \piso.data_li [2010];
      \piso.data_r_2009_sv2v_reg  <= \piso.data_li [2009];
      \piso.data_r_2008_sv2v_reg  <= \piso.data_li [2008];
      \piso.data_r_2007_sv2v_reg  <= \piso.data_li [2007];
      \piso.data_r_2006_sv2v_reg  <= \piso.data_li [2006];
      \piso.data_r_2005_sv2v_reg  <= \piso.data_li [2005];
      \piso.data_r_2004_sv2v_reg  <= \piso.data_li [2004];
      \piso.data_r_2003_sv2v_reg  <= \piso.data_li [2003];
      \piso.data_r_2002_sv2v_reg  <= \piso.data_li [2002];
      \piso.data_r_2001_sv2v_reg  <= \piso.data_li [2001];
      \piso.data_r_2000_sv2v_reg  <= \piso.data_li [2000];
      \piso.data_r_1999_sv2v_reg  <= \piso.data_li [1999];
      \piso.data_r_1998_sv2v_reg  <= \piso.data_li [1998];
      \piso.data_r_1997_sv2v_reg  <= \piso.data_li [1997];
      \piso.data_r_1996_sv2v_reg  <= \piso.data_li [1996];
      \piso.data_r_1995_sv2v_reg  <= \piso.data_li [1995];
      \piso.data_r_1994_sv2v_reg  <= \piso.data_li [1994];
      \piso.data_r_1993_sv2v_reg  <= \piso.data_li [1993];
      \piso.data_r_1992_sv2v_reg  <= \piso.data_li [1992];
      \piso.data_r_1991_sv2v_reg  <= \piso.data_li [1991];
      \piso.data_r_1990_sv2v_reg  <= \piso.data_li [1990];
      \piso.data_r_1989_sv2v_reg  <= \piso.data_li [1989];
      \piso.data_r_1988_sv2v_reg  <= \piso.data_li [1988];
      \piso.data_r_1987_sv2v_reg  <= \piso.data_li [1987];
      \piso.data_r_1986_sv2v_reg  <= \piso.data_li [1986];
      \piso.data_r_1985_sv2v_reg  <= \piso.data_li [1985];
      \piso.data_r_1984_sv2v_reg  <= \piso.data_li [1984];
      \piso.data_r_1983_sv2v_reg  <= \piso.data_li [1983];
      \piso.data_r_1982_sv2v_reg  <= \piso.data_li [1982];
      \piso.data_r_1981_sv2v_reg  <= \piso.data_li [1981];
      \piso.data_r_1980_sv2v_reg  <= \piso.data_li [1980];
      \piso.data_r_1979_sv2v_reg  <= \piso.data_li [1979];
      \piso.data_r_1978_sv2v_reg  <= \piso.data_li [1978];
      \piso.data_r_1977_sv2v_reg  <= \piso.data_li [1977];
      \piso.data_r_1976_sv2v_reg  <= \piso.data_li [1976];
      \piso.data_r_1975_sv2v_reg  <= \piso.data_li [1975];
      \piso.data_r_1974_sv2v_reg  <= \piso.data_li [1974];
      \piso.data_r_1973_sv2v_reg  <= \piso.data_li [1973];
      \piso.data_r_1972_sv2v_reg  <= \piso.data_li [1972];
      \piso.data_r_1971_sv2v_reg  <= \piso.data_li [1971];
      \piso.data_r_1970_sv2v_reg  <= \piso.data_li [1970];
      \piso.data_r_1969_sv2v_reg  <= \piso.data_li [1969];
      \piso.data_r_1968_sv2v_reg  <= \piso.data_li [1968];
      \piso.data_r_1967_sv2v_reg  <= \piso.data_li [1967];
      \piso.data_r_1966_sv2v_reg  <= \piso.data_li [1966];
      \piso.data_r_1965_sv2v_reg  <= \piso.data_li [1965];
      \piso.data_r_1964_sv2v_reg  <= \piso.data_li [1964];
      \piso.data_r_1963_sv2v_reg  <= \piso.data_li [1963];
      \piso.data_r_1962_sv2v_reg  <= \piso.data_li [1962];
      \piso.data_r_1961_sv2v_reg  <= \piso.data_li [1961];
      \piso.data_r_1960_sv2v_reg  <= \piso.data_li [1960];
      \piso.data_r_1959_sv2v_reg  <= \piso.data_li [1959];
      \piso.data_r_1958_sv2v_reg  <= \piso.data_li [1958];
      \piso.data_r_1957_sv2v_reg  <= \piso.data_li [1957];
      \piso.data_r_1956_sv2v_reg  <= \piso.data_li [1956];
      \piso.data_r_1955_sv2v_reg  <= \piso.data_li [1955];
      \piso.data_r_1954_sv2v_reg  <= \piso.data_li [1954];
      \piso.data_r_1953_sv2v_reg  <= \piso.data_li [1953];
      \piso.data_r_1952_sv2v_reg  <= \piso.data_li [1952];
      \piso.data_r_1951_sv2v_reg  <= \piso.data_li [1951];
      \piso.data_r_1950_sv2v_reg  <= \piso.data_li [1950];
      \piso.data_r_1949_sv2v_reg  <= \piso.data_li [1949];
      \piso.data_r_1948_sv2v_reg  <= \piso.data_li [1948];
      \piso.data_r_1947_sv2v_reg  <= \piso.data_li [1947];
      \piso.data_r_1946_sv2v_reg  <= \piso.data_li [1946];
      \piso.data_r_1945_sv2v_reg  <= \piso.data_li [1945];
      \piso.data_r_1944_sv2v_reg  <= \piso.data_li [1944];
      \piso.data_r_1943_sv2v_reg  <= \piso.data_li [1943];
      \piso.data_r_1942_sv2v_reg  <= \piso.data_li [1942];
      \piso.data_r_1941_sv2v_reg  <= \piso.data_li [1941];
      \piso.data_r_1940_sv2v_reg  <= \piso.data_li [1940];
      \piso.data_r_1939_sv2v_reg  <= \piso.data_li [1939];
      \piso.data_r_1938_sv2v_reg  <= \piso.data_li [1938];
      \piso.data_r_1937_sv2v_reg  <= \piso.data_li [1937];
      \piso.data_r_1936_sv2v_reg  <= \piso.data_li [1936];
      \piso.data_r_1935_sv2v_reg  <= \piso.data_li [1935];
      \piso.data_r_1934_sv2v_reg  <= \piso.data_li [1934];
      \piso.data_r_1933_sv2v_reg  <= \piso.data_li [1933];
      \piso.data_r_1932_sv2v_reg  <= \piso.data_li [1932];
      \piso.data_r_1931_sv2v_reg  <= \piso.data_li [1931];
      \piso.data_r_1930_sv2v_reg  <= \piso.data_li [1930];
      \piso.data_r_1929_sv2v_reg  <= \piso.data_li [1929];
      \piso.data_r_1928_sv2v_reg  <= \piso.data_li [1928];
      \piso.data_r_1927_sv2v_reg  <= \piso.data_li [1927];
      \piso.data_r_1926_sv2v_reg  <= \piso.data_li [1926];
      \piso.data_r_1925_sv2v_reg  <= \piso.data_li [1925];
      \piso.data_r_1924_sv2v_reg  <= \piso.data_li [1924];
      \piso.data_r_1923_sv2v_reg  <= \piso.data_li [1923];
      \piso.data_r_1922_sv2v_reg  <= \piso.data_li [1922];
      \piso.data_r_1921_sv2v_reg  <= \piso.data_li [1921];
      \piso.data_r_1920_sv2v_reg  <= \piso.data_li [1920];
      \piso.data_r_1919_sv2v_reg  <= \piso.data_li [1919];
      \piso.data_r_1918_sv2v_reg  <= \piso.data_li [1918];
      \piso.data_r_1917_sv2v_reg  <= \piso.data_li [1917];
      \piso.data_r_1916_sv2v_reg  <= \piso.data_li [1916];
      \piso.data_r_1915_sv2v_reg  <= \piso.data_li [1915];
      \piso.data_r_1914_sv2v_reg  <= \piso.data_li [1914];
      \piso.data_r_1913_sv2v_reg  <= \piso.data_li [1913];
      \piso.data_r_1912_sv2v_reg  <= \piso.data_li [1912];
      \piso.data_r_1911_sv2v_reg  <= \piso.data_li [1911];
      \piso.data_r_1910_sv2v_reg  <= \piso.data_li [1910];
      \piso.data_r_1909_sv2v_reg  <= \piso.data_li [1909];
      \piso.data_r_1908_sv2v_reg  <= \piso.data_li [1908];
      \piso.data_r_1907_sv2v_reg  <= \piso.data_li [1907];
      \piso.data_r_1906_sv2v_reg  <= \piso.data_li [1906];
      \piso.data_r_1905_sv2v_reg  <= \piso.data_li [1905];
      \piso.data_r_1904_sv2v_reg  <= \piso.data_li [1904];
      \piso.data_r_1903_sv2v_reg  <= \piso.data_li [1903];
      \piso.data_r_1902_sv2v_reg  <= \piso.data_li [1902];
      \piso.data_r_1901_sv2v_reg  <= \piso.data_li [1901];
      \piso.data_r_1900_sv2v_reg  <= \piso.data_li [1900];
      \piso.data_r_1899_sv2v_reg  <= \piso.data_li [1899];
      \piso.data_r_1898_sv2v_reg  <= \piso.data_li [1898];
      \piso.data_r_1897_sv2v_reg  <= \piso.data_li [1897];
      \piso.data_r_1896_sv2v_reg  <= \piso.data_li [1896];
      \piso.data_r_1895_sv2v_reg  <= \piso.data_li [1895];
      \piso.data_r_1894_sv2v_reg  <= \piso.data_li [1894];
      \piso.data_r_1893_sv2v_reg  <= \piso.data_li [1893];
      \piso.data_r_1892_sv2v_reg  <= \piso.data_li [1892];
      \piso.data_r_1891_sv2v_reg  <= \piso.data_li [1891];
      \piso.data_r_1890_sv2v_reg  <= \piso.data_li [1890];
      \piso.data_r_1889_sv2v_reg  <= \piso.data_li [1889];
      \piso.data_r_1888_sv2v_reg  <= \piso.data_li [1888];
      \piso.data_r_1887_sv2v_reg  <= \piso.data_li [1887];
      \piso.data_r_1886_sv2v_reg  <= \piso.data_li [1886];
      \piso.data_r_1885_sv2v_reg  <= \piso.data_li [1885];
      \piso.data_r_1884_sv2v_reg  <= \piso.data_li [1884];
      \piso.data_r_1883_sv2v_reg  <= \piso.data_li [1883];
      \piso.data_r_1882_sv2v_reg  <= \piso.data_li [1882];
      \piso.data_r_1881_sv2v_reg  <= \piso.data_li [1881];
      \piso.data_r_1880_sv2v_reg  <= \piso.data_li [1880];
      \piso.data_r_1879_sv2v_reg  <= \piso.data_li [1879];
      \piso.data_r_1878_sv2v_reg  <= \piso.data_li [1878];
      \piso.data_r_1877_sv2v_reg  <= \piso.data_li [1877];
      \piso.data_r_1876_sv2v_reg  <= \piso.data_li [1876];
      \piso.data_r_1875_sv2v_reg  <= \piso.data_li [1875];
      \piso.data_r_1874_sv2v_reg  <= \piso.data_li [1874];
      \piso.data_r_1873_sv2v_reg  <= \piso.data_li [1873];
      \piso.data_r_1872_sv2v_reg  <= \piso.data_li [1872];
      \piso.data_r_1871_sv2v_reg  <= \piso.data_li [1871];
      \piso.data_r_1870_sv2v_reg  <= \piso.data_li [1870];
      \piso.data_r_1869_sv2v_reg  <= \piso.data_li [1869];
      \piso.data_r_1868_sv2v_reg  <= \piso.data_li [1868];
      \piso.data_r_1867_sv2v_reg  <= \piso.data_li [1867];
      \piso.data_r_1866_sv2v_reg  <= \piso.data_li [1866];
      \piso.data_r_1865_sv2v_reg  <= \piso.data_li [1865];
      \piso.data_r_1864_sv2v_reg  <= \piso.data_li [1864];
      \piso.data_r_1863_sv2v_reg  <= \piso.data_li [1863];
      \piso.data_r_1862_sv2v_reg  <= \piso.data_li [1862];
      \piso.data_r_1861_sv2v_reg  <= \piso.data_li [1861];
      \piso.data_r_1860_sv2v_reg  <= \piso.data_li [1860];
      \piso.data_r_1859_sv2v_reg  <= \piso.data_li [1859];
      \piso.data_r_1858_sv2v_reg  <= \piso.data_li [1858];
      \piso.data_r_1857_sv2v_reg  <= \piso.data_li [1857];
      \piso.data_r_1856_sv2v_reg  <= \piso.data_li [1856];
      \piso.data_r_1855_sv2v_reg  <= \piso.data_li [1855];
      \piso.data_r_1854_sv2v_reg  <= \piso.data_li [1854];
      \piso.data_r_1853_sv2v_reg  <= \piso.data_li [1853];
      \piso.data_r_1852_sv2v_reg  <= \piso.data_li [1852];
      \piso.data_r_1851_sv2v_reg  <= \piso.data_li [1851];
      \piso.data_r_1850_sv2v_reg  <= \piso.data_li [1850];
      \piso.data_r_1849_sv2v_reg  <= \piso.data_li [1849];
      \piso.data_r_1848_sv2v_reg  <= \piso.data_li [1848];
      \piso.data_r_1847_sv2v_reg  <= \piso.data_li [1847];
      \piso.data_r_1846_sv2v_reg  <= \piso.data_li [1846];
      \piso.data_r_1845_sv2v_reg  <= \piso.data_li [1845];
      \piso.data_r_1844_sv2v_reg  <= \piso.data_li [1844];
      \piso.data_r_1843_sv2v_reg  <= \piso.data_li [1843];
      \piso.data_r_1842_sv2v_reg  <= \piso.data_li [1842];
      \piso.data_r_1841_sv2v_reg  <= \piso.data_li [1841];
      \piso.data_r_1840_sv2v_reg  <= \piso.data_li [1840];
      \piso.data_r_1839_sv2v_reg  <= \piso.data_li [1839];
      \piso.data_r_1838_sv2v_reg  <= \piso.data_li [1838];
      \piso.data_r_1837_sv2v_reg  <= \piso.data_li [1837];
      \piso.data_r_1836_sv2v_reg  <= \piso.data_li [1836];
      \piso.data_r_1835_sv2v_reg  <= \piso.data_li [1835];
      \piso.data_r_1834_sv2v_reg  <= \piso.data_li [1834];
      \piso.data_r_1833_sv2v_reg  <= \piso.data_li [1833];
      \piso.data_r_1832_sv2v_reg  <= \piso.data_li [1832];
      \piso.data_r_1831_sv2v_reg  <= \piso.data_li [1831];
      \piso.data_r_1830_sv2v_reg  <= \piso.data_li [1830];
      \piso.data_r_1829_sv2v_reg  <= \piso.data_li [1829];
      \piso.data_r_1828_sv2v_reg  <= \piso.data_li [1828];
      \piso.data_r_1827_sv2v_reg  <= \piso.data_li [1827];
      \piso.data_r_1826_sv2v_reg  <= \piso.data_li [1826];
      \piso.data_r_1825_sv2v_reg  <= \piso.data_li [1825];
      \piso.data_r_1824_sv2v_reg  <= \piso.data_li [1824];
      \piso.data_r_1823_sv2v_reg  <= \piso.data_li [1823];
      \piso.data_r_1822_sv2v_reg  <= \piso.data_li [1822];
      \piso.data_r_1821_sv2v_reg  <= \piso.data_li [1821];
      \piso.data_r_1820_sv2v_reg  <= \piso.data_li [1820];
      \piso.data_r_1819_sv2v_reg  <= \piso.data_li [1819];
      \piso.data_r_1818_sv2v_reg  <= \piso.data_li [1818];
      \piso.data_r_1817_sv2v_reg  <= \piso.data_li [1817];
      \piso.data_r_1816_sv2v_reg  <= \piso.data_li [1816];
      \piso.data_r_1815_sv2v_reg  <= \piso.data_li [1815];
      \piso.data_r_1814_sv2v_reg  <= \piso.data_li [1814];
      \piso.data_r_1813_sv2v_reg  <= \piso.data_li [1813];
      \piso.data_r_1812_sv2v_reg  <= \piso.data_li [1812];
      \piso.data_r_1811_sv2v_reg  <= \piso.data_li [1811];
      \piso.data_r_1810_sv2v_reg  <= \piso.data_li [1810];
      \piso.data_r_1809_sv2v_reg  <= \piso.data_li [1809];
      \piso.data_r_1808_sv2v_reg  <= \piso.data_li [1808];
      \piso.data_r_1807_sv2v_reg  <= \piso.data_li [1807];
      \piso.data_r_1806_sv2v_reg  <= \piso.data_li [1806];
      \piso.data_r_1805_sv2v_reg  <= \piso.data_li [1805];
      \piso.data_r_1804_sv2v_reg  <= \piso.data_li [1804];
      \piso.data_r_1803_sv2v_reg  <= \piso.data_li [1803];
      \piso.data_r_1802_sv2v_reg  <= \piso.data_li [1802];
      \piso.data_r_1801_sv2v_reg  <= \piso.data_li [1801];
      \piso.data_r_1800_sv2v_reg  <= \piso.data_li [1800];
      \piso.data_r_1799_sv2v_reg  <= \piso.data_li [1799];
      \piso.data_r_1798_sv2v_reg  <= \piso.data_li [1798];
      \piso.data_r_1797_sv2v_reg  <= \piso.data_li [1797];
      \piso.data_r_1796_sv2v_reg  <= \piso.data_li [1796];
      \piso.data_r_1795_sv2v_reg  <= \piso.data_li [1795];
      \piso.data_r_1794_sv2v_reg  <= \piso.data_li [1794];
      \piso.data_r_1793_sv2v_reg  <= \piso.data_li [1793];
      \piso.data_r_1792_sv2v_reg  <= \piso.data_li [1792];
      \piso.data_r_1791_sv2v_reg  <= \piso.data_li [1791];
      \piso.data_r_1790_sv2v_reg  <= \piso.data_li [1790];
      \piso.data_r_1789_sv2v_reg  <= \piso.data_li [1789];
      \piso.data_r_1788_sv2v_reg  <= \piso.data_li [1788];
      \piso.data_r_1787_sv2v_reg  <= \piso.data_li [1787];
      \piso.data_r_1786_sv2v_reg  <= \piso.data_li [1786];
      \piso.data_r_1785_sv2v_reg  <= \piso.data_li [1785];
      \piso.data_r_1784_sv2v_reg  <= \piso.data_li [1784];
      \piso.data_r_1783_sv2v_reg  <= \piso.data_li [1783];
      \piso.data_r_1782_sv2v_reg  <= \piso.data_li [1782];
      \piso.data_r_1781_sv2v_reg  <= \piso.data_li [1781];
      \piso.data_r_1780_sv2v_reg  <= \piso.data_li [1780];
      \piso.data_r_1779_sv2v_reg  <= \piso.data_li [1779];
      \piso.data_r_1778_sv2v_reg  <= \piso.data_li [1778];
      \piso.data_r_1777_sv2v_reg  <= \piso.data_li [1777];
      \piso.data_r_1776_sv2v_reg  <= \piso.data_li [1776];
      \piso.data_r_1775_sv2v_reg  <= \piso.data_li [1775];
      \piso.data_r_1774_sv2v_reg  <= \piso.data_li [1774];
      \piso.data_r_1773_sv2v_reg  <= \piso.data_li [1773];
      \piso.data_r_1772_sv2v_reg  <= \piso.data_li [1772];
      \piso.data_r_1771_sv2v_reg  <= \piso.data_li [1771];
      \piso.data_r_1770_sv2v_reg  <= \piso.data_li [1770];
      \piso.data_r_1769_sv2v_reg  <= \piso.data_li [1769];
      \piso.data_r_1768_sv2v_reg  <= \piso.data_li [1768];
      \piso.data_r_1767_sv2v_reg  <= \piso.data_li [1767];
      \piso.data_r_1766_sv2v_reg  <= \piso.data_li [1766];
      \piso.data_r_1765_sv2v_reg  <= \piso.data_li [1765];
      \piso.data_r_1764_sv2v_reg  <= \piso.data_li [1764];
      \piso.data_r_1763_sv2v_reg  <= \piso.data_li [1763];
      \piso.data_r_1762_sv2v_reg  <= \piso.data_li [1762];
      \piso.data_r_1761_sv2v_reg  <= \piso.data_li [1761];
      \piso.data_r_1760_sv2v_reg  <= \piso.data_li [1760];
      \piso.data_r_1759_sv2v_reg  <= \piso.data_li [1759];
      \piso.data_r_1758_sv2v_reg  <= \piso.data_li [1758];
      \piso.data_r_1757_sv2v_reg  <= \piso.data_li [1757];
      \piso.data_r_1756_sv2v_reg  <= \piso.data_li [1756];
      \piso.data_r_1755_sv2v_reg  <= \piso.data_li [1755];
      \piso.data_r_1754_sv2v_reg  <= \piso.data_li [1754];
      \piso.data_r_1753_sv2v_reg  <= \piso.data_li [1753];
      \piso.data_r_1752_sv2v_reg  <= \piso.data_li [1752];
      \piso.data_r_1751_sv2v_reg  <= \piso.data_li [1751];
      \piso.data_r_1750_sv2v_reg  <= \piso.data_li [1750];
      \piso.data_r_1749_sv2v_reg  <= \piso.data_li [1749];
      \piso.data_r_1748_sv2v_reg  <= \piso.data_li [1748];
      \piso.data_r_1747_sv2v_reg  <= \piso.data_li [1747];
      \piso.data_r_1746_sv2v_reg  <= \piso.data_li [1746];
      \piso.data_r_1745_sv2v_reg  <= \piso.data_li [1745];
      \piso.data_r_1744_sv2v_reg  <= \piso.data_li [1744];
      \piso.data_r_1743_sv2v_reg  <= \piso.data_li [1743];
      \piso.data_r_1742_sv2v_reg  <= \piso.data_li [1742];
      \piso.data_r_1741_sv2v_reg  <= \piso.data_li [1741];
      \piso.data_r_1740_sv2v_reg  <= \piso.data_li [1740];
      \piso.data_r_1739_sv2v_reg  <= \piso.data_li [1739];
      \piso.data_r_1738_sv2v_reg  <= \piso.data_li [1738];
      \piso.data_r_1737_sv2v_reg  <= \piso.data_li [1737];
      \piso.data_r_1736_sv2v_reg  <= \piso.data_li [1736];
      \piso.data_r_1735_sv2v_reg  <= \piso.data_li [1735];
      \piso.data_r_1734_sv2v_reg  <= \piso.data_li [1734];
      \piso.data_r_1733_sv2v_reg  <= \piso.data_li [1733];
      \piso.data_r_1732_sv2v_reg  <= \piso.data_li [1732];
      \piso.data_r_1731_sv2v_reg  <= \piso.data_li [1731];
      \piso.data_r_1730_sv2v_reg  <= \piso.data_li [1730];
      \piso.data_r_1729_sv2v_reg  <= \piso.data_li [1729];
      \piso.data_r_1728_sv2v_reg  <= \piso.data_li [1728];
      \piso.data_r_1727_sv2v_reg  <= \piso.data_li [1727];
      \piso.data_r_1726_sv2v_reg  <= \piso.data_li [1726];
      \piso.data_r_1725_sv2v_reg  <= \piso.data_li [1725];
      \piso.data_r_1724_sv2v_reg  <= \piso.data_li [1724];
      \piso.data_r_1723_sv2v_reg  <= \piso.data_li [1723];
      \piso.data_r_1722_sv2v_reg  <= \piso.data_li [1722];
      \piso.data_r_1721_sv2v_reg  <= \piso.data_li [1721];
      \piso.data_r_1720_sv2v_reg  <= \piso.data_li [1720];
      \piso.data_r_1719_sv2v_reg  <= \piso.data_li [1719];
      \piso.data_r_1718_sv2v_reg  <= \piso.data_li [1718];
      \piso.data_r_1717_sv2v_reg  <= \piso.data_li [1717];
      \piso.data_r_1716_sv2v_reg  <= \piso.data_li [1716];
      \piso.data_r_1715_sv2v_reg  <= \piso.data_li [1715];
      \piso.data_r_1714_sv2v_reg  <= \piso.data_li [1714];
      \piso.data_r_1713_sv2v_reg  <= \piso.data_li [1713];
      \piso.data_r_1712_sv2v_reg  <= \piso.data_li [1712];
      \piso.data_r_1711_sv2v_reg  <= \piso.data_li [1711];
      \piso.data_r_1710_sv2v_reg  <= \piso.data_li [1710];
      \piso.data_r_1709_sv2v_reg  <= \piso.data_li [1709];
      \piso.data_r_1708_sv2v_reg  <= \piso.data_li [1708];
      \piso.data_r_1707_sv2v_reg  <= \piso.data_li [1707];
      \piso.data_r_1706_sv2v_reg  <= \piso.data_li [1706];
      \piso.data_r_1705_sv2v_reg  <= \piso.data_li [1705];
      \piso.data_r_1704_sv2v_reg  <= \piso.data_li [1704];
      \piso.data_r_1703_sv2v_reg  <= \piso.data_li [1703];
      \piso.data_r_1702_sv2v_reg  <= \piso.data_li [1702];
      \piso.data_r_1701_sv2v_reg  <= \piso.data_li [1701];
      \piso.data_r_1700_sv2v_reg  <= \piso.data_li [1700];
      \piso.data_r_1699_sv2v_reg  <= \piso.data_li [1699];
      \piso.data_r_1698_sv2v_reg  <= \piso.data_li [1698];
      \piso.data_r_1697_sv2v_reg  <= \piso.data_li [1697];
      \piso.data_r_1696_sv2v_reg  <= \piso.data_li [1696];
      \piso.data_r_1695_sv2v_reg  <= \piso.data_li [1695];
      \piso.data_r_1694_sv2v_reg  <= \piso.data_li [1694];
      \piso.data_r_1693_sv2v_reg  <= \piso.data_li [1693];
      \piso.data_r_1692_sv2v_reg  <= \piso.data_li [1692];
      \piso.data_r_1691_sv2v_reg  <= \piso.data_li [1691];
      \piso.data_r_1690_sv2v_reg  <= \piso.data_li [1690];
      \piso.data_r_1689_sv2v_reg  <= \piso.data_li [1689];
      \piso.data_r_1688_sv2v_reg  <= \piso.data_li [1688];
      \piso.data_r_1687_sv2v_reg  <= \piso.data_li [1687];
      \piso.data_r_1686_sv2v_reg  <= \piso.data_li [1686];
      \piso.data_r_1685_sv2v_reg  <= \piso.data_li [1685];
      \piso.data_r_1684_sv2v_reg  <= \piso.data_li [1684];
      \piso.data_r_1683_sv2v_reg  <= \piso.data_li [1683];
      \piso.data_r_1682_sv2v_reg  <= \piso.data_li [1682];
      \piso.data_r_1681_sv2v_reg  <= \piso.data_li [1681];
      \piso.data_r_1680_sv2v_reg  <= \piso.data_li [1680];
      \piso.data_r_1679_sv2v_reg  <= \piso.data_li [1679];
      \piso.data_r_1678_sv2v_reg  <= \piso.data_li [1678];
      \piso.data_r_1677_sv2v_reg  <= \piso.data_li [1677];
      \piso.data_r_1676_sv2v_reg  <= \piso.data_li [1676];
      \piso.data_r_1675_sv2v_reg  <= \piso.data_li [1675];
      \piso.data_r_1674_sv2v_reg  <= \piso.data_li [1674];
      \piso.data_r_1673_sv2v_reg  <= \piso.data_li [1673];
      \piso.data_r_1672_sv2v_reg  <= \piso.data_li [1672];
      \piso.data_r_1671_sv2v_reg  <= \piso.data_li [1671];
      \piso.data_r_1670_sv2v_reg  <= \piso.data_li [1670];
      \piso.data_r_1669_sv2v_reg  <= \piso.data_li [1669];
      \piso.data_r_1668_sv2v_reg  <= \piso.data_li [1668];
      \piso.data_r_1667_sv2v_reg  <= \piso.data_li [1667];
      \piso.data_r_1666_sv2v_reg  <= \piso.data_li [1666];
      \piso.data_r_1665_sv2v_reg  <= \piso.data_li [1665];
      \piso.data_r_1664_sv2v_reg  <= \piso.data_li [1664];
      \piso.data_r_1663_sv2v_reg  <= \piso.data_li [1663];
      \piso.data_r_1662_sv2v_reg  <= \piso.data_li [1662];
      \piso.data_r_1661_sv2v_reg  <= \piso.data_li [1661];
      \piso.data_r_1660_sv2v_reg  <= \piso.data_li [1660];
      \piso.data_r_1659_sv2v_reg  <= \piso.data_li [1659];
      \piso.data_r_1658_sv2v_reg  <= \piso.data_li [1658];
      \piso.data_r_1657_sv2v_reg  <= \piso.data_li [1657];
      \piso.data_r_1656_sv2v_reg  <= \piso.data_li [1656];
      \piso.data_r_1655_sv2v_reg  <= \piso.data_li [1655];
      \piso.data_r_1654_sv2v_reg  <= \piso.data_li [1654];
      \piso.data_r_1653_sv2v_reg  <= \piso.data_li [1653];
      \piso.data_r_1652_sv2v_reg  <= \piso.data_li [1652];
      \piso.data_r_1651_sv2v_reg  <= \piso.data_li [1651];
      \piso.data_r_1650_sv2v_reg  <= \piso.data_li [1650];
      \piso.data_r_1649_sv2v_reg  <= \piso.data_li [1649];
      \piso.data_r_1648_sv2v_reg  <= \piso.data_li [1648];
      \piso.data_r_1647_sv2v_reg  <= \piso.data_li [1647];
      \piso.data_r_1646_sv2v_reg  <= \piso.data_li [1646];
      \piso.data_r_1645_sv2v_reg  <= \piso.data_li [1645];
      \piso.data_r_1644_sv2v_reg  <= \piso.data_li [1644];
      \piso.data_r_1643_sv2v_reg  <= \piso.data_li [1643];
      \piso.data_r_1642_sv2v_reg  <= \piso.data_li [1642];
      \piso.data_r_1641_sv2v_reg  <= \piso.data_li [1641];
      \piso.data_r_1640_sv2v_reg  <= \piso.data_li [1640];
      \piso.data_r_1639_sv2v_reg  <= \piso.data_li [1639];
      \piso.data_r_1638_sv2v_reg  <= \piso.data_li [1638];
      \piso.data_r_1637_sv2v_reg  <= \piso.data_li [1637];
      \piso.data_r_1636_sv2v_reg  <= \piso.data_li [1636];
      \piso.data_r_1635_sv2v_reg  <= \piso.data_li [1635];
      \piso.data_r_1634_sv2v_reg  <= \piso.data_li [1634];
      \piso.data_r_1633_sv2v_reg  <= \piso.data_li [1633];
      \piso.data_r_1632_sv2v_reg  <= \piso.data_li [1632];
      \piso.data_r_1631_sv2v_reg  <= \piso.data_li [1631];
      \piso.data_r_1630_sv2v_reg  <= \piso.data_li [1630];
      \piso.data_r_1629_sv2v_reg  <= \piso.data_li [1629];
      \piso.data_r_1628_sv2v_reg  <= \piso.data_li [1628];
      \piso.data_r_1627_sv2v_reg  <= \piso.data_li [1627];
      \piso.data_r_1626_sv2v_reg  <= \piso.data_li [1626];
      \piso.data_r_1625_sv2v_reg  <= \piso.data_li [1625];
      \piso.data_r_1624_sv2v_reg  <= \piso.data_li [1624];
      \piso.data_r_1623_sv2v_reg  <= \piso.data_li [1623];
      \piso.data_r_1622_sv2v_reg  <= \piso.data_li [1622];
      \piso.data_r_1621_sv2v_reg  <= \piso.data_li [1621];
      \piso.data_r_1620_sv2v_reg  <= \piso.data_li [1620];
      \piso.data_r_1619_sv2v_reg  <= \piso.data_li [1619];
      \piso.data_r_1618_sv2v_reg  <= \piso.data_li [1618];
      \piso.data_r_1617_sv2v_reg  <= \piso.data_li [1617];
      \piso.data_r_1616_sv2v_reg  <= \piso.data_li [1616];
      \piso.data_r_1615_sv2v_reg  <= \piso.data_li [1615];
      \piso.data_r_1614_sv2v_reg  <= \piso.data_li [1614];
      \piso.data_r_1613_sv2v_reg  <= \piso.data_li [1613];
      \piso.data_r_1612_sv2v_reg  <= \piso.data_li [1612];
      \piso.data_r_1611_sv2v_reg  <= \piso.data_li [1611];
      \piso.data_r_1610_sv2v_reg  <= \piso.data_li [1610];
      \piso.data_r_1609_sv2v_reg  <= \piso.data_li [1609];
      \piso.data_r_1608_sv2v_reg  <= \piso.data_li [1608];
      \piso.data_r_1607_sv2v_reg  <= \piso.data_li [1607];
      \piso.data_r_1606_sv2v_reg  <= \piso.data_li [1606];
      \piso.data_r_1605_sv2v_reg  <= \piso.data_li [1605];
      \piso.data_r_1604_sv2v_reg  <= \piso.data_li [1604];
      \piso.data_r_1603_sv2v_reg  <= \piso.data_li [1603];
      \piso.data_r_1602_sv2v_reg  <= \piso.data_li [1602];
      \piso.data_r_1601_sv2v_reg  <= \piso.data_li [1601];
      \piso.data_r_1600_sv2v_reg  <= \piso.data_li [1600];
      \piso.data_r_1599_sv2v_reg  <= \piso.data_li [1599];
      \piso.data_r_1598_sv2v_reg  <= \piso.data_li [1598];
      \piso.data_r_1597_sv2v_reg  <= \piso.data_li [1597];
      \piso.data_r_1596_sv2v_reg  <= \piso.data_li [1596];
      \piso.data_r_1595_sv2v_reg  <= \piso.data_li [1595];
      \piso.data_r_1594_sv2v_reg  <= \piso.data_li [1594];
      \piso.data_r_1593_sv2v_reg  <= \piso.data_li [1593];
      \piso.data_r_1592_sv2v_reg  <= \piso.data_li [1592];
      \piso.data_r_1591_sv2v_reg  <= \piso.data_li [1591];
      \piso.data_r_1590_sv2v_reg  <= \piso.data_li [1590];
      \piso.data_r_1589_sv2v_reg  <= \piso.data_li [1589];
      \piso.data_r_1588_sv2v_reg  <= \piso.data_li [1588];
      \piso.data_r_1587_sv2v_reg  <= \piso.data_li [1587];
      \piso.data_r_1586_sv2v_reg  <= \piso.data_li [1586];
      \piso.data_r_1585_sv2v_reg  <= \piso.data_li [1585];
      \piso.data_r_1584_sv2v_reg  <= \piso.data_li [1584];
      \piso.data_r_1583_sv2v_reg  <= \piso.data_li [1583];
      \piso.data_r_1582_sv2v_reg  <= \piso.data_li [1582];
      \piso.data_r_1581_sv2v_reg  <= \piso.data_li [1581];
      \piso.data_r_1580_sv2v_reg  <= \piso.data_li [1580];
      \piso.data_r_1579_sv2v_reg  <= \piso.data_li [1579];
      \piso.data_r_1578_sv2v_reg  <= \piso.data_li [1578];
      \piso.data_r_1577_sv2v_reg  <= \piso.data_li [1577];
      \piso.data_r_1576_sv2v_reg  <= \piso.data_li [1576];
      \piso.data_r_1575_sv2v_reg  <= \piso.data_li [1575];
      \piso.data_r_1574_sv2v_reg  <= \piso.data_li [1574];
      \piso.data_r_1573_sv2v_reg  <= \piso.data_li [1573];
      \piso.data_r_1572_sv2v_reg  <= \piso.data_li [1572];
      \piso.data_r_1571_sv2v_reg  <= \piso.data_li [1571];
      \piso.data_r_1570_sv2v_reg  <= \piso.data_li [1570];
      \piso.data_r_1569_sv2v_reg  <= \piso.data_li [1569];
      \piso.data_r_1568_sv2v_reg  <= \piso.data_li [1568];
      \piso.data_r_1567_sv2v_reg  <= \piso.data_li [1567];
      \piso.data_r_1566_sv2v_reg  <= \piso.data_li [1566];
      \piso.data_r_1565_sv2v_reg  <= \piso.data_li [1565];
      \piso.data_r_1564_sv2v_reg  <= \piso.data_li [1564];
      \piso.data_r_1563_sv2v_reg  <= \piso.data_li [1563];
      \piso.data_r_1562_sv2v_reg  <= \piso.data_li [1562];
      \piso.data_r_1561_sv2v_reg  <= \piso.data_li [1561];
      \piso.data_r_1560_sv2v_reg  <= \piso.data_li [1560];
      \piso.data_r_1559_sv2v_reg  <= \piso.data_li [1559];
      \piso.data_r_1558_sv2v_reg  <= \piso.data_li [1558];
      \piso.data_r_1557_sv2v_reg  <= \piso.data_li [1557];
      \piso.data_r_1556_sv2v_reg  <= \piso.data_li [1556];
      \piso.data_r_1555_sv2v_reg  <= \piso.data_li [1555];
      \piso.data_r_1554_sv2v_reg  <= \piso.data_li [1554];
      \piso.data_r_1553_sv2v_reg  <= \piso.data_li [1553];
      \piso.data_r_1552_sv2v_reg  <= \piso.data_li [1552];
      \piso.data_r_1551_sv2v_reg  <= \piso.data_li [1551];
      \piso.data_r_1550_sv2v_reg  <= \piso.data_li [1550];
      \piso.data_r_1549_sv2v_reg  <= \piso.data_li [1549];
      \piso.data_r_1548_sv2v_reg  <= \piso.data_li [1548];
      \piso.data_r_1547_sv2v_reg  <= \piso.data_li [1547];
      \piso.data_r_1546_sv2v_reg  <= \piso.data_li [1546];
      \piso.data_r_1545_sv2v_reg  <= \piso.data_li [1545];
      \piso.data_r_1544_sv2v_reg  <= \piso.data_li [1544];
      \piso.data_r_1543_sv2v_reg  <= \piso.data_li [1543];
      \piso.data_r_1542_sv2v_reg  <= \piso.data_li [1542];
      \piso.data_r_1541_sv2v_reg  <= \piso.data_li [1541];
      \piso.data_r_1540_sv2v_reg  <= \piso.data_li [1540];
      \piso.data_r_1539_sv2v_reg  <= \piso.data_li [1539];
      \piso.data_r_1538_sv2v_reg  <= \piso.data_li [1538];
      \piso.data_r_1537_sv2v_reg  <= \piso.data_li [1537];
      \piso.data_r_1536_sv2v_reg  <= \piso.data_li [1536];
      \piso.data_r_1535_sv2v_reg  <= \piso.data_li [1535];
      \piso.data_r_1534_sv2v_reg  <= \piso.data_li [1534];
      \piso.data_r_1533_sv2v_reg  <= \piso.data_li [1533];
      \piso.data_r_1532_sv2v_reg  <= \piso.data_li [1532];
      \piso.data_r_1531_sv2v_reg  <= \piso.data_li [1531];
      \piso.data_r_1530_sv2v_reg  <= \piso.data_li [1530];
      \piso.data_r_1529_sv2v_reg  <= \piso.data_li [1529];
      \piso.data_r_1528_sv2v_reg  <= \piso.data_li [1528];
      \piso.data_r_1527_sv2v_reg  <= \piso.data_li [1527];
      \piso.data_r_1526_sv2v_reg  <= \piso.data_li [1526];
      \piso.data_r_1525_sv2v_reg  <= \piso.data_li [1525];
      \piso.data_r_1524_sv2v_reg  <= \piso.data_li [1524];
      \piso.data_r_1523_sv2v_reg  <= \piso.data_li [1523];
      \piso.data_r_1522_sv2v_reg  <= \piso.data_li [1522];
      \piso.data_r_1521_sv2v_reg  <= \piso.data_li [1521];
      \piso.data_r_1520_sv2v_reg  <= \piso.data_li [1520];
      \piso.data_r_1519_sv2v_reg  <= \piso.data_li [1519];
      \piso.data_r_1518_sv2v_reg  <= \piso.data_li [1518];
      \piso.data_r_1517_sv2v_reg  <= \piso.data_li [1517];
      \piso.data_r_1516_sv2v_reg  <= \piso.data_li [1516];
      \piso.data_r_1515_sv2v_reg  <= \piso.data_li [1515];
      \piso.data_r_1514_sv2v_reg  <= \piso.data_li [1514];
      \piso.data_r_1513_sv2v_reg  <= \piso.data_li [1513];
      \piso.data_r_1512_sv2v_reg  <= \piso.data_li [1512];
      \piso.data_r_1511_sv2v_reg  <= \piso.data_li [1511];
      \piso.data_r_1510_sv2v_reg  <= \piso.data_li [1510];
      \piso.data_r_1509_sv2v_reg  <= \piso.data_li [1509];
      \piso.data_r_1508_sv2v_reg  <= \piso.data_li [1508];
      \piso.data_r_1507_sv2v_reg  <= \piso.data_li [1507];
      \piso.data_r_1506_sv2v_reg  <= \piso.data_li [1506];
      \piso.data_r_1505_sv2v_reg  <= \piso.data_li [1505];
      \piso.data_r_1504_sv2v_reg  <= \piso.data_li [1504];
      \piso.data_r_1503_sv2v_reg  <= \piso.data_li [1503];
      \piso.data_r_1502_sv2v_reg  <= \piso.data_li [1502];
      \piso.data_r_1501_sv2v_reg  <= \piso.data_li [1501];
      \piso.data_r_1500_sv2v_reg  <= \piso.data_li [1500];
      \piso.data_r_1499_sv2v_reg  <= \piso.data_li [1499];
      \piso.data_r_1498_sv2v_reg  <= \piso.data_li [1498];
      \piso.data_r_1497_sv2v_reg  <= \piso.data_li [1497];
      \piso.data_r_1496_sv2v_reg  <= \piso.data_li [1496];
      \piso.data_r_1495_sv2v_reg  <= \piso.data_li [1495];
      \piso.data_r_1494_sv2v_reg  <= \piso.data_li [1494];
      \piso.data_r_1493_sv2v_reg  <= \piso.data_li [1493];
      \piso.data_r_1492_sv2v_reg  <= \piso.data_li [1492];
      \piso.data_r_1491_sv2v_reg  <= \piso.data_li [1491];
      \piso.data_r_1490_sv2v_reg  <= \piso.data_li [1490];
      \piso.data_r_1489_sv2v_reg  <= \piso.data_li [1489];
      \piso.data_r_1488_sv2v_reg  <= \piso.data_li [1488];
      \piso.data_r_1487_sv2v_reg  <= \piso.data_li [1487];
      \piso.data_r_1486_sv2v_reg  <= \piso.data_li [1486];
      \piso.data_r_1485_sv2v_reg  <= \piso.data_li [1485];
      \piso.data_r_1484_sv2v_reg  <= \piso.data_li [1484];
      \piso.data_r_1483_sv2v_reg  <= \piso.data_li [1483];
      \piso.data_r_1482_sv2v_reg  <= \piso.data_li [1482];
      \piso.data_r_1481_sv2v_reg  <= \piso.data_li [1481];
      \piso.data_r_1480_sv2v_reg  <= \piso.data_li [1480];
      \piso.data_r_1479_sv2v_reg  <= \piso.data_li [1479];
      \piso.data_r_1478_sv2v_reg  <= \piso.data_li [1478];
      \piso.data_r_1477_sv2v_reg  <= \piso.data_li [1477];
      \piso.data_r_1476_sv2v_reg  <= \piso.data_li [1476];
      \piso.data_r_1475_sv2v_reg  <= \piso.data_li [1475];
      \piso.data_r_1474_sv2v_reg  <= \piso.data_li [1474];
      \piso.data_r_1473_sv2v_reg  <= \piso.data_li [1473];
      \piso.data_r_1472_sv2v_reg  <= \piso.data_li [1472];
      \piso.data_r_1471_sv2v_reg  <= \piso.data_li [1471];
      \piso.data_r_1470_sv2v_reg  <= \piso.data_li [1470];
      \piso.data_r_1469_sv2v_reg  <= \piso.data_li [1469];
      \piso.data_r_1468_sv2v_reg  <= \piso.data_li [1468];
      \piso.data_r_1467_sv2v_reg  <= \piso.data_li [1467];
      \piso.data_r_1466_sv2v_reg  <= \piso.data_li [1466];
      \piso.data_r_1465_sv2v_reg  <= \piso.data_li [1465];
      \piso.data_r_1464_sv2v_reg  <= \piso.data_li [1464];
      \piso.data_r_1463_sv2v_reg  <= \piso.data_li [1463];
      \piso.data_r_1462_sv2v_reg  <= \piso.data_li [1462];
      \piso.data_r_1461_sv2v_reg  <= \piso.data_li [1461];
      \piso.data_r_1460_sv2v_reg  <= \piso.data_li [1460];
      \piso.data_r_1459_sv2v_reg  <= \piso.data_li [1459];
      \piso.data_r_1458_sv2v_reg  <= \piso.data_li [1458];
      \piso.data_r_1457_sv2v_reg  <= \piso.data_li [1457];
      \piso.data_r_1456_sv2v_reg  <= \piso.data_li [1456];
      \piso.data_r_1455_sv2v_reg  <= \piso.data_li [1455];
      \piso.data_r_1454_sv2v_reg  <= \piso.data_li [1454];
      \piso.data_r_1453_sv2v_reg  <= \piso.data_li [1453];
      \piso.data_r_1452_sv2v_reg  <= \piso.data_li [1452];
      \piso.data_r_1451_sv2v_reg  <= \piso.data_li [1451];
      \piso.data_r_1450_sv2v_reg  <= \piso.data_li [1450];
      \piso.data_r_1449_sv2v_reg  <= \piso.data_li [1449];
      \piso.data_r_1448_sv2v_reg  <= \piso.data_li [1448];
      \piso.data_r_1447_sv2v_reg  <= \piso.data_li [1447];
      \piso.data_r_1446_sv2v_reg  <= \piso.data_li [1446];
      \piso.data_r_1445_sv2v_reg  <= \piso.data_li [1445];
      \piso.data_r_1444_sv2v_reg  <= \piso.data_li [1444];
      \piso.data_r_1443_sv2v_reg  <= \piso.data_li [1443];
      \piso.data_r_1442_sv2v_reg  <= \piso.data_li [1442];
      \piso.data_r_1441_sv2v_reg  <= \piso.data_li [1441];
      \piso.data_r_1440_sv2v_reg  <= \piso.data_li [1440];
      \piso.data_r_1439_sv2v_reg  <= \piso.data_li [1439];
      \piso.data_r_1438_sv2v_reg  <= \piso.data_li [1438];
      \piso.data_r_1437_sv2v_reg  <= \piso.data_li [1437];
      \piso.data_r_1436_sv2v_reg  <= \piso.data_li [1436];
      \piso.data_r_1435_sv2v_reg  <= \piso.data_li [1435];
      \piso.data_r_1434_sv2v_reg  <= \piso.data_li [1434];
      \piso.data_r_1433_sv2v_reg  <= \piso.data_li [1433];
      \piso.data_r_1432_sv2v_reg  <= \piso.data_li [1432];
      \piso.data_r_1431_sv2v_reg  <= \piso.data_li [1431];
      \piso.data_r_1430_sv2v_reg  <= \piso.data_li [1430];
      \piso.data_r_1429_sv2v_reg  <= \piso.data_li [1429];
      \piso.data_r_1428_sv2v_reg  <= \piso.data_li [1428];
      \piso.data_r_1427_sv2v_reg  <= \piso.data_li [1427];
      \piso.data_r_1426_sv2v_reg  <= \piso.data_li [1426];
      \piso.data_r_1425_sv2v_reg  <= \piso.data_li [1425];
      \piso.data_r_1424_sv2v_reg  <= \piso.data_li [1424];
      \piso.data_r_1423_sv2v_reg  <= \piso.data_li [1423];
      \piso.data_r_1422_sv2v_reg  <= \piso.data_li [1422];
      \piso.data_r_1421_sv2v_reg  <= \piso.data_li [1421];
      \piso.data_r_1420_sv2v_reg  <= \piso.data_li [1420];
      \piso.data_r_1419_sv2v_reg  <= \piso.data_li [1419];
      \piso.data_r_1418_sv2v_reg  <= \piso.data_li [1418];
      \piso.data_r_1417_sv2v_reg  <= \piso.data_li [1417];
      \piso.data_r_1416_sv2v_reg  <= \piso.data_li [1416];
      \piso.data_r_1415_sv2v_reg  <= \piso.data_li [1415];
      \piso.data_r_1414_sv2v_reg  <= \piso.data_li [1414];
      \piso.data_r_1413_sv2v_reg  <= \piso.data_li [1413];
      \piso.data_r_1412_sv2v_reg  <= \piso.data_li [1412];
      \piso.data_r_1411_sv2v_reg  <= \piso.data_li [1411];
      \piso.data_r_1410_sv2v_reg  <= \piso.data_li [1410];
      \piso.data_r_1409_sv2v_reg  <= \piso.data_li [1409];
      \piso.data_r_1408_sv2v_reg  <= \piso.data_li [1408];
      \piso.data_r_1407_sv2v_reg  <= \piso.data_li [1407];
      \piso.data_r_1406_sv2v_reg  <= \piso.data_li [1406];
      \piso.data_r_1405_sv2v_reg  <= \piso.data_li [1405];
      \piso.data_r_1404_sv2v_reg  <= \piso.data_li [1404];
      \piso.data_r_1403_sv2v_reg  <= \piso.data_li [1403];
      \piso.data_r_1402_sv2v_reg  <= \piso.data_li [1402];
      \piso.data_r_1401_sv2v_reg  <= \piso.data_li [1401];
      \piso.data_r_1400_sv2v_reg  <= \piso.data_li [1400];
      \piso.data_r_1399_sv2v_reg  <= \piso.data_li [1399];
      \piso.data_r_1398_sv2v_reg  <= \piso.data_li [1398];
      \piso.data_r_1397_sv2v_reg  <= \piso.data_li [1397];
      \piso.data_r_1396_sv2v_reg  <= \piso.data_li [1396];
      \piso.data_r_1395_sv2v_reg  <= \piso.data_li [1395];
      \piso.data_r_1394_sv2v_reg  <= \piso.data_li [1394];
      \piso.data_r_1393_sv2v_reg  <= \piso.data_li [1393];
      \piso.data_r_1392_sv2v_reg  <= \piso.data_li [1392];
      \piso.data_r_1391_sv2v_reg  <= \piso.data_li [1391];
      \piso.data_r_1390_sv2v_reg  <= \piso.data_li [1390];
      \piso.data_r_1389_sv2v_reg  <= \piso.data_li [1389];
      \piso.data_r_1388_sv2v_reg  <= \piso.data_li [1388];
      \piso.data_r_1387_sv2v_reg  <= \piso.data_li [1387];
      \piso.data_r_1386_sv2v_reg  <= \piso.data_li [1386];
      \piso.data_r_1385_sv2v_reg  <= \piso.data_li [1385];
      \piso.data_r_1384_sv2v_reg  <= \piso.data_li [1384];
      \piso.data_r_1383_sv2v_reg  <= \piso.data_li [1383];
      \piso.data_r_1382_sv2v_reg  <= \piso.data_li [1382];
      \piso.data_r_1381_sv2v_reg  <= \piso.data_li [1381];
      \piso.data_r_1380_sv2v_reg  <= \piso.data_li [1380];
      \piso.data_r_1379_sv2v_reg  <= \piso.data_li [1379];
      \piso.data_r_1378_sv2v_reg  <= \piso.data_li [1378];
      \piso.data_r_1377_sv2v_reg  <= \piso.data_li [1377];
      \piso.data_r_1376_sv2v_reg  <= \piso.data_li [1376];
      \piso.data_r_1375_sv2v_reg  <= \piso.data_li [1375];
      \piso.data_r_1374_sv2v_reg  <= \piso.data_li [1374];
      \piso.data_r_1373_sv2v_reg  <= \piso.data_li [1373];
      \piso.data_r_1372_sv2v_reg  <= \piso.data_li [1372];
      \piso.data_r_1371_sv2v_reg  <= \piso.data_li [1371];
      \piso.data_r_1370_sv2v_reg  <= \piso.data_li [1370];
      \piso.data_r_1369_sv2v_reg  <= \piso.data_li [1369];
      \piso.data_r_1368_sv2v_reg  <= \piso.data_li [1368];
      \piso.data_r_1367_sv2v_reg  <= \piso.data_li [1367];
      \piso.data_r_1366_sv2v_reg  <= \piso.data_li [1366];
      \piso.data_r_1365_sv2v_reg  <= \piso.data_li [1365];
      \piso.data_r_1364_sv2v_reg  <= \piso.data_li [1364];
      \piso.data_r_1363_sv2v_reg  <= \piso.data_li [1363];
      \piso.data_r_1362_sv2v_reg  <= \piso.data_li [1362];
      \piso.data_r_1361_sv2v_reg  <= \piso.data_li [1361];
      \piso.data_r_1360_sv2v_reg  <= \piso.data_li [1360];
      \piso.data_r_1359_sv2v_reg  <= \piso.data_li [1359];
      \piso.data_r_1358_sv2v_reg  <= \piso.data_li [1358];
      \piso.data_r_1357_sv2v_reg  <= \piso.data_li [1357];
      \piso.data_r_1356_sv2v_reg  <= \piso.data_li [1356];
      \piso.data_r_1355_sv2v_reg  <= \piso.data_li [1355];
      \piso.data_r_1354_sv2v_reg  <= \piso.data_li [1354];
      \piso.data_r_1353_sv2v_reg  <= \piso.data_li [1353];
      \piso.data_r_1352_sv2v_reg  <= \piso.data_li [1352];
      \piso.data_r_1351_sv2v_reg  <= \piso.data_li [1351];
      \piso.data_r_1350_sv2v_reg  <= \piso.data_li [1350];
      \piso.data_r_1349_sv2v_reg  <= \piso.data_li [1349];
      \piso.data_r_1348_sv2v_reg  <= \piso.data_li [1348];
      \piso.data_r_1347_sv2v_reg  <= \piso.data_li [1347];
      \piso.data_r_1346_sv2v_reg  <= \piso.data_li [1346];
      \piso.data_r_1345_sv2v_reg  <= \piso.data_li [1345];
      \piso.data_r_1344_sv2v_reg  <= \piso.data_li [1344];
      \piso.data_r_1343_sv2v_reg  <= \piso.data_li [1343];
      \piso.data_r_1342_sv2v_reg  <= \piso.data_li [1342];
      \piso.data_r_1341_sv2v_reg  <= \piso.data_li [1341];
      \piso.data_r_1340_sv2v_reg  <= \piso.data_li [1340];
      \piso.data_r_1339_sv2v_reg  <= \piso.data_li [1339];
      \piso.data_r_1338_sv2v_reg  <= \piso.data_li [1338];
      \piso.data_r_1337_sv2v_reg  <= \piso.data_li [1337];
      \piso.data_r_1336_sv2v_reg  <= \piso.data_li [1336];
      \piso.data_r_1335_sv2v_reg  <= \piso.data_li [1335];
      \piso.data_r_1334_sv2v_reg  <= \piso.data_li [1334];
      \piso.data_r_1333_sv2v_reg  <= \piso.data_li [1333];
      \piso.data_r_1332_sv2v_reg  <= \piso.data_li [1332];
      \piso.data_r_1331_sv2v_reg  <= \piso.data_li [1331];
      \piso.data_r_1330_sv2v_reg  <= \piso.data_li [1330];
      \piso.data_r_1329_sv2v_reg  <= \piso.data_li [1329];
      \piso.data_r_1328_sv2v_reg  <= \piso.data_li [1328];
      \piso.data_r_1327_sv2v_reg  <= \piso.data_li [1327];
      \piso.data_r_1326_sv2v_reg  <= \piso.data_li [1326];
      \piso.data_r_1325_sv2v_reg  <= \piso.data_li [1325];
      \piso.data_r_1324_sv2v_reg  <= \piso.data_li [1324];
      \piso.data_r_1323_sv2v_reg  <= \piso.data_li [1323];
      \piso.data_r_1322_sv2v_reg  <= \piso.data_li [1322];
      \piso.data_r_1321_sv2v_reg  <= \piso.data_li [1321];
      \piso.data_r_1320_sv2v_reg  <= \piso.data_li [1320];
      \piso.data_r_1319_sv2v_reg  <= \piso.data_li [1319];
      \piso.data_r_1318_sv2v_reg  <= \piso.data_li [1318];
      \piso.data_r_1317_sv2v_reg  <= \piso.data_li [1317];
      \piso.data_r_1316_sv2v_reg  <= \piso.data_li [1316];
      \piso.data_r_1315_sv2v_reg  <= \piso.data_li [1315];
      \piso.data_r_1314_sv2v_reg  <= \piso.data_li [1314];
      \piso.data_r_1313_sv2v_reg  <= \piso.data_li [1313];
      \piso.data_r_1312_sv2v_reg  <= \piso.data_li [1312];
      \piso.data_r_1311_sv2v_reg  <= \piso.data_li [1311];
      \piso.data_r_1310_sv2v_reg  <= \piso.data_li [1310];
      \piso.data_r_1309_sv2v_reg  <= \piso.data_li [1309];
      \piso.data_r_1308_sv2v_reg  <= \piso.data_li [1308];
      \piso.data_r_1307_sv2v_reg  <= \piso.data_li [1307];
      \piso.data_r_1306_sv2v_reg  <= \piso.data_li [1306];
      \piso.data_r_1305_sv2v_reg  <= \piso.data_li [1305];
      \piso.data_r_1304_sv2v_reg  <= \piso.data_li [1304];
      \piso.data_r_1303_sv2v_reg  <= \piso.data_li [1303];
      \piso.data_r_1302_sv2v_reg  <= \piso.data_li [1302];
      \piso.data_r_1301_sv2v_reg  <= \piso.data_li [1301];
      \piso.data_r_1300_sv2v_reg  <= \piso.data_li [1300];
      \piso.data_r_1299_sv2v_reg  <= \piso.data_li [1299];
      \piso.data_r_1298_sv2v_reg  <= \piso.data_li [1298];
      \piso.data_r_1297_sv2v_reg  <= \piso.data_li [1297];
      \piso.data_r_1296_sv2v_reg  <= \piso.data_li [1296];
      \piso.data_r_1295_sv2v_reg  <= \piso.data_li [1295];
      \piso.data_r_1294_sv2v_reg  <= \piso.data_li [1294];
      \piso.data_r_1293_sv2v_reg  <= \piso.data_li [1293];
      \piso.data_r_1292_sv2v_reg  <= \piso.data_li [1292];
      \piso.data_r_1291_sv2v_reg  <= \piso.data_li [1291];
      \piso.data_r_1290_sv2v_reg  <= \piso.data_li [1290];
      \piso.data_r_1289_sv2v_reg  <= \piso.data_li [1289];
      \piso.data_r_1288_sv2v_reg  <= \piso.data_li [1288];
      \piso.data_r_1287_sv2v_reg  <= \piso.data_li [1287];
      \piso.data_r_1286_sv2v_reg  <= \piso.data_li [1286];
      \piso.data_r_1285_sv2v_reg  <= \piso.data_li [1285];
      \piso.data_r_1284_sv2v_reg  <= \piso.data_li [1284];
      \piso.data_r_1283_sv2v_reg  <= \piso.data_li [1283];
      \piso.data_r_1282_sv2v_reg  <= \piso.data_li [1282];
      \piso.data_r_1281_sv2v_reg  <= \piso.data_li [1281];
      \piso.data_r_1280_sv2v_reg  <= \piso.data_li [1280];
      \piso.data_r_1279_sv2v_reg  <= \piso.data_li [1279];
      \piso.data_r_1278_sv2v_reg  <= \piso.data_li [1278];
      \piso.data_r_1277_sv2v_reg  <= \piso.data_li [1277];
      \piso.data_r_1276_sv2v_reg  <= \piso.data_li [1276];
      \piso.data_r_1275_sv2v_reg  <= \piso.data_li [1275];
      \piso.data_r_1274_sv2v_reg  <= \piso.data_li [1274];
      \piso.data_r_1273_sv2v_reg  <= \piso.data_li [1273];
      \piso.data_r_1272_sv2v_reg  <= \piso.data_li [1272];
      \piso.data_r_1271_sv2v_reg  <= \piso.data_li [1271];
      \piso.data_r_1270_sv2v_reg  <= \piso.data_li [1270];
      \piso.data_r_1269_sv2v_reg  <= \piso.data_li [1269];
      \piso.data_r_1268_sv2v_reg  <= \piso.data_li [1268];
      \piso.data_r_1267_sv2v_reg  <= \piso.data_li [1267];
      \piso.data_r_1266_sv2v_reg  <= \piso.data_li [1266];
      \piso.data_r_1265_sv2v_reg  <= \piso.data_li [1265];
      \piso.data_r_1264_sv2v_reg  <= \piso.data_li [1264];
      \piso.data_r_1263_sv2v_reg  <= \piso.data_li [1263];
      \piso.data_r_1262_sv2v_reg  <= \piso.data_li [1262];
      \piso.data_r_1261_sv2v_reg  <= \piso.data_li [1261];
      \piso.data_r_1260_sv2v_reg  <= \piso.data_li [1260];
      \piso.data_r_1259_sv2v_reg  <= \piso.data_li [1259];
      \piso.data_r_1258_sv2v_reg  <= \piso.data_li [1258];
      \piso.data_r_1257_sv2v_reg  <= \piso.data_li [1257];
      \piso.data_r_1256_sv2v_reg  <= \piso.data_li [1256];
      \piso.data_r_1255_sv2v_reg  <= \piso.data_li [1255];
      \piso.data_r_1254_sv2v_reg  <= \piso.data_li [1254];
      \piso.data_r_1253_sv2v_reg  <= \piso.data_li [1253];
      \piso.data_r_1252_sv2v_reg  <= \piso.data_li [1252];
      \piso.data_r_1251_sv2v_reg  <= \piso.data_li [1251];
      \piso.data_r_1250_sv2v_reg  <= \piso.data_li [1250];
      \piso.data_r_1249_sv2v_reg  <= \piso.data_li [1249];
      \piso.data_r_1248_sv2v_reg  <= \piso.data_li [1248];
      \piso.data_r_1247_sv2v_reg  <= \piso.data_li [1247];
      \piso.data_r_1246_sv2v_reg  <= \piso.data_li [1246];
      \piso.data_r_1245_sv2v_reg  <= \piso.data_li [1245];
      \piso.data_r_1244_sv2v_reg  <= \piso.data_li [1244];
      \piso.data_r_1243_sv2v_reg  <= \piso.data_li [1243];
      \piso.data_r_1242_sv2v_reg  <= \piso.data_li [1242];
      \piso.data_r_1241_sv2v_reg  <= \piso.data_li [1241];
      \piso.data_r_1240_sv2v_reg  <= \piso.data_li [1240];
      \piso.data_r_1239_sv2v_reg  <= \piso.data_li [1239];
      \piso.data_r_1238_sv2v_reg  <= \piso.data_li [1238];
      \piso.data_r_1237_sv2v_reg  <= \piso.data_li [1237];
      \piso.data_r_1236_sv2v_reg  <= \piso.data_li [1236];
      \piso.data_r_1235_sv2v_reg  <= \piso.data_li [1235];
      \piso.data_r_1234_sv2v_reg  <= \piso.data_li [1234];
      \piso.data_r_1233_sv2v_reg  <= \piso.data_li [1233];
      \piso.data_r_1232_sv2v_reg  <= \piso.data_li [1232];
      \piso.data_r_1231_sv2v_reg  <= \piso.data_li [1231];
      \piso.data_r_1230_sv2v_reg  <= \piso.data_li [1230];
      \piso.data_r_1229_sv2v_reg  <= \piso.data_li [1229];
      \piso.data_r_1228_sv2v_reg  <= \piso.data_li [1228];
      \piso.data_r_1227_sv2v_reg  <= \piso.data_li [1227];
      \piso.data_r_1226_sv2v_reg  <= \piso.data_li [1226];
      \piso.data_r_1225_sv2v_reg  <= \piso.data_li [1225];
      \piso.data_r_1224_sv2v_reg  <= \piso.data_li [1224];
      \piso.data_r_1223_sv2v_reg  <= \piso.data_li [1223];
      \piso.data_r_1222_sv2v_reg  <= \piso.data_li [1222];
      \piso.data_r_1221_sv2v_reg  <= \piso.data_li [1221];
      \piso.data_r_1220_sv2v_reg  <= \piso.data_li [1220];
      \piso.data_r_1219_sv2v_reg  <= \piso.data_li [1219];
      \piso.data_r_1218_sv2v_reg  <= \piso.data_li [1218];
      \piso.data_r_1217_sv2v_reg  <= \piso.data_li [1217];
      \piso.data_r_1216_sv2v_reg  <= \piso.data_li [1216];
      \piso.data_r_1215_sv2v_reg  <= \piso.data_li [1215];
      \piso.data_r_1214_sv2v_reg  <= \piso.data_li [1214];
      \piso.data_r_1213_sv2v_reg  <= \piso.data_li [1213];
      \piso.data_r_1212_sv2v_reg  <= \piso.data_li [1212];
      \piso.data_r_1211_sv2v_reg  <= \piso.data_li [1211];
      \piso.data_r_1210_sv2v_reg  <= \piso.data_li [1210];
      \piso.data_r_1209_sv2v_reg  <= \piso.data_li [1209];
      \piso.data_r_1208_sv2v_reg  <= \piso.data_li [1208];
      \piso.data_r_1207_sv2v_reg  <= \piso.data_li [1207];
      \piso.data_r_1206_sv2v_reg  <= \piso.data_li [1206];
      \piso.data_r_1205_sv2v_reg  <= \piso.data_li [1205];
      \piso.data_r_1204_sv2v_reg  <= \piso.data_li [1204];
      \piso.data_r_1203_sv2v_reg  <= \piso.data_li [1203];
      \piso.data_r_1202_sv2v_reg  <= \piso.data_li [1202];
      \piso.data_r_1201_sv2v_reg  <= \piso.data_li [1201];
      \piso.data_r_1200_sv2v_reg  <= \piso.data_li [1200];
      \piso.data_r_1199_sv2v_reg  <= \piso.data_li [1199];
      \piso.data_r_1198_sv2v_reg  <= \piso.data_li [1198];
      \piso.data_r_1197_sv2v_reg  <= \piso.data_li [1197];
      \piso.data_r_1196_sv2v_reg  <= \piso.data_li [1196];
      \piso.data_r_1195_sv2v_reg  <= \piso.data_li [1195];
      \piso.data_r_1194_sv2v_reg  <= \piso.data_li [1194];
      \piso.data_r_1193_sv2v_reg  <= \piso.data_li [1193];
      \piso.data_r_1192_sv2v_reg  <= \piso.data_li [1192];
      \piso.data_r_1191_sv2v_reg  <= \piso.data_li [1191];
      \piso.data_r_1190_sv2v_reg  <= \piso.data_li [1190];
      \piso.data_r_1189_sv2v_reg  <= \piso.data_li [1189];
      \piso.data_r_1188_sv2v_reg  <= \piso.data_li [1188];
      \piso.data_r_1187_sv2v_reg  <= \piso.data_li [1187];
      \piso.data_r_1186_sv2v_reg  <= \piso.data_li [1186];
      \piso.data_r_1185_sv2v_reg  <= \piso.data_li [1185];
      \piso.data_r_1184_sv2v_reg  <= \piso.data_li [1184];
      \piso.data_r_1183_sv2v_reg  <= \piso.data_li [1183];
      \piso.data_r_1182_sv2v_reg  <= \piso.data_li [1182];
      \piso.data_r_1181_sv2v_reg  <= \piso.data_li [1181];
      \piso.data_r_1180_sv2v_reg  <= \piso.data_li [1180];
      \piso.data_r_1179_sv2v_reg  <= \piso.data_li [1179];
      \piso.data_r_1178_sv2v_reg  <= \piso.data_li [1178];
      \piso.data_r_1177_sv2v_reg  <= \piso.data_li [1177];
      \piso.data_r_1176_sv2v_reg  <= \piso.data_li [1176];
      \piso.data_r_1175_sv2v_reg  <= \piso.data_li [1175];
      \piso.data_r_1174_sv2v_reg  <= \piso.data_li [1174];
      \piso.data_r_1173_sv2v_reg  <= \piso.data_li [1173];
      \piso.data_r_1172_sv2v_reg  <= \piso.data_li [1172];
      \piso.data_r_1171_sv2v_reg  <= \piso.data_li [1171];
      \piso.data_r_1170_sv2v_reg  <= \piso.data_li [1170];
      \piso.data_r_1169_sv2v_reg  <= \piso.data_li [1169];
      \piso.data_r_1168_sv2v_reg  <= \piso.data_li [1168];
      \piso.data_r_1167_sv2v_reg  <= \piso.data_li [1167];
      \piso.data_r_1166_sv2v_reg  <= \piso.data_li [1166];
      \piso.data_r_1165_sv2v_reg  <= \piso.data_li [1165];
      \piso.data_r_1164_sv2v_reg  <= \piso.data_li [1164];
      \piso.data_r_1163_sv2v_reg  <= \piso.data_li [1163];
      \piso.data_r_1162_sv2v_reg  <= \piso.data_li [1162];
      \piso.data_r_1161_sv2v_reg  <= \piso.data_li [1161];
      \piso.data_r_1160_sv2v_reg  <= \piso.data_li [1160];
      \piso.data_r_1159_sv2v_reg  <= \piso.data_li [1159];
      \piso.data_r_1158_sv2v_reg  <= \piso.data_li [1158];
      \piso.data_r_1157_sv2v_reg  <= \piso.data_li [1157];
      \piso.data_r_1156_sv2v_reg  <= \piso.data_li [1156];
      \piso.data_r_1155_sv2v_reg  <= \piso.data_li [1155];
      \piso.data_r_1154_sv2v_reg  <= \piso.data_li [1154];
      \piso.data_r_1153_sv2v_reg  <= \piso.data_li [1153];
      \piso.data_r_1152_sv2v_reg  <= \piso.data_li [1152];
      \piso.data_r_1151_sv2v_reg  <= \piso.data_li [1151];
      \piso.data_r_1150_sv2v_reg  <= \piso.data_li [1150];
      \piso.data_r_1149_sv2v_reg  <= \piso.data_li [1149];
      \piso.data_r_1148_sv2v_reg  <= \piso.data_li [1148];
      \piso.data_r_1147_sv2v_reg  <= \piso.data_li [1147];
      \piso.data_r_1146_sv2v_reg  <= \piso.data_li [1146];
      \piso.data_r_1145_sv2v_reg  <= \piso.data_li [1145];
      \piso.data_r_1144_sv2v_reg  <= \piso.data_li [1144];
      \piso.data_r_1143_sv2v_reg  <= \piso.data_li [1143];
      \piso.data_r_1142_sv2v_reg  <= \piso.data_li [1142];
      \piso.data_r_1141_sv2v_reg  <= \piso.data_li [1141];
      \piso.data_r_1140_sv2v_reg  <= \piso.data_li [1140];
      \piso.data_r_1139_sv2v_reg  <= \piso.data_li [1139];
      \piso.data_r_1138_sv2v_reg  <= \piso.data_li [1138];
      \piso.data_r_1137_sv2v_reg  <= \piso.data_li [1137];
      \piso.data_r_1136_sv2v_reg  <= \piso.data_li [1136];
      \piso.data_r_1135_sv2v_reg  <= \piso.data_li [1135];
      \piso.data_r_1134_sv2v_reg  <= \piso.data_li [1134];
      \piso.data_r_1133_sv2v_reg  <= \piso.data_li [1133];
      \piso.data_r_1132_sv2v_reg  <= \piso.data_li [1132];
      \piso.data_r_1131_sv2v_reg  <= \piso.data_li [1131];
      \piso.data_r_1130_sv2v_reg  <= \piso.data_li [1130];
      \piso.data_r_1129_sv2v_reg  <= \piso.data_li [1129];
      \piso.data_r_1128_sv2v_reg  <= \piso.data_li [1128];
      \piso.data_r_1127_sv2v_reg  <= \piso.data_li [1127];
      \piso.data_r_1126_sv2v_reg  <= \piso.data_li [1126];
      \piso.data_r_1125_sv2v_reg  <= \piso.data_li [1125];
      \piso.data_r_1124_sv2v_reg  <= \piso.data_li [1124];
      \piso.data_r_1123_sv2v_reg  <= \piso.data_li [1123];
      \piso.data_r_1122_sv2v_reg  <= \piso.data_li [1122];
      \piso.data_r_1121_sv2v_reg  <= \piso.data_li [1121];
      \piso.data_r_1120_sv2v_reg  <= \piso.data_li [1120];
      \piso.data_r_1119_sv2v_reg  <= \piso.data_li [1119];
      \piso.data_r_1118_sv2v_reg  <= \piso.data_li [1118];
      \piso.data_r_1117_sv2v_reg  <= \piso.data_li [1117];
      \piso.data_r_1116_sv2v_reg  <= \piso.data_li [1116];
      \piso.data_r_1115_sv2v_reg  <= \piso.data_li [1115];
      \piso.data_r_1114_sv2v_reg  <= \piso.data_li [1114];
      \piso.data_r_1113_sv2v_reg  <= \piso.data_li [1113];
      \piso.data_r_1112_sv2v_reg  <= \piso.data_li [1112];
      \piso.data_r_1111_sv2v_reg  <= \piso.data_li [1111];
      \piso.data_r_1110_sv2v_reg  <= \piso.data_li [1110];
      \piso.data_r_1109_sv2v_reg  <= \piso.data_li [1109];
      \piso.data_r_1108_sv2v_reg  <= \piso.data_li [1108];
      \piso.data_r_1107_sv2v_reg  <= \piso.data_li [1107];
      \piso.data_r_1106_sv2v_reg  <= \piso.data_li [1106];
      \piso.data_r_1105_sv2v_reg  <= \piso.data_li [1105];
      \piso.data_r_1104_sv2v_reg  <= \piso.data_li [1104];
      \piso.data_r_1103_sv2v_reg  <= \piso.data_li [1103];
      \piso.data_r_1102_sv2v_reg  <= \piso.data_li [1102];
      \piso.data_r_1101_sv2v_reg  <= \piso.data_li [1101];
      \piso.data_r_1100_sv2v_reg  <= \piso.data_li [1100];
      \piso.data_r_1099_sv2v_reg  <= \piso.data_li [1099];
      \piso.data_r_1098_sv2v_reg  <= \piso.data_li [1098];
      \piso.data_r_1097_sv2v_reg  <= \piso.data_li [1097];
      \piso.data_r_1096_sv2v_reg  <= \piso.data_li [1096];
      \piso.data_r_1095_sv2v_reg  <= \piso.data_li [1095];
      \piso.data_r_1094_sv2v_reg  <= \piso.data_li [1094];
      \piso.data_r_1093_sv2v_reg  <= \piso.data_li [1093];
      \piso.data_r_1092_sv2v_reg  <= \piso.data_li [1092];
      \piso.data_r_1091_sv2v_reg  <= \piso.data_li [1091];
      \piso.data_r_1090_sv2v_reg  <= \piso.data_li [1090];
      \piso.data_r_1089_sv2v_reg  <= \piso.data_li [1089];
      \piso.data_r_1088_sv2v_reg  <= \piso.data_li [1088];
      \piso.data_r_1087_sv2v_reg  <= \piso.data_li [1087];
      \piso.data_r_1086_sv2v_reg  <= \piso.data_li [1086];
      \piso.data_r_1085_sv2v_reg  <= \piso.data_li [1085];
      \piso.data_r_1084_sv2v_reg  <= \piso.data_li [1084];
      \piso.data_r_1083_sv2v_reg  <= \piso.data_li [1083];
      \piso.data_r_1082_sv2v_reg  <= \piso.data_li [1082];
      \piso.data_r_1081_sv2v_reg  <= \piso.data_li [1081];
      \piso.data_r_1080_sv2v_reg  <= \piso.data_li [1080];
      \piso.data_r_1079_sv2v_reg  <= \piso.data_li [1079];
      \piso.data_r_1078_sv2v_reg  <= \piso.data_li [1078];
      \piso.data_r_1077_sv2v_reg  <= \piso.data_li [1077];
      \piso.data_r_1076_sv2v_reg  <= \piso.data_li [1076];
      \piso.data_r_1075_sv2v_reg  <= \piso.data_li [1075];
      \piso.data_r_1074_sv2v_reg  <= \piso.data_li [1074];
      \piso.data_r_1073_sv2v_reg  <= \piso.data_li [1073];
      \piso.data_r_1072_sv2v_reg  <= \piso.data_li [1072];
      \piso.data_r_1071_sv2v_reg  <= \piso.data_li [1071];
      \piso.data_r_1070_sv2v_reg  <= \piso.data_li [1070];
      \piso.data_r_1069_sv2v_reg  <= \piso.data_li [1069];
      \piso.data_r_1068_sv2v_reg  <= \piso.data_li [1068];
      \piso.data_r_1067_sv2v_reg  <= \piso.data_li [1067];
      \piso.data_r_1066_sv2v_reg  <= \piso.data_li [1066];
      \piso.data_r_1065_sv2v_reg  <= \piso.data_li [1065];
      \piso.data_r_1064_sv2v_reg  <= \piso.data_li [1064];
      \piso.data_r_1063_sv2v_reg  <= \piso.data_li [1063];
      \piso.data_r_1062_sv2v_reg  <= \piso.data_li [1062];
      \piso.data_r_1061_sv2v_reg  <= \piso.data_li [1061];
      \piso.data_r_1060_sv2v_reg  <= \piso.data_li [1060];
      \piso.data_r_1059_sv2v_reg  <= \piso.data_li [1059];
      \piso.data_r_1058_sv2v_reg  <= \piso.data_li [1058];
      \piso.data_r_1057_sv2v_reg  <= \piso.data_li [1057];
      \piso.data_r_1056_sv2v_reg  <= \piso.data_li [1056];
      \piso.data_r_1055_sv2v_reg  <= \piso.data_li [1055];
      \piso.data_r_1054_sv2v_reg  <= \piso.data_li [1054];
      \piso.data_r_1053_sv2v_reg  <= \piso.data_li [1053];
      \piso.data_r_1052_sv2v_reg  <= \piso.data_li [1052];
      \piso.data_r_1051_sv2v_reg  <= \piso.data_li [1051];
      \piso.data_r_1050_sv2v_reg  <= \piso.data_li [1050];
      \piso.data_r_1049_sv2v_reg  <= \piso.data_li [1049];
      \piso.data_r_1048_sv2v_reg  <= \piso.data_li [1048];
      \piso.data_r_1047_sv2v_reg  <= \piso.data_li [1047];
      \piso.data_r_1046_sv2v_reg  <= \piso.data_li [1046];
      \piso.data_r_1045_sv2v_reg  <= \piso.data_li [1045];
      \piso.data_r_1044_sv2v_reg  <= \piso.data_li [1044];
      \piso.data_r_1043_sv2v_reg  <= \piso.data_li [1043];
      \piso.data_r_1042_sv2v_reg  <= \piso.data_li [1042];
      \piso.data_r_1041_sv2v_reg  <= \piso.data_li [1041];
      \piso.data_r_1040_sv2v_reg  <= \piso.data_li [1040];
      \piso.data_r_1039_sv2v_reg  <= \piso.data_li [1039];
      \piso.data_r_1038_sv2v_reg  <= \piso.data_li [1038];
      \piso.data_r_1037_sv2v_reg  <= \piso.data_li [1037];
      \piso.data_r_1036_sv2v_reg  <= \piso.data_li [1036];
      \piso.data_r_1035_sv2v_reg  <= \piso.data_li [1035];
      \piso.data_r_1034_sv2v_reg  <= \piso.data_li [1034];
      \piso.data_r_1033_sv2v_reg  <= \piso.data_li [1033];
      \piso.data_r_1032_sv2v_reg  <= \piso.data_li [1032];
      \piso.data_r_1031_sv2v_reg  <= \piso.data_li [1031];
      \piso.data_r_1030_sv2v_reg  <= \piso.data_li [1030];
      \piso.data_r_1029_sv2v_reg  <= \piso.data_li [1029];
      \piso.data_r_1028_sv2v_reg  <= \piso.data_li [1028];
      \piso.data_r_1027_sv2v_reg  <= \piso.data_li [1027];
      \piso.data_r_1026_sv2v_reg  <= \piso.data_li [1026];
      \piso.data_r_1025_sv2v_reg  <= \piso.data_li [1025];
      \piso.data_r_1024_sv2v_reg  <= \piso.data_li [1024];
      \piso.data_r_1023_sv2v_reg  <= \piso.data_li [1023];
      \piso.data_r_1022_sv2v_reg  <= \piso.data_li [1022];
      \piso.data_r_1021_sv2v_reg  <= \piso.data_li [1021];
      \piso.data_r_1020_sv2v_reg  <= \piso.data_li [1020];
      \piso.data_r_1019_sv2v_reg  <= \piso.data_li [1019];
      \piso.data_r_1018_sv2v_reg  <= \piso.data_li [1018];
      \piso.data_r_1017_sv2v_reg  <= \piso.data_li [1017];
      \piso.data_r_1016_sv2v_reg  <= \piso.data_li [1016];
      \piso.data_r_1015_sv2v_reg  <= \piso.data_li [1015];
      \piso.data_r_1014_sv2v_reg  <= \piso.data_li [1014];
      \piso.data_r_1013_sv2v_reg  <= \piso.data_li [1013];
      \piso.data_r_1012_sv2v_reg  <= \piso.data_li [1012];
      \piso.data_r_1011_sv2v_reg  <= \piso.data_li [1011];
      \piso.data_r_1010_sv2v_reg  <= \piso.data_li [1010];
      \piso.data_r_1009_sv2v_reg  <= \piso.data_li [1009];
      \piso.data_r_1008_sv2v_reg  <= \piso.data_li [1008];
      \piso.data_r_1007_sv2v_reg  <= \piso.data_li [1007];
      \piso.data_r_1006_sv2v_reg  <= \piso.data_li [1006];
      \piso.data_r_1005_sv2v_reg  <= \piso.data_li [1005];
      \piso.data_r_1004_sv2v_reg  <= \piso.data_li [1004];
      \piso.data_r_1003_sv2v_reg  <= \piso.data_li [1003];
      \piso.data_r_1002_sv2v_reg  <= \piso.data_li [1002];
      \piso.data_r_1001_sv2v_reg  <= \piso.data_li [1001];
      \piso.data_r_1000_sv2v_reg  <= \piso.data_li [1000];
      \piso.data_r_999_sv2v_reg  <= \piso.data_li [999];
      \piso.data_r_998_sv2v_reg  <= \piso.data_li [998];
      \piso.data_r_997_sv2v_reg  <= \piso.data_li [997];
      \piso.data_r_996_sv2v_reg  <= \piso.data_li [996];
      \piso.data_r_995_sv2v_reg  <= \piso.data_li [995];
      \piso.data_r_994_sv2v_reg  <= \piso.data_li [994];
      \piso.data_r_993_sv2v_reg  <= \piso.data_li [993];
      \piso.data_r_992_sv2v_reg  <= \piso.data_li [992];
      \piso.data_r_991_sv2v_reg  <= \piso.data_li [991];
      \piso.data_r_990_sv2v_reg  <= \piso.data_li [990];
      \piso.data_r_989_sv2v_reg  <= \piso.data_li [989];
      \piso.data_r_988_sv2v_reg  <= \piso.data_li [988];
      \piso.data_r_987_sv2v_reg  <= \piso.data_li [987];
      \piso.data_r_986_sv2v_reg  <= \piso.data_li [986];
      \piso.data_r_985_sv2v_reg  <= \piso.data_li [985];
      \piso.data_r_984_sv2v_reg  <= \piso.data_li [984];
      \piso.data_r_983_sv2v_reg  <= \piso.data_li [983];
      \piso.data_r_982_sv2v_reg  <= \piso.data_li [982];
      \piso.data_r_981_sv2v_reg  <= \piso.data_li [981];
      \piso.data_r_980_sv2v_reg  <= \piso.data_li [980];
      \piso.data_r_979_sv2v_reg  <= \piso.data_li [979];
      \piso.data_r_978_sv2v_reg  <= \piso.data_li [978];
      \piso.data_r_977_sv2v_reg  <= \piso.data_li [977];
      \piso.data_r_976_sv2v_reg  <= \piso.data_li [976];
      \piso.data_r_975_sv2v_reg  <= \piso.data_li [975];
      \piso.data_r_974_sv2v_reg  <= \piso.data_li [974];
      \piso.data_r_973_sv2v_reg  <= \piso.data_li [973];
      \piso.data_r_972_sv2v_reg  <= \piso.data_li [972];
      \piso.data_r_971_sv2v_reg  <= \piso.data_li [971];
      \piso.data_r_970_sv2v_reg  <= \piso.data_li [970];
      \piso.data_r_969_sv2v_reg  <= \piso.data_li [969];
      \piso.data_r_968_sv2v_reg  <= \piso.data_li [968];
      \piso.data_r_967_sv2v_reg  <= \piso.data_li [967];
      \piso.data_r_966_sv2v_reg  <= \piso.data_li [966];
      \piso.data_r_965_sv2v_reg  <= \piso.data_li [965];
      \piso.data_r_964_sv2v_reg  <= \piso.data_li [964];
      \piso.data_r_963_sv2v_reg  <= \piso.data_li [963];
      \piso.data_r_962_sv2v_reg  <= \piso.data_li [962];
      \piso.data_r_961_sv2v_reg  <= \piso.data_li [961];
      \piso.data_r_960_sv2v_reg  <= \piso.data_li [960];
      \piso.data_r_959_sv2v_reg  <= \piso.data_li [959];
      \piso.data_r_958_sv2v_reg  <= \piso.data_li [958];
      \piso.data_r_957_sv2v_reg  <= \piso.data_li [957];
      \piso.data_r_956_sv2v_reg  <= \piso.data_li [956];
      \piso.data_r_955_sv2v_reg  <= \piso.data_li [955];
      \piso.data_r_954_sv2v_reg  <= \piso.data_li [954];
      \piso.data_r_953_sv2v_reg  <= \piso.data_li [953];
      \piso.data_r_952_sv2v_reg  <= \piso.data_li [952];
      \piso.data_r_951_sv2v_reg  <= \piso.data_li [951];
      \piso.data_r_950_sv2v_reg  <= \piso.data_li [950];
      \piso.data_r_949_sv2v_reg  <= \piso.data_li [949];
      \piso.data_r_948_sv2v_reg  <= \piso.data_li [948];
      \piso.data_r_947_sv2v_reg  <= \piso.data_li [947];
      \piso.data_r_946_sv2v_reg  <= \piso.data_li [946];
      \piso.data_r_945_sv2v_reg  <= \piso.data_li [945];
      \piso.data_r_944_sv2v_reg  <= \piso.data_li [944];
      \piso.data_r_943_sv2v_reg  <= \piso.data_li [943];
      \piso.data_r_942_sv2v_reg  <= \piso.data_li [942];
      \piso.data_r_941_sv2v_reg  <= \piso.data_li [941];
      \piso.data_r_940_sv2v_reg  <= \piso.data_li [940];
      \piso.data_r_939_sv2v_reg  <= \piso.data_li [939];
      \piso.data_r_938_sv2v_reg  <= \piso.data_li [938];
      \piso.data_r_937_sv2v_reg  <= \piso.data_li [937];
      \piso.data_r_936_sv2v_reg  <= \piso.data_li [936];
      \piso.data_r_935_sv2v_reg  <= \piso.data_li [935];
      \piso.data_r_934_sv2v_reg  <= \piso.data_li [934];
      \piso.data_r_933_sv2v_reg  <= \piso.data_li [933];
      \piso.data_r_932_sv2v_reg  <= \piso.data_li [932];
      \piso.data_r_931_sv2v_reg  <= \piso.data_li [931];
      \piso.data_r_930_sv2v_reg  <= \piso.data_li [930];
      \piso.data_r_929_sv2v_reg  <= \piso.data_li [929];
      \piso.data_r_928_sv2v_reg  <= \piso.data_li [928];
      \piso.data_r_927_sv2v_reg  <= \piso.data_li [927];
      \piso.data_r_926_sv2v_reg  <= \piso.data_li [926];
      \piso.data_r_925_sv2v_reg  <= \piso.data_li [925];
      \piso.data_r_924_sv2v_reg  <= \piso.data_li [924];
      \piso.data_r_923_sv2v_reg  <= \piso.data_li [923];
      \piso.data_r_922_sv2v_reg  <= \piso.data_li [922];
      \piso.data_r_921_sv2v_reg  <= \piso.data_li [921];
      \piso.data_r_920_sv2v_reg  <= \piso.data_li [920];
      \piso.data_r_919_sv2v_reg  <= \piso.data_li [919];
      \piso.data_r_918_sv2v_reg  <= \piso.data_li [918];
      \piso.data_r_917_sv2v_reg  <= \piso.data_li [917];
      \piso.data_r_916_sv2v_reg  <= \piso.data_li [916];
      \piso.data_r_915_sv2v_reg  <= \piso.data_li [915];
      \piso.data_r_914_sv2v_reg  <= \piso.data_li [914];
      \piso.data_r_913_sv2v_reg  <= \piso.data_li [913];
      \piso.data_r_912_sv2v_reg  <= \piso.data_li [912];
      \piso.data_r_911_sv2v_reg  <= \piso.data_li [911];
      \piso.data_r_910_sv2v_reg  <= \piso.data_li [910];
      \piso.data_r_909_sv2v_reg  <= \piso.data_li [909];
      \piso.data_r_908_sv2v_reg  <= \piso.data_li [908];
      \piso.data_r_907_sv2v_reg  <= \piso.data_li [907];
      \piso.data_r_906_sv2v_reg  <= \piso.data_li [906];
      \piso.data_r_905_sv2v_reg  <= \piso.data_li [905];
      \piso.data_r_904_sv2v_reg  <= \piso.data_li [904];
      \piso.data_r_903_sv2v_reg  <= \piso.data_li [903];
      \piso.data_r_902_sv2v_reg  <= \piso.data_li [902];
      \piso.data_r_901_sv2v_reg  <= \piso.data_li [901];
      \piso.data_r_900_sv2v_reg  <= \piso.data_li [900];
      \piso.data_r_899_sv2v_reg  <= \piso.data_li [899];
      \piso.data_r_898_sv2v_reg  <= \piso.data_li [898];
      \piso.data_r_897_sv2v_reg  <= \piso.data_li [897];
      \piso.data_r_896_sv2v_reg  <= \piso.data_li [896];
      \piso.data_r_895_sv2v_reg  <= \piso.data_li [895];
      \piso.data_r_894_sv2v_reg  <= \piso.data_li [894];
      \piso.data_r_893_sv2v_reg  <= \piso.data_li [893];
      \piso.data_r_892_sv2v_reg  <= \piso.data_li [892];
      \piso.data_r_891_sv2v_reg  <= \piso.data_li [891];
      \piso.data_r_890_sv2v_reg  <= \piso.data_li [890];
      \piso.data_r_889_sv2v_reg  <= \piso.data_li [889];
      \piso.data_r_888_sv2v_reg  <= \piso.data_li [888];
      \piso.data_r_887_sv2v_reg  <= \piso.data_li [887];
      \piso.data_r_886_sv2v_reg  <= \piso.data_li [886];
      \piso.data_r_885_sv2v_reg  <= \piso.data_li [885];
      \piso.data_r_884_sv2v_reg  <= \piso.data_li [884];
      \piso.data_r_883_sv2v_reg  <= \piso.data_li [883];
      \piso.data_r_882_sv2v_reg  <= \piso.data_li [882];
      \piso.data_r_881_sv2v_reg  <= \piso.data_li [881];
      \piso.data_r_880_sv2v_reg  <= \piso.data_li [880];
      \piso.data_r_879_sv2v_reg  <= \piso.data_li [879];
      \piso.data_r_878_sv2v_reg  <= \piso.data_li [878];
      \piso.data_r_877_sv2v_reg  <= \piso.data_li [877];
      \piso.data_r_876_sv2v_reg  <= \piso.data_li [876];
      \piso.data_r_875_sv2v_reg  <= \piso.data_li [875];
      \piso.data_r_874_sv2v_reg  <= \piso.data_li [874];
      \piso.data_r_873_sv2v_reg  <= \piso.data_li [873];
      \piso.data_r_872_sv2v_reg  <= \piso.data_li [872];
      \piso.data_r_871_sv2v_reg  <= \piso.data_li [871];
      \piso.data_r_870_sv2v_reg  <= \piso.data_li [870];
      \piso.data_r_869_sv2v_reg  <= \piso.data_li [869];
      \piso.data_r_868_sv2v_reg  <= \piso.data_li [868];
      \piso.data_r_867_sv2v_reg  <= \piso.data_li [867];
      \piso.data_r_866_sv2v_reg  <= \piso.data_li [866];
      \piso.data_r_865_sv2v_reg  <= \piso.data_li [865];
      \piso.data_r_864_sv2v_reg  <= \piso.data_li [864];
      \piso.data_r_863_sv2v_reg  <= \piso.data_li [863];
      \piso.data_r_862_sv2v_reg  <= \piso.data_li [862];
      \piso.data_r_861_sv2v_reg  <= \piso.data_li [861];
      \piso.data_r_860_sv2v_reg  <= \piso.data_li [860];
      \piso.data_r_859_sv2v_reg  <= \piso.data_li [859];
      \piso.data_r_858_sv2v_reg  <= \piso.data_li [858];
      \piso.data_r_857_sv2v_reg  <= \piso.data_li [857];
      \piso.data_r_856_sv2v_reg  <= \piso.data_li [856];
      \piso.data_r_855_sv2v_reg  <= \piso.data_li [855];
      \piso.data_r_854_sv2v_reg  <= \piso.data_li [854];
      \piso.data_r_853_sv2v_reg  <= \piso.data_li [853];
      \piso.data_r_852_sv2v_reg  <= \piso.data_li [852];
      \piso.data_r_851_sv2v_reg  <= \piso.data_li [851];
      \piso.data_r_850_sv2v_reg  <= \piso.data_li [850];
      \piso.data_r_849_sv2v_reg  <= \piso.data_li [849];
      \piso.data_r_848_sv2v_reg  <= \piso.data_li [848];
      \piso.data_r_847_sv2v_reg  <= \piso.data_li [847];
      \piso.data_r_846_sv2v_reg  <= \piso.data_li [846];
      \piso.data_r_845_sv2v_reg  <= \piso.data_li [845];
      \piso.data_r_844_sv2v_reg  <= \piso.data_li [844];
      \piso.data_r_843_sv2v_reg  <= \piso.data_li [843];
      \piso.data_r_842_sv2v_reg  <= \piso.data_li [842];
      \piso.data_r_841_sv2v_reg  <= \piso.data_li [841];
      \piso.data_r_840_sv2v_reg  <= \piso.data_li [840];
      \piso.data_r_839_sv2v_reg  <= \piso.data_li [839];
      \piso.data_r_838_sv2v_reg  <= \piso.data_li [838];
      \piso.data_r_837_sv2v_reg  <= \piso.data_li [837];
      \piso.data_r_836_sv2v_reg  <= \piso.data_li [836];
      \piso.data_r_835_sv2v_reg  <= \piso.data_li [835];
      \piso.data_r_834_sv2v_reg  <= \piso.data_li [834];
      \piso.data_r_833_sv2v_reg  <= \piso.data_li [833];
      \piso.data_r_832_sv2v_reg  <= \piso.data_li [832];
      \piso.data_r_831_sv2v_reg  <= \piso.data_li [831];
      \piso.data_r_830_sv2v_reg  <= \piso.data_li [830];
      \piso.data_r_829_sv2v_reg  <= \piso.data_li [829];
      \piso.data_r_828_sv2v_reg  <= \piso.data_li [828];
      \piso.data_r_827_sv2v_reg  <= \piso.data_li [827];
      \piso.data_r_826_sv2v_reg  <= \piso.data_li [826];
      \piso.data_r_825_sv2v_reg  <= \piso.data_li [825];
      \piso.data_r_824_sv2v_reg  <= \piso.data_li [824];
      \piso.data_r_823_sv2v_reg  <= \piso.data_li [823];
      \piso.data_r_822_sv2v_reg  <= \piso.data_li [822];
      \piso.data_r_821_sv2v_reg  <= \piso.data_li [821];
      \piso.data_r_820_sv2v_reg  <= \piso.data_li [820];
      \piso.data_r_819_sv2v_reg  <= \piso.data_li [819];
      \piso.data_r_818_sv2v_reg  <= \piso.data_li [818];
      \piso.data_r_817_sv2v_reg  <= \piso.data_li [817];
      \piso.data_r_816_sv2v_reg  <= \piso.data_li [816];
      \piso.data_r_815_sv2v_reg  <= \piso.data_li [815];
      \piso.data_r_814_sv2v_reg  <= \piso.data_li [814];
      \piso.data_r_813_sv2v_reg  <= \piso.data_li [813];
      \piso.data_r_812_sv2v_reg  <= \piso.data_li [812];
      \piso.data_r_811_sv2v_reg  <= \piso.data_li [811];
      \piso.data_r_810_sv2v_reg  <= \piso.data_li [810];
      \piso.data_r_809_sv2v_reg  <= \piso.data_li [809];
      \piso.data_r_808_sv2v_reg  <= \piso.data_li [808];
      \piso.data_r_807_sv2v_reg  <= \piso.data_li [807];
      \piso.data_r_806_sv2v_reg  <= \piso.data_li [806];
      \piso.data_r_805_sv2v_reg  <= \piso.data_li [805];
      \piso.data_r_804_sv2v_reg  <= \piso.data_li [804];
      \piso.data_r_803_sv2v_reg  <= \piso.data_li [803];
      \piso.data_r_802_sv2v_reg  <= \piso.data_li [802];
      \piso.data_r_801_sv2v_reg  <= \piso.data_li [801];
      \piso.data_r_800_sv2v_reg  <= \piso.data_li [800];
      \piso.data_r_799_sv2v_reg  <= \piso.data_li [799];
      \piso.data_r_798_sv2v_reg  <= \piso.data_li [798];
      \piso.data_r_797_sv2v_reg  <= \piso.data_li [797];
      \piso.data_r_796_sv2v_reg  <= \piso.data_li [796];
      \piso.data_r_795_sv2v_reg  <= \piso.data_li [795];
      \piso.data_r_794_sv2v_reg  <= \piso.data_li [794];
      \piso.data_r_793_sv2v_reg  <= \piso.data_li [793];
      \piso.data_r_792_sv2v_reg  <= \piso.data_li [792];
      \piso.data_r_791_sv2v_reg  <= \piso.data_li [791];
      \piso.data_r_790_sv2v_reg  <= \piso.data_li [790];
      \piso.data_r_789_sv2v_reg  <= \piso.data_li [789];
      \piso.data_r_788_sv2v_reg  <= \piso.data_li [788];
      \piso.data_r_787_sv2v_reg  <= \piso.data_li [787];
      \piso.data_r_786_sv2v_reg  <= \piso.data_li [786];
      \piso.data_r_785_sv2v_reg  <= \piso.data_li [785];
      \piso.data_r_784_sv2v_reg  <= \piso.data_li [784];
      \piso.data_r_783_sv2v_reg  <= \piso.data_li [783];
      \piso.data_r_782_sv2v_reg  <= \piso.data_li [782];
      \piso.data_r_781_sv2v_reg  <= \piso.data_li [781];
      \piso.data_r_780_sv2v_reg  <= \piso.data_li [780];
      \piso.data_r_779_sv2v_reg  <= \piso.data_li [779];
      \piso.data_r_778_sv2v_reg  <= \piso.data_li [778];
      \piso.data_r_777_sv2v_reg  <= \piso.data_li [777];
      \piso.data_r_776_sv2v_reg  <= \piso.data_li [776];
      \piso.data_r_775_sv2v_reg  <= \piso.data_li [775];
      \piso.data_r_774_sv2v_reg  <= \piso.data_li [774];
      \piso.data_r_773_sv2v_reg  <= \piso.data_li [773];
      \piso.data_r_772_sv2v_reg  <= \piso.data_li [772];
      \piso.data_r_771_sv2v_reg  <= \piso.data_li [771];
      \piso.data_r_770_sv2v_reg  <= \piso.data_li [770];
      \piso.data_r_769_sv2v_reg  <= \piso.data_li [769];
      \piso.data_r_768_sv2v_reg  <= \piso.data_li [768];
      \piso.data_r_767_sv2v_reg  <= \piso.data_li [767];
      \piso.data_r_766_sv2v_reg  <= \piso.data_li [766];
      \piso.data_r_765_sv2v_reg  <= \piso.data_li [765];
      \piso.data_r_764_sv2v_reg  <= \piso.data_li [764];
      \piso.data_r_763_sv2v_reg  <= \piso.data_li [763];
      \piso.data_r_762_sv2v_reg  <= \piso.data_li [762];
      \piso.data_r_761_sv2v_reg  <= \piso.data_li [761];
      \piso.data_r_760_sv2v_reg  <= \piso.data_li [760];
      \piso.data_r_759_sv2v_reg  <= \piso.data_li [759];
      \piso.data_r_758_sv2v_reg  <= \piso.data_li [758];
      \piso.data_r_757_sv2v_reg  <= \piso.data_li [757];
      \piso.data_r_756_sv2v_reg  <= \piso.data_li [756];
      \piso.data_r_755_sv2v_reg  <= \piso.data_li [755];
      \piso.data_r_754_sv2v_reg  <= \piso.data_li [754];
      \piso.data_r_753_sv2v_reg  <= \piso.data_li [753];
      \piso.data_r_752_sv2v_reg  <= \piso.data_li [752];
      \piso.data_r_751_sv2v_reg  <= \piso.data_li [751];
      \piso.data_r_750_sv2v_reg  <= \piso.data_li [750];
      \piso.data_r_749_sv2v_reg  <= \piso.data_li [749];
      \piso.data_r_748_sv2v_reg  <= \piso.data_li [748];
      \piso.data_r_747_sv2v_reg  <= \piso.data_li [747];
      \piso.data_r_746_sv2v_reg  <= \piso.data_li [746];
      \piso.data_r_745_sv2v_reg  <= \piso.data_li [745];
      \piso.data_r_744_sv2v_reg  <= \piso.data_li [744];
      \piso.data_r_743_sv2v_reg  <= \piso.data_li [743];
      \piso.data_r_742_sv2v_reg  <= \piso.data_li [742];
      \piso.data_r_741_sv2v_reg  <= \piso.data_li [741];
      \piso.data_r_740_sv2v_reg  <= \piso.data_li [740];
      \piso.data_r_739_sv2v_reg  <= \piso.data_li [739];
      \piso.data_r_738_sv2v_reg  <= \piso.data_li [738];
      \piso.data_r_737_sv2v_reg  <= \piso.data_li [737];
      \piso.data_r_736_sv2v_reg  <= \piso.data_li [736];
      \piso.data_r_735_sv2v_reg  <= \piso.data_li [735];
      \piso.data_r_734_sv2v_reg  <= \piso.data_li [734];
      \piso.data_r_733_sv2v_reg  <= \piso.data_li [733];
      \piso.data_r_732_sv2v_reg  <= \piso.data_li [732];
      \piso.data_r_731_sv2v_reg  <= \piso.data_li [731];
      \piso.data_r_730_sv2v_reg  <= \piso.data_li [730];
      \piso.data_r_729_sv2v_reg  <= \piso.data_li [729];
      \piso.data_r_728_sv2v_reg  <= \piso.data_li [728];
      \piso.data_r_727_sv2v_reg  <= \piso.data_li [727];
      \piso.data_r_726_sv2v_reg  <= \piso.data_li [726];
      \piso.data_r_725_sv2v_reg  <= \piso.data_li [725];
      \piso.data_r_724_sv2v_reg  <= \piso.data_li [724];
      \piso.data_r_723_sv2v_reg  <= \piso.data_li [723];
      \piso.data_r_722_sv2v_reg  <= \piso.data_li [722];
      \piso.data_r_721_sv2v_reg  <= \piso.data_li [721];
      \piso.data_r_720_sv2v_reg  <= \piso.data_li [720];
      \piso.data_r_719_sv2v_reg  <= \piso.data_li [719];
      \piso.data_r_718_sv2v_reg  <= \piso.data_li [718];
      \piso.data_r_717_sv2v_reg  <= \piso.data_li [717];
      \piso.data_r_716_sv2v_reg  <= \piso.data_li [716];
      \piso.data_r_715_sv2v_reg  <= \piso.data_li [715];
      \piso.data_r_714_sv2v_reg  <= \piso.data_li [714];
      \piso.data_r_713_sv2v_reg  <= \piso.data_li [713];
      \piso.data_r_712_sv2v_reg  <= \piso.data_li [712];
      \piso.data_r_711_sv2v_reg  <= \piso.data_li [711];
      \piso.data_r_710_sv2v_reg  <= \piso.data_li [710];
      \piso.data_r_709_sv2v_reg  <= \piso.data_li [709];
      \piso.data_r_708_sv2v_reg  <= \piso.data_li [708];
      \piso.data_r_707_sv2v_reg  <= \piso.data_li [707];
      \piso.data_r_706_sv2v_reg  <= \piso.data_li [706];
      \piso.data_r_705_sv2v_reg  <= \piso.data_li [705];
      \piso.data_r_704_sv2v_reg  <= \piso.data_li [704];
      \piso.data_r_703_sv2v_reg  <= \piso.data_li [703];
      \piso.data_r_702_sv2v_reg  <= \piso.data_li [702];
      \piso.data_r_701_sv2v_reg  <= \piso.data_li [701];
      \piso.data_r_700_sv2v_reg  <= \piso.data_li [700];
      \piso.data_r_699_sv2v_reg  <= \piso.data_li [699];
      \piso.data_r_698_sv2v_reg  <= \piso.data_li [698];
      \piso.data_r_697_sv2v_reg  <= \piso.data_li [697];
      \piso.data_r_696_sv2v_reg  <= \piso.data_li [696];
      \piso.data_r_695_sv2v_reg  <= \piso.data_li [695];
      \piso.data_r_694_sv2v_reg  <= \piso.data_li [694];
      \piso.data_r_693_sv2v_reg  <= \piso.data_li [693];
      \piso.data_r_692_sv2v_reg  <= \piso.data_li [692];
      \piso.data_r_691_sv2v_reg  <= \piso.data_li [691];
      \piso.data_r_690_sv2v_reg  <= \piso.data_li [690];
      \piso.data_r_689_sv2v_reg  <= \piso.data_li [689];
      \piso.data_r_688_sv2v_reg  <= \piso.data_li [688];
      \piso.data_r_687_sv2v_reg  <= \piso.data_li [687];
      \piso.data_r_686_sv2v_reg  <= \piso.data_li [686];
      \piso.data_r_685_sv2v_reg  <= \piso.data_li [685];
      \piso.data_r_684_sv2v_reg  <= \piso.data_li [684];
      \piso.data_r_683_sv2v_reg  <= \piso.data_li [683];
      \piso.data_r_682_sv2v_reg  <= \piso.data_li [682];
      \piso.data_r_681_sv2v_reg  <= \piso.data_li [681];
      \piso.data_r_680_sv2v_reg  <= \piso.data_li [680];
      \piso.data_r_679_sv2v_reg  <= \piso.data_li [679];
      \piso.data_r_678_sv2v_reg  <= \piso.data_li [678];
      \piso.data_r_677_sv2v_reg  <= \piso.data_li [677];
      \piso.data_r_676_sv2v_reg  <= \piso.data_li [676];
      \piso.data_r_675_sv2v_reg  <= \piso.data_li [675];
      \piso.data_r_674_sv2v_reg  <= \piso.data_li [674];
      \piso.data_r_673_sv2v_reg  <= \piso.data_li [673];
      \piso.data_r_672_sv2v_reg  <= \piso.data_li [672];
      \piso.data_r_671_sv2v_reg  <= \piso.data_li [671];
      \piso.data_r_670_sv2v_reg  <= \piso.data_li [670];
      \piso.data_r_669_sv2v_reg  <= \piso.data_li [669];
      \piso.data_r_668_sv2v_reg  <= \piso.data_li [668];
      \piso.data_r_667_sv2v_reg  <= \piso.data_li [667];
      \piso.data_r_666_sv2v_reg  <= \piso.data_li [666];
      \piso.data_r_665_sv2v_reg  <= \piso.data_li [665];
      \piso.data_r_664_sv2v_reg  <= \piso.data_li [664];
      \piso.data_r_663_sv2v_reg  <= \piso.data_li [663];
      \piso.data_r_662_sv2v_reg  <= \piso.data_li [662];
      \piso.data_r_661_sv2v_reg  <= \piso.data_li [661];
      \piso.data_r_660_sv2v_reg  <= \piso.data_li [660];
      \piso.data_r_659_sv2v_reg  <= \piso.data_li [659];
      \piso.data_r_658_sv2v_reg  <= \piso.data_li [658];
      \piso.data_r_657_sv2v_reg  <= \piso.data_li [657];
      \piso.data_r_656_sv2v_reg  <= \piso.data_li [656];
      \piso.data_r_655_sv2v_reg  <= \piso.data_li [655];
      \piso.data_r_654_sv2v_reg  <= \piso.data_li [654];
      \piso.data_r_653_sv2v_reg  <= \piso.data_li [653];
      \piso.data_r_652_sv2v_reg  <= \piso.data_li [652];
      \piso.data_r_651_sv2v_reg  <= \piso.data_li [651];
      \piso.data_r_650_sv2v_reg  <= \piso.data_li [650];
      \piso.data_r_649_sv2v_reg  <= \piso.data_li [649];
      \piso.data_r_648_sv2v_reg  <= \piso.data_li [648];
      \piso.data_r_647_sv2v_reg  <= \piso.data_li [647];
      \piso.data_r_646_sv2v_reg  <= \piso.data_li [646];
      \piso.data_r_645_sv2v_reg  <= \piso.data_li [645];
      \piso.data_r_644_sv2v_reg  <= \piso.data_li [644];
      \piso.data_r_643_sv2v_reg  <= \piso.data_li [643];
      \piso.data_r_642_sv2v_reg  <= \piso.data_li [642];
      \piso.data_r_641_sv2v_reg  <= \piso.data_li [641];
      \piso.data_r_640_sv2v_reg  <= \piso.data_li [640];
      \piso.data_r_639_sv2v_reg  <= \piso.data_li [639];
      \piso.data_r_638_sv2v_reg  <= \piso.data_li [638];
      \piso.data_r_637_sv2v_reg  <= \piso.data_li [637];
      \piso.data_r_636_sv2v_reg  <= \piso.data_li [636];
      \piso.data_r_635_sv2v_reg  <= \piso.data_li [635];
      \piso.data_r_634_sv2v_reg  <= \piso.data_li [634];
      \piso.data_r_633_sv2v_reg  <= \piso.data_li [633];
      \piso.data_r_632_sv2v_reg  <= \piso.data_li [632];
      \piso.data_r_631_sv2v_reg  <= \piso.data_li [631];
      \piso.data_r_630_sv2v_reg  <= \piso.data_li [630];
      \piso.data_r_629_sv2v_reg  <= \piso.data_li [629];
      \piso.data_r_628_sv2v_reg  <= \piso.data_li [628];
      \piso.data_r_627_sv2v_reg  <= \piso.data_li [627];
      \piso.data_r_626_sv2v_reg  <= \piso.data_li [626];
      \piso.data_r_625_sv2v_reg  <= \piso.data_li [625];
      \piso.data_r_624_sv2v_reg  <= \piso.data_li [624];
      \piso.data_r_623_sv2v_reg  <= \piso.data_li [623];
      \piso.data_r_622_sv2v_reg  <= \piso.data_li [622];
      \piso.data_r_621_sv2v_reg  <= \piso.data_li [621];
      \piso.data_r_620_sv2v_reg  <= \piso.data_li [620];
      \piso.data_r_619_sv2v_reg  <= \piso.data_li [619];
      \piso.data_r_618_sv2v_reg  <= \piso.data_li [618];
      \piso.data_r_617_sv2v_reg  <= \piso.data_li [617];
      \piso.data_r_616_sv2v_reg  <= \piso.data_li [616];
      \piso.data_r_615_sv2v_reg  <= \piso.data_li [615];
      \piso.data_r_614_sv2v_reg  <= \piso.data_li [614];
      \piso.data_r_613_sv2v_reg  <= \piso.data_li [613];
      \piso.data_r_612_sv2v_reg  <= \piso.data_li [612];
      \piso.data_r_611_sv2v_reg  <= \piso.data_li [611];
      \piso.data_r_610_sv2v_reg  <= \piso.data_li [610];
      \piso.data_r_609_sv2v_reg  <= \piso.data_li [609];
      \piso.data_r_608_sv2v_reg  <= \piso.data_li [608];
      \piso.data_r_607_sv2v_reg  <= \piso.data_li [607];
      \piso.data_r_606_sv2v_reg  <= \piso.data_li [606];
      \piso.data_r_605_sv2v_reg  <= \piso.data_li [605];
      \piso.data_r_604_sv2v_reg  <= \piso.data_li [604];
      \piso.data_r_603_sv2v_reg  <= \piso.data_li [603];
      \piso.data_r_602_sv2v_reg  <= \piso.data_li [602];
      \piso.data_r_601_sv2v_reg  <= \piso.data_li [601];
      \piso.data_r_600_sv2v_reg  <= \piso.data_li [600];
      \piso.data_r_599_sv2v_reg  <= \piso.data_li [599];
      \piso.data_r_598_sv2v_reg  <= \piso.data_li [598];
      \piso.data_r_597_sv2v_reg  <= \piso.data_li [597];
      \piso.data_r_596_sv2v_reg  <= \piso.data_li [596];
      \piso.data_r_595_sv2v_reg  <= \piso.data_li [595];
      \piso.data_r_594_sv2v_reg  <= \piso.data_li [594];
      \piso.data_r_593_sv2v_reg  <= \piso.data_li [593];
      \piso.data_r_592_sv2v_reg  <= \piso.data_li [592];
      \piso.data_r_591_sv2v_reg  <= \piso.data_li [591];
      \piso.data_r_590_sv2v_reg  <= \piso.data_li [590];
      \piso.data_r_589_sv2v_reg  <= \piso.data_li [589];
      \piso.data_r_588_sv2v_reg  <= \piso.data_li [588];
      \piso.data_r_587_sv2v_reg  <= \piso.data_li [587];
      \piso.data_r_586_sv2v_reg  <= \piso.data_li [586];
      \piso.data_r_585_sv2v_reg  <= \piso.data_li [585];
      \piso.data_r_584_sv2v_reg  <= \piso.data_li [584];
      \piso.data_r_583_sv2v_reg  <= \piso.data_li [583];
      \piso.data_r_582_sv2v_reg  <= \piso.data_li [582];
      \piso.data_r_581_sv2v_reg  <= \piso.data_li [581];
      \piso.data_r_580_sv2v_reg  <= \piso.data_li [580];
      \piso.data_r_579_sv2v_reg  <= \piso.data_li [579];
      \piso.data_r_578_sv2v_reg  <= \piso.data_li [578];
      \piso.data_r_577_sv2v_reg  <= \piso.data_li [577];
      \piso.data_r_576_sv2v_reg  <= \piso.data_li [576];
      \piso.data_r_575_sv2v_reg  <= \piso.data_li [575];
      \piso.data_r_574_sv2v_reg  <= \piso.data_li [574];
      \piso.data_r_573_sv2v_reg  <= \piso.data_li [573];
      \piso.data_r_572_sv2v_reg  <= \piso.data_li [572];
      \piso.data_r_571_sv2v_reg  <= \piso.data_li [571];
      \piso.data_r_570_sv2v_reg  <= \piso.data_li [570];
      \piso.data_r_569_sv2v_reg  <= \piso.data_li [569];
      \piso.data_r_568_sv2v_reg  <= \piso.data_li [568];
      \piso.data_r_567_sv2v_reg  <= \piso.data_li [567];
      \piso.data_r_566_sv2v_reg  <= \piso.data_li [566];
      \piso.data_r_565_sv2v_reg  <= \piso.data_li [565];
      \piso.data_r_564_sv2v_reg  <= \piso.data_li [564];
      \piso.data_r_563_sv2v_reg  <= \piso.data_li [563];
      \piso.data_r_562_sv2v_reg  <= \piso.data_li [562];
      \piso.data_r_561_sv2v_reg  <= \piso.data_li [561];
      \piso.data_r_560_sv2v_reg  <= \piso.data_li [560];
      \piso.data_r_559_sv2v_reg  <= \piso.data_li [559];
      \piso.data_r_558_sv2v_reg  <= \piso.data_li [558];
      \piso.data_r_557_sv2v_reg  <= \piso.data_li [557];
      \piso.data_r_556_sv2v_reg  <= \piso.data_li [556];
      \piso.data_r_555_sv2v_reg  <= \piso.data_li [555];
      \piso.data_r_554_sv2v_reg  <= \piso.data_li [554];
      \piso.data_r_553_sv2v_reg  <= \piso.data_li [553];
      \piso.data_r_552_sv2v_reg  <= \piso.data_li [552];
      \piso.data_r_551_sv2v_reg  <= \piso.data_li [551];
      \piso.data_r_550_sv2v_reg  <= \piso.data_li [550];
      \piso.data_r_549_sv2v_reg  <= \piso.data_li [549];
      \piso.data_r_548_sv2v_reg  <= \piso.data_li [548];
      \piso.data_r_547_sv2v_reg  <= \piso.data_li [547];
      \piso.data_r_546_sv2v_reg  <= \piso.data_li [546];
      \piso.data_r_545_sv2v_reg  <= \piso.data_li [545];
      \piso.data_r_544_sv2v_reg  <= \piso.data_li [544];
      \piso.data_r_543_sv2v_reg  <= \piso.data_li [543];
      \piso.data_r_542_sv2v_reg  <= \piso.data_li [542];
      \piso.data_r_541_sv2v_reg  <= \piso.data_li [541];
      \piso.data_r_540_sv2v_reg  <= \piso.data_li [540];
      \piso.data_r_539_sv2v_reg  <= \piso.data_li [539];
      \piso.data_r_538_sv2v_reg  <= \piso.data_li [538];
      \piso.data_r_537_sv2v_reg  <= \piso.data_li [537];
      \piso.data_r_536_sv2v_reg  <= \piso.data_li [536];
      \piso.data_r_535_sv2v_reg  <= \piso.data_li [535];
      \piso.data_r_534_sv2v_reg  <= \piso.data_li [534];
      \piso.data_r_533_sv2v_reg  <= \piso.data_li [533];
      \piso.data_r_532_sv2v_reg  <= \piso.data_li [532];
      \piso.data_r_531_sv2v_reg  <= \piso.data_li [531];
      \piso.data_r_530_sv2v_reg  <= \piso.data_li [530];
      \piso.data_r_529_sv2v_reg  <= \piso.data_li [529];
      \piso.data_r_528_sv2v_reg  <= \piso.data_li [528];
      \piso.data_r_527_sv2v_reg  <= \piso.data_li [527];
      \piso.data_r_526_sv2v_reg  <= \piso.data_li [526];
      \piso.data_r_525_sv2v_reg  <= \piso.data_li [525];
      \piso.data_r_524_sv2v_reg  <= \piso.data_li [524];
      \piso.data_r_523_sv2v_reg  <= \piso.data_li [523];
      \piso.data_r_522_sv2v_reg  <= \piso.data_li [522];
      \piso.data_r_521_sv2v_reg  <= \piso.data_li [521];
      \piso.data_r_520_sv2v_reg  <= \piso.data_li [520];
      \piso.data_r_519_sv2v_reg  <= \piso.data_li [519];
      \piso.data_r_518_sv2v_reg  <= \piso.data_li [518];
      \piso.data_r_517_sv2v_reg  <= \piso.data_li [517];
      \piso.data_r_516_sv2v_reg  <= \piso.data_li [516];
      \piso.data_r_515_sv2v_reg  <= \piso.data_li [515];
      \piso.data_r_514_sv2v_reg  <= \piso.data_li [514];
      \piso.data_r_513_sv2v_reg  <= \piso.data_li [513];
      \piso.data_r_512_sv2v_reg  <= \piso.data_li [512];
      \piso.data_r_511_sv2v_reg  <= \piso.data_li [511];
      \piso.data_r_510_sv2v_reg  <= \piso.data_li [510];
      \piso.data_r_509_sv2v_reg  <= \piso.data_li [509];
      \piso.data_r_508_sv2v_reg  <= \piso.data_li [508];
      \piso.data_r_507_sv2v_reg  <= \piso.data_li [507];
      \piso.data_r_506_sv2v_reg  <= \piso.data_li [506];
      \piso.data_r_505_sv2v_reg  <= \piso.data_li [505];
      \piso.data_r_504_sv2v_reg  <= \piso.data_li [504];
      \piso.data_r_503_sv2v_reg  <= \piso.data_li [503];
      \piso.data_r_502_sv2v_reg  <= \piso.data_li [502];
      \piso.data_r_501_sv2v_reg  <= \piso.data_li [501];
      \piso.data_r_500_sv2v_reg  <= \piso.data_li [500];
      \piso.data_r_499_sv2v_reg  <= \piso.data_li [499];
      \piso.data_r_498_sv2v_reg  <= \piso.data_li [498];
      \piso.data_r_497_sv2v_reg  <= \piso.data_li [497];
      \piso.data_r_496_sv2v_reg  <= \piso.data_li [496];
      \piso.data_r_495_sv2v_reg  <= \piso.data_li [495];
      \piso.data_r_494_sv2v_reg  <= \piso.data_li [494];
      \piso.data_r_493_sv2v_reg  <= \piso.data_li [493];
      \piso.data_r_492_sv2v_reg  <= \piso.data_li [492];
      \piso.data_r_491_sv2v_reg  <= \piso.data_li [491];
      \piso.data_r_490_sv2v_reg  <= \piso.data_li [490];
      \piso.data_r_489_sv2v_reg  <= \piso.data_li [489];
      \piso.data_r_488_sv2v_reg  <= \piso.data_li [488];
      \piso.data_r_487_sv2v_reg  <= \piso.data_li [487];
      \piso.data_r_486_sv2v_reg  <= \piso.data_li [486];
      \piso.data_r_485_sv2v_reg  <= \piso.data_li [485];
      \piso.data_r_484_sv2v_reg  <= \piso.data_li [484];
      \piso.data_r_483_sv2v_reg  <= \piso.data_li [483];
      \piso.data_r_482_sv2v_reg  <= \piso.data_li [482];
      \piso.data_r_481_sv2v_reg  <= \piso.data_li [481];
      \piso.data_r_480_sv2v_reg  <= \piso.data_li [480];
      \piso.data_r_479_sv2v_reg  <= \piso.data_li [479];
      \piso.data_r_478_sv2v_reg  <= \piso.data_li [478];
      \piso.data_r_477_sv2v_reg  <= \piso.data_li [477];
      \piso.data_r_476_sv2v_reg  <= \piso.data_li [476];
      \piso.data_r_475_sv2v_reg  <= \piso.data_li [475];
      \piso.data_r_474_sv2v_reg  <= \piso.data_li [474];
      \piso.data_r_473_sv2v_reg  <= \piso.data_li [473];
      \piso.data_r_472_sv2v_reg  <= \piso.data_li [472];
      \piso.data_r_471_sv2v_reg  <= \piso.data_li [471];
      \piso.data_r_470_sv2v_reg  <= \piso.data_li [470];
      \piso.data_r_469_sv2v_reg  <= \piso.data_li [469];
      \piso.data_r_468_sv2v_reg  <= \piso.data_li [468];
      \piso.data_r_467_sv2v_reg  <= \piso.data_li [467];
      \piso.data_r_466_sv2v_reg  <= \piso.data_li [466];
      \piso.data_r_465_sv2v_reg  <= \piso.data_li [465];
      \piso.data_r_464_sv2v_reg  <= \piso.data_li [464];
      \piso.data_r_463_sv2v_reg  <= \piso.data_li [463];
      \piso.data_r_462_sv2v_reg  <= \piso.data_li [462];
      \piso.data_r_461_sv2v_reg  <= \piso.data_li [461];
      \piso.data_r_460_sv2v_reg  <= \piso.data_li [460];
      \piso.data_r_459_sv2v_reg  <= \piso.data_li [459];
      \piso.data_r_458_sv2v_reg  <= \piso.data_li [458];
      \piso.data_r_457_sv2v_reg  <= \piso.data_li [457];
      \piso.data_r_456_sv2v_reg  <= \piso.data_li [456];
      \piso.data_r_455_sv2v_reg  <= \piso.data_li [455];
      \piso.data_r_454_sv2v_reg  <= \piso.data_li [454];
      \piso.data_r_453_sv2v_reg  <= \piso.data_li [453];
      \piso.data_r_452_sv2v_reg  <= \piso.data_li [452];
      \piso.data_r_451_sv2v_reg  <= \piso.data_li [451];
      \piso.data_r_450_sv2v_reg  <= \piso.data_li [450];
      \piso.data_r_449_sv2v_reg  <= \piso.data_li [449];
      \piso.data_r_448_sv2v_reg  <= \piso.data_li [448];
      \piso.data_r_447_sv2v_reg  <= \piso.data_li [447];
      \piso.data_r_446_sv2v_reg  <= \piso.data_li [446];
      \piso.data_r_445_sv2v_reg  <= \piso.data_li [445];
      \piso.data_r_444_sv2v_reg  <= \piso.data_li [444];
      \piso.data_r_443_sv2v_reg  <= \piso.data_li [443];
      \piso.data_r_442_sv2v_reg  <= \piso.data_li [442];
      \piso.data_r_441_sv2v_reg  <= \piso.data_li [441];
      \piso.data_r_440_sv2v_reg  <= \piso.data_li [440];
      \piso.data_r_439_sv2v_reg  <= \piso.data_li [439];
      \piso.data_r_438_sv2v_reg  <= \piso.data_li [438];
      \piso.data_r_437_sv2v_reg  <= \piso.data_li [437];
      \piso.data_r_436_sv2v_reg  <= \piso.data_li [436];
      \piso.data_r_435_sv2v_reg  <= \piso.data_li [435];
      \piso.data_r_434_sv2v_reg  <= \piso.data_li [434];
      \piso.data_r_433_sv2v_reg  <= \piso.data_li [433];
      \piso.data_r_432_sv2v_reg  <= \piso.data_li [432];
      \piso.data_r_431_sv2v_reg  <= \piso.data_li [431];
      \piso.data_r_430_sv2v_reg  <= \piso.data_li [430];
      \piso.data_r_429_sv2v_reg  <= \piso.data_li [429];
      \piso.data_r_428_sv2v_reg  <= \piso.data_li [428];
      \piso.data_r_427_sv2v_reg  <= \piso.data_li [427];
      \piso.data_r_426_sv2v_reg  <= \piso.data_li [426];
      \piso.data_r_425_sv2v_reg  <= \piso.data_li [425];
      \piso.data_r_424_sv2v_reg  <= \piso.data_li [424];
      \piso.data_r_423_sv2v_reg  <= \piso.data_li [423];
      \piso.data_r_422_sv2v_reg  <= \piso.data_li [422];
      \piso.data_r_421_sv2v_reg  <= \piso.data_li [421];
      \piso.data_r_420_sv2v_reg  <= \piso.data_li [420];
      \piso.data_r_419_sv2v_reg  <= \piso.data_li [419];
      \piso.data_r_418_sv2v_reg  <= \piso.data_li [418];
      \piso.data_r_417_sv2v_reg  <= \piso.data_li [417];
      \piso.data_r_416_sv2v_reg  <= \piso.data_li [416];
      \piso.data_r_415_sv2v_reg  <= \piso.data_li [415];
      \piso.data_r_414_sv2v_reg  <= \piso.data_li [414];
      \piso.data_r_413_sv2v_reg  <= \piso.data_li [413];
      \piso.data_r_412_sv2v_reg  <= \piso.data_li [412];
      \piso.data_r_411_sv2v_reg  <= \piso.data_li [411];
      \piso.data_r_410_sv2v_reg  <= \piso.data_li [410];
      \piso.data_r_409_sv2v_reg  <= \piso.data_li [409];
      \piso.data_r_408_sv2v_reg  <= \piso.data_li [408];
      \piso.data_r_407_sv2v_reg  <= \piso.data_li [407];
      \piso.data_r_406_sv2v_reg  <= \piso.data_li [406];
      \piso.data_r_405_sv2v_reg  <= \piso.data_li [405];
      \piso.data_r_404_sv2v_reg  <= \piso.data_li [404];
      \piso.data_r_403_sv2v_reg  <= \piso.data_li [403];
      \piso.data_r_402_sv2v_reg  <= \piso.data_li [402];
      \piso.data_r_401_sv2v_reg  <= \piso.data_li [401];
      \piso.data_r_400_sv2v_reg  <= \piso.data_li [400];
      \piso.data_r_399_sv2v_reg  <= \piso.data_li [399];
      \piso.data_r_398_sv2v_reg  <= \piso.data_li [398];
      \piso.data_r_397_sv2v_reg  <= \piso.data_li [397];
      \piso.data_r_396_sv2v_reg  <= \piso.data_li [396];
      \piso.data_r_395_sv2v_reg  <= \piso.data_li [395];
      \piso.data_r_394_sv2v_reg  <= \piso.data_li [394];
      \piso.data_r_393_sv2v_reg  <= \piso.data_li [393];
      \piso.data_r_392_sv2v_reg  <= \piso.data_li [392];
      \piso.data_r_391_sv2v_reg  <= \piso.data_li [391];
      \piso.data_r_390_sv2v_reg  <= \piso.data_li [390];
      \piso.data_r_389_sv2v_reg  <= \piso.data_li [389];
      \piso.data_r_388_sv2v_reg  <= \piso.data_li [388];
      \piso.data_r_387_sv2v_reg  <= \piso.data_li [387];
      \piso.data_r_386_sv2v_reg  <= \piso.data_li [386];
      \piso.data_r_385_sv2v_reg  <= \piso.data_li [385];
      \piso.data_r_384_sv2v_reg  <= \piso.data_li [384];
      \piso.data_r_383_sv2v_reg  <= \piso.data_li [383];
      \piso.data_r_382_sv2v_reg  <= \piso.data_li [382];
      \piso.data_r_381_sv2v_reg  <= \piso.data_li [381];
      \piso.data_r_380_sv2v_reg  <= \piso.data_li [380];
      \piso.data_r_379_sv2v_reg  <= \piso.data_li [379];
      \piso.data_r_378_sv2v_reg  <= \piso.data_li [378];
      \piso.data_r_377_sv2v_reg  <= \piso.data_li [377];
      \piso.data_r_376_sv2v_reg  <= \piso.data_li [376];
      \piso.data_r_375_sv2v_reg  <= \piso.data_li [375];
      \piso.data_r_374_sv2v_reg  <= \piso.data_li [374];
      \piso.data_r_373_sv2v_reg  <= \piso.data_li [373];
      \piso.data_r_372_sv2v_reg  <= \piso.data_li [372];
      \piso.data_r_371_sv2v_reg  <= \piso.data_li [371];
      \piso.data_r_370_sv2v_reg  <= \piso.data_li [370];
      \piso.data_r_369_sv2v_reg  <= \piso.data_li [369];
      \piso.data_r_368_sv2v_reg  <= \piso.data_li [368];
      \piso.data_r_367_sv2v_reg  <= \piso.data_li [367];
      \piso.data_r_366_sv2v_reg  <= \piso.data_li [366];
      \piso.data_r_365_sv2v_reg  <= \piso.data_li [365];
      \piso.data_r_364_sv2v_reg  <= \piso.data_li [364];
      \piso.data_r_363_sv2v_reg  <= \piso.data_li [363];
      \piso.data_r_362_sv2v_reg  <= \piso.data_li [362];
      \piso.data_r_361_sv2v_reg  <= \piso.data_li [361];
      \piso.data_r_360_sv2v_reg  <= \piso.data_li [360];
      \piso.data_r_359_sv2v_reg  <= \piso.data_li [359];
      \piso.data_r_358_sv2v_reg  <= \piso.data_li [358];
      \piso.data_r_357_sv2v_reg  <= \piso.data_li [357];
      \piso.data_r_356_sv2v_reg  <= \piso.data_li [356];
      \piso.data_r_355_sv2v_reg  <= \piso.data_li [355];
      \piso.data_r_354_sv2v_reg  <= \piso.data_li [354];
      \piso.data_r_353_sv2v_reg  <= \piso.data_li [353];
      \piso.data_r_352_sv2v_reg  <= \piso.data_li [352];
      \piso.data_r_351_sv2v_reg  <= \piso.data_li [351];
      \piso.data_r_350_sv2v_reg  <= \piso.data_li [350];
      \piso.data_r_349_sv2v_reg  <= \piso.data_li [349];
      \piso.data_r_348_sv2v_reg  <= \piso.data_li [348];
      \piso.data_r_347_sv2v_reg  <= \piso.data_li [347];
      \piso.data_r_346_sv2v_reg  <= \piso.data_li [346];
      \piso.data_r_345_sv2v_reg  <= \piso.data_li [345];
      \piso.data_r_344_sv2v_reg  <= \piso.data_li [344];
      \piso.data_r_343_sv2v_reg  <= \piso.data_li [343];
      \piso.data_r_342_sv2v_reg  <= \piso.data_li [342];
      \piso.data_r_341_sv2v_reg  <= \piso.data_li [341];
      \piso.data_r_340_sv2v_reg  <= \piso.data_li [340];
      \piso.data_r_339_sv2v_reg  <= \piso.data_li [339];
      \piso.data_r_338_sv2v_reg  <= \piso.data_li [338];
      \piso.data_r_337_sv2v_reg  <= \piso.data_li [337];
      \piso.data_r_336_sv2v_reg  <= \piso.data_li [336];
      \piso.data_r_335_sv2v_reg  <= \piso.data_li [335];
      \piso.data_r_334_sv2v_reg  <= \piso.data_li [334];
      \piso.data_r_333_sv2v_reg  <= \piso.data_li [333];
      \piso.data_r_332_sv2v_reg  <= \piso.data_li [332];
      \piso.data_r_331_sv2v_reg  <= \piso.data_li [331];
      \piso.data_r_330_sv2v_reg  <= \piso.data_li [330];
      \piso.data_r_329_sv2v_reg  <= \piso.data_li [329];
      \piso.data_r_328_sv2v_reg  <= \piso.data_li [328];
      \piso.data_r_327_sv2v_reg  <= \piso.data_li [327];
      \piso.data_r_326_sv2v_reg  <= \piso.data_li [326];
      \piso.data_r_325_sv2v_reg  <= \piso.data_li [325];
      \piso.data_r_324_sv2v_reg  <= \piso.data_li [324];
      \piso.data_r_323_sv2v_reg  <= \piso.data_li [323];
      \piso.data_r_322_sv2v_reg  <= \piso.data_li [322];
      \piso.data_r_321_sv2v_reg  <= \piso.data_li [321];
      \piso.data_r_320_sv2v_reg  <= \piso.data_li [320];
      \piso.data_r_319_sv2v_reg  <= \piso.data_li [319];
      \piso.data_r_318_sv2v_reg  <= \piso.data_li [318];
      \piso.data_r_317_sv2v_reg  <= \piso.data_li [317];
      \piso.data_r_316_sv2v_reg  <= \piso.data_li [316];
      \piso.data_r_315_sv2v_reg  <= \piso.data_li [315];
      \piso.data_r_314_sv2v_reg  <= \piso.data_li [314];
      \piso.data_r_313_sv2v_reg  <= \piso.data_li [313];
      \piso.data_r_312_sv2v_reg  <= \piso.data_li [312];
      \piso.data_r_311_sv2v_reg  <= \piso.data_li [311];
      \piso.data_r_310_sv2v_reg  <= \piso.data_li [310];
      \piso.data_r_309_sv2v_reg  <= \piso.data_li [309];
      \piso.data_r_308_sv2v_reg  <= \piso.data_li [308];
      \piso.data_r_307_sv2v_reg  <= \piso.data_li [307];
      \piso.data_r_306_sv2v_reg  <= \piso.data_li [306];
      \piso.data_r_305_sv2v_reg  <= \piso.data_li [305];
      \piso.data_r_304_sv2v_reg  <= \piso.data_li [304];
      \piso.data_r_303_sv2v_reg  <= \piso.data_li [303];
      \piso.data_r_302_sv2v_reg  <= \piso.data_li [302];
      \piso.data_r_301_sv2v_reg  <= \piso.data_li [301];
      \piso.data_r_300_sv2v_reg  <= \piso.data_li [300];
      \piso.data_r_299_sv2v_reg  <= \piso.data_li [299];
      \piso.data_r_298_sv2v_reg  <= \piso.data_li [298];
      \piso.data_r_297_sv2v_reg  <= \piso.data_li [297];
      \piso.data_r_296_sv2v_reg  <= \piso.data_li [296];
      \piso.data_r_295_sv2v_reg  <= \piso.data_li [295];
      \piso.data_r_294_sv2v_reg  <= \piso.data_li [294];
      \piso.data_r_293_sv2v_reg  <= \piso.data_li [293];
      \piso.data_r_292_sv2v_reg  <= \piso.data_li [292];
      \piso.data_r_291_sv2v_reg  <= \piso.data_li [291];
      \piso.data_r_290_sv2v_reg  <= \piso.data_li [290];
      \piso.data_r_289_sv2v_reg  <= \piso.data_li [289];
      \piso.data_r_288_sv2v_reg  <= \piso.data_li [288];
      \piso.data_r_287_sv2v_reg  <= \piso.data_li [287];
      \piso.data_r_286_sv2v_reg  <= \piso.data_li [286];
      \piso.data_r_285_sv2v_reg  <= \piso.data_li [285];
      \piso.data_r_284_sv2v_reg  <= \piso.data_li [284];
      \piso.data_r_283_sv2v_reg  <= \piso.data_li [283];
      \piso.data_r_282_sv2v_reg  <= \piso.data_li [282];
      \piso.data_r_281_sv2v_reg  <= \piso.data_li [281];
      \piso.data_r_280_sv2v_reg  <= \piso.data_li [280];
      \piso.data_r_279_sv2v_reg  <= \piso.data_li [279];
      \piso.data_r_278_sv2v_reg  <= \piso.data_li [278];
      \piso.data_r_277_sv2v_reg  <= \piso.data_li [277];
      \piso.data_r_276_sv2v_reg  <= \piso.data_li [276];
      \piso.data_r_275_sv2v_reg  <= \piso.data_li [275];
      \piso.data_r_274_sv2v_reg  <= \piso.data_li [274];
      \piso.data_r_273_sv2v_reg  <= \piso.data_li [273];
      \piso.data_r_272_sv2v_reg  <= \piso.data_li [272];
      \piso.data_r_271_sv2v_reg  <= \piso.data_li [271];
      \piso.data_r_270_sv2v_reg  <= \piso.data_li [270];
      \piso.data_r_269_sv2v_reg  <= \piso.data_li [269];
      \piso.data_r_268_sv2v_reg  <= \piso.data_li [268];
      \piso.data_r_267_sv2v_reg  <= \piso.data_li [267];
      \piso.data_r_266_sv2v_reg  <= \piso.data_li [266];
      \piso.data_r_265_sv2v_reg  <= \piso.data_li [265];
      \piso.data_r_264_sv2v_reg  <= \piso.data_li [264];
      \piso.data_r_263_sv2v_reg  <= \piso.data_li [263];
      \piso.data_r_262_sv2v_reg  <= \piso.data_li [262];
      \piso.data_r_261_sv2v_reg  <= \piso.data_li [261];
      \piso.data_r_260_sv2v_reg  <= \piso.data_li [260];
      \piso.data_r_259_sv2v_reg  <= \piso.data_li [259];
      \piso.data_r_258_sv2v_reg  <= \piso.data_li [258];
      \piso.data_r_257_sv2v_reg  <= \piso.data_li [257];
      \piso.data_r_256_sv2v_reg  <= \piso.data_li [256];
      \piso.data_r_255_sv2v_reg  <= \piso.data_li [255];
      \piso.data_r_254_sv2v_reg  <= \piso.data_li [254];
      \piso.data_r_253_sv2v_reg  <= \piso.data_li [253];
      \piso.data_r_252_sv2v_reg  <= \piso.data_li [252];
      \piso.data_r_251_sv2v_reg  <= \piso.data_li [251];
      \piso.data_r_250_sv2v_reg  <= \piso.data_li [250];
      \piso.data_r_249_sv2v_reg  <= \piso.data_li [249];
      \piso.data_r_248_sv2v_reg  <= \piso.data_li [248];
      \piso.data_r_247_sv2v_reg  <= \piso.data_li [247];
      \piso.data_r_246_sv2v_reg  <= \piso.data_li [246];
      \piso.data_r_245_sv2v_reg  <= \piso.data_li [245];
      \piso.data_r_244_sv2v_reg  <= \piso.data_li [244];
      \piso.data_r_243_sv2v_reg  <= \piso.data_li [243];
      \piso.data_r_242_sv2v_reg  <= \piso.data_li [242];
      \piso.data_r_241_sv2v_reg  <= \piso.data_li [241];
      \piso.data_r_240_sv2v_reg  <= \piso.data_li [240];
      \piso.data_r_239_sv2v_reg  <= \piso.data_li [239];
      \piso.data_r_238_sv2v_reg  <= \piso.data_li [238];
      \piso.data_r_237_sv2v_reg  <= \piso.data_li [237];
      \piso.data_r_236_sv2v_reg  <= \piso.data_li [236];
      \piso.data_r_235_sv2v_reg  <= \piso.data_li [235];
      \piso.data_r_234_sv2v_reg  <= \piso.data_li [234];
      \piso.data_r_233_sv2v_reg  <= \piso.data_li [233];
      \piso.data_r_232_sv2v_reg  <= \piso.data_li [232];
      \piso.data_r_231_sv2v_reg  <= \piso.data_li [231];
      \piso.data_r_230_sv2v_reg  <= \piso.data_li [230];
      \piso.data_r_229_sv2v_reg  <= \piso.data_li [229];
      \piso.data_r_228_sv2v_reg  <= \piso.data_li [228];
      \piso.data_r_227_sv2v_reg  <= \piso.data_li [227];
      \piso.data_r_226_sv2v_reg  <= \piso.data_li [226];
      \piso.data_r_225_sv2v_reg  <= \piso.data_li [225];
      \piso.data_r_224_sv2v_reg  <= \piso.data_li [224];
      \piso.data_r_223_sv2v_reg  <= \piso.data_li [223];
      \piso.data_r_222_sv2v_reg  <= \piso.data_li [222];
      \piso.data_r_221_sv2v_reg  <= \piso.data_li [221];
      \piso.data_r_220_sv2v_reg  <= \piso.data_li [220];
      \piso.data_r_219_sv2v_reg  <= \piso.data_li [219];
      \piso.data_r_218_sv2v_reg  <= \piso.data_li [218];
      \piso.data_r_217_sv2v_reg  <= \piso.data_li [217];
      \piso.data_r_216_sv2v_reg  <= \piso.data_li [216];
      \piso.data_r_215_sv2v_reg  <= \piso.data_li [215];
      \piso.data_r_214_sv2v_reg  <= \piso.data_li [214];
      \piso.data_r_213_sv2v_reg  <= \piso.data_li [213];
      \piso.data_r_212_sv2v_reg  <= \piso.data_li [212];
      \piso.data_r_211_sv2v_reg  <= \piso.data_li [211];
      \piso.data_r_210_sv2v_reg  <= \piso.data_li [210];
      \piso.data_r_209_sv2v_reg  <= \piso.data_li [209];
      \piso.data_r_208_sv2v_reg  <= \piso.data_li [208];
      \piso.data_r_207_sv2v_reg  <= \piso.data_li [207];
      \piso.data_r_206_sv2v_reg  <= \piso.data_li [206];
      \piso.data_r_205_sv2v_reg  <= \piso.data_li [205];
      \piso.data_r_204_sv2v_reg  <= \piso.data_li [204];
      \piso.data_r_203_sv2v_reg  <= \piso.data_li [203];
      \piso.data_r_202_sv2v_reg  <= \piso.data_li [202];
      \piso.data_r_201_sv2v_reg  <= \piso.data_li [201];
      \piso.data_r_200_sv2v_reg  <= \piso.data_li [200];
      \piso.data_r_199_sv2v_reg  <= \piso.data_li [199];
      \piso.data_r_198_sv2v_reg  <= \piso.data_li [198];
      \piso.data_r_197_sv2v_reg  <= \piso.data_li [197];
      \piso.data_r_196_sv2v_reg  <= \piso.data_li [196];
      \piso.data_r_195_sv2v_reg  <= \piso.data_li [195];
      \piso.data_r_194_sv2v_reg  <= \piso.data_li [194];
      \piso.data_r_193_sv2v_reg  <= \piso.data_li [193];
      \piso.data_r_192_sv2v_reg  <= \piso.data_li [192];
      \piso.data_r_191_sv2v_reg  <= \piso.data_li [191];
      \piso.data_r_190_sv2v_reg  <= \piso.data_li [190];
      \piso.data_r_189_sv2v_reg  <= \piso.data_li [189];
      \piso.data_r_188_sv2v_reg  <= \piso.data_li [188];
      \piso.data_r_187_sv2v_reg  <= \piso.data_li [187];
      \piso.data_r_186_sv2v_reg  <= \piso.data_li [186];
      \piso.data_r_185_sv2v_reg  <= \piso.data_li [185];
      \piso.data_r_184_sv2v_reg  <= \piso.data_li [184];
      \piso.data_r_183_sv2v_reg  <= \piso.data_li [183];
      \piso.data_r_182_sv2v_reg  <= \piso.data_li [182];
      \piso.data_r_181_sv2v_reg  <= \piso.data_li [181];
      \piso.data_r_180_sv2v_reg  <= \piso.data_li [180];
      \piso.data_r_179_sv2v_reg  <= \piso.data_li [179];
      \piso.data_r_178_sv2v_reg  <= \piso.data_li [178];
      \piso.data_r_177_sv2v_reg  <= \piso.data_li [177];
      \piso.data_r_176_sv2v_reg  <= \piso.data_li [176];
      \piso.data_r_175_sv2v_reg  <= \piso.data_li [175];
      \piso.data_r_174_sv2v_reg  <= \piso.data_li [174];
      \piso.data_r_173_sv2v_reg  <= \piso.data_li [173];
      \piso.data_r_172_sv2v_reg  <= \piso.data_li [172];
      \piso.data_r_171_sv2v_reg  <= \piso.data_li [171];
      \piso.data_r_170_sv2v_reg  <= \piso.data_li [170];
      \piso.data_r_169_sv2v_reg  <= \piso.data_li [169];
      \piso.data_r_168_sv2v_reg  <= \piso.data_li [168];
      \piso.data_r_167_sv2v_reg  <= \piso.data_li [167];
      \piso.data_r_166_sv2v_reg  <= \piso.data_li [166];
      \piso.data_r_165_sv2v_reg  <= \piso.data_li [165];
      \piso.data_r_164_sv2v_reg  <= \piso.data_li [164];
      \piso.data_r_163_sv2v_reg  <= \piso.data_li [163];
      \piso.data_r_162_sv2v_reg  <= \piso.data_li [162];
      \piso.data_r_161_sv2v_reg  <= \piso.data_li [161];
      \piso.data_r_160_sv2v_reg  <= \piso.data_li [160];
      \piso.data_r_159_sv2v_reg  <= \piso.data_li [159];
      \piso.data_r_158_sv2v_reg  <= \piso.data_li [158];
      \piso.data_r_157_sv2v_reg  <= \piso.data_li [157];
      \piso.data_r_156_sv2v_reg  <= \piso.data_li [156];
      \piso.data_r_155_sv2v_reg  <= \piso.data_li [155];
      \piso.data_r_154_sv2v_reg  <= \piso.data_li [154];
      \piso.data_r_153_sv2v_reg  <= \piso.data_li [153];
      \piso.data_r_152_sv2v_reg  <= \piso.data_li [152];
      \piso.data_r_151_sv2v_reg  <= \piso.data_li [151];
      \piso.data_r_150_sv2v_reg  <= \piso.data_li [150];
      \piso.data_r_149_sv2v_reg  <= \piso.data_li [149];
      \piso.data_r_148_sv2v_reg  <= \piso.data_li [148];
      \piso.data_r_147_sv2v_reg  <= \piso.data_li [147];
      \piso.data_r_146_sv2v_reg  <= \piso.data_li [146];
      \piso.data_r_145_sv2v_reg  <= \piso.data_li [145];
      \piso.data_r_144_sv2v_reg  <= \piso.data_li [144];
      \piso.data_r_143_sv2v_reg  <= \piso.data_li [143];
      \piso.data_r_142_sv2v_reg  <= \piso.data_li [142];
      \piso.data_r_141_sv2v_reg  <= \piso.data_li [141];
      \piso.data_r_140_sv2v_reg  <= \piso.data_li [140];
      \piso.data_r_139_sv2v_reg  <= \piso.data_li [139];
      \piso.data_r_138_sv2v_reg  <= \piso.data_li [138];
      \piso.data_r_137_sv2v_reg  <= \piso.data_li [137];
      \piso.data_r_136_sv2v_reg  <= \piso.data_li [136];
      \piso.data_r_135_sv2v_reg  <= \piso.data_li [135];
      \piso.data_r_134_sv2v_reg  <= \piso.data_li [134];
      \piso.data_r_133_sv2v_reg  <= \piso.data_li [133];
      \piso.data_r_132_sv2v_reg  <= \piso.data_li [132];
      \piso.data_r_131_sv2v_reg  <= \piso.data_li [131];
      \piso.data_r_130_sv2v_reg  <= \piso.data_li [130];
      \piso.data_r_129_sv2v_reg  <= \piso.data_li [129];
      \piso.data_r_128_sv2v_reg  <= \piso.data_li [128];
      \piso.data_r_127_sv2v_reg  <= \piso.data_li [127];
      \piso.data_r_126_sv2v_reg  <= \piso.data_li [126];
      \piso.data_r_125_sv2v_reg  <= \piso.data_li [125];
      \piso.data_r_124_sv2v_reg  <= \piso.data_li [124];
      \piso.data_r_123_sv2v_reg  <= \piso.data_li [123];
      \piso.data_r_122_sv2v_reg  <= \piso.data_li [122];
      \piso.data_r_121_sv2v_reg  <= \piso.data_li [121];
      \piso.data_r_120_sv2v_reg  <= \piso.data_li [120];
      \piso.data_r_119_sv2v_reg  <= \piso.data_li [119];
      \piso.data_r_118_sv2v_reg  <= \piso.data_li [118];
      \piso.data_r_117_sv2v_reg  <= \piso.data_li [117];
      \piso.data_r_116_sv2v_reg  <= \piso.data_li [116];
      \piso.data_r_115_sv2v_reg  <= \piso.data_li [115];
      \piso.data_r_114_sv2v_reg  <= \piso.data_li [114];
      \piso.data_r_113_sv2v_reg  <= \piso.data_li [113];
      \piso.data_r_112_sv2v_reg  <= \piso.data_li [112];
      \piso.data_r_111_sv2v_reg  <= \piso.data_li [111];
      \piso.data_r_110_sv2v_reg  <= \piso.data_li [110];
      \piso.data_r_109_sv2v_reg  <= \piso.data_li [109];
      \piso.data_r_108_sv2v_reg  <= \piso.data_li [108];
      \piso.data_r_107_sv2v_reg  <= \piso.data_li [107];
      \piso.data_r_106_sv2v_reg  <= \piso.data_li [106];
      \piso.data_r_105_sv2v_reg  <= \piso.data_li [105];
      \piso.data_r_104_sv2v_reg  <= \piso.data_li [104];
      \piso.data_r_103_sv2v_reg  <= \piso.data_li [103];
      \piso.data_r_102_sv2v_reg  <= \piso.data_li [102];
      \piso.data_r_101_sv2v_reg  <= \piso.data_li [101];
      \piso.data_r_100_sv2v_reg  <= \piso.data_li [100];
      \piso.data_r_99_sv2v_reg  <= \piso.data_li [99];
      \piso.data_r_98_sv2v_reg  <= \piso.data_li [98];
      \piso.data_r_97_sv2v_reg  <= \piso.data_li [97];
      \piso.data_r_96_sv2v_reg  <= \piso.data_li [96];
      \piso.data_r_95_sv2v_reg  <= \piso.data_li [95];
      \piso.data_r_94_sv2v_reg  <= \piso.data_li [94];
      \piso.data_r_93_sv2v_reg  <= \piso.data_li [93];
      \piso.data_r_92_sv2v_reg  <= \piso.data_li [92];
      \piso.data_r_91_sv2v_reg  <= \piso.data_li [91];
      \piso.data_r_90_sv2v_reg  <= \piso.data_li [90];
      \piso.data_r_89_sv2v_reg  <= \piso.data_li [89];
      \piso.data_r_88_sv2v_reg  <= \piso.data_li [88];
      \piso.data_r_87_sv2v_reg  <= \piso.data_li [87];
      \piso.data_r_86_sv2v_reg  <= \piso.data_li [86];
      \piso.data_r_85_sv2v_reg  <= \piso.data_li [85];
      \piso.data_r_84_sv2v_reg  <= \piso.data_li [84];
      \piso.data_r_83_sv2v_reg  <= \piso.data_li [83];
      \piso.data_r_82_sv2v_reg  <= \piso.data_li [82];
      \piso.data_r_81_sv2v_reg  <= \piso.data_li [81];
      \piso.data_r_80_sv2v_reg  <= \piso.data_li [80];
      \piso.data_r_79_sv2v_reg  <= \piso.data_li [79];
      \piso.data_r_78_sv2v_reg  <= \piso.data_li [78];
      \piso.data_r_77_sv2v_reg  <= \piso.data_li [77];
      \piso.data_r_76_sv2v_reg  <= \piso.data_li [76];
      \piso.data_r_75_sv2v_reg  <= \piso.data_li [75];
      \piso.data_r_74_sv2v_reg  <= \piso.data_li [74];
      \piso.data_r_73_sv2v_reg  <= \piso.data_li [73];
      \piso.data_r_72_sv2v_reg  <= \piso.data_li [72];
      \piso.data_r_71_sv2v_reg  <= \piso.data_li [71];
      \piso.data_r_70_sv2v_reg  <= \piso.data_li [70];
      \piso.data_r_69_sv2v_reg  <= \piso.data_li [69];
      \piso.data_r_68_sv2v_reg  <= \piso.data_li [68];
      \piso.data_r_67_sv2v_reg  <= \piso.data_li [67];
      \piso.data_r_66_sv2v_reg  <= \piso.data_li [66];
      \piso.data_r_65_sv2v_reg  <= \piso.data_li [65];
      \piso.data_r_64_sv2v_reg  <= \piso.data_li [64];
      \piso.data_r_63_sv2v_reg  <= \piso.data_li [63];
      \piso.data_r_62_sv2v_reg  <= \piso.data_li [62];
      \piso.data_r_61_sv2v_reg  <= \piso.data_li [61];
      \piso.data_r_60_sv2v_reg  <= \piso.data_li [60];
      \piso.data_r_59_sv2v_reg  <= \piso.data_li [59];
      \piso.data_r_58_sv2v_reg  <= \piso.data_li [58];
      \piso.data_r_57_sv2v_reg  <= \piso.data_li [57];
      \piso.data_r_56_sv2v_reg  <= \piso.data_li [56];
      \piso.data_r_55_sv2v_reg  <= \piso.data_li [55];
      \piso.data_r_54_sv2v_reg  <= \piso.data_li [54];
      \piso.data_r_53_sv2v_reg  <= \piso.data_li [53];
      \piso.data_r_52_sv2v_reg  <= \piso.data_li [52];
      \piso.data_r_51_sv2v_reg  <= \piso.data_li [51];
      \piso.data_r_50_sv2v_reg  <= \piso.data_li [50];
      \piso.data_r_49_sv2v_reg  <= \piso.data_li [49];
      \piso.data_r_48_sv2v_reg  <= \piso.data_li [48];
      \piso.data_r_47_sv2v_reg  <= \piso.data_li [47];
      \piso.data_r_46_sv2v_reg  <= \piso.data_li [46];
      \piso.data_r_45_sv2v_reg  <= \piso.data_li [45];
      \piso.data_r_44_sv2v_reg  <= \piso.data_li [44];
      \piso.data_r_43_sv2v_reg  <= \piso.data_li [43];
      \piso.data_r_42_sv2v_reg  <= \piso.data_li [42];
      \piso.data_r_41_sv2v_reg  <= \piso.data_li [41];
      \piso.data_r_40_sv2v_reg  <= \piso.data_li [40];
      \piso.data_r_39_sv2v_reg  <= \piso.data_li [39];
      \piso.data_r_38_sv2v_reg  <= \piso.data_li [38];
      \piso.data_r_37_sv2v_reg  <= \piso.data_li [37];
      \piso.data_r_36_sv2v_reg  <= \piso.data_li [36];
      \piso.data_r_35_sv2v_reg  <= \piso.data_li [35];
      \piso.data_r_34_sv2v_reg  <= \piso.data_li [34];
      \piso.data_r_33_sv2v_reg  <= \piso.data_li [33];
      \piso.data_r_32_sv2v_reg  <= \piso.data_li [32];
      \piso.data_r_31_sv2v_reg  <= \piso.data_li [31];
      \piso.data_r_30_sv2v_reg  <= \piso.data_li [30];
      \piso.data_r_29_sv2v_reg  <= \piso.data_li [29];
      \piso.data_r_28_sv2v_reg  <= \piso.data_li [28];
      \piso.data_r_27_sv2v_reg  <= \piso.data_li [27];
      \piso.data_r_26_sv2v_reg  <= \piso.data_li [26];
      \piso.data_r_25_sv2v_reg  <= \piso.data_li [25];
      \piso.data_r_24_sv2v_reg  <= \piso.data_li [24];
      \piso.data_r_23_sv2v_reg  <= \piso.data_li [23];
      \piso.data_r_22_sv2v_reg  <= \piso.data_li [22];
      \piso.data_r_21_sv2v_reg  <= \piso.data_li [21];
      \piso.data_r_20_sv2v_reg  <= \piso.data_li [20];
      \piso.data_r_19_sv2v_reg  <= \piso.data_li [19];
      \piso.data_r_18_sv2v_reg  <= \piso.data_li [18];
      \piso.data_r_17_sv2v_reg  <= \piso.data_li [17];
      \piso.data_r_16_sv2v_reg  <= \piso.data_li [16];
      \piso.data_r_15_sv2v_reg  <= \piso.data_li [15];
      \piso.data_r_14_sv2v_reg  <= \piso.data_li [14];
      \piso.data_r_13_sv2v_reg  <= \piso.data_li [13];
      \piso.data_r_12_sv2v_reg  <= \piso.data_li [12];
      \piso.data_r_11_sv2v_reg  <= \piso.data_li [11];
      \piso.data_r_10_sv2v_reg  <= \piso.data_li [10];
      \piso.data_r_9_sv2v_reg  <= \piso.data_li [9];
      \piso.data_r_8_sv2v_reg  <= \piso.data_li [8];
      \piso.data_r_7_sv2v_reg  <= \piso.data_li [7];
      \piso.data_r_6_sv2v_reg  <= \piso.data_li [6];
      \piso.data_r_5_sv2v_reg  <= \piso.data_li [5];
      \piso.data_r_4_sv2v_reg  <= \piso.data_li [4];
      \piso.data_r_3_sv2v_reg  <= \piso.data_li [3];
      \piso.data_r_2_sv2v_reg  <= \piso.data_li [2];
      \piso.data_r_1_sv2v_reg  <= \piso.data_li [1];
      \piso.data_r_0_sv2v_reg  <= \piso.data_li [0];
    end 
    if(reset_i) begin
      \piso.shift_ctr_r_5_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_4_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_3_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_2_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_1_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_0_sv2v_reg  <= 1'b0;
    end else if(N154) begin
      \piso.shift_ctr_r_5_sv2v_reg  <= N14;
      \piso.shift_ctr_r_4_sv2v_reg  <= N13;
      \piso.shift_ctr_r_3_sv2v_reg  <= N12;
      \piso.shift_ctr_r_2_sv2v_reg  <= N11;
      \piso.shift_ctr_r_1_sv2v_reg  <= N10;
      \piso.shift_ctr_r_0_sv2v_reg  <= N9;
    end 
  end


endmodule

