

module top
(
  clk_i,
  reset_i,
  ready_o,
  v_i,
  data_i,
  v_o,
  data_o,
  ready_i
);

  input [31:0] data_i;
  output [49:0] v_o;
  output [1599:0] data_o;
  input [49:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output ready_o;

  bsg_front_side_bus_hop_in
  wrapper
  (
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .ready_i(ready_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [63:0] \nz.mem ;
  reg \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [62] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [61] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [60] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [59] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [58] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [57] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [56] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [55] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [54] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [53] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [52] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [51] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [50] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [49] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [48] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [47] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [46] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [45] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [44] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [43] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [42] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [41] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [40] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [39] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [38] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [37] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [36] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [35] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [34] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [33] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_63_sv2v_reg  <= w_data_i[31];
      \nz.mem_62_sv2v_reg  <= w_data_i[30];
      \nz.mem_61_sv2v_reg  <= w_data_i[29];
      \nz.mem_60_sv2v_reg  <= w_data_i[28];
      \nz.mem_59_sv2v_reg  <= w_data_i[27];
      \nz.mem_58_sv2v_reg  <= w_data_i[26];
      \nz.mem_57_sv2v_reg  <= w_data_i[25];
      \nz.mem_56_sv2v_reg  <= w_data_i[24];
      \nz.mem_55_sv2v_reg  <= w_data_i[23];
      \nz.mem_54_sv2v_reg  <= w_data_i[22];
      \nz.mem_53_sv2v_reg  <= w_data_i[21];
      \nz.mem_52_sv2v_reg  <= w_data_i[20];
      \nz.mem_51_sv2v_reg  <= w_data_i[19];
      \nz.mem_50_sv2v_reg  <= w_data_i[18];
      \nz.mem_49_sv2v_reg  <= w_data_i[17];
      \nz.mem_48_sv2v_reg  <= w_data_i[16];
      \nz.mem_47_sv2v_reg  <= w_data_i[15];
      \nz.mem_46_sv2v_reg  <= w_data_i[14];
      \nz.mem_45_sv2v_reg  <= w_data_i[13];
      \nz.mem_44_sv2v_reg  <= w_data_i[12];
      \nz.mem_43_sv2v_reg  <= w_data_i[11];
      \nz.mem_42_sv2v_reg  <= w_data_i[10];
      \nz.mem_41_sv2v_reg  <= w_data_i[9];
      \nz.mem_40_sv2v_reg  <= w_data_i[8];
      \nz.mem_39_sv2v_reg  <= w_data_i[7];
      \nz.mem_38_sv2v_reg  <= w_data_i[6];
      \nz.mem_37_sv2v_reg  <= w_data_i[5];
      \nz.mem_36_sv2v_reg  <= w_data_i[4];
      \nz.mem_35_sv2v_reg  <= w_data_i[3];
      \nz.mem_34_sv2v_reg  <= w_data_i[2];
      \nz.mem_33_sv2v_reg  <= w_data_i[1];
      \nz.mem_32_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_front_side_bus_hop_in
(
  clk_i,
  reset_i,
  ready_o,
  v_i,
  data_i,
  v_o,
  data_o,
  ready_i
);

  input [31:0] data_i;
  output [49:0] v_o;
  output [1599:0] data_o;
  input [49:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output ready_o;
  wire [49:0] v_o,sent_r,sent_n;
  wire [1599:0] data_o;
  wire ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,data_o_0__31_,data_o_0__30_,data_o_0__29_,
  data_o_0__28_,data_o_0__27_,data_o_0__26_,data_o_0__25_,data_o_0__24_,
  data_o_0__23_,data_o_0__22_,data_o_0__21_,data_o_0__20_,data_o_0__19_,data_o_0__18_,
  data_o_0__17_,data_o_0__16_,data_o_0__15_,data_o_0__14_,data_o_0__13_,data_o_0__12_,
  data_o_0__11_,data_o_0__10_,data_o_0__9_,data_o_0__8_,data_o_0__7_,data_o_0__6_,
  data_o_0__5_,data_o_0__4_,data_o_0__3_,data_o_0__2_,data_o_0__1_,data_o_0__0_,
  fifo_v,fifo_yumi,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,
  N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,
  N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,
  N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,
  N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,
  N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,
  N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,
  N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,
  N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,
  N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
  N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,
  N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,
  N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,
  N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,
  N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,
  N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,
  N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
  N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,
  N345,N346,N347;
  reg sent_r_0_sv2v_reg,sent_r_1_sv2v_reg,sent_r_2_sv2v_reg,sent_r_3_sv2v_reg,
  sent_r_4_sv2v_reg,sent_r_5_sv2v_reg,sent_r_6_sv2v_reg,sent_r_7_sv2v_reg,
  sent_r_8_sv2v_reg,sent_r_9_sv2v_reg,sent_r_10_sv2v_reg,sent_r_11_sv2v_reg,sent_r_12_sv2v_reg,
  sent_r_13_sv2v_reg,sent_r_14_sv2v_reg,sent_r_15_sv2v_reg,sent_r_16_sv2v_reg,
  sent_r_17_sv2v_reg,sent_r_18_sv2v_reg,sent_r_19_sv2v_reg,sent_r_20_sv2v_reg,
  sent_r_21_sv2v_reg,sent_r_22_sv2v_reg,sent_r_23_sv2v_reg,sent_r_24_sv2v_reg,
  sent_r_25_sv2v_reg,sent_r_26_sv2v_reg,sent_r_27_sv2v_reg,sent_r_28_sv2v_reg,sent_r_29_sv2v_reg,
  sent_r_30_sv2v_reg,sent_r_31_sv2v_reg,sent_r_32_sv2v_reg,sent_r_33_sv2v_reg,
  sent_r_34_sv2v_reg,sent_r_35_sv2v_reg,sent_r_36_sv2v_reg,sent_r_37_sv2v_reg,
  sent_r_38_sv2v_reg,sent_r_39_sv2v_reg,sent_r_40_sv2v_reg,sent_r_41_sv2v_reg,
  sent_r_42_sv2v_reg,sent_r_43_sv2v_reg,sent_r_44_sv2v_reg,sent_r_45_sv2v_reg,
  sent_r_46_sv2v_reg,sent_r_47_sv2v_reg,sent_r_48_sv2v_reg,sent_r_49_sv2v_reg;
  assign sent_r[0] = sent_r_0_sv2v_reg;
  assign sent_r[1] = sent_r_1_sv2v_reg;
  assign sent_r[2] = sent_r_2_sv2v_reg;
  assign sent_r[3] = sent_r_3_sv2v_reg;
  assign sent_r[4] = sent_r_4_sv2v_reg;
  assign sent_r[5] = sent_r_5_sv2v_reg;
  assign sent_r[6] = sent_r_6_sv2v_reg;
  assign sent_r[7] = sent_r_7_sv2v_reg;
  assign sent_r[8] = sent_r_8_sv2v_reg;
  assign sent_r[9] = sent_r_9_sv2v_reg;
  assign sent_r[10] = sent_r_10_sv2v_reg;
  assign sent_r[11] = sent_r_11_sv2v_reg;
  assign sent_r[12] = sent_r_12_sv2v_reg;
  assign sent_r[13] = sent_r_13_sv2v_reg;
  assign sent_r[14] = sent_r_14_sv2v_reg;
  assign sent_r[15] = sent_r_15_sv2v_reg;
  assign sent_r[16] = sent_r_16_sv2v_reg;
  assign sent_r[17] = sent_r_17_sv2v_reg;
  assign sent_r[18] = sent_r_18_sv2v_reg;
  assign sent_r[19] = sent_r_19_sv2v_reg;
  assign sent_r[20] = sent_r_20_sv2v_reg;
  assign sent_r[21] = sent_r_21_sv2v_reg;
  assign sent_r[22] = sent_r_22_sv2v_reg;
  assign sent_r[23] = sent_r_23_sv2v_reg;
  assign sent_r[24] = sent_r_24_sv2v_reg;
  assign sent_r[25] = sent_r_25_sv2v_reg;
  assign sent_r[26] = sent_r_26_sv2v_reg;
  assign sent_r[27] = sent_r_27_sv2v_reg;
  assign sent_r[28] = sent_r_28_sv2v_reg;
  assign sent_r[29] = sent_r_29_sv2v_reg;
  assign sent_r[30] = sent_r_30_sv2v_reg;
  assign sent_r[31] = sent_r_31_sv2v_reg;
  assign sent_r[32] = sent_r_32_sv2v_reg;
  assign sent_r[33] = sent_r_33_sv2v_reg;
  assign sent_r[34] = sent_r_34_sv2v_reg;
  assign sent_r[35] = sent_r_35_sv2v_reg;
  assign sent_r[36] = sent_r_36_sv2v_reg;
  assign sent_r[37] = sent_r_37_sv2v_reg;
  assign sent_r[38] = sent_r_38_sv2v_reg;
  assign sent_r[39] = sent_r_39_sv2v_reg;
  assign sent_r[40] = sent_r_40_sv2v_reg;
  assign sent_r[41] = sent_r_41_sv2v_reg;
  assign sent_r[42] = sent_r_42_sv2v_reg;
  assign sent_r[43] = sent_r_43_sv2v_reg;
  assign sent_r[44] = sent_r_44_sv2v_reg;
  assign sent_r[45] = sent_r_45_sv2v_reg;
  assign sent_r[46] = sent_r_46_sv2v_reg;
  assign sent_r[47] = sent_r_47_sv2v_reg;
  assign sent_r[48] = sent_r_48_sv2v_reg;
  assign sent_r[49] = sent_r_49_sv2v_reg;
  assign data_o[31] = data_o_0__31_;
  assign data_o[63] = data_o_0__31_;
  assign data_o[95] = data_o_0__31_;
  assign data_o[127] = data_o_0__31_;
  assign data_o[159] = data_o_0__31_;
  assign data_o[191] = data_o_0__31_;
  assign data_o[223] = data_o_0__31_;
  assign data_o[255] = data_o_0__31_;
  assign data_o[287] = data_o_0__31_;
  assign data_o[319] = data_o_0__31_;
  assign data_o[351] = data_o_0__31_;
  assign data_o[383] = data_o_0__31_;
  assign data_o[415] = data_o_0__31_;
  assign data_o[447] = data_o_0__31_;
  assign data_o[479] = data_o_0__31_;
  assign data_o[511] = data_o_0__31_;
  assign data_o[543] = data_o_0__31_;
  assign data_o[575] = data_o_0__31_;
  assign data_o[607] = data_o_0__31_;
  assign data_o[639] = data_o_0__31_;
  assign data_o[671] = data_o_0__31_;
  assign data_o[703] = data_o_0__31_;
  assign data_o[735] = data_o_0__31_;
  assign data_o[767] = data_o_0__31_;
  assign data_o[799] = data_o_0__31_;
  assign data_o[831] = data_o_0__31_;
  assign data_o[863] = data_o_0__31_;
  assign data_o[895] = data_o_0__31_;
  assign data_o[927] = data_o_0__31_;
  assign data_o[959] = data_o_0__31_;
  assign data_o[991] = data_o_0__31_;
  assign data_o[1023] = data_o_0__31_;
  assign data_o[1055] = data_o_0__31_;
  assign data_o[1087] = data_o_0__31_;
  assign data_o[1119] = data_o_0__31_;
  assign data_o[1151] = data_o_0__31_;
  assign data_o[1183] = data_o_0__31_;
  assign data_o[1215] = data_o_0__31_;
  assign data_o[1247] = data_o_0__31_;
  assign data_o[1279] = data_o_0__31_;
  assign data_o[1311] = data_o_0__31_;
  assign data_o[1343] = data_o_0__31_;
  assign data_o[1375] = data_o_0__31_;
  assign data_o[1407] = data_o_0__31_;
  assign data_o[1439] = data_o_0__31_;
  assign data_o[1471] = data_o_0__31_;
  assign data_o[1503] = data_o_0__31_;
  assign data_o[1535] = data_o_0__31_;
  assign data_o[1567] = data_o_0__31_;
  assign data_o[1599] = data_o_0__31_;
  assign data_o[30] = data_o_0__30_;
  assign data_o[62] = data_o_0__30_;
  assign data_o[94] = data_o_0__30_;
  assign data_o[126] = data_o_0__30_;
  assign data_o[158] = data_o_0__30_;
  assign data_o[190] = data_o_0__30_;
  assign data_o[222] = data_o_0__30_;
  assign data_o[254] = data_o_0__30_;
  assign data_o[286] = data_o_0__30_;
  assign data_o[318] = data_o_0__30_;
  assign data_o[350] = data_o_0__30_;
  assign data_o[382] = data_o_0__30_;
  assign data_o[414] = data_o_0__30_;
  assign data_o[446] = data_o_0__30_;
  assign data_o[478] = data_o_0__30_;
  assign data_o[510] = data_o_0__30_;
  assign data_o[542] = data_o_0__30_;
  assign data_o[574] = data_o_0__30_;
  assign data_o[606] = data_o_0__30_;
  assign data_o[638] = data_o_0__30_;
  assign data_o[670] = data_o_0__30_;
  assign data_o[702] = data_o_0__30_;
  assign data_o[734] = data_o_0__30_;
  assign data_o[766] = data_o_0__30_;
  assign data_o[798] = data_o_0__30_;
  assign data_o[830] = data_o_0__30_;
  assign data_o[862] = data_o_0__30_;
  assign data_o[894] = data_o_0__30_;
  assign data_o[926] = data_o_0__30_;
  assign data_o[958] = data_o_0__30_;
  assign data_o[990] = data_o_0__30_;
  assign data_o[1022] = data_o_0__30_;
  assign data_o[1054] = data_o_0__30_;
  assign data_o[1086] = data_o_0__30_;
  assign data_o[1118] = data_o_0__30_;
  assign data_o[1150] = data_o_0__30_;
  assign data_o[1182] = data_o_0__30_;
  assign data_o[1214] = data_o_0__30_;
  assign data_o[1246] = data_o_0__30_;
  assign data_o[1278] = data_o_0__30_;
  assign data_o[1310] = data_o_0__30_;
  assign data_o[1342] = data_o_0__30_;
  assign data_o[1374] = data_o_0__30_;
  assign data_o[1406] = data_o_0__30_;
  assign data_o[1438] = data_o_0__30_;
  assign data_o[1470] = data_o_0__30_;
  assign data_o[1502] = data_o_0__30_;
  assign data_o[1534] = data_o_0__30_;
  assign data_o[1566] = data_o_0__30_;
  assign data_o[1598] = data_o_0__30_;
  assign data_o[29] = data_o_0__29_;
  assign data_o[61] = data_o_0__29_;
  assign data_o[93] = data_o_0__29_;
  assign data_o[125] = data_o_0__29_;
  assign data_o[157] = data_o_0__29_;
  assign data_o[189] = data_o_0__29_;
  assign data_o[221] = data_o_0__29_;
  assign data_o[253] = data_o_0__29_;
  assign data_o[285] = data_o_0__29_;
  assign data_o[317] = data_o_0__29_;
  assign data_o[349] = data_o_0__29_;
  assign data_o[381] = data_o_0__29_;
  assign data_o[413] = data_o_0__29_;
  assign data_o[445] = data_o_0__29_;
  assign data_o[477] = data_o_0__29_;
  assign data_o[509] = data_o_0__29_;
  assign data_o[541] = data_o_0__29_;
  assign data_o[573] = data_o_0__29_;
  assign data_o[605] = data_o_0__29_;
  assign data_o[637] = data_o_0__29_;
  assign data_o[669] = data_o_0__29_;
  assign data_o[701] = data_o_0__29_;
  assign data_o[733] = data_o_0__29_;
  assign data_o[765] = data_o_0__29_;
  assign data_o[797] = data_o_0__29_;
  assign data_o[829] = data_o_0__29_;
  assign data_o[861] = data_o_0__29_;
  assign data_o[893] = data_o_0__29_;
  assign data_o[925] = data_o_0__29_;
  assign data_o[957] = data_o_0__29_;
  assign data_o[989] = data_o_0__29_;
  assign data_o[1021] = data_o_0__29_;
  assign data_o[1053] = data_o_0__29_;
  assign data_o[1085] = data_o_0__29_;
  assign data_o[1117] = data_o_0__29_;
  assign data_o[1149] = data_o_0__29_;
  assign data_o[1181] = data_o_0__29_;
  assign data_o[1213] = data_o_0__29_;
  assign data_o[1245] = data_o_0__29_;
  assign data_o[1277] = data_o_0__29_;
  assign data_o[1309] = data_o_0__29_;
  assign data_o[1341] = data_o_0__29_;
  assign data_o[1373] = data_o_0__29_;
  assign data_o[1405] = data_o_0__29_;
  assign data_o[1437] = data_o_0__29_;
  assign data_o[1469] = data_o_0__29_;
  assign data_o[1501] = data_o_0__29_;
  assign data_o[1533] = data_o_0__29_;
  assign data_o[1565] = data_o_0__29_;
  assign data_o[1597] = data_o_0__29_;
  assign data_o[28] = data_o_0__28_;
  assign data_o[60] = data_o_0__28_;
  assign data_o[92] = data_o_0__28_;
  assign data_o[124] = data_o_0__28_;
  assign data_o[156] = data_o_0__28_;
  assign data_o[188] = data_o_0__28_;
  assign data_o[220] = data_o_0__28_;
  assign data_o[252] = data_o_0__28_;
  assign data_o[284] = data_o_0__28_;
  assign data_o[316] = data_o_0__28_;
  assign data_o[348] = data_o_0__28_;
  assign data_o[380] = data_o_0__28_;
  assign data_o[412] = data_o_0__28_;
  assign data_o[444] = data_o_0__28_;
  assign data_o[476] = data_o_0__28_;
  assign data_o[508] = data_o_0__28_;
  assign data_o[540] = data_o_0__28_;
  assign data_o[572] = data_o_0__28_;
  assign data_o[604] = data_o_0__28_;
  assign data_o[636] = data_o_0__28_;
  assign data_o[668] = data_o_0__28_;
  assign data_o[700] = data_o_0__28_;
  assign data_o[732] = data_o_0__28_;
  assign data_o[764] = data_o_0__28_;
  assign data_o[796] = data_o_0__28_;
  assign data_o[828] = data_o_0__28_;
  assign data_o[860] = data_o_0__28_;
  assign data_o[892] = data_o_0__28_;
  assign data_o[924] = data_o_0__28_;
  assign data_o[956] = data_o_0__28_;
  assign data_o[988] = data_o_0__28_;
  assign data_o[1020] = data_o_0__28_;
  assign data_o[1052] = data_o_0__28_;
  assign data_o[1084] = data_o_0__28_;
  assign data_o[1116] = data_o_0__28_;
  assign data_o[1148] = data_o_0__28_;
  assign data_o[1180] = data_o_0__28_;
  assign data_o[1212] = data_o_0__28_;
  assign data_o[1244] = data_o_0__28_;
  assign data_o[1276] = data_o_0__28_;
  assign data_o[1308] = data_o_0__28_;
  assign data_o[1340] = data_o_0__28_;
  assign data_o[1372] = data_o_0__28_;
  assign data_o[1404] = data_o_0__28_;
  assign data_o[1436] = data_o_0__28_;
  assign data_o[1468] = data_o_0__28_;
  assign data_o[1500] = data_o_0__28_;
  assign data_o[1532] = data_o_0__28_;
  assign data_o[1564] = data_o_0__28_;
  assign data_o[1596] = data_o_0__28_;
  assign data_o[27] = data_o_0__27_;
  assign data_o[59] = data_o_0__27_;
  assign data_o[91] = data_o_0__27_;
  assign data_o[123] = data_o_0__27_;
  assign data_o[155] = data_o_0__27_;
  assign data_o[187] = data_o_0__27_;
  assign data_o[219] = data_o_0__27_;
  assign data_o[251] = data_o_0__27_;
  assign data_o[283] = data_o_0__27_;
  assign data_o[315] = data_o_0__27_;
  assign data_o[347] = data_o_0__27_;
  assign data_o[379] = data_o_0__27_;
  assign data_o[411] = data_o_0__27_;
  assign data_o[443] = data_o_0__27_;
  assign data_o[475] = data_o_0__27_;
  assign data_o[507] = data_o_0__27_;
  assign data_o[539] = data_o_0__27_;
  assign data_o[571] = data_o_0__27_;
  assign data_o[603] = data_o_0__27_;
  assign data_o[635] = data_o_0__27_;
  assign data_o[667] = data_o_0__27_;
  assign data_o[699] = data_o_0__27_;
  assign data_o[731] = data_o_0__27_;
  assign data_o[763] = data_o_0__27_;
  assign data_o[795] = data_o_0__27_;
  assign data_o[827] = data_o_0__27_;
  assign data_o[859] = data_o_0__27_;
  assign data_o[891] = data_o_0__27_;
  assign data_o[923] = data_o_0__27_;
  assign data_o[955] = data_o_0__27_;
  assign data_o[987] = data_o_0__27_;
  assign data_o[1019] = data_o_0__27_;
  assign data_o[1051] = data_o_0__27_;
  assign data_o[1083] = data_o_0__27_;
  assign data_o[1115] = data_o_0__27_;
  assign data_o[1147] = data_o_0__27_;
  assign data_o[1179] = data_o_0__27_;
  assign data_o[1211] = data_o_0__27_;
  assign data_o[1243] = data_o_0__27_;
  assign data_o[1275] = data_o_0__27_;
  assign data_o[1307] = data_o_0__27_;
  assign data_o[1339] = data_o_0__27_;
  assign data_o[1371] = data_o_0__27_;
  assign data_o[1403] = data_o_0__27_;
  assign data_o[1435] = data_o_0__27_;
  assign data_o[1467] = data_o_0__27_;
  assign data_o[1499] = data_o_0__27_;
  assign data_o[1531] = data_o_0__27_;
  assign data_o[1563] = data_o_0__27_;
  assign data_o[1595] = data_o_0__27_;
  assign data_o[26] = data_o_0__26_;
  assign data_o[58] = data_o_0__26_;
  assign data_o[90] = data_o_0__26_;
  assign data_o[122] = data_o_0__26_;
  assign data_o[154] = data_o_0__26_;
  assign data_o[186] = data_o_0__26_;
  assign data_o[218] = data_o_0__26_;
  assign data_o[250] = data_o_0__26_;
  assign data_o[282] = data_o_0__26_;
  assign data_o[314] = data_o_0__26_;
  assign data_o[346] = data_o_0__26_;
  assign data_o[378] = data_o_0__26_;
  assign data_o[410] = data_o_0__26_;
  assign data_o[442] = data_o_0__26_;
  assign data_o[474] = data_o_0__26_;
  assign data_o[506] = data_o_0__26_;
  assign data_o[538] = data_o_0__26_;
  assign data_o[570] = data_o_0__26_;
  assign data_o[602] = data_o_0__26_;
  assign data_o[634] = data_o_0__26_;
  assign data_o[666] = data_o_0__26_;
  assign data_o[698] = data_o_0__26_;
  assign data_o[730] = data_o_0__26_;
  assign data_o[762] = data_o_0__26_;
  assign data_o[794] = data_o_0__26_;
  assign data_o[826] = data_o_0__26_;
  assign data_o[858] = data_o_0__26_;
  assign data_o[890] = data_o_0__26_;
  assign data_o[922] = data_o_0__26_;
  assign data_o[954] = data_o_0__26_;
  assign data_o[986] = data_o_0__26_;
  assign data_o[1018] = data_o_0__26_;
  assign data_o[1050] = data_o_0__26_;
  assign data_o[1082] = data_o_0__26_;
  assign data_o[1114] = data_o_0__26_;
  assign data_o[1146] = data_o_0__26_;
  assign data_o[1178] = data_o_0__26_;
  assign data_o[1210] = data_o_0__26_;
  assign data_o[1242] = data_o_0__26_;
  assign data_o[1274] = data_o_0__26_;
  assign data_o[1306] = data_o_0__26_;
  assign data_o[1338] = data_o_0__26_;
  assign data_o[1370] = data_o_0__26_;
  assign data_o[1402] = data_o_0__26_;
  assign data_o[1434] = data_o_0__26_;
  assign data_o[1466] = data_o_0__26_;
  assign data_o[1498] = data_o_0__26_;
  assign data_o[1530] = data_o_0__26_;
  assign data_o[1562] = data_o_0__26_;
  assign data_o[1594] = data_o_0__26_;
  assign data_o[25] = data_o_0__25_;
  assign data_o[57] = data_o_0__25_;
  assign data_o[89] = data_o_0__25_;
  assign data_o[121] = data_o_0__25_;
  assign data_o[153] = data_o_0__25_;
  assign data_o[185] = data_o_0__25_;
  assign data_o[217] = data_o_0__25_;
  assign data_o[249] = data_o_0__25_;
  assign data_o[281] = data_o_0__25_;
  assign data_o[313] = data_o_0__25_;
  assign data_o[345] = data_o_0__25_;
  assign data_o[377] = data_o_0__25_;
  assign data_o[409] = data_o_0__25_;
  assign data_o[441] = data_o_0__25_;
  assign data_o[473] = data_o_0__25_;
  assign data_o[505] = data_o_0__25_;
  assign data_o[537] = data_o_0__25_;
  assign data_o[569] = data_o_0__25_;
  assign data_o[601] = data_o_0__25_;
  assign data_o[633] = data_o_0__25_;
  assign data_o[665] = data_o_0__25_;
  assign data_o[697] = data_o_0__25_;
  assign data_o[729] = data_o_0__25_;
  assign data_o[761] = data_o_0__25_;
  assign data_o[793] = data_o_0__25_;
  assign data_o[825] = data_o_0__25_;
  assign data_o[857] = data_o_0__25_;
  assign data_o[889] = data_o_0__25_;
  assign data_o[921] = data_o_0__25_;
  assign data_o[953] = data_o_0__25_;
  assign data_o[985] = data_o_0__25_;
  assign data_o[1017] = data_o_0__25_;
  assign data_o[1049] = data_o_0__25_;
  assign data_o[1081] = data_o_0__25_;
  assign data_o[1113] = data_o_0__25_;
  assign data_o[1145] = data_o_0__25_;
  assign data_o[1177] = data_o_0__25_;
  assign data_o[1209] = data_o_0__25_;
  assign data_o[1241] = data_o_0__25_;
  assign data_o[1273] = data_o_0__25_;
  assign data_o[1305] = data_o_0__25_;
  assign data_o[1337] = data_o_0__25_;
  assign data_o[1369] = data_o_0__25_;
  assign data_o[1401] = data_o_0__25_;
  assign data_o[1433] = data_o_0__25_;
  assign data_o[1465] = data_o_0__25_;
  assign data_o[1497] = data_o_0__25_;
  assign data_o[1529] = data_o_0__25_;
  assign data_o[1561] = data_o_0__25_;
  assign data_o[1593] = data_o_0__25_;
  assign data_o[24] = data_o_0__24_;
  assign data_o[56] = data_o_0__24_;
  assign data_o[88] = data_o_0__24_;
  assign data_o[120] = data_o_0__24_;
  assign data_o[152] = data_o_0__24_;
  assign data_o[184] = data_o_0__24_;
  assign data_o[216] = data_o_0__24_;
  assign data_o[248] = data_o_0__24_;
  assign data_o[280] = data_o_0__24_;
  assign data_o[312] = data_o_0__24_;
  assign data_o[344] = data_o_0__24_;
  assign data_o[376] = data_o_0__24_;
  assign data_o[408] = data_o_0__24_;
  assign data_o[440] = data_o_0__24_;
  assign data_o[472] = data_o_0__24_;
  assign data_o[504] = data_o_0__24_;
  assign data_o[536] = data_o_0__24_;
  assign data_o[568] = data_o_0__24_;
  assign data_o[600] = data_o_0__24_;
  assign data_o[632] = data_o_0__24_;
  assign data_o[664] = data_o_0__24_;
  assign data_o[696] = data_o_0__24_;
  assign data_o[728] = data_o_0__24_;
  assign data_o[760] = data_o_0__24_;
  assign data_o[792] = data_o_0__24_;
  assign data_o[824] = data_o_0__24_;
  assign data_o[856] = data_o_0__24_;
  assign data_o[888] = data_o_0__24_;
  assign data_o[920] = data_o_0__24_;
  assign data_o[952] = data_o_0__24_;
  assign data_o[984] = data_o_0__24_;
  assign data_o[1016] = data_o_0__24_;
  assign data_o[1048] = data_o_0__24_;
  assign data_o[1080] = data_o_0__24_;
  assign data_o[1112] = data_o_0__24_;
  assign data_o[1144] = data_o_0__24_;
  assign data_o[1176] = data_o_0__24_;
  assign data_o[1208] = data_o_0__24_;
  assign data_o[1240] = data_o_0__24_;
  assign data_o[1272] = data_o_0__24_;
  assign data_o[1304] = data_o_0__24_;
  assign data_o[1336] = data_o_0__24_;
  assign data_o[1368] = data_o_0__24_;
  assign data_o[1400] = data_o_0__24_;
  assign data_o[1432] = data_o_0__24_;
  assign data_o[1464] = data_o_0__24_;
  assign data_o[1496] = data_o_0__24_;
  assign data_o[1528] = data_o_0__24_;
  assign data_o[1560] = data_o_0__24_;
  assign data_o[1592] = data_o_0__24_;
  assign data_o[23] = data_o_0__23_;
  assign data_o[55] = data_o_0__23_;
  assign data_o[87] = data_o_0__23_;
  assign data_o[119] = data_o_0__23_;
  assign data_o[151] = data_o_0__23_;
  assign data_o[183] = data_o_0__23_;
  assign data_o[215] = data_o_0__23_;
  assign data_o[247] = data_o_0__23_;
  assign data_o[279] = data_o_0__23_;
  assign data_o[311] = data_o_0__23_;
  assign data_o[343] = data_o_0__23_;
  assign data_o[375] = data_o_0__23_;
  assign data_o[407] = data_o_0__23_;
  assign data_o[439] = data_o_0__23_;
  assign data_o[471] = data_o_0__23_;
  assign data_o[503] = data_o_0__23_;
  assign data_o[535] = data_o_0__23_;
  assign data_o[567] = data_o_0__23_;
  assign data_o[599] = data_o_0__23_;
  assign data_o[631] = data_o_0__23_;
  assign data_o[663] = data_o_0__23_;
  assign data_o[695] = data_o_0__23_;
  assign data_o[727] = data_o_0__23_;
  assign data_o[759] = data_o_0__23_;
  assign data_o[791] = data_o_0__23_;
  assign data_o[823] = data_o_0__23_;
  assign data_o[855] = data_o_0__23_;
  assign data_o[887] = data_o_0__23_;
  assign data_o[919] = data_o_0__23_;
  assign data_o[951] = data_o_0__23_;
  assign data_o[983] = data_o_0__23_;
  assign data_o[1015] = data_o_0__23_;
  assign data_o[1047] = data_o_0__23_;
  assign data_o[1079] = data_o_0__23_;
  assign data_o[1111] = data_o_0__23_;
  assign data_o[1143] = data_o_0__23_;
  assign data_o[1175] = data_o_0__23_;
  assign data_o[1207] = data_o_0__23_;
  assign data_o[1239] = data_o_0__23_;
  assign data_o[1271] = data_o_0__23_;
  assign data_o[1303] = data_o_0__23_;
  assign data_o[1335] = data_o_0__23_;
  assign data_o[1367] = data_o_0__23_;
  assign data_o[1399] = data_o_0__23_;
  assign data_o[1431] = data_o_0__23_;
  assign data_o[1463] = data_o_0__23_;
  assign data_o[1495] = data_o_0__23_;
  assign data_o[1527] = data_o_0__23_;
  assign data_o[1559] = data_o_0__23_;
  assign data_o[1591] = data_o_0__23_;
  assign data_o[22] = data_o_0__22_;
  assign data_o[54] = data_o_0__22_;
  assign data_o[86] = data_o_0__22_;
  assign data_o[118] = data_o_0__22_;
  assign data_o[150] = data_o_0__22_;
  assign data_o[182] = data_o_0__22_;
  assign data_o[214] = data_o_0__22_;
  assign data_o[246] = data_o_0__22_;
  assign data_o[278] = data_o_0__22_;
  assign data_o[310] = data_o_0__22_;
  assign data_o[342] = data_o_0__22_;
  assign data_o[374] = data_o_0__22_;
  assign data_o[406] = data_o_0__22_;
  assign data_o[438] = data_o_0__22_;
  assign data_o[470] = data_o_0__22_;
  assign data_o[502] = data_o_0__22_;
  assign data_o[534] = data_o_0__22_;
  assign data_o[566] = data_o_0__22_;
  assign data_o[598] = data_o_0__22_;
  assign data_o[630] = data_o_0__22_;
  assign data_o[662] = data_o_0__22_;
  assign data_o[694] = data_o_0__22_;
  assign data_o[726] = data_o_0__22_;
  assign data_o[758] = data_o_0__22_;
  assign data_o[790] = data_o_0__22_;
  assign data_o[822] = data_o_0__22_;
  assign data_o[854] = data_o_0__22_;
  assign data_o[886] = data_o_0__22_;
  assign data_o[918] = data_o_0__22_;
  assign data_o[950] = data_o_0__22_;
  assign data_o[982] = data_o_0__22_;
  assign data_o[1014] = data_o_0__22_;
  assign data_o[1046] = data_o_0__22_;
  assign data_o[1078] = data_o_0__22_;
  assign data_o[1110] = data_o_0__22_;
  assign data_o[1142] = data_o_0__22_;
  assign data_o[1174] = data_o_0__22_;
  assign data_o[1206] = data_o_0__22_;
  assign data_o[1238] = data_o_0__22_;
  assign data_o[1270] = data_o_0__22_;
  assign data_o[1302] = data_o_0__22_;
  assign data_o[1334] = data_o_0__22_;
  assign data_o[1366] = data_o_0__22_;
  assign data_o[1398] = data_o_0__22_;
  assign data_o[1430] = data_o_0__22_;
  assign data_o[1462] = data_o_0__22_;
  assign data_o[1494] = data_o_0__22_;
  assign data_o[1526] = data_o_0__22_;
  assign data_o[1558] = data_o_0__22_;
  assign data_o[1590] = data_o_0__22_;
  assign data_o[21] = data_o_0__21_;
  assign data_o[53] = data_o_0__21_;
  assign data_o[85] = data_o_0__21_;
  assign data_o[117] = data_o_0__21_;
  assign data_o[149] = data_o_0__21_;
  assign data_o[181] = data_o_0__21_;
  assign data_o[213] = data_o_0__21_;
  assign data_o[245] = data_o_0__21_;
  assign data_o[277] = data_o_0__21_;
  assign data_o[309] = data_o_0__21_;
  assign data_o[341] = data_o_0__21_;
  assign data_o[373] = data_o_0__21_;
  assign data_o[405] = data_o_0__21_;
  assign data_o[437] = data_o_0__21_;
  assign data_o[469] = data_o_0__21_;
  assign data_o[501] = data_o_0__21_;
  assign data_o[533] = data_o_0__21_;
  assign data_o[565] = data_o_0__21_;
  assign data_o[597] = data_o_0__21_;
  assign data_o[629] = data_o_0__21_;
  assign data_o[661] = data_o_0__21_;
  assign data_o[693] = data_o_0__21_;
  assign data_o[725] = data_o_0__21_;
  assign data_o[757] = data_o_0__21_;
  assign data_o[789] = data_o_0__21_;
  assign data_o[821] = data_o_0__21_;
  assign data_o[853] = data_o_0__21_;
  assign data_o[885] = data_o_0__21_;
  assign data_o[917] = data_o_0__21_;
  assign data_o[949] = data_o_0__21_;
  assign data_o[981] = data_o_0__21_;
  assign data_o[1013] = data_o_0__21_;
  assign data_o[1045] = data_o_0__21_;
  assign data_o[1077] = data_o_0__21_;
  assign data_o[1109] = data_o_0__21_;
  assign data_o[1141] = data_o_0__21_;
  assign data_o[1173] = data_o_0__21_;
  assign data_o[1205] = data_o_0__21_;
  assign data_o[1237] = data_o_0__21_;
  assign data_o[1269] = data_o_0__21_;
  assign data_o[1301] = data_o_0__21_;
  assign data_o[1333] = data_o_0__21_;
  assign data_o[1365] = data_o_0__21_;
  assign data_o[1397] = data_o_0__21_;
  assign data_o[1429] = data_o_0__21_;
  assign data_o[1461] = data_o_0__21_;
  assign data_o[1493] = data_o_0__21_;
  assign data_o[1525] = data_o_0__21_;
  assign data_o[1557] = data_o_0__21_;
  assign data_o[1589] = data_o_0__21_;
  assign data_o[20] = data_o_0__20_;
  assign data_o[52] = data_o_0__20_;
  assign data_o[84] = data_o_0__20_;
  assign data_o[116] = data_o_0__20_;
  assign data_o[148] = data_o_0__20_;
  assign data_o[180] = data_o_0__20_;
  assign data_o[212] = data_o_0__20_;
  assign data_o[244] = data_o_0__20_;
  assign data_o[276] = data_o_0__20_;
  assign data_o[308] = data_o_0__20_;
  assign data_o[340] = data_o_0__20_;
  assign data_o[372] = data_o_0__20_;
  assign data_o[404] = data_o_0__20_;
  assign data_o[436] = data_o_0__20_;
  assign data_o[468] = data_o_0__20_;
  assign data_o[500] = data_o_0__20_;
  assign data_o[532] = data_o_0__20_;
  assign data_o[564] = data_o_0__20_;
  assign data_o[596] = data_o_0__20_;
  assign data_o[628] = data_o_0__20_;
  assign data_o[660] = data_o_0__20_;
  assign data_o[692] = data_o_0__20_;
  assign data_o[724] = data_o_0__20_;
  assign data_o[756] = data_o_0__20_;
  assign data_o[788] = data_o_0__20_;
  assign data_o[820] = data_o_0__20_;
  assign data_o[852] = data_o_0__20_;
  assign data_o[884] = data_o_0__20_;
  assign data_o[916] = data_o_0__20_;
  assign data_o[948] = data_o_0__20_;
  assign data_o[980] = data_o_0__20_;
  assign data_o[1012] = data_o_0__20_;
  assign data_o[1044] = data_o_0__20_;
  assign data_o[1076] = data_o_0__20_;
  assign data_o[1108] = data_o_0__20_;
  assign data_o[1140] = data_o_0__20_;
  assign data_o[1172] = data_o_0__20_;
  assign data_o[1204] = data_o_0__20_;
  assign data_o[1236] = data_o_0__20_;
  assign data_o[1268] = data_o_0__20_;
  assign data_o[1300] = data_o_0__20_;
  assign data_o[1332] = data_o_0__20_;
  assign data_o[1364] = data_o_0__20_;
  assign data_o[1396] = data_o_0__20_;
  assign data_o[1428] = data_o_0__20_;
  assign data_o[1460] = data_o_0__20_;
  assign data_o[1492] = data_o_0__20_;
  assign data_o[1524] = data_o_0__20_;
  assign data_o[1556] = data_o_0__20_;
  assign data_o[1588] = data_o_0__20_;
  assign data_o[19] = data_o_0__19_;
  assign data_o[51] = data_o_0__19_;
  assign data_o[83] = data_o_0__19_;
  assign data_o[115] = data_o_0__19_;
  assign data_o[147] = data_o_0__19_;
  assign data_o[179] = data_o_0__19_;
  assign data_o[211] = data_o_0__19_;
  assign data_o[243] = data_o_0__19_;
  assign data_o[275] = data_o_0__19_;
  assign data_o[307] = data_o_0__19_;
  assign data_o[339] = data_o_0__19_;
  assign data_o[371] = data_o_0__19_;
  assign data_o[403] = data_o_0__19_;
  assign data_o[435] = data_o_0__19_;
  assign data_o[467] = data_o_0__19_;
  assign data_o[499] = data_o_0__19_;
  assign data_o[531] = data_o_0__19_;
  assign data_o[563] = data_o_0__19_;
  assign data_o[595] = data_o_0__19_;
  assign data_o[627] = data_o_0__19_;
  assign data_o[659] = data_o_0__19_;
  assign data_o[691] = data_o_0__19_;
  assign data_o[723] = data_o_0__19_;
  assign data_o[755] = data_o_0__19_;
  assign data_o[787] = data_o_0__19_;
  assign data_o[819] = data_o_0__19_;
  assign data_o[851] = data_o_0__19_;
  assign data_o[883] = data_o_0__19_;
  assign data_o[915] = data_o_0__19_;
  assign data_o[947] = data_o_0__19_;
  assign data_o[979] = data_o_0__19_;
  assign data_o[1011] = data_o_0__19_;
  assign data_o[1043] = data_o_0__19_;
  assign data_o[1075] = data_o_0__19_;
  assign data_o[1107] = data_o_0__19_;
  assign data_o[1139] = data_o_0__19_;
  assign data_o[1171] = data_o_0__19_;
  assign data_o[1203] = data_o_0__19_;
  assign data_o[1235] = data_o_0__19_;
  assign data_o[1267] = data_o_0__19_;
  assign data_o[1299] = data_o_0__19_;
  assign data_o[1331] = data_o_0__19_;
  assign data_o[1363] = data_o_0__19_;
  assign data_o[1395] = data_o_0__19_;
  assign data_o[1427] = data_o_0__19_;
  assign data_o[1459] = data_o_0__19_;
  assign data_o[1491] = data_o_0__19_;
  assign data_o[1523] = data_o_0__19_;
  assign data_o[1555] = data_o_0__19_;
  assign data_o[1587] = data_o_0__19_;
  assign data_o[18] = data_o_0__18_;
  assign data_o[50] = data_o_0__18_;
  assign data_o[82] = data_o_0__18_;
  assign data_o[114] = data_o_0__18_;
  assign data_o[146] = data_o_0__18_;
  assign data_o[178] = data_o_0__18_;
  assign data_o[210] = data_o_0__18_;
  assign data_o[242] = data_o_0__18_;
  assign data_o[274] = data_o_0__18_;
  assign data_o[306] = data_o_0__18_;
  assign data_o[338] = data_o_0__18_;
  assign data_o[370] = data_o_0__18_;
  assign data_o[402] = data_o_0__18_;
  assign data_o[434] = data_o_0__18_;
  assign data_o[466] = data_o_0__18_;
  assign data_o[498] = data_o_0__18_;
  assign data_o[530] = data_o_0__18_;
  assign data_o[562] = data_o_0__18_;
  assign data_o[594] = data_o_0__18_;
  assign data_o[626] = data_o_0__18_;
  assign data_o[658] = data_o_0__18_;
  assign data_o[690] = data_o_0__18_;
  assign data_o[722] = data_o_0__18_;
  assign data_o[754] = data_o_0__18_;
  assign data_o[786] = data_o_0__18_;
  assign data_o[818] = data_o_0__18_;
  assign data_o[850] = data_o_0__18_;
  assign data_o[882] = data_o_0__18_;
  assign data_o[914] = data_o_0__18_;
  assign data_o[946] = data_o_0__18_;
  assign data_o[978] = data_o_0__18_;
  assign data_o[1010] = data_o_0__18_;
  assign data_o[1042] = data_o_0__18_;
  assign data_o[1074] = data_o_0__18_;
  assign data_o[1106] = data_o_0__18_;
  assign data_o[1138] = data_o_0__18_;
  assign data_o[1170] = data_o_0__18_;
  assign data_o[1202] = data_o_0__18_;
  assign data_o[1234] = data_o_0__18_;
  assign data_o[1266] = data_o_0__18_;
  assign data_o[1298] = data_o_0__18_;
  assign data_o[1330] = data_o_0__18_;
  assign data_o[1362] = data_o_0__18_;
  assign data_o[1394] = data_o_0__18_;
  assign data_o[1426] = data_o_0__18_;
  assign data_o[1458] = data_o_0__18_;
  assign data_o[1490] = data_o_0__18_;
  assign data_o[1522] = data_o_0__18_;
  assign data_o[1554] = data_o_0__18_;
  assign data_o[1586] = data_o_0__18_;
  assign data_o[17] = data_o_0__17_;
  assign data_o[49] = data_o_0__17_;
  assign data_o[81] = data_o_0__17_;
  assign data_o[113] = data_o_0__17_;
  assign data_o[145] = data_o_0__17_;
  assign data_o[177] = data_o_0__17_;
  assign data_o[209] = data_o_0__17_;
  assign data_o[241] = data_o_0__17_;
  assign data_o[273] = data_o_0__17_;
  assign data_o[305] = data_o_0__17_;
  assign data_o[337] = data_o_0__17_;
  assign data_o[369] = data_o_0__17_;
  assign data_o[401] = data_o_0__17_;
  assign data_o[433] = data_o_0__17_;
  assign data_o[465] = data_o_0__17_;
  assign data_o[497] = data_o_0__17_;
  assign data_o[529] = data_o_0__17_;
  assign data_o[561] = data_o_0__17_;
  assign data_o[593] = data_o_0__17_;
  assign data_o[625] = data_o_0__17_;
  assign data_o[657] = data_o_0__17_;
  assign data_o[689] = data_o_0__17_;
  assign data_o[721] = data_o_0__17_;
  assign data_o[753] = data_o_0__17_;
  assign data_o[785] = data_o_0__17_;
  assign data_o[817] = data_o_0__17_;
  assign data_o[849] = data_o_0__17_;
  assign data_o[881] = data_o_0__17_;
  assign data_o[913] = data_o_0__17_;
  assign data_o[945] = data_o_0__17_;
  assign data_o[977] = data_o_0__17_;
  assign data_o[1009] = data_o_0__17_;
  assign data_o[1041] = data_o_0__17_;
  assign data_o[1073] = data_o_0__17_;
  assign data_o[1105] = data_o_0__17_;
  assign data_o[1137] = data_o_0__17_;
  assign data_o[1169] = data_o_0__17_;
  assign data_o[1201] = data_o_0__17_;
  assign data_o[1233] = data_o_0__17_;
  assign data_o[1265] = data_o_0__17_;
  assign data_o[1297] = data_o_0__17_;
  assign data_o[1329] = data_o_0__17_;
  assign data_o[1361] = data_o_0__17_;
  assign data_o[1393] = data_o_0__17_;
  assign data_o[1425] = data_o_0__17_;
  assign data_o[1457] = data_o_0__17_;
  assign data_o[1489] = data_o_0__17_;
  assign data_o[1521] = data_o_0__17_;
  assign data_o[1553] = data_o_0__17_;
  assign data_o[1585] = data_o_0__17_;
  assign data_o[16] = data_o_0__16_;
  assign data_o[48] = data_o_0__16_;
  assign data_o[80] = data_o_0__16_;
  assign data_o[112] = data_o_0__16_;
  assign data_o[144] = data_o_0__16_;
  assign data_o[176] = data_o_0__16_;
  assign data_o[208] = data_o_0__16_;
  assign data_o[240] = data_o_0__16_;
  assign data_o[272] = data_o_0__16_;
  assign data_o[304] = data_o_0__16_;
  assign data_o[336] = data_o_0__16_;
  assign data_o[368] = data_o_0__16_;
  assign data_o[400] = data_o_0__16_;
  assign data_o[432] = data_o_0__16_;
  assign data_o[464] = data_o_0__16_;
  assign data_o[496] = data_o_0__16_;
  assign data_o[528] = data_o_0__16_;
  assign data_o[560] = data_o_0__16_;
  assign data_o[592] = data_o_0__16_;
  assign data_o[624] = data_o_0__16_;
  assign data_o[656] = data_o_0__16_;
  assign data_o[688] = data_o_0__16_;
  assign data_o[720] = data_o_0__16_;
  assign data_o[752] = data_o_0__16_;
  assign data_o[784] = data_o_0__16_;
  assign data_o[816] = data_o_0__16_;
  assign data_o[848] = data_o_0__16_;
  assign data_o[880] = data_o_0__16_;
  assign data_o[912] = data_o_0__16_;
  assign data_o[944] = data_o_0__16_;
  assign data_o[976] = data_o_0__16_;
  assign data_o[1008] = data_o_0__16_;
  assign data_o[1040] = data_o_0__16_;
  assign data_o[1072] = data_o_0__16_;
  assign data_o[1104] = data_o_0__16_;
  assign data_o[1136] = data_o_0__16_;
  assign data_o[1168] = data_o_0__16_;
  assign data_o[1200] = data_o_0__16_;
  assign data_o[1232] = data_o_0__16_;
  assign data_o[1264] = data_o_0__16_;
  assign data_o[1296] = data_o_0__16_;
  assign data_o[1328] = data_o_0__16_;
  assign data_o[1360] = data_o_0__16_;
  assign data_o[1392] = data_o_0__16_;
  assign data_o[1424] = data_o_0__16_;
  assign data_o[1456] = data_o_0__16_;
  assign data_o[1488] = data_o_0__16_;
  assign data_o[1520] = data_o_0__16_;
  assign data_o[1552] = data_o_0__16_;
  assign data_o[1584] = data_o_0__16_;
  assign data_o[15] = data_o_0__15_;
  assign data_o[47] = data_o_0__15_;
  assign data_o[79] = data_o_0__15_;
  assign data_o[111] = data_o_0__15_;
  assign data_o[143] = data_o_0__15_;
  assign data_o[175] = data_o_0__15_;
  assign data_o[207] = data_o_0__15_;
  assign data_o[239] = data_o_0__15_;
  assign data_o[271] = data_o_0__15_;
  assign data_o[303] = data_o_0__15_;
  assign data_o[335] = data_o_0__15_;
  assign data_o[367] = data_o_0__15_;
  assign data_o[399] = data_o_0__15_;
  assign data_o[431] = data_o_0__15_;
  assign data_o[463] = data_o_0__15_;
  assign data_o[495] = data_o_0__15_;
  assign data_o[527] = data_o_0__15_;
  assign data_o[559] = data_o_0__15_;
  assign data_o[591] = data_o_0__15_;
  assign data_o[623] = data_o_0__15_;
  assign data_o[655] = data_o_0__15_;
  assign data_o[687] = data_o_0__15_;
  assign data_o[719] = data_o_0__15_;
  assign data_o[751] = data_o_0__15_;
  assign data_o[783] = data_o_0__15_;
  assign data_o[815] = data_o_0__15_;
  assign data_o[847] = data_o_0__15_;
  assign data_o[879] = data_o_0__15_;
  assign data_o[911] = data_o_0__15_;
  assign data_o[943] = data_o_0__15_;
  assign data_o[975] = data_o_0__15_;
  assign data_o[1007] = data_o_0__15_;
  assign data_o[1039] = data_o_0__15_;
  assign data_o[1071] = data_o_0__15_;
  assign data_o[1103] = data_o_0__15_;
  assign data_o[1135] = data_o_0__15_;
  assign data_o[1167] = data_o_0__15_;
  assign data_o[1199] = data_o_0__15_;
  assign data_o[1231] = data_o_0__15_;
  assign data_o[1263] = data_o_0__15_;
  assign data_o[1295] = data_o_0__15_;
  assign data_o[1327] = data_o_0__15_;
  assign data_o[1359] = data_o_0__15_;
  assign data_o[1391] = data_o_0__15_;
  assign data_o[1423] = data_o_0__15_;
  assign data_o[1455] = data_o_0__15_;
  assign data_o[1487] = data_o_0__15_;
  assign data_o[1519] = data_o_0__15_;
  assign data_o[1551] = data_o_0__15_;
  assign data_o[1583] = data_o_0__15_;
  assign data_o[14] = data_o_0__14_;
  assign data_o[46] = data_o_0__14_;
  assign data_o[78] = data_o_0__14_;
  assign data_o[110] = data_o_0__14_;
  assign data_o[142] = data_o_0__14_;
  assign data_o[174] = data_o_0__14_;
  assign data_o[206] = data_o_0__14_;
  assign data_o[238] = data_o_0__14_;
  assign data_o[270] = data_o_0__14_;
  assign data_o[302] = data_o_0__14_;
  assign data_o[334] = data_o_0__14_;
  assign data_o[366] = data_o_0__14_;
  assign data_o[398] = data_o_0__14_;
  assign data_o[430] = data_o_0__14_;
  assign data_o[462] = data_o_0__14_;
  assign data_o[494] = data_o_0__14_;
  assign data_o[526] = data_o_0__14_;
  assign data_o[558] = data_o_0__14_;
  assign data_o[590] = data_o_0__14_;
  assign data_o[622] = data_o_0__14_;
  assign data_o[654] = data_o_0__14_;
  assign data_o[686] = data_o_0__14_;
  assign data_o[718] = data_o_0__14_;
  assign data_o[750] = data_o_0__14_;
  assign data_o[782] = data_o_0__14_;
  assign data_o[814] = data_o_0__14_;
  assign data_o[846] = data_o_0__14_;
  assign data_o[878] = data_o_0__14_;
  assign data_o[910] = data_o_0__14_;
  assign data_o[942] = data_o_0__14_;
  assign data_o[974] = data_o_0__14_;
  assign data_o[1006] = data_o_0__14_;
  assign data_o[1038] = data_o_0__14_;
  assign data_o[1070] = data_o_0__14_;
  assign data_o[1102] = data_o_0__14_;
  assign data_o[1134] = data_o_0__14_;
  assign data_o[1166] = data_o_0__14_;
  assign data_o[1198] = data_o_0__14_;
  assign data_o[1230] = data_o_0__14_;
  assign data_o[1262] = data_o_0__14_;
  assign data_o[1294] = data_o_0__14_;
  assign data_o[1326] = data_o_0__14_;
  assign data_o[1358] = data_o_0__14_;
  assign data_o[1390] = data_o_0__14_;
  assign data_o[1422] = data_o_0__14_;
  assign data_o[1454] = data_o_0__14_;
  assign data_o[1486] = data_o_0__14_;
  assign data_o[1518] = data_o_0__14_;
  assign data_o[1550] = data_o_0__14_;
  assign data_o[1582] = data_o_0__14_;
  assign data_o[13] = data_o_0__13_;
  assign data_o[45] = data_o_0__13_;
  assign data_o[77] = data_o_0__13_;
  assign data_o[109] = data_o_0__13_;
  assign data_o[141] = data_o_0__13_;
  assign data_o[173] = data_o_0__13_;
  assign data_o[205] = data_o_0__13_;
  assign data_o[237] = data_o_0__13_;
  assign data_o[269] = data_o_0__13_;
  assign data_o[301] = data_o_0__13_;
  assign data_o[333] = data_o_0__13_;
  assign data_o[365] = data_o_0__13_;
  assign data_o[397] = data_o_0__13_;
  assign data_o[429] = data_o_0__13_;
  assign data_o[461] = data_o_0__13_;
  assign data_o[493] = data_o_0__13_;
  assign data_o[525] = data_o_0__13_;
  assign data_o[557] = data_o_0__13_;
  assign data_o[589] = data_o_0__13_;
  assign data_o[621] = data_o_0__13_;
  assign data_o[653] = data_o_0__13_;
  assign data_o[685] = data_o_0__13_;
  assign data_o[717] = data_o_0__13_;
  assign data_o[749] = data_o_0__13_;
  assign data_o[781] = data_o_0__13_;
  assign data_o[813] = data_o_0__13_;
  assign data_o[845] = data_o_0__13_;
  assign data_o[877] = data_o_0__13_;
  assign data_o[909] = data_o_0__13_;
  assign data_o[941] = data_o_0__13_;
  assign data_o[973] = data_o_0__13_;
  assign data_o[1005] = data_o_0__13_;
  assign data_o[1037] = data_o_0__13_;
  assign data_o[1069] = data_o_0__13_;
  assign data_o[1101] = data_o_0__13_;
  assign data_o[1133] = data_o_0__13_;
  assign data_o[1165] = data_o_0__13_;
  assign data_o[1197] = data_o_0__13_;
  assign data_o[1229] = data_o_0__13_;
  assign data_o[1261] = data_o_0__13_;
  assign data_o[1293] = data_o_0__13_;
  assign data_o[1325] = data_o_0__13_;
  assign data_o[1357] = data_o_0__13_;
  assign data_o[1389] = data_o_0__13_;
  assign data_o[1421] = data_o_0__13_;
  assign data_o[1453] = data_o_0__13_;
  assign data_o[1485] = data_o_0__13_;
  assign data_o[1517] = data_o_0__13_;
  assign data_o[1549] = data_o_0__13_;
  assign data_o[1581] = data_o_0__13_;
  assign data_o[12] = data_o_0__12_;
  assign data_o[44] = data_o_0__12_;
  assign data_o[76] = data_o_0__12_;
  assign data_o[108] = data_o_0__12_;
  assign data_o[140] = data_o_0__12_;
  assign data_o[172] = data_o_0__12_;
  assign data_o[204] = data_o_0__12_;
  assign data_o[236] = data_o_0__12_;
  assign data_o[268] = data_o_0__12_;
  assign data_o[300] = data_o_0__12_;
  assign data_o[332] = data_o_0__12_;
  assign data_o[364] = data_o_0__12_;
  assign data_o[396] = data_o_0__12_;
  assign data_o[428] = data_o_0__12_;
  assign data_o[460] = data_o_0__12_;
  assign data_o[492] = data_o_0__12_;
  assign data_o[524] = data_o_0__12_;
  assign data_o[556] = data_o_0__12_;
  assign data_o[588] = data_o_0__12_;
  assign data_o[620] = data_o_0__12_;
  assign data_o[652] = data_o_0__12_;
  assign data_o[684] = data_o_0__12_;
  assign data_o[716] = data_o_0__12_;
  assign data_o[748] = data_o_0__12_;
  assign data_o[780] = data_o_0__12_;
  assign data_o[812] = data_o_0__12_;
  assign data_o[844] = data_o_0__12_;
  assign data_o[876] = data_o_0__12_;
  assign data_o[908] = data_o_0__12_;
  assign data_o[940] = data_o_0__12_;
  assign data_o[972] = data_o_0__12_;
  assign data_o[1004] = data_o_0__12_;
  assign data_o[1036] = data_o_0__12_;
  assign data_o[1068] = data_o_0__12_;
  assign data_o[1100] = data_o_0__12_;
  assign data_o[1132] = data_o_0__12_;
  assign data_o[1164] = data_o_0__12_;
  assign data_o[1196] = data_o_0__12_;
  assign data_o[1228] = data_o_0__12_;
  assign data_o[1260] = data_o_0__12_;
  assign data_o[1292] = data_o_0__12_;
  assign data_o[1324] = data_o_0__12_;
  assign data_o[1356] = data_o_0__12_;
  assign data_o[1388] = data_o_0__12_;
  assign data_o[1420] = data_o_0__12_;
  assign data_o[1452] = data_o_0__12_;
  assign data_o[1484] = data_o_0__12_;
  assign data_o[1516] = data_o_0__12_;
  assign data_o[1548] = data_o_0__12_;
  assign data_o[1580] = data_o_0__12_;
  assign data_o[11] = data_o_0__11_;
  assign data_o[43] = data_o_0__11_;
  assign data_o[75] = data_o_0__11_;
  assign data_o[107] = data_o_0__11_;
  assign data_o[139] = data_o_0__11_;
  assign data_o[171] = data_o_0__11_;
  assign data_o[203] = data_o_0__11_;
  assign data_o[235] = data_o_0__11_;
  assign data_o[267] = data_o_0__11_;
  assign data_o[299] = data_o_0__11_;
  assign data_o[331] = data_o_0__11_;
  assign data_o[363] = data_o_0__11_;
  assign data_o[395] = data_o_0__11_;
  assign data_o[427] = data_o_0__11_;
  assign data_o[459] = data_o_0__11_;
  assign data_o[491] = data_o_0__11_;
  assign data_o[523] = data_o_0__11_;
  assign data_o[555] = data_o_0__11_;
  assign data_o[587] = data_o_0__11_;
  assign data_o[619] = data_o_0__11_;
  assign data_o[651] = data_o_0__11_;
  assign data_o[683] = data_o_0__11_;
  assign data_o[715] = data_o_0__11_;
  assign data_o[747] = data_o_0__11_;
  assign data_o[779] = data_o_0__11_;
  assign data_o[811] = data_o_0__11_;
  assign data_o[843] = data_o_0__11_;
  assign data_o[875] = data_o_0__11_;
  assign data_o[907] = data_o_0__11_;
  assign data_o[939] = data_o_0__11_;
  assign data_o[971] = data_o_0__11_;
  assign data_o[1003] = data_o_0__11_;
  assign data_o[1035] = data_o_0__11_;
  assign data_o[1067] = data_o_0__11_;
  assign data_o[1099] = data_o_0__11_;
  assign data_o[1131] = data_o_0__11_;
  assign data_o[1163] = data_o_0__11_;
  assign data_o[1195] = data_o_0__11_;
  assign data_o[1227] = data_o_0__11_;
  assign data_o[1259] = data_o_0__11_;
  assign data_o[1291] = data_o_0__11_;
  assign data_o[1323] = data_o_0__11_;
  assign data_o[1355] = data_o_0__11_;
  assign data_o[1387] = data_o_0__11_;
  assign data_o[1419] = data_o_0__11_;
  assign data_o[1451] = data_o_0__11_;
  assign data_o[1483] = data_o_0__11_;
  assign data_o[1515] = data_o_0__11_;
  assign data_o[1547] = data_o_0__11_;
  assign data_o[1579] = data_o_0__11_;
  assign data_o[10] = data_o_0__10_;
  assign data_o[42] = data_o_0__10_;
  assign data_o[74] = data_o_0__10_;
  assign data_o[106] = data_o_0__10_;
  assign data_o[138] = data_o_0__10_;
  assign data_o[170] = data_o_0__10_;
  assign data_o[202] = data_o_0__10_;
  assign data_o[234] = data_o_0__10_;
  assign data_o[266] = data_o_0__10_;
  assign data_o[298] = data_o_0__10_;
  assign data_o[330] = data_o_0__10_;
  assign data_o[362] = data_o_0__10_;
  assign data_o[394] = data_o_0__10_;
  assign data_o[426] = data_o_0__10_;
  assign data_o[458] = data_o_0__10_;
  assign data_o[490] = data_o_0__10_;
  assign data_o[522] = data_o_0__10_;
  assign data_o[554] = data_o_0__10_;
  assign data_o[586] = data_o_0__10_;
  assign data_o[618] = data_o_0__10_;
  assign data_o[650] = data_o_0__10_;
  assign data_o[682] = data_o_0__10_;
  assign data_o[714] = data_o_0__10_;
  assign data_o[746] = data_o_0__10_;
  assign data_o[778] = data_o_0__10_;
  assign data_o[810] = data_o_0__10_;
  assign data_o[842] = data_o_0__10_;
  assign data_o[874] = data_o_0__10_;
  assign data_o[906] = data_o_0__10_;
  assign data_o[938] = data_o_0__10_;
  assign data_o[970] = data_o_0__10_;
  assign data_o[1002] = data_o_0__10_;
  assign data_o[1034] = data_o_0__10_;
  assign data_o[1066] = data_o_0__10_;
  assign data_o[1098] = data_o_0__10_;
  assign data_o[1130] = data_o_0__10_;
  assign data_o[1162] = data_o_0__10_;
  assign data_o[1194] = data_o_0__10_;
  assign data_o[1226] = data_o_0__10_;
  assign data_o[1258] = data_o_0__10_;
  assign data_o[1290] = data_o_0__10_;
  assign data_o[1322] = data_o_0__10_;
  assign data_o[1354] = data_o_0__10_;
  assign data_o[1386] = data_o_0__10_;
  assign data_o[1418] = data_o_0__10_;
  assign data_o[1450] = data_o_0__10_;
  assign data_o[1482] = data_o_0__10_;
  assign data_o[1514] = data_o_0__10_;
  assign data_o[1546] = data_o_0__10_;
  assign data_o[1578] = data_o_0__10_;
  assign data_o[9] = data_o_0__9_;
  assign data_o[41] = data_o_0__9_;
  assign data_o[73] = data_o_0__9_;
  assign data_o[105] = data_o_0__9_;
  assign data_o[137] = data_o_0__9_;
  assign data_o[169] = data_o_0__9_;
  assign data_o[201] = data_o_0__9_;
  assign data_o[233] = data_o_0__9_;
  assign data_o[265] = data_o_0__9_;
  assign data_o[297] = data_o_0__9_;
  assign data_o[329] = data_o_0__9_;
  assign data_o[361] = data_o_0__9_;
  assign data_o[393] = data_o_0__9_;
  assign data_o[425] = data_o_0__9_;
  assign data_o[457] = data_o_0__9_;
  assign data_o[489] = data_o_0__9_;
  assign data_o[521] = data_o_0__9_;
  assign data_o[553] = data_o_0__9_;
  assign data_o[585] = data_o_0__9_;
  assign data_o[617] = data_o_0__9_;
  assign data_o[649] = data_o_0__9_;
  assign data_o[681] = data_o_0__9_;
  assign data_o[713] = data_o_0__9_;
  assign data_o[745] = data_o_0__9_;
  assign data_o[777] = data_o_0__9_;
  assign data_o[809] = data_o_0__9_;
  assign data_o[841] = data_o_0__9_;
  assign data_o[873] = data_o_0__9_;
  assign data_o[905] = data_o_0__9_;
  assign data_o[937] = data_o_0__9_;
  assign data_o[969] = data_o_0__9_;
  assign data_o[1001] = data_o_0__9_;
  assign data_o[1033] = data_o_0__9_;
  assign data_o[1065] = data_o_0__9_;
  assign data_o[1097] = data_o_0__9_;
  assign data_o[1129] = data_o_0__9_;
  assign data_o[1161] = data_o_0__9_;
  assign data_o[1193] = data_o_0__9_;
  assign data_o[1225] = data_o_0__9_;
  assign data_o[1257] = data_o_0__9_;
  assign data_o[1289] = data_o_0__9_;
  assign data_o[1321] = data_o_0__9_;
  assign data_o[1353] = data_o_0__9_;
  assign data_o[1385] = data_o_0__9_;
  assign data_o[1417] = data_o_0__9_;
  assign data_o[1449] = data_o_0__9_;
  assign data_o[1481] = data_o_0__9_;
  assign data_o[1513] = data_o_0__9_;
  assign data_o[1545] = data_o_0__9_;
  assign data_o[1577] = data_o_0__9_;
  assign data_o[8] = data_o_0__8_;
  assign data_o[40] = data_o_0__8_;
  assign data_o[72] = data_o_0__8_;
  assign data_o[104] = data_o_0__8_;
  assign data_o[136] = data_o_0__8_;
  assign data_o[168] = data_o_0__8_;
  assign data_o[200] = data_o_0__8_;
  assign data_o[232] = data_o_0__8_;
  assign data_o[264] = data_o_0__8_;
  assign data_o[296] = data_o_0__8_;
  assign data_o[328] = data_o_0__8_;
  assign data_o[360] = data_o_0__8_;
  assign data_o[392] = data_o_0__8_;
  assign data_o[424] = data_o_0__8_;
  assign data_o[456] = data_o_0__8_;
  assign data_o[488] = data_o_0__8_;
  assign data_o[520] = data_o_0__8_;
  assign data_o[552] = data_o_0__8_;
  assign data_o[584] = data_o_0__8_;
  assign data_o[616] = data_o_0__8_;
  assign data_o[648] = data_o_0__8_;
  assign data_o[680] = data_o_0__8_;
  assign data_o[712] = data_o_0__8_;
  assign data_o[744] = data_o_0__8_;
  assign data_o[776] = data_o_0__8_;
  assign data_o[808] = data_o_0__8_;
  assign data_o[840] = data_o_0__8_;
  assign data_o[872] = data_o_0__8_;
  assign data_o[904] = data_o_0__8_;
  assign data_o[936] = data_o_0__8_;
  assign data_o[968] = data_o_0__8_;
  assign data_o[1000] = data_o_0__8_;
  assign data_o[1032] = data_o_0__8_;
  assign data_o[1064] = data_o_0__8_;
  assign data_o[1096] = data_o_0__8_;
  assign data_o[1128] = data_o_0__8_;
  assign data_o[1160] = data_o_0__8_;
  assign data_o[1192] = data_o_0__8_;
  assign data_o[1224] = data_o_0__8_;
  assign data_o[1256] = data_o_0__8_;
  assign data_o[1288] = data_o_0__8_;
  assign data_o[1320] = data_o_0__8_;
  assign data_o[1352] = data_o_0__8_;
  assign data_o[1384] = data_o_0__8_;
  assign data_o[1416] = data_o_0__8_;
  assign data_o[1448] = data_o_0__8_;
  assign data_o[1480] = data_o_0__8_;
  assign data_o[1512] = data_o_0__8_;
  assign data_o[1544] = data_o_0__8_;
  assign data_o[1576] = data_o_0__8_;
  assign data_o[7] = data_o_0__7_;
  assign data_o[39] = data_o_0__7_;
  assign data_o[71] = data_o_0__7_;
  assign data_o[103] = data_o_0__7_;
  assign data_o[135] = data_o_0__7_;
  assign data_o[167] = data_o_0__7_;
  assign data_o[199] = data_o_0__7_;
  assign data_o[231] = data_o_0__7_;
  assign data_o[263] = data_o_0__7_;
  assign data_o[295] = data_o_0__7_;
  assign data_o[327] = data_o_0__7_;
  assign data_o[359] = data_o_0__7_;
  assign data_o[391] = data_o_0__7_;
  assign data_o[423] = data_o_0__7_;
  assign data_o[455] = data_o_0__7_;
  assign data_o[487] = data_o_0__7_;
  assign data_o[519] = data_o_0__7_;
  assign data_o[551] = data_o_0__7_;
  assign data_o[583] = data_o_0__7_;
  assign data_o[615] = data_o_0__7_;
  assign data_o[647] = data_o_0__7_;
  assign data_o[679] = data_o_0__7_;
  assign data_o[711] = data_o_0__7_;
  assign data_o[743] = data_o_0__7_;
  assign data_o[775] = data_o_0__7_;
  assign data_o[807] = data_o_0__7_;
  assign data_o[839] = data_o_0__7_;
  assign data_o[871] = data_o_0__7_;
  assign data_o[903] = data_o_0__7_;
  assign data_o[935] = data_o_0__7_;
  assign data_o[967] = data_o_0__7_;
  assign data_o[999] = data_o_0__7_;
  assign data_o[1031] = data_o_0__7_;
  assign data_o[1063] = data_o_0__7_;
  assign data_o[1095] = data_o_0__7_;
  assign data_o[1127] = data_o_0__7_;
  assign data_o[1159] = data_o_0__7_;
  assign data_o[1191] = data_o_0__7_;
  assign data_o[1223] = data_o_0__7_;
  assign data_o[1255] = data_o_0__7_;
  assign data_o[1287] = data_o_0__7_;
  assign data_o[1319] = data_o_0__7_;
  assign data_o[1351] = data_o_0__7_;
  assign data_o[1383] = data_o_0__7_;
  assign data_o[1415] = data_o_0__7_;
  assign data_o[1447] = data_o_0__7_;
  assign data_o[1479] = data_o_0__7_;
  assign data_o[1511] = data_o_0__7_;
  assign data_o[1543] = data_o_0__7_;
  assign data_o[1575] = data_o_0__7_;
  assign data_o[6] = data_o_0__6_;
  assign data_o[38] = data_o_0__6_;
  assign data_o[70] = data_o_0__6_;
  assign data_o[102] = data_o_0__6_;
  assign data_o[134] = data_o_0__6_;
  assign data_o[166] = data_o_0__6_;
  assign data_o[198] = data_o_0__6_;
  assign data_o[230] = data_o_0__6_;
  assign data_o[262] = data_o_0__6_;
  assign data_o[294] = data_o_0__6_;
  assign data_o[326] = data_o_0__6_;
  assign data_o[358] = data_o_0__6_;
  assign data_o[390] = data_o_0__6_;
  assign data_o[422] = data_o_0__6_;
  assign data_o[454] = data_o_0__6_;
  assign data_o[486] = data_o_0__6_;
  assign data_o[518] = data_o_0__6_;
  assign data_o[550] = data_o_0__6_;
  assign data_o[582] = data_o_0__6_;
  assign data_o[614] = data_o_0__6_;
  assign data_o[646] = data_o_0__6_;
  assign data_o[678] = data_o_0__6_;
  assign data_o[710] = data_o_0__6_;
  assign data_o[742] = data_o_0__6_;
  assign data_o[774] = data_o_0__6_;
  assign data_o[806] = data_o_0__6_;
  assign data_o[838] = data_o_0__6_;
  assign data_o[870] = data_o_0__6_;
  assign data_o[902] = data_o_0__6_;
  assign data_o[934] = data_o_0__6_;
  assign data_o[966] = data_o_0__6_;
  assign data_o[998] = data_o_0__6_;
  assign data_o[1030] = data_o_0__6_;
  assign data_o[1062] = data_o_0__6_;
  assign data_o[1094] = data_o_0__6_;
  assign data_o[1126] = data_o_0__6_;
  assign data_o[1158] = data_o_0__6_;
  assign data_o[1190] = data_o_0__6_;
  assign data_o[1222] = data_o_0__6_;
  assign data_o[1254] = data_o_0__6_;
  assign data_o[1286] = data_o_0__6_;
  assign data_o[1318] = data_o_0__6_;
  assign data_o[1350] = data_o_0__6_;
  assign data_o[1382] = data_o_0__6_;
  assign data_o[1414] = data_o_0__6_;
  assign data_o[1446] = data_o_0__6_;
  assign data_o[1478] = data_o_0__6_;
  assign data_o[1510] = data_o_0__6_;
  assign data_o[1542] = data_o_0__6_;
  assign data_o[1574] = data_o_0__6_;
  assign data_o[5] = data_o_0__5_;
  assign data_o[37] = data_o_0__5_;
  assign data_o[69] = data_o_0__5_;
  assign data_o[101] = data_o_0__5_;
  assign data_o[133] = data_o_0__5_;
  assign data_o[165] = data_o_0__5_;
  assign data_o[197] = data_o_0__5_;
  assign data_o[229] = data_o_0__5_;
  assign data_o[261] = data_o_0__5_;
  assign data_o[293] = data_o_0__5_;
  assign data_o[325] = data_o_0__5_;
  assign data_o[357] = data_o_0__5_;
  assign data_o[389] = data_o_0__5_;
  assign data_o[421] = data_o_0__5_;
  assign data_o[453] = data_o_0__5_;
  assign data_o[485] = data_o_0__5_;
  assign data_o[517] = data_o_0__5_;
  assign data_o[549] = data_o_0__5_;
  assign data_o[581] = data_o_0__5_;
  assign data_o[613] = data_o_0__5_;
  assign data_o[645] = data_o_0__5_;
  assign data_o[677] = data_o_0__5_;
  assign data_o[709] = data_o_0__5_;
  assign data_o[741] = data_o_0__5_;
  assign data_o[773] = data_o_0__5_;
  assign data_o[805] = data_o_0__5_;
  assign data_o[837] = data_o_0__5_;
  assign data_o[869] = data_o_0__5_;
  assign data_o[901] = data_o_0__5_;
  assign data_o[933] = data_o_0__5_;
  assign data_o[965] = data_o_0__5_;
  assign data_o[997] = data_o_0__5_;
  assign data_o[1029] = data_o_0__5_;
  assign data_o[1061] = data_o_0__5_;
  assign data_o[1093] = data_o_0__5_;
  assign data_o[1125] = data_o_0__5_;
  assign data_o[1157] = data_o_0__5_;
  assign data_o[1189] = data_o_0__5_;
  assign data_o[1221] = data_o_0__5_;
  assign data_o[1253] = data_o_0__5_;
  assign data_o[1285] = data_o_0__5_;
  assign data_o[1317] = data_o_0__5_;
  assign data_o[1349] = data_o_0__5_;
  assign data_o[1381] = data_o_0__5_;
  assign data_o[1413] = data_o_0__5_;
  assign data_o[1445] = data_o_0__5_;
  assign data_o[1477] = data_o_0__5_;
  assign data_o[1509] = data_o_0__5_;
  assign data_o[1541] = data_o_0__5_;
  assign data_o[1573] = data_o_0__5_;
  assign data_o[4] = data_o_0__4_;
  assign data_o[36] = data_o_0__4_;
  assign data_o[68] = data_o_0__4_;
  assign data_o[100] = data_o_0__4_;
  assign data_o[132] = data_o_0__4_;
  assign data_o[164] = data_o_0__4_;
  assign data_o[196] = data_o_0__4_;
  assign data_o[228] = data_o_0__4_;
  assign data_o[260] = data_o_0__4_;
  assign data_o[292] = data_o_0__4_;
  assign data_o[324] = data_o_0__4_;
  assign data_o[356] = data_o_0__4_;
  assign data_o[388] = data_o_0__4_;
  assign data_o[420] = data_o_0__4_;
  assign data_o[452] = data_o_0__4_;
  assign data_o[484] = data_o_0__4_;
  assign data_o[516] = data_o_0__4_;
  assign data_o[548] = data_o_0__4_;
  assign data_o[580] = data_o_0__4_;
  assign data_o[612] = data_o_0__4_;
  assign data_o[644] = data_o_0__4_;
  assign data_o[676] = data_o_0__4_;
  assign data_o[708] = data_o_0__4_;
  assign data_o[740] = data_o_0__4_;
  assign data_o[772] = data_o_0__4_;
  assign data_o[804] = data_o_0__4_;
  assign data_o[836] = data_o_0__4_;
  assign data_o[868] = data_o_0__4_;
  assign data_o[900] = data_o_0__4_;
  assign data_o[932] = data_o_0__4_;
  assign data_o[964] = data_o_0__4_;
  assign data_o[996] = data_o_0__4_;
  assign data_o[1028] = data_o_0__4_;
  assign data_o[1060] = data_o_0__4_;
  assign data_o[1092] = data_o_0__4_;
  assign data_o[1124] = data_o_0__4_;
  assign data_o[1156] = data_o_0__4_;
  assign data_o[1188] = data_o_0__4_;
  assign data_o[1220] = data_o_0__4_;
  assign data_o[1252] = data_o_0__4_;
  assign data_o[1284] = data_o_0__4_;
  assign data_o[1316] = data_o_0__4_;
  assign data_o[1348] = data_o_0__4_;
  assign data_o[1380] = data_o_0__4_;
  assign data_o[1412] = data_o_0__4_;
  assign data_o[1444] = data_o_0__4_;
  assign data_o[1476] = data_o_0__4_;
  assign data_o[1508] = data_o_0__4_;
  assign data_o[1540] = data_o_0__4_;
  assign data_o[1572] = data_o_0__4_;
  assign data_o[3] = data_o_0__3_;
  assign data_o[35] = data_o_0__3_;
  assign data_o[67] = data_o_0__3_;
  assign data_o[99] = data_o_0__3_;
  assign data_o[131] = data_o_0__3_;
  assign data_o[163] = data_o_0__3_;
  assign data_o[195] = data_o_0__3_;
  assign data_o[227] = data_o_0__3_;
  assign data_o[259] = data_o_0__3_;
  assign data_o[291] = data_o_0__3_;
  assign data_o[323] = data_o_0__3_;
  assign data_o[355] = data_o_0__3_;
  assign data_o[387] = data_o_0__3_;
  assign data_o[419] = data_o_0__3_;
  assign data_o[451] = data_o_0__3_;
  assign data_o[483] = data_o_0__3_;
  assign data_o[515] = data_o_0__3_;
  assign data_o[547] = data_o_0__3_;
  assign data_o[579] = data_o_0__3_;
  assign data_o[611] = data_o_0__3_;
  assign data_o[643] = data_o_0__3_;
  assign data_o[675] = data_o_0__3_;
  assign data_o[707] = data_o_0__3_;
  assign data_o[739] = data_o_0__3_;
  assign data_o[771] = data_o_0__3_;
  assign data_o[803] = data_o_0__3_;
  assign data_o[835] = data_o_0__3_;
  assign data_o[867] = data_o_0__3_;
  assign data_o[899] = data_o_0__3_;
  assign data_o[931] = data_o_0__3_;
  assign data_o[963] = data_o_0__3_;
  assign data_o[995] = data_o_0__3_;
  assign data_o[1027] = data_o_0__3_;
  assign data_o[1059] = data_o_0__3_;
  assign data_o[1091] = data_o_0__3_;
  assign data_o[1123] = data_o_0__3_;
  assign data_o[1155] = data_o_0__3_;
  assign data_o[1187] = data_o_0__3_;
  assign data_o[1219] = data_o_0__3_;
  assign data_o[1251] = data_o_0__3_;
  assign data_o[1283] = data_o_0__3_;
  assign data_o[1315] = data_o_0__3_;
  assign data_o[1347] = data_o_0__3_;
  assign data_o[1379] = data_o_0__3_;
  assign data_o[1411] = data_o_0__3_;
  assign data_o[1443] = data_o_0__3_;
  assign data_o[1475] = data_o_0__3_;
  assign data_o[1507] = data_o_0__3_;
  assign data_o[1539] = data_o_0__3_;
  assign data_o[1571] = data_o_0__3_;
  assign data_o[2] = data_o_0__2_;
  assign data_o[34] = data_o_0__2_;
  assign data_o[66] = data_o_0__2_;
  assign data_o[98] = data_o_0__2_;
  assign data_o[130] = data_o_0__2_;
  assign data_o[162] = data_o_0__2_;
  assign data_o[194] = data_o_0__2_;
  assign data_o[226] = data_o_0__2_;
  assign data_o[258] = data_o_0__2_;
  assign data_o[290] = data_o_0__2_;
  assign data_o[322] = data_o_0__2_;
  assign data_o[354] = data_o_0__2_;
  assign data_o[386] = data_o_0__2_;
  assign data_o[418] = data_o_0__2_;
  assign data_o[450] = data_o_0__2_;
  assign data_o[482] = data_o_0__2_;
  assign data_o[514] = data_o_0__2_;
  assign data_o[546] = data_o_0__2_;
  assign data_o[578] = data_o_0__2_;
  assign data_o[610] = data_o_0__2_;
  assign data_o[642] = data_o_0__2_;
  assign data_o[674] = data_o_0__2_;
  assign data_o[706] = data_o_0__2_;
  assign data_o[738] = data_o_0__2_;
  assign data_o[770] = data_o_0__2_;
  assign data_o[802] = data_o_0__2_;
  assign data_o[834] = data_o_0__2_;
  assign data_o[866] = data_o_0__2_;
  assign data_o[898] = data_o_0__2_;
  assign data_o[930] = data_o_0__2_;
  assign data_o[962] = data_o_0__2_;
  assign data_o[994] = data_o_0__2_;
  assign data_o[1026] = data_o_0__2_;
  assign data_o[1058] = data_o_0__2_;
  assign data_o[1090] = data_o_0__2_;
  assign data_o[1122] = data_o_0__2_;
  assign data_o[1154] = data_o_0__2_;
  assign data_o[1186] = data_o_0__2_;
  assign data_o[1218] = data_o_0__2_;
  assign data_o[1250] = data_o_0__2_;
  assign data_o[1282] = data_o_0__2_;
  assign data_o[1314] = data_o_0__2_;
  assign data_o[1346] = data_o_0__2_;
  assign data_o[1378] = data_o_0__2_;
  assign data_o[1410] = data_o_0__2_;
  assign data_o[1442] = data_o_0__2_;
  assign data_o[1474] = data_o_0__2_;
  assign data_o[1506] = data_o_0__2_;
  assign data_o[1538] = data_o_0__2_;
  assign data_o[1570] = data_o_0__2_;
  assign data_o[1] = data_o_0__1_;
  assign data_o[33] = data_o_0__1_;
  assign data_o[65] = data_o_0__1_;
  assign data_o[97] = data_o_0__1_;
  assign data_o[129] = data_o_0__1_;
  assign data_o[161] = data_o_0__1_;
  assign data_o[193] = data_o_0__1_;
  assign data_o[225] = data_o_0__1_;
  assign data_o[257] = data_o_0__1_;
  assign data_o[289] = data_o_0__1_;
  assign data_o[321] = data_o_0__1_;
  assign data_o[353] = data_o_0__1_;
  assign data_o[385] = data_o_0__1_;
  assign data_o[417] = data_o_0__1_;
  assign data_o[449] = data_o_0__1_;
  assign data_o[481] = data_o_0__1_;
  assign data_o[513] = data_o_0__1_;
  assign data_o[545] = data_o_0__1_;
  assign data_o[577] = data_o_0__1_;
  assign data_o[609] = data_o_0__1_;
  assign data_o[641] = data_o_0__1_;
  assign data_o[673] = data_o_0__1_;
  assign data_o[705] = data_o_0__1_;
  assign data_o[737] = data_o_0__1_;
  assign data_o[769] = data_o_0__1_;
  assign data_o[801] = data_o_0__1_;
  assign data_o[833] = data_o_0__1_;
  assign data_o[865] = data_o_0__1_;
  assign data_o[897] = data_o_0__1_;
  assign data_o[929] = data_o_0__1_;
  assign data_o[961] = data_o_0__1_;
  assign data_o[993] = data_o_0__1_;
  assign data_o[1025] = data_o_0__1_;
  assign data_o[1057] = data_o_0__1_;
  assign data_o[1089] = data_o_0__1_;
  assign data_o[1121] = data_o_0__1_;
  assign data_o[1153] = data_o_0__1_;
  assign data_o[1185] = data_o_0__1_;
  assign data_o[1217] = data_o_0__1_;
  assign data_o[1249] = data_o_0__1_;
  assign data_o[1281] = data_o_0__1_;
  assign data_o[1313] = data_o_0__1_;
  assign data_o[1345] = data_o_0__1_;
  assign data_o[1377] = data_o_0__1_;
  assign data_o[1409] = data_o_0__1_;
  assign data_o[1441] = data_o_0__1_;
  assign data_o[1473] = data_o_0__1_;
  assign data_o[1505] = data_o_0__1_;
  assign data_o[1537] = data_o_0__1_;
  assign data_o[1569] = data_o_0__1_;
  assign data_o[0] = data_o_0__0_;
  assign data_o[32] = data_o_0__0_;
  assign data_o[64] = data_o_0__0_;
  assign data_o[96] = data_o_0__0_;
  assign data_o[128] = data_o_0__0_;
  assign data_o[160] = data_o_0__0_;
  assign data_o[192] = data_o_0__0_;
  assign data_o[224] = data_o_0__0_;
  assign data_o[256] = data_o_0__0_;
  assign data_o[288] = data_o_0__0_;
  assign data_o[320] = data_o_0__0_;
  assign data_o[352] = data_o_0__0_;
  assign data_o[384] = data_o_0__0_;
  assign data_o[416] = data_o_0__0_;
  assign data_o[448] = data_o_0__0_;
  assign data_o[480] = data_o_0__0_;
  assign data_o[512] = data_o_0__0_;
  assign data_o[544] = data_o_0__0_;
  assign data_o[576] = data_o_0__0_;
  assign data_o[608] = data_o_0__0_;
  assign data_o[640] = data_o_0__0_;
  assign data_o[672] = data_o_0__0_;
  assign data_o[704] = data_o_0__0_;
  assign data_o[736] = data_o_0__0_;
  assign data_o[768] = data_o_0__0_;
  assign data_o[800] = data_o_0__0_;
  assign data_o[832] = data_o_0__0_;
  assign data_o[864] = data_o_0__0_;
  assign data_o[896] = data_o_0__0_;
  assign data_o[928] = data_o_0__0_;
  assign data_o[960] = data_o_0__0_;
  assign data_o[992] = data_o_0__0_;
  assign data_o[1024] = data_o_0__0_;
  assign data_o[1056] = data_o_0__0_;
  assign data_o[1088] = data_o_0__0_;
  assign data_o[1120] = data_o_0__0_;
  assign data_o[1152] = data_o_0__0_;
  assign data_o[1184] = data_o_0__0_;
  assign data_o[1216] = data_o_0__0_;
  assign data_o[1248] = data_o_0__0_;
  assign data_o[1280] = data_o_0__0_;
  assign data_o[1312] = data_o_0__0_;
  assign data_o[1344] = data_o_0__0_;
  assign data_o[1376] = data_o_0__0_;
  assign data_o[1408] = data_o_0__0_;
  assign data_o[1440] = data_o_0__0_;
  assign data_o[1472] = data_o_0__0_;
  assign data_o[1504] = data_o_0__0_;
  assign data_o[1536] = data_o_0__0_;
  assign data_o[1568] = data_o_0__0_;

  bsg_two_fifo_width_p32
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_i(v_i),
    .v_o(fifo_v),
    .data_o({ data_o_0__31_, data_o_0__30_, data_o_0__29_, data_o_0__28_, data_o_0__27_, data_o_0__26_, data_o_0__25_, data_o_0__24_, data_o_0__23_, data_o_0__22_, data_o_0__21_, data_o_0__20_, data_o_0__19_, data_o_0__18_, data_o_0__17_, data_o_0__16_, data_o_0__15_, data_o_0__14_, data_o_0__13_, data_o_0__12_, data_o_0__11_, data_o_0__10_, data_o_0__9_, data_o_0__8_, data_o_0__7_, data_o_0__6_, data_o_0__5_, data_o_0__4_, data_o_0__3_, data_o_0__2_, data_o_0__1_, data_o_0__0_ }),
    .yumi_i(fifo_yumi)
  );

  assign sent_n[0] = (N0)? 1'b1 : 
                     (N52)? sent_r[0] : 1'b0;
  assign N0 = N51;
  assign sent_n[1] = (N1)? 1'b1 : 
                     (N55)? sent_r[1] : 1'b0;
  assign N1 = N54;
  assign sent_n[2] = (N2)? 1'b1 : 
                     (N58)? sent_r[2] : 1'b0;
  assign N2 = N57;
  assign sent_n[3] = (N3)? 1'b1 : 
                     (N61)? sent_r[3] : 1'b0;
  assign N3 = N60;
  assign sent_n[4] = (N4)? 1'b1 : 
                     (N64)? sent_r[4] : 1'b0;
  assign N4 = N63;
  assign sent_n[5] = (N5)? 1'b1 : 
                     (N67)? sent_r[5] : 1'b0;
  assign N5 = N66;
  assign sent_n[6] = (N6)? 1'b1 : 
                     (N70)? sent_r[6] : 1'b0;
  assign N6 = N69;
  assign sent_n[7] = (N7)? 1'b1 : 
                     (N73)? sent_r[7] : 1'b0;
  assign N7 = N72;
  assign sent_n[8] = (N8)? 1'b1 : 
                     (N76)? sent_r[8] : 1'b0;
  assign N8 = N75;
  assign sent_n[9] = (N9)? 1'b1 : 
                     (N79)? sent_r[9] : 1'b0;
  assign N9 = N78;
  assign sent_n[10] = (N10)? 1'b1 : 
                      (N82)? sent_r[10] : 1'b0;
  assign N10 = N81;
  assign sent_n[11] = (N11)? 1'b1 : 
                      (N85)? sent_r[11] : 1'b0;
  assign N11 = N84;
  assign sent_n[12] = (N12)? 1'b1 : 
                      (N88)? sent_r[12] : 1'b0;
  assign N12 = N87;
  assign sent_n[13] = (N13)? 1'b1 : 
                      (N91)? sent_r[13] : 1'b0;
  assign N13 = N90;
  assign sent_n[14] = (N14)? 1'b1 : 
                      (N94)? sent_r[14] : 1'b0;
  assign N14 = N93;
  assign sent_n[15] = (N15)? 1'b1 : 
                      (N97)? sent_r[15] : 1'b0;
  assign N15 = N96;
  assign sent_n[16] = (N16)? 1'b1 : 
                      (N100)? sent_r[16] : 1'b0;
  assign N16 = N99;
  assign sent_n[17] = (N17)? 1'b1 : 
                      (N103)? sent_r[17] : 1'b0;
  assign N17 = N102;
  assign sent_n[18] = (N18)? 1'b1 : 
                      (N106)? sent_r[18] : 1'b0;
  assign N18 = N105;
  assign sent_n[19] = (N19)? 1'b1 : 
                      (N109)? sent_r[19] : 1'b0;
  assign N19 = N108;
  assign sent_n[20] = (N20)? 1'b1 : 
                      (N112)? sent_r[20] : 1'b0;
  assign N20 = N111;
  assign sent_n[21] = (N21)? 1'b1 : 
                      (N115)? sent_r[21] : 1'b0;
  assign N21 = N114;
  assign sent_n[22] = (N22)? 1'b1 : 
                      (N118)? sent_r[22] : 1'b0;
  assign N22 = N117;
  assign sent_n[23] = (N23)? 1'b1 : 
                      (N121)? sent_r[23] : 1'b0;
  assign N23 = N120;
  assign sent_n[24] = (N24)? 1'b1 : 
                      (N124)? sent_r[24] : 1'b0;
  assign N24 = N123;
  assign sent_n[25] = (N25)? 1'b1 : 
                      (N127)? sent_r[25] : 1'b0;
  assign N25 = N126;
  assign sent_n[26] = (N26)? 1'b1 : 
                      (N130)? sent_r[26] : 1'b0;
  assign N26 = N129;
  assign sent_n[27] = (N27)? 1'b1 : 
                      (N133)? sent_r[27] : 1'b0;
  assign N27 = N132;
  assign sent_n[28] = (N28)? 1'b1 : 
                      (N136)? sent_r[28] : 1'b0;
  assign N28 = N135;
  assign sent_n[29] = (N29)? 1'b1 : 
                      (N139)? sent_r[29] : 1'b0;
  assign N29 = N138;
  assign sent_n[30] = (N30)? 1'b1 : 
                      (N142)? sent_r[30] : 1'b0;
  assign N30 = N141;
  assign sent_n[31] = (N31)? 1'b1 : 
                      (N145)? sent_r[31] : 1'b0;
  assign N31 = N144;
  assign sent_n[32] = (N32)? 1'b1 : 
                      (N148)? sent_r[32] : 1'b0;
  assign N32 = N147;
  assign sent_n[33] = (N33)? 1'b1 : 
                      (N151)? sent_r[33] : 1'b0;
  assign N33 = N150;
  assign sent_n[34] = (N34)? 1'b1 : 
                      (N154)? sent_r[34] : 1'b0;
  assign N34 = N153;
  assign sent_n[35] = (N35)? 1'b1 : 
                      (N157)? sent_r[35] : 1'b0;
  assign N35 = N156;
  assign sent_n[36] = (N36)? 1'b1 : 
                      (N160)? sent_r[36] : 1'b0;
  assign N36 = N159;
  assign sent_n[37] = (N37)? 1'b1 : 
                      (N163)? sent_r[37] : 1'b0;
  assign N37 = N162;
  assign sent_n[38] = (N38)? 1'b1 : 
                      (N166)? sent_r[38] : 1'b0;
  assign N38 = N165;
  assign sent_n[39] = (N39)? 1'b1 : 
                      (N169)? sent_r[39] : 1'b0;
  assign N39 = N168;
  assign sent_n[40] = (N40)? 1'b1 : 
                      (N172)? sent_r[40] : 1'b0;
  assign N40 = N171;
  assign sent_n[41] = (N41)? 1'b1 : 
                      (N175)? sent_r[41] : 1'b0;
  assign N41 = N174;
  assign sent_n[42] = (N42)? 1'b1 : 
                      (N178)? sent_r[42] : 1'b0;
  assign N42 = N177;
  assign sent_n[43] = (N43)? 1'b1 : 
                      (N181)? sent_r[43] : 1'b0;
  assign N43 = N180;
  assign sent_n[44] = (N44)? 1'b1 : 
                      (N184)? sent_r[44] : 1'b0;
  assign N44 = N183;
  assign sent_n[45] = (N45)? 1'b1 : 
                      (N187)? sent_r[45] : 1'b0;
  assign N45 = N186;
  assign sent_n[46] = (N46)? 1'b1 : 
                      (N190)? sent_r[46] : 1'b0;
  assign N46 = N189;
  assign sent_n[47] = (N47)? 1'b1 : 
                      (N193)? sent_r[47] : 1'b0;
  assign N47 = N192;
  assign sent_n[48] = (N48)? 1'b1 : 
                      (N196)? sent_r[48] : 1'b0;
  assign N48 = N195;
  assign sent_n[49] = (N49)? 1'b1 : 
                      (N199)? sent_r[49] : 1'b0;
  assign N49 = N198;
  assign v_o[0] = fifo_v & N200;
  assign N200 = ~sent_r[0];
  assign N50 = sent_n[0] & N201;
  assign N201 = ~fifo_yumi;
  assign N51 = v_o[0] & ready_i[0];
  assign N52 = ~N51;
  assign v_o[1] = fifo_v & N202;
  assign N202 = ~sent_r[1];
  assign N53 = sent_n[1] & N203;
  assign N203 = ~fifo_yumi;
  assign N54 = v_o[1] & ready_i[1];
  assign N55 = ~N54;
  assign v_o[2] = fifo_v & N204;
  assign N204 = ~sent_r[2];
  assign N56 = sent_n[2] & N205;
  assign N205 = ~fifo_yumi;
  assign N57 = v_o[2] & ready_i[2];
  assign N58 = ~N57;
  assign v_o[3] = fifo_v & N206;
  assign N206 = ~sent_r[3];
  assign N59 = sent_n[3] & N207;
  assign N207 = ~fifo_yumi;
  assign N60 = v_o[3] & ready_i[3];
  assign N61 = ~N60;
  assign v_o[4] = fifo_v & N208;
  assign N208 = ~sent_r[4];
  assign N62 = sent_n[4] & N209;
  assign N209 = ~fifo_yumi;
  assign N63 = v_o[4] & ready_i[4];
  assign N64 = ~N63;
  assign v_o[5] = fifo_v & N210;
  assign N210 = ~sent_r[5];
  assign N65 = sent_n[5] & N211;
  assign N211 = ~fifo_yumi;
  assign N66 = v_o[5] & ready_i[5];
  assign N67 = ~N66;
  assign v_o[6] = fifo_v & N212;
  assign N212 = ~sent_r[6];
  assign N68 = sent_n[6] & N213;
  assign N213 = ~fifo_yumi;
  assign N69 = v_o[6] & ready_i[6];
  assign N70 = ~N69;
  assign v_o[7] = fifo_v & N214;
  assign N214 = ~sent_r[7];
  assign N71 = sent_n[7] & N215;
  assign N215 = ~fifo_yumi;
  assign N72 = v_o[7] & ready_i[7];
  assign N73 = ~N72;
  assign v_o[8] = fifo_v & N216;
  assign N216 = ~sent_r[8];
  assign N74 = sent_n[8] & N217;
  assign N217 = ~fifo_yumi;
  assign N75 = v_o[8] & ready_i[8];
  assign N76 = ~N75;
  assign v_o[9] = fifo_v & N218;
  assign N218 = ~sent_r[9];
  assign N77 = sent_n[9] & N219;
  assign N219 = ~fifo_yumi;
  assign N78 = v_o[9] & ready_i[9];
  assign N79 = ~N78;
  assign v_o[10] = fifo_v & N220;
  assign N220 = ~sent_r[10];
  assign N80 = sent_n[10] & N221;
  assign N221 = ~fifo_yumi;
  assign N81 = v_o[10] & ready_i[10];
  assign N82 = ~N81;
  assign v_o[11] = fifo_v & N222;
  assign N222 = ~sent_r[11];
  assign N83 = sent_n[11] & N223;
  assign N223 = ~fifo_yumi;
  assign N84 = v_o[11] & ready_i[11];
  assign N85 = ~N84;
  assign v_o[12] = fifo_v & N224;
  assign N224 = ~sent_r[12];
  assign N86 = sent_n[12] & N225;
  assign N225 = ~fifo_yumi;
  assign N87 = v_o[12] & ready_i[12];
  assign N88 = ~N87;
  assign v_o[13] = fifo_v & N226;
  assign N226 = ~sent_r[13];
  assign N89 = sent_n[13] & N227;
  assign N227 = ~fifo_yumi;
  assign N90 = v_o[13] & ready_i[13];
  assign N91 = ~N90;
  assign v_o[14] = fifo_v & N228;
  assign N228 = ~sent_r[14];
  assign N92 = sent_n[14] & N229;
  assign N229 = ~fifo_yumi;
  assign N93 = v_o[14] & ready_i[14];
  assign N94 = ~N93;
  assign v_o[15] = fifo_v & N230;
  assign N230 = ~sent_r[15];
  assign N95 = sent_n[15] & N231;
  assign N231 = ~fifo_yumi;
  assign N96 = v_o[15] & ready_i[15];
  assign N97 = ~N96;
  assign v_o[16] = fifo_v & N232;
  assign N232 = ~sent_r[16];
  assign N98 = sent_n[16] & N233;
  assign N233 = ~fifo_yumi;
  assign N99 = v_o[16] & ready_i[16];
  assign N100 = ~N99;
  assign v_o[17] = fifo_v & N234;
  assign N234 = ~sent_r[17];
  assign N101 = sent_n[17] & N235;
  assign N235 = ~fifo_yumi;
  assign N102 = v_o[17] & ready_i[17];
  assign N103 = ~N102;
  assign v_o[18] = fifo_v & N236;
  assign N236 = ~sent_r[18];
  assign N104 = sent_n[18] & N237;
  assign N237 = ~fifo_yumi;
  assign N105 = v_o[18] & ready_i[18];
  assign N106 = ~N105;
  assign v_o[19] = fifo_v & N238;
  assign N238 = ~sent_r[19];
  assign N107 = sent_n[19] & N239;
  assign N239 = ~fifo_yumi;
  assign N108 = v_o[19] & ready_i[19];
  assign N109 = ~N108;
  assign v_o[20] = fifo_v & N240;
  assign N240 = ~sent_r[20];
  assign N110 = sent_n[20] & N241;
  assign N241 = ~fifo_yumi;
  assign N111 = v_o[20] & ready_i[20];
  assign N112 = ~N111;
  assign v_o[21] = fifo_v & N242;
  assign N242 = ~sent_r[21];
  assign N113 = sent_n[21] & N243;
  assign N243 = ~fifo_yumi;
  assign N114 = v_o[21] & ready_i[21];
  assign N115 = ~N114;
  assign v_o[22] = fifo_v & N244;
  assign N244 = ~sent_r[22];
  assign N116 = sent_n[22] & N245;
  assign N245 = ~fifo_yumi;
  assign N117 = v_o[22] & ready_i[22];
  assign N118 = ~N117;
  assign v_o[23] = fifo_v & N246;
  assign N246 = ~sent_r[23];
  assign N119 = sent_n[23] & N247;
  assign N247 = ~fifo_yumi;
  assign N120 = v_o[23] & ready_i[23];
  assign N121 = ~N120;
  assign v_o[24] = fifo_v & N248;
  assign N248 = ~sent_r[24];
  assign N122 = sent_n[24] & N249;
  assign N249 = ~fifo_yumi;
  assign N123 = v_o[24] & ready_i[24];
  assign N124 = ~N123;
  assign v_o[25] = fifo_v & N250;
  assign N250 = ~sent_r[25];
  assign N125 = sent_n[25] & N251;
  assign N251 = ~fifo_yumi;
  assign N126 = v_o[25] & ready_i[25];
  assign N127 = ~N126;
  assign v_o[26] = fifo_v & N252;
  assign N252 = ~sent_r[26];
  assign N128 = sent_n[26] & N253;
  assign N253 = ~fifo_yumi;
  assign N129 = v_o[26] & ready_i[26];
  assign N130 = ~N129;
  assign v_o[27] = fifo_v & N254;
  assign N254 = ~sent_r[27];
  assign N131 = sent_n[27] & N255;
  assign N255 = ~fifo_yumi;
  assign N132 = v_o[27] & ready_i[27];
  assign N133 = ~N132;
  assign v_o[28] = fifo_v & N256;
  assign N256 = ~sent_r[28];
  assign N134 = sent_n[28] & N257;
  assign N257 = ~fifo_yumi;
  assign N135 = v_o[28] & ready_i[28];
  assign N136 = ~N135;
  assign v_o[29] = fifo_v & N258;
  assign N258 = ~sent_r[29];
  assign N137 = sent_n[29] & N259;
  assign N259 = ~fifo_yumi;
  assign N138 = v_o[29] & ready_i[29];
  assign N139 = ~N138;
  assign v_o[30] = fifo_v & N260;
  assign N260 = ~sent_r[30];
  assign N140 = sent_n[30] & N261;
  assign N261 = ~fifo_yumi;
  assign N141 = v_o[30] & ready_i[30];
  assign N142 = ~N141;
  assign v_o[31] = fifo_v & N262;
  assign N262 = ~sent_r[31];
  assign N143 = sent_n[31] & N263;
  assign N263 = ~fifo_yumi;
  assign N144 = v_o[31] & ready_i[31];
  assign N145 = ~N144;
  assign v_o[32] = fifo_v & N264;
  assign N264 = ~sent_r[32];
  assign N146 = sent_n[32] & N265;
  assign N265 = ~fifo_yumi;
  assign N147 = v_o[32] & ready_i[32];
  assign N148 = ~N147;
  assign v_o[33] = fifo_v & N266;
  assign N266 = ~sent_r[33];
  assign N149 = sent_n[33] & N267;
  assign N267 = ~fifo_yumi;
  assign N150 = v_o[33] & ready_i[33];
  assign N151 = ~N150;
  assign v_o[34] = fifo_v & N268;
  assign N268 = ~sent_r[34];
  assign N152 = sent_n[34] & N269;
  assign N269 = ~fifo_yumi;
  assign N153 = v_o[34] & ready_i[34];
  assign N154 = ~N153;
  assign v_o[35] = fifo_v & N270;
  assign N270 = ~sent_r[35];
  assign N155 = sent_n[35] & N271;
  assign N271 = ~fifo_yumi;
  assign N156 = v_o[35] & ready_i[35];
  assign N157 = ~N156;
  assign v_o[36] = fifo_v & N272;
  assign N272 = ~sent_r[36];
  assign N158 = sent_n[36] & N273;
  assign N273 = ~fifo_yumi;
  assign N159 = v_o[36] & ready_i[36];
  assign N160 = ~N159;
  assign v_o[37] = fifo_v & N274;
  assign N274 = ~sent_r[37];
  assign N161 = sent_n[37] & N275;
  assign N275 = ~fifo_yumi;
  assign N162 = v_o[37] & ready_i[37];
  assign N163 = ~N162;
  assign v_o[38] = fifo_v & N276;
  assign N276 = ~sent_r[38];
  assign N164 = sent_n[38] & N277;
  assign N277 = ~fifo_yumi;
  assign N165 = v_o[38] & ready_i[38];
  assign N166 = ~N165;
  assign v_o[39] = fifo_v & N278;
  assign N278 = ~sent_r[39];
  assign N167 = sent_n[39] & N279;
  assign N279 = ~fifo_yumi;
  assign N168 = v_o[39] & ready_i[39];
  assign N169 = ~N168;
  assign v_o[40] = fifo_v & N280;
  assign N280 = ~sent_r[40];
  assign N170 = sent_n[40] & N281;
  assign N281 = ~fifo_yumi;
  assign N171 = v_o[40] & ready_i[40];
  assign N172 = ~N171;
  assign v_o[41] = fifo_v & N282;
  assign N282 = ~sent_r[41];
  assign N173 = sent_n[41] & N283;
  assign N283 = ~fifo_yumi;
  assign N174 = v_o[41] & ready_i[41];
  assign N175 = ~N174;
  assign v_o[42] = fifo_v & N284;
  assign N284 = ~sent_r[42];
  assign N176 = sent_n[42] & N285;
  assign N285 = ~fifo_yumi;
  assign N177 = v_o[42] & ready_i[42];
  assign N178 = ~N177;
  assign v_o[43] = fifo_v & N286;
  assign N286 = ~sent_r[43];
  assign N179 = sent_n[43] & N287;
  assign N287 = ~fifo_yumi;
  assign N180 = v_o[43] & ready_i[43];
  assign N181 = ~N180;
  assign v_o[44] = fifo_v & N288;
  assign N288 = ~sent_r[44];
  assign N182 = sent_n[44] & N289;
  assign N289 = ~fifo_yumi;
  assign N183 = v_o[44] & ready_i[44];
  assign N184 = ~N183;
  assign v_o[45] = fifo_v & N290;
  assign N290 = ~sent_r[45];
  assign N185 = sent_n[45] & N291;
  assign N291 = ~fifo_yumi;
  assign N186 = v_o[45] & ready_i[45];
  assign N187 = ~N186;
  assign v_o[46] = fifo_v & N292;
  assign N292 = ~sent_r[46];
  assign N188 = sent_n[46] & N293;
  assign N293 = ~fifo_yumi;
  assign N189 = v_o[46] & ready_i[46];
  assign N190 = ~N189;
  assign v_o[47] = fifo_v & N294;
  assign N294 = ~sent_r[47];
  assign N191 = sent_n[47] & N295;
  assign N295 = ~fifo_yumi;
  assign N192 = v_o[47] & ready_i[47];
  assign N193 = ~N192;
  assign v_o[48] = fifo_v & N296;
  assign N296 = ~sent_r[48];
  assign N194 = sent_n[48] & N297;
  assign N297 = ~fifo_yumi;
  assign N195 = v_o[48] & ready_i[48];
  assign N196 = ~N195;
  assign v_o[49] = fifo_v & N298;
  assign N298 = ~sent_r[49];
  assign N197 = sent_n[49] & N299;
  assign N299 = ~fifo_yumi;
  assign N198 = v_o[49] & ready_i[49];
  assign N199 = ~N198;
  assign fifo_yumi = N347 & sent_n[0];
  assign N347 = N346 & sent_n[1];
  assign N346 = N345 & sent_n[2];
  assign N345 = N344 & sent_n[3];
  assign N344 = N343 & sent_n[4];
  assign N343 = N342 & sent_n[5];
  assign N342 = N341 & sent_n[6];
  assign N341 = N340 & sent_n[7];
  assign N340 = N339 & sent_n[8];
  assign N339 = N338 & sent_n[9];
  assign N338 = N337 & sent_n[10];
  assign N337 = N336 & sent_n[11];
  assign N336 = N335 & sent_n[12];
  assign N335 = N334 & sent_n[13];
  assign N334 = N333 & sent_n[14];
  assign N333 = N332 & sent_n[15];
  assign N332 = N331 & sent_n[16];
  assign N331 = N330 & sent_n[17];
  assign N330 = N329 & sent_n[18];
  assign N329 = N328 & sent_n[19];
  assign N328 = N327 & sent_n[20];
  assign N327 = N326 & sent_n[21];
  assign N326 = N325 & sent_n[22];
  assign N325 = N324 & sent_n[23];
  assign N324 = N323 & sent_n[24];
  assign N323 = N322 & sent_n[25];
  assign N322 = N321 & sent_n[26];
  assign N321 = N320 & sent_n[27];
  assign N320 = N319 & sent_n[28];
  assign N319 = N318 & sent_n[29];
  assign N318 = N317 & sent_n[30];
  assign N317 = N316 & sent_n[31];
  assign N316 = N315 & sent_n[32];
  assign N315 = N314 & sent_n[33];
  assign N314 = N313 & sent_n[34];
  assign N313 = N312 & sent_n[35];
  assign N312 = N311 & sent_n[36];
  assign N311 = N310 & sent_n[37];
  assign N310 = N309 & sent_n[38];
  assign N309 = N308 & sent_n[39];
  assign N308 = N307 & sent_n[40];
  assign N307 = N306 & sent_n[41];
  assign N306 = N305 & sent_n[42];
  assign N305 = N304 & sent_n[43];
  assign N304 = N303 & sent_n[44];
  assign N303 = N302 & sent_n[45];
  assign N302 = N301 & sent_n[46];
  assign N301 = N300 & sent_n[47];
  assign N300 = sent_n[49] & sent_n[48];

  always @(posedge clk_i) begin
    if(reset_i) begin
      sent_r_0_sv2v_reg <= 1'b0;
      sent_r_1_sv2v_reg <= 1'b0;
      sent_r_2_sv2v_reg <= 1'b0;
      sent_r_3_sv2v_reg <= 1'b0;
      sent_r_4_sv2v_reg <= 1'b0;
      sent_r_5_sv2v_reg <= 1'b0;
      sent_r_6_sv2v_reg <= 1'b0;
      sent_r_7_sv2v_reg <= 1'b0;
      sent_r_8_sv2v_reg <= 1'b0;
      sent_r_9_sv2v_reg <= 1'b0;
      sent_r_10_sv2v_reg <= 1'b0;
      sent_r_11_sv2v_reg <= 1'b0;
      sent_r_12_sv2v_reg <= 1'b0;
      sent_r_13_sv2v_reg <= 1'b0;
      sent_r_14_sv2v_reg <= 1'b0;
      sent_r_15_sv2v_reg <= 1'b0;
      sent_r_16_sv2v_reg <= 1'b0;
      sent_r_17_sv2v_reg <= 1'b0;
      sent_r_18_sv2v_reg <= 1'b0;
      sent_r_19_sv2v_reg <= 1'b0;
      sent_r_20_sv2v_reg <= 1'b0;
      sent_r_21_sv2v_reg <= 1'b0;
      sent_r_22_sv2v_reg <= 1'b0;
      sent_r_23_sv2v_reg <= 1'b0;
      sent_r_24_sv2v_reg <= 1'b0;
      sent_r_25_sv2v_reg <= 1'b0;
      sent_r_26_sv2v_reg <= 1'b0;
      sent_r_27_sv2v_reg <= 1'b0;
      sent_r_28_sv2v_reg <= 1'b0;
      sent_r_29_sv2v_reg <= 1'b0;
      sent_r_30_sv2v_reg <= 1'b0;
      sent_r_31_sv2v_reg <= 1'b0;
      sent_r_32_sv2v_reg <= 1'b0;
      sent_r_33_sv2v_reg <= 1'b0;
      sent_r_34_sv2v_reg <= 1'b0;
      sent_r_35_sv2v_reg <= 1'b0;
      sent_r_36_sv2v_reg <= 1'b0;
      sent_r_37_sv2v_reg <= 1'b0;
      sent_r_38_sv2v_reg <= 1'b0;
      sent_r_39_sv2v_reg <= 1'b0;
      sent_r_40_sv2v_reg <= 1'b0;
      sent_r_41_sv2v_reg <= 1'b0;
      sent_r_42_sv2v_reg <= 1'b0;
      sent_r_43_sv2v_reg <= 1'b0;
      sent_r_44_sv2v_reg <= 1'b0;
      sent_r_45_sv2v_reg <= 1'b0;
      sent_r_46_sv2v_reg <= 1'b0;
      sent_r_47_sv2v_reg <= 1'b0;
      sent_r_48_sv2v_reg <= 1'b0;
      sent_r_49_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      sent_r_0_sv2v_reg <= N50;
      sent_r_1_sv2v_reg <= N53;
      sent_r_2_sv2v_reg <= N56;
      sent_r_3_sv2v_reg <= N59;
      sent_r_4_sv2v_reg <= N62;
      sent_r_5_sv2v_reg <= N65;
      sent_r_6_sv2v_reg <= N68;
      sent_r_7_sv2v_reg <= N71;
      sent_r_8_sv2v_reg <= N74;
      sent_r_9_sv2v_reg <= N77;
      sent_r_10_sv2v_reg <= N80;
      sent_r_11_sv2v_reg <= N83;
      sent_r_12_sv2v_reg <= N86;
      sent_r_13_sv2v_reg <= N89;
      sent_r_14_sv2v_reg <= N92;
      sent_r_15_sv2v_reg <= N95;
      sent_r_16_sv2v_reg <= N98;
      sent_r_17_sv2v_reg <= N101;
      sent_r_18_sv2v_reg <= N104;
      sent_r_19_sv2v_reg <= N107;
      sent_r_20_sv2v_reg <= N110;
      sent_r_21_sv2v_reg <= N113;
      sent_r_22_sv2v_reg <= N116;
      sent_r_23_sv2v_reg <= N119;
      sent_r_24_sv2v_reg <= N122;
      sent_r_25_sv2v_reg <= N125;
      sent_r_26_sv2v_reg <= N128;
      sent_r_27_sv2v_reg <= N131;
      sent_r_28_sv2v_reg <= N134;
      sent_r_29_sv2v_reg <= N137;
      sent_r_30_sv2v_reg <= N140;
      sent_r_31_sv2v_reg <= N143;
      sent_r_32_sv2v_reg <= N146;
      sent_r_33_sv2v_reg <= N149;
      sent_r_34_sv2v_reg <= N152;
      sent_r_35_sv2v_reg <= N155;
      sent_r_36_sv2v_reg <= N158;
      sent_r_37_sv2v_reg <= N161;
      sent_r_38_sv2v_reg <= N164;
      sent_r_39_sv2v_reg <= N167;
      sent_r_40_sv2v_reg <= N170;
      sent_r_41_sv2v_reg <= N173;
      sent_r_42_sv2v_reg <= N176;
      sent_r_43_sv2v_reg <= N179;
      sent_r_44_sv2v_reg <= N182;
      sent_r_45_sv2v_reg <= N185;
      sent_r_46_sv2v_reg <= N188;
      sent_r_47_sv2v_reg <= N191;
      sent_r_48_sv2v_reg <= N194;
      sent_r_49_sv2v_reg <= N197;
    end 
  end


endmodule

