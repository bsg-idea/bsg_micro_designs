

module top
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  credit_o,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output credit_o;
  output v_o;

  bsg_fifo_1r1w_small_credit_on_input
  wrapper
  (
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .credit_o(credit_o),
    .v_o(v_o)
  );


endmodule



module bsg_circular_ptr_slots_p50_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [5:0] o;
  output [5:0] n_o;
  input clk;
  input reset_i;
  wire [5:0] o,n_o,ptr_nowrap;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9;
  wire [6:0] ptr_wrap;
  reg o_5_sv2v_reg,o_4_sv2v_reg,o_3_sv2v_reg,o_2_sv2v_reg,o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[5] = o_5_sv2v_reg;
  assign o[4] = o_4_sv2v_reg;
  assign o[3] = o_3_sv2v_reg;
  assign o[2] = o_2_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign ptr_nowrap = o + add_i[0];
  assign { N8, N7, N6, N5, N4, N3, N2 } = o - { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 };
  assign ptr_wrap = { N8, N7, N6, N5, N4, N3, N2 } + add_i[0];
  assign n_o = (N0)? ptr_wrap[5:0] : 
               (N1)? ptr_nowrap : 1'b0;
  assign N0 = N9;
  assign N1 = ptr_wrap[6];
  assign N9 = ~ptr_wrap[6];

  always @(posedge clk) begin
    if(reset_i) begin
      o_5_sv2v_reg <= 1'b0;
      o_4_sv2v_reg <= 1'b0;
      o_3_sv2v_reg <= 1'b0;
      o_2_sv2v_reg <= 1'b0;
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_5_sv2v_reg <= n_o[5];
      o_4_sv2v_reg <= n_o[4];
      o_3_sv2v_reg <= n_o[3];
      o_2_sv2v_reg <= n_o[2];
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_els_p50
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [5:0] wptr_r_o;
  output [5:0] rptr_r_o;
  output [5:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [5:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,enq_r,deq_r,N0,equal_ptrs,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,
  sv2v_dc_4,sv2v_dc_5,sv2v_dc_6;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_slots_p50_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p50_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N0 = enq_i | deq_i;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N0) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p50_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [31:0] w_data_i;
  input [5:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448;
  wire [1599:0] \nz.mem ;
  reg \nz.mem_1599_sv2v_reg ,\nz.mem_1598_sv2v_reg ,\nz.mem_1597_sv2v_reg ,
  \nz.mem_1596_sv2v_reg ,\nz.mem_1595_sv2v_reg ,\nz.mem_1594_sv2v_reg ,
  \nz.mem_1593_sv2v_reg ,\nz.mem_1592_sv2v_reg ,\nz.mem_1591_sv2v_reg ,\nz.mem_1590_sv2v_reg ,
  \nz.mem_1589_sv2v_reg ,\nz.mem_1588_sv2v_reg ,\nz.mem_1587_sv2v_reg ,
  \nz.mem_1586_sv2v_reg ,\nz.mem_1585_sv2v_reg ,\nz.mem_1584_sv2v_reg ,\nz.mem_1583_sv2v_reg ,
  \nz.mem_1582_sv2v_reg ,\nz.mem_1581_sv2v_reg ,\nz.mem_1580_sv2v_reg ,
  \nz.mem_1579_sv2v_reg ,\nz.mem_1578_sv2v_reg ,\nz.mem_1577_sv2v_reg ,\nz.mem_1576_sv2v_reg ,
  \nz.mem_1575_sv2v_reg ,\nz.mem_1574_sv2v_reg ,\nz.mem_1573_sv2v_reg ,
  \nz.mem_1572_sv2v_reg ,\nz.mem_1571_sv2v_reg ,\nz.mem_1570_sv2v_reg ,\nz.mem_1569_sv2v_reg ,
  \nz.mem_1568_sv2v_reg ,\nz.mem_1567_sv2v_reg ,\nz.mem_1566_sv2v_reg ,
  \nz.mem_1565_sv2v_reg ,\nz.mem_1564_sv2v_reg ,\nz.mem_1563_sv2v_reg ,\nz.mem_1562_sv2v_reg ,
  \nz.mem_1561_sv2v_reg ,\nz.mem_1560_sv2v_reg ,\nz.mem_1559_sv2v_reg ,
  \nz.mem_1558_sv2v_reg ,\nz.mem_1557_sv2v_reg ,\nz.mem_1556_sv2v_reg ,\nz.mem_1555_sv2v_reg ,
  \nz.mem_1554_sv2v_reg ,\nz.mem_1553_sv2v_reg ,\nz.mem_1552_sv2v_reg ,
  \nz.mem_1551_sv2v_reg ,\nz.mem_1550_sv2v_reg ,\nz.mem_1549_sv2v_reg ,\nz.mem_1548_sv2v_reg ,
  \nz.mem_1547_sv2v_reg ,\nz.mem_1546_sv2v_reg ,\nz.mem_1545_sv2v_reg ,
  \nz.mem_1544_sv2v_reg ,\nz.mem_1543_sv2v_reg ,\nz.mem_1542_sv2v_reg ,\nz.mem_1541_sv2v_reg ,
  \nz.mem_1540_sv2v_reg ,\nz.mem_1539_sv2v_reg ,\nz.mem_1538_sv2v_reg ,
  \nz.mem_1537_sv2v_reg ,\nz.mem_1536_sv2v_reg ,\nz.mem_1535_sv2v_reg ,\nz.mem_1534_sv2v_reg ,
  \nz.mem_1533_sv2v_reg ,\nz.mem_1532_sv2v_reg ,\nz.mem_1531_sv2v_reg ,
  \nz.mem_1530_sv2v_reg ,\nz.mem_1529_sv2v_reg ,\nz.mem_1528_sv2v_reg ,\nz.mem_1527_sv2v_reg ,
  \nz.mem_1526_sv2v_reg ,\nz.mem_1525_sv2v_reg ,\nz.mem_1524_sv2v_reg ,
  \nz.mem_1523_sv2v_reg ,\nz.mem_1522_sv2v_reg ,\nz.mem_1521_sv2v_reg ,\nz.mem_1520_sv2v_reg ,
  \nz.mem_1519_sv2v_reg ,\nz.mem_1518_sv2v_reg ,\nz.mem_1517_sv2v_reg ,
  \nz.mem_1516_sv2v_reg ,\nz.mem_1515_sv2v_reg ,\nz.mem_1514_sv2v_reg ,
  \nz.mem_1513_sv2v_reg ,\nz.mem_1512_sv2v_reg ,\nz.mem_1511_sv2v_reg ,\nz.mem_1510_sv2v_reg ,
  \nz.mem_1509_sv2v_reg ,\nz.mem_1508_sv2v_reg ,\nz.mem_1507_sv2v_reg ,
  \nz.mem_1506_sv2v_reg ,\nz.mem_1505_sv2v_reg ,\nz.mem_1504_sv2v_reg ,\nz.mem_1503_sv2v_reg ,
  \nz.mem_1502_sv2v_reg ,\nz.mem_1501_sv2v_reg ,\nz.mem_1500_sv2v_reg ,
  \nz.mem_1499_sv2v_reg ,\nz.mem_1498_sv2v_reg ,\nz.mem_1497_sv2v_reg ,\nz.mem_1496_sv2v_reg ,
  \nz.mem_1495_sv2v_reg ,\nz.mem_1494_sv2v_reg ,\nz.mem_1493_sv2v_reg ,
  \nz.mem_1492_sv2v_reg ,\nz.mem_1491_sv2v_reg ,\nz.mem_1490_sv2v_reg ,\nz.mem_1489_sv2v_reg ,
  \nz.mem_1488_sv2v_reg ,\nz.mem_1487_sv2v_reg ,\nz.mem_1486_sv2v_reg ,
  \nz.mem_1485_sv2v_reg ,\nz.mem_1484_sv2v_reg ,\nz.mem_1483_sv2v_reg ,\nz.mem_1482_sv2v_reg ,
  \nz.mem_1481_sv2v_reg ,\nz.mem_1480_sv2v_reg ,\nz.mem_1479_sv2v_reg ,
  \nz.mem_1478_sv2v_reg ,\nz.mem_1477_sv2v_reg ,\nz.mem_1476_sv2v_reg ,\nz.mem_1475_sv2v_reg ,
  \nz.mem_1474_sv2v_reg ,\nz.mem_1473_sv2v_reg ,\nz.mem_1472_sv2v_reg ,
  \nz.mem_1471_sv2v_reg ,\nz.mem_1470_sv2v_reg ,\nz.mem_1469_sv2v_reg ,\nz.mem_1468_sv2v_reg ,
  \nz.mem_1467_sv2v_reg ,\nz.mem_1466_sv2v_reg ,\nz.mem_1465_sv2v_reg ,
  \nz.mem_1464_sv2v_reg ,\nz.mem_1463_sv2v_reg ,\nz.mem_1462_sv2v_reg ,\nz.mem_1461_sv2v_reg ,
  \nz.mem_1460_sv2v_reg ,\nz.mem_1459_sv2v_reg ,\nz.mem_1458_sv2v_reg ,
  \nz.mem_1457_sv2v_reg ,\nz.mem_1456_sv2v_reg ,\nz.mem_1455_sv2v_reg ,\nz.mem_1454_sv2v_reg ,
  \nz.mem_1453_sv2v_reg ,\nz.mem_1452_sv2v_reg ,\nz.mem_1451_sv2v_reg ,
  \nz.mem_1450_sv2v_reg ,\nz.mem_1449_sv2v_reg ,\nz.mem_1448_sv2v_reg ,\nz.mem_1447_sv2v_reg ,
  \nz.mem_1446_sv2v_reg ,\nz.mem_1445_sv2v_reg ,\nz.mem_1444_sv2v_reg ,
  \nz.mem_1443_sv2v_reg ,\nz.mem_1442_sv2v_reg ,\nz.mem_1441_sv2v_reg ,\nz.mem_1440_sv2v_reg ,
  \nz.mem_1439_sv2v_reg ,\nz.mem_1438_sv2v_reg ,\nz.mem_1437_sv2v_reg ,
  \nz.mem_1436_sv2v_reg ,\nz.mem_1435_sv2v_reg ,\nz.mem_1434_sv2v_reg ,
  \nz.mem_1433_sv2v_reg ,\nz.mem_1432_sv2v_reg ,\nz.mem_1431_sv2v_reg ,\nz.mem_1430_sv2v_reg ,
  \nz.mem_1429_sv2v_reg ,\nz.mem_1428_sv2v_reg ,\nz.mem_1427_sv2v_reg ,
  \nz.mem_1426_sv2v_reg ,\nz.mem_1425_sv2v_reg ,\nz.mem_1424_sv2v_reg ,\nz.mem_1423_sv2v_reg ,
  \nz.mem_1422_sv2v_reg ,\nz.mem_1421_sv2v_reg ,\nz.mem_1420_sv2v_reg ,
  \nz.mem_1419_sv2v_reg ,\nz.mem_1418_sv2v_reg ,\nz.mem_1417_sv2v_reg ,\nz.mem_1416_sv2v_reg ,
  \nz.mem_1415_sv2v_reg ,\nz.mem_1414_sv2v_reg ,\nz.mem_1413_sv2v_reg ,
  \nz.mem_1412_sv2v_reg ,\nz.mem_1411_sv2v_reg ,\nz.mem_1410_sv2v_reg ,\nz.mem_1409_sv2v_reg ,
  \nz.mem_1408_sv2v_reg ,\nz.mem_1407_sv2v_reg ,\nz.mem_1406_sv2v_reg ,
  \nz.mem_1405_sv2v_reg ,\nz.mem_1404_sv2v_reg ,\nz.mem_1403_sv2v_reg ,\nz.mem_1402_sv2v_reg ,
  \nz.mem_1401_sv2v_reg ,\nz.mem_1400_sv2v_reg ,\nz.mem_1399_sv2v_reg ,
  \nz.mem_1398_sv2v_reg ,\nz.mem_1397_sv2v_reg ,\nz.mem_1396_sv2v_reg ,\nz.mem_1395_sv2v_reg ,
  \nz.mem_1394_sv2v_reg ,\nz.mem_1393_sv2v_reg ,\nz.mem_1392_sv2v_reg ,
  \nz.mem_1391_sv2v_reg ,\nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,\nz.mem_1388_sv2v_reg ,
  \nz.mem_1387_sv2v_reg ,\nz.mem_1386_sv2v_reg ,\nz.mem_1385_sv2v_reg ,
  \nz.mem_1384_sv2v_reg ,\nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,\nz.mem_1381_sv2v_reg ,
  \nz.mem_1380_sv2v_reg ,\nz.mem_1379_sv2v_reg ,\nz.mem_1378_sv2v_reg ,
  \nz.mem_1377_sv2v_reg ,\nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,\nz.mem_1374_sv2v_reg ,
  \nz.mem_1373_sv2v_reg ,\nz.mem_1372_sv2v_reg ,\nz.mem_1371_sv2v_reg ,
  \nz.mem_1370_sv2v_reg ,\nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,\nz.mem_1367_sv2v_reg ,
  \nz.mem_1366_sv2v_reg ,\nz.mem_1365_sv2v_reg ,\nz.mem_1364_sv2v_reg ,
  \nz.mem_1363_sv2v_reg ,\nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,\nz.mem_1360_sv2v_reg ,
  \nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,\nz.mem_1357_sv2v_reg ,
  \nz.mem_1356_sv2v_reg ,\nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,
  \nz.mem_1353_sv2v_reg ,\nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,\nz.mem_1350_sv2v_reg ,
  \nz.mem_1349_sv2v_reg ,\nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,
  \nz.mem_1346_sv2v_reg ,\nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,\nz.mem_1343_sv2v_reg ,
  \nz.mem_1342_sv2v_reg ,\nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,
  \nz.mem_1339_sv2v_reg ,\nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,\nz.mem_1336_sv2v_reg ,
  \nz.mem_1335_sv2v_reg ,\nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,
  \nz.mem_1332_sv2v_reg ,\nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,\nz.mem_1329_sv2v_reg ,
  \nz.mem_1328_sv2v_reg ,\nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,
  \nz.mem_1325_sv2v_reg ,\nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,\nz.mem_1322_sv2v_reg ,
  \nz.mem_1321_sv2v_reg ,\nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,
  \nz.mem_1318_sv2v_reg ,\nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,\nz.mem_1315_sv2v_reg ,
  \nz.mem_1314_sv2v_reg ,\nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,
  \nz.mem_1311_sv2v_reg ,\nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,\nz.mem_1308_sv2v_reg ,
  \nz.mem_1307_sv2v_reg ,\nz.mem_1306_sv2v_reg ,\nz.mem_1305_sv2v_reg ,
  \nz.mem_1304_sv2v_reg ,\nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,\nz.mem_1301_sv2v_reg ,
  \nz.mem_1300_sv2v_reg ,\nz.mem_1299_sv2v_reg ,\nz.mem_1298_sv2v_reg ,
  \nz.mem_1297_sv2v_reg ,\nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,\nz.mem_1294_sv2v_reg ,
  \nz.mem_1293_sv2v_reg ,\nz.mem_1292_sv2v_reg ,\nz.mem_1291_sv2v_reg ,
  \nz.mem_1290_sv2v_reg ,\nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,\nz.mem_1287_sv2v_reg ,
  \nz.mem_1286_sv2v_reg ,\nz.mem_1285_sv2v_reg ,\nz.mem_1284_sv2v_reg ,
  \nz.mem_1283_sv2v_reg ,\nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,\nz.mem_1280_sv2v_reg ,
  \nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,\nz.mem_1277_sv2v_reg ,
  \nz.mem_1276_sv2v_reg ,\nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,
  \nz.mem_1273_sv2v_reg ,\nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,\nz.mem_1270_sv2v_reg ,
  \nz.mem_1269_sv2v_reg ,\nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,
  \nz.mem_1266_sv2v_reg ,\nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,\nz.mem_1263_sv2v_reg ,
  \nz.mem_1262_sv2v_reg ,\nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,
  \nz.mem_1259_sv2v_reg ,\nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,\nz.mem_1256_sv2v_reg ,
  \nz.mem_1255_sv2v_reg ,\nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,
  \nz.mem_1252_sv2v_reg ,\nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,\nz.mem_1249_sv2v_reg ,
  \nz.mem_1248_sv2v_reg ,\nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,
  \nz.mem_1245_sv2v_reg ,\nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,\nz.mem_1242_sv2v_reg ,
  \nz.mem_1241_sv2v_reg ,\nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,
  \nz.mem_1238_sv2v_reg ,\nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,\nz.mem_1235_sv2v_reg ,
  \nz.mem_1234_sv2v_reg ,\nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,
  \nz.mem_1231_sv2v_reg ,\nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,\nz.mem_1228_sv2v_reg ,
  \nz.mem_1227_sv2v_reg ,\nz.mem_1226_sv2v_reg ,\nz.mem_1225_sv2v_reg ,
  \nz.mem_1224_sv2v_reg ,\nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,\nz.mem_1221_sv2v_reg ,
  \nz.mem_1220_sv2v_reg ,\nz.mem_1219_sv2v_reg ,\nz.mem_1218_sv2v_reg ,
  \nz.mem_1217_sv2v_reg ,\nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,\nz.mem_1214_sv2v_reg ,
  \nz.mem_1213_sv2v_reg ,\nz.mem_1212_sv2v_reg ,\nz.mem_1211_sv2v_reg ,
  \nz.mem_1210_sv2v_reg ,\nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,\nz.mem_1207_sv2v_reg ,
  \nz.mem_1206_sv2v_reg ,\nz.mem_1205_sv2v_reg ,\nz.mem_1204_sv2v_reg ,
  \nz.mem_1203_sv2v_reg ,\nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,\nz.mem_1200_sv2v_reg ,
  \nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,\nz.mem_1197_sv2v_reg ,
  \nz.mem_1196_sv2v_reg ,\nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,
  \nz.mem_1193_sv2v_reg ,\nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,\nz.mem_1190_sv2v_reg ,
  \nz.mem_1189_sv2v_reg ,\nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,
  \nz.mem_1186_sv2v_reg ,\nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,\nz.mem_1183_sv2v_reg ,
  \nz.mem_1182_sv2v_reg ,\nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,
  \nz.mem_1179_sv2v_reg ,\nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,\nz.mem_1176_sv2v_reg ,
  \nz.mem_1175_sv2v_reg ,\nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,
  \nz.mem_1172_sv2v_reg ,\nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,\nz.mem_1169_sv2v_reg ,
  \nz.mem_1168_sv2v_reg ,\nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,
  \nz.mem_1165_sv2v_reg ,\nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,\nz.mem_1162_sv2v_reg ,
  \nz.mem_1161_sv2v_reg ,\nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,
  \nz.mem_1158_sv2v_reg ,\nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,\nz.mem_1155_sv2v_reg ,
  \nz.mem_1154_sv2v_reg ,\nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,
  \nz.mem_1151_sv2v_reg ,\nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,\nz.mem_1148_sv2v_reg ,
  \nz.mem_1147_sv2v_reg ,\nz.mem_1146_sv2v_reg ,\nz.mem_1145_sv2v_reg ,
  \nz.mem_1144_sv2v_reg ,\nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,\nz.mem_1141_sv2v_reg ,
  \nz.mem_1140_sv2v_reg ,\nz.mem_1139_sv2v_reg ,\nz.mem_1138_sv2v_reg ,
  \nz.mem_1137_sv2v_reg ,\nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,\nz.mem_1134_sv2v_reg ,
  \nz.mem_1133_sv2v_reg ,\nz.mem_1132_sv2v_reg ,\nz.mem_1131_sv2v_reg ,
  \nz.mem_1130_sv2v_reg ,\nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,\nz.mem_1127_sv2v_reg ,
  \nz.mem_1126_sv2v_reg ,\nz.mem_1125_sv2v_reg ,\nz.mem_1124_sv2v_reg ,
  \nz.mem_1123_sv2v_reg ,\nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,\nz.mem_1120_sv2v_reg ,
  \nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,\nz.mem_1117_sv2v_reg ,
  \nz.mem_1116_sv2v_reg ,\nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,
  \nz.mem_1113_sv2v_reg ,\nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,\nz.mem_1110_sv2v_reg ,
  \nz.mem_1109_sv2v_reg ,\nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,
  \nz.mem_1106_sv2v_reg ,\nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,\nz.mem_1103_sv2v_reg ,
  \nz.mem_1102_sv2v_reg ,\nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,
  \nz.mem_1099_sv2v_reg ,\nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,\nz.mem_1096_sv2v_reg ,
  \nz.mem_1095_sv2v_reg ,\nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,
  \nz.mem_1092_sv2v_reg ,\nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,\nz.mem_1089_sv2v_reg ,
  \nz.mem_1088_sv2v_reg ,\nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,
  \nz.mem_1085_sv2v_reg ,\nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,\nz.mem_1082_sv2v_reg ,
  \nz.mem_1081_sv2v_reg ,\nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,
  \nz.mem_1078_sv2v_reg ,\nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,\nz.mem_1075_sv2v_reg ,
  \nz.mem_1074_sv2v_reg ,\nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,
  \nz.mem_1071_sv2v_reg ,\nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,\nz.mem_1068_sv2v_reg ,
  \nz.mem_1067_sv2v_reg ,\nz.mem_1066_sv2v_reg ,\nz.mem_1065_sv2v_reg ,
  \nz.mem_1064_sv2v_reg ,\nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,\nz.mem_1061_sv2v_reg ,
  \nz.mem_1060_sv2v_reg ,\nz.mem_1059_sv2v_reg ,\nz.mem_1058_sv2v_reg ,
  \nz.mem_1057_sv2v_reg ,\nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,\nz.mem_1054_sv2v_reg ,
  \nz.mem_1053_sv2v_reg ,\nz.mem_1052_sv2v_reg ,\nz.mem_1051_sv2v_reg ,
  \nz.mem_1050_sv2v_reg ,\nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,\nz.mem_1047_sv2v_reg ,
  \nz.mem_1046_sv2v_reg ,\nz.mem_1045_sv2v_reg ,\nz.mem_1044_sv2v_reg ,
  \nz.mem_1043_sv2v_reg ,\nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,\nz.mem_1040_sv2v_reg ,
  \nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,\nz.mem_1037_sv2v_reg ,
  \nz.mem_1036_sv2v_reg ,\nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,
  \nz.mem_1033_sv2v_reg ,\nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,\nz.mem_1030_sv2v_reg ,
  \nz.mem_1029_sv2v_reg ,\nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,
  \nz.mem_1026_sv2v_reg ,\nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,\nz.mem_1023_sv2v_reg ,
  \nz.mem_1022_sv2v_reg ,\nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,
  \nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,\nz.mem_1016_sv2v_reg ,
  \nz.mem_1015_sv2v_reg ,\nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,
  \nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,\nz.mem_1009_sv2v_reg ,
  \nz.mem_1008_sv2v_reg ,\nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,
  \nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,\nz.mem_1002_sv2v_reg ,
  \nz.mem_1001_sv2v_reg ,\nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,
  \nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,
  \nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,\nz.mem_991_sv2v_reg ,
  \nz.mem_990_sv2v_reg ,\nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,
  \nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,\nz.mem_984_sv2v_reg ,
  \nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,\nz.mem_980_sv2v_reg ,
  \nz.mem_979_sv2v_reg ,\nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,
  \nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,\nz.mem_973_sv2v_reg ,
  \nz.mem_972_sv2v_reg ,\nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,
  \nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,
  \nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,\nz.mem_962_sv2v_reg ,
  \nz.mem_961_sv2v_reg ,\nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,
  \nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,
  \nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,\nz.mem_951_sv2v_reg ,
  \nz.mem_950_sv2v_reg ,\nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,
  \nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,\nz.mem_944_sv2v_reg ,
  \nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,\nz.mem_940_sv2v_reg ,
  \nz.mem_939_sv2v_reg ,\nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,
  \nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,\nz.mem_933_sv2v_reg ,
  \nz.mem_932_sv2v_reg ,\nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,
  \nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,
  \nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,\nz.mem_922_sv2v_reg ,
  \nz.mem_921_sv2v_reg ,\nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,
  \nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,
  \nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,\nz.mem_911_sv2v_reg ,
  \nz.mem_910_sv2v_reg ,\nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,
  \nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,\nz.mem_904_sv2v_reg ,
  \nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,\nz.mem_900_sv2v_reg ,
  \nz.mem_899_sv2v_reg ,\nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,
  \nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,\nz.mem_893_sv2v_reg ,
  \nz.mem_892_sv2v_reg ,\nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,
  \nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,
  \nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,\nz.mem_882_sv2v_reg ,
  \nz.mem_881_sv2v_reg ,\nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,
  \nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,
  \nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,\nz.mem_871_sv2v_reg ,
  \nz.mem_870_sv2v_reg ,\nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,
  \nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,\nz.mem_864_sv2v_reg ,
  \nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,\nz.mem_860_sv2v_reg ,
  \nz.mem_859_sv2v_reg ,\nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,
  \nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,\nz.mem_853_sv2v_reg ,
  \nz.mem_852_sv2v_reg ,\nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,
  \nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,
  \nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,\nz.mem_842_sv2v_reg ,
  \nz.mem_841_sv2v_reg ,\nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,
  \nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,
  \nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,\nz.mem_831_sv2v_reg ,
  \nz.mem_830_sv2v_reg ,\nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,
  \nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,\nz.mem_824_sv2v_reg ,
  \nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,\nz.mem_820_sv2v_reg ,
  \nz.mem_819_sv2v_reg ,\nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,
  \nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,\nz.mem_813_sv2v_reg ,
  \nz.mem_812_sv2v_reg ,\nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,
  \nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,
  \nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,\nz.mem_802_sv2v_reg ,
  \nz.mem_801_sv2v_reg ,\nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,
  \nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,
  \nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,\nz.mem_791_sv2v_reg ,
  \nz.mem_790_sv2v_reg ,\nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,
  \nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,\nz.mem_784_sv2v_reg ,
  \nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,\nz.mem_780_sv2v_reg ,
  \nz.mem_779_sv2v_reg ,\nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,
  \nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,\nz.mem_773_sv2v_reg ,
  \nz.mem_772_sv2v_reg ,\nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,
  \nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,
  \nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,\nz.mem_762_sv2v_reg ,
  \nz.mem_761_sv2v_reg ,\nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,
  \nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,
  \nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,\nz.mem_751_sv2v_reg ,
  \nz.mem_750_sv2v_reg ,\nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,
  \nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,\nz.mem_744_sv2v_reg ,
  \nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,\nz.mem_740_sv2v_reg ,
  \nz.mem_739_sv2v_reg ,\nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,
  \nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,\nz.mem_733_sv2v_reg ,
  \nz.mem_732_sv2v_reg ,\nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,
  \nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,
  \nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,\nz.mem_722_sv2v_reg ,
  \nz.mem_721_sv2v_reg ,\nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,
  \nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,
  \nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,\nz.mem_711_sv2v_reg ,
  \nz.mem_710_sv2v_reg ,\nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,
  \nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,\nz.mem_704_sv2v_reg ,
  \nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,\nz.mem_700_sv2v_reg ,
  \nz.mem_699_sv2v_reg ,\nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,
  \nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,\nz.mem_693_sv2v_reg ,
  \nz.mem_692_sv2v_reg ,\nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,
  \nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,
  \nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,\nz.mem_682_sv2v_reg ,
  \nz.mem_681_sv2v_reg ,\nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,
  \nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,
  \nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,\nz.mem_671_sv2v_reg ,
  \nz.mem_670_sv2v_reg ,\nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,
  \nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,
  \nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,\nz.mem_660_sv2v_reg ,
  \nz.mem_659_sv2v_reg ,\nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,
  \nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,\nz.mem_653_sv2v_reg ,
  \nz.mem_652_sv2v_reg ,\nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,
  \nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,
  \nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,\nz.mem_642_sv2v_reg ,
  \nz.mem_641_sv2v_reg ,\nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,
  \nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,
  \nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,
  \nz.mem_630_sv2v_reg ,\nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,
  \nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,
  \nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,
  \nz.mem_619_sv2v_reg ,\nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,
  \nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,
  \nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,
  \nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,
  \nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,
  \nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,
  \nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,
  \nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,
  \nz.mem_590_sv2v_reg ,\nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,
  \nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,
  \nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,
  \nz.mem_579_sv2v_reg ,\nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,
  \nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,
  \nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,
  \nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,
  \nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,
  \nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,
  \nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,
  \nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,
  \nz.mem_550_sv2v_reg ,\nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,
  \nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,
  \nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,
  \nz.mem_539_sv2v_reg ,\nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,
  \nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,
  \nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,
  \nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,
  \nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,
  \nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,
  \nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,
  \nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,
  \nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,
  \nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,
  \nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,
  \nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,
  \nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,
  \nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,
  \nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,
  \nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,
  \nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,
  \nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,
  \nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,
  \nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,
  \nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,
  \nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,
  \nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,
  \nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,
  \nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,
  \nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,
  \nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,
  \nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,
  \nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,
  \nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,
  \nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,
  \nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,
  \nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,
  \nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,
  \nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,
  \nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,
  \nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,
  \nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,
  \nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,
  \nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,
  \nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,
  \nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,
  \nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,
  \nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,
  \nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,
  \nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,
  \nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,
  \nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,
  \nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,
  \nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,
  \nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,
  \nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,
  \nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,
  \nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,
  \nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,
  \nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,
  \nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,
  \nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,
  \nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,
  \nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,
  \nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,
  \nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,
  \nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,
  \nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,
  \nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,
  \nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,
  \nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,
  \nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,
  \nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,
  \nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,
  \nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,
  \nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,
  \nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,
  \nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,
  \nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,
  \nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,
  \nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,
  \nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,
  \nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,
  \nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,
  \nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,
  \nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,
  \nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,
  \nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,
  \nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,
  \nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,
  \nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,
  \nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,
  \nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,
  \nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,
  \nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,
  \nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,
  \nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,
  \nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,
  \nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,
  \nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,
  \nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.mem [1599] = \nz.mem_1599_sv2v_reg ;
  assign \nz.mem [1598] = \nz.mem_1598_sv2v_reg ;
  assign \nz.mem [1597] = \nz.mem_1597_sv2v_reg ;
  assign \nz.mem [1596] = \nz.mem_1596_sv2v_reg ;
  assign \nz.mem [1595] = \nz.mem_1595_sv2v_reg ;
  assign \nz.mem [1594] = \nz.mem_1594_sv2v_reg ;
  assign \nz.mem [1593] = \nz.mem_1593_sv2v_reg ;
  assign \nz.mem [1592] = \nz.mem_1592_sv2v_reg ;
  assign \nz.mem [1591] = \nz.mem_1591_sv2v_reg ;
  assign \nz.mem [1590] = \nz.mem_1590_sv2v_reg ;
  assign \nz.mem [1589] = \nz.mem_1589_sv2v_reg ;
  assign \nz.mem [1588] = \nz.mem_1588_sv2v_reg ;
  assign \nz.mem [1587] = \nz.mem_1587_sv2v_reg ;
  assign \nz.mem [1586] = \nz.mem_1586_sv2v_reg ;
  assign \nz.mem [1585] = \nz.mem_1585_sv2v_reg ;
  assign \nz.mem [1584] = \nz.mem_1584_sv2v_reg ;
  assign \nz.mem [1583] = \nz.mem_1583_sv2v_reg ;
  assign \nz.mem [1582] = \nz.mem_1582_sv2v_reg ;
  assign \nz.mem [1581] = \nz.mem_1581_sv2v_reg ;
  assign \nz.mem [1580] = \nz.mem_1580_sv2v_reg ;
  assign \nz.mem [1579] = \nz.mem_1579_sv2v_reg ;
  assign \nz.mem [1578] = \nz.mem_1578_sv2v_reg ;
  assign \nz.mem [1577] = \nz.mem_1577_sv2v_reg ;
  assign \nz.mem [1576] = \nz.mem_1576_sv2v_reg ;
  assign \nz.mem [1575] = \nz.mem_1575_sv2v_reg ;
  assign \nz.mem [1574] = \nz.mem_1574_sv2v_reg ;
  assign \nz.mem [1573] = \nz.mem_1573_sv2v_reg ;
  assign \nz.mem [1572] = \nz.mem_1572_sv2v_reg ;
  assign \nz.mem [1571] = \nz.mem_1571_sv2v_reg ;
  assign \nz.mem [1570] = \nz.mem_1570_sv2v_reg ;
  assign \nz.mem [1569] = \nz.mem_1569_sv2v_reg ;
  assign \nz.mem [1568] = \nz.mem_1568_sv2v_reg ;
  assign \nz.mem [1567] = \nz.mem_1567_sv2v_reg ;
  assign \nz.mem [1566] = \nz.mem_1566_sv2v_reg ;
  assign \nz.mem [1565] = \nz.mem_1565_sv2v_reg ;
  assign \nz.mem [1564] = \nz.mem_1564_sv2v_reg ;
  assign \nz.mem [1563] = \nz.mem_1563_sv2v_reg ;
  assign \nz.mem [1562] = \nz.mem_1562_sv2v_reg ;
  assign \nz.mem [1561] = \nz.mem_1561_sv2v_reg ;
  assign \nz.mem [1560] = \nz.mem_1560_sv2v_reg ;
  assign \nz.mem [1559] = \nz.mem_1559_sv2v_reg ;
  assign \nz.mem [1558] = \nz.mem_1558_sv2v_reg ;
  assign \nz.mem [1557] = \nz.mem_1557_sv2v_reg ;
  assign \nz.mem [1556] = \nz.mem_1556_sv2v_reg ;
  assign \nz.mem [1555] = \nz.mem_1555_sv2v_reg ;
  assign \nz.mem [1554] = \nz.mem_1554_sv2v_reg ;
  assign \nz.mem [1553] = \nz.mem_1553_sv2v_reg ;
  assign \nz.mem [1552] = \nz.mem_1552_sv2v_reg ;
  assign \nz.mem [1551] = \nz.mem_1551_sv2v_reg ;
  assign \nz.mem [1550] = \nz.mem_1550_sv2v_reg ;
  assign \nz.mem [1549] = \nz.mem_1549_sv2v_reg ;
  assign \nz.mem [1548] = \nz.mem_1548_sv2v_reg ;
  assign \nz.mem [1547] = \nz.mem_1547_sv2v_reg ;
  assign \nz.mem [1546] = \nz.mem_1546_sv2v_reg ;
  assign \nz.mem [1545] = \nz.mem_1545_sv2v_reg ;
  assign \nz.mem [1544] = \nz.mem_1544_sv2v_reg ;
  assign \nz.mem [1543] = \nz.mem_1543_sv2v_reg ;
  assign \nz.mem [1542] = \nz.mem_1542_sv2v_reg ;
  assign \nz.mem [1541] = \nz.mem_1541_sv2v_reg ;
  assign \nz.mem [1540] = \nz.mem_1540_sv2v_reg ;
  assign \nz.mem [1539] = \nz.mem_1539_sv2v_reg ;
  assign \nz.mem [1538] = \nz.mem_1538_sv2v_reg ;
  assign \nz.mem [1537] = \nz.mem_1537_sv2v_reg ;
  assign \nz.mem [1536] = \nz.mem_1536_sv2v_reg ;
  assign \nz.mem [1535] = \nz.mem_1535_sv2v_reg ;
  assign \nz.mem [1534] = \nz.mem_1534_sv2v_reg ;
  assign \nz.mem [1533] = \nz.mem_1533_sv2v_reg ;
  assign \nz.mem [1532] = \nz.mem_1532_sv2v_reg ;
  assign \nz.mem [1531] = \nz.mem_1531_sv2v_reg ;
  assign \nz.mem [1530] = \nz.mem_1530_sv2v_reg ;
  assign \nz.mem [1529] = \nz.mem_1529_sv2v_reg ;
  assign \nz.mem [1528] = \nz.mem_1528_sv2v_reg ;
  assign \nz.mem [1527] = \nz.mem_1527_sv2v_reg ;
  assign \nz.mem [1526] = \nz.mem_1526_sv2v_reg ;
  assign \nz.mem [1525] = \nz.mem_1525_sv2v_reg ;
  assign \nz.mem [1524] = \nz.mem_1524_sv2v_reg ;
  assign \nz.mem [1523] = \nz.mem_1523_sv2v_reg ;
  assign \nz.mem [1522] = \nz.mem_1522_sv2v_reg ;
  assign \nz.mem [1521] = \nz.mem_1521_sv2v_reg ;
  assign \nz.mem [1520] = \nz.mem_1520_sv2v_reg ;
  assign \nz.mem [1519] = \nz.mem_1519_sv2v_reg ;
  assign \nz.mem [1518] = \nz.mem_1518_sv2v_reg ;
  assign \nz.mem [1517] = \nz.mem_1517_sv2v_reg ;
  assign \nz.mem [1516] = \nz.mem_1516_sv2v_reg ;
  assign \nz.mem [1515] = \nz.mem_1515_sv2v_reg ;
  assign \nz.mem [1514] = \nz.mem_1514_sv2v_reg ;
  assign \nz.mem [1513] = \nz.mem_1513_sv2v_reg ;
  assign \nz.mem [1512] = \nz.mem_1512_sv2v_reg ;
  assign \nz.mem [1511] = \nz.mem_1511_sv2v_reg ;
  assign \nz.mem [1510] = \nz.mem_1510_sv2v_reg ;
  assign \nz.mem [1509] = \nz.mem_1509_sv2v_reg ;
  assign \nz.mem [1508] = \nz.mem_1508_sv2v_reg ;
  assign \nz.mem [1507] = \nz.mem_1507_sv2v_reg ;
  assign \nz.mem [1506] = \nz.mem_1506_sv2v_reg ;
  assign \nz.mem [1505] = \nz.mem_1505_sv2v_reg ;
  assign \nz.mem [1504] = \nz.mem_1504_sv2v_reg ;
  assign \nz.mem [1503] = \nz.mem_1503_sv2v_reg ;
  assign \nz.mem [1502] = \nz.mem_1502_sv2v_reg ;
  assign \nz.mem [1501] = \nz.mem_1501_sv2v_reg ;
  assign \nz.mem [1500] = \nz.mem_1500_sv2v_reg ;
  assign \nz.mem [1499] = \nz.mem_1499_sv2v_reg ;
  assign \nz.mem [1498] = \nz.mem_1498_sv2v_reg ;
  assign \nz.mem [1497] = \nz.mem_1497_sv2v_reg ;
  assign \nz.mem [1496] = \nz.mem_1496_sv2v_reg ;
  assign \nz.mem [1495] = \nz.mem_1495_sv2v_reg ;
  assign \nz.mem [1494] = \nz.mem_1494_sv2v_reg ;
  assign \nz.mem [1493] = \nz.mem_1493_sv2v_reg ;
  assign \nz.mem [1492] = \nz.mem_1492_sv2v_reg ;
  assign \nz.mem [1491] = \nz.mem_1491_sv2v_reg ;
  assign \nz.mem [1490] = \nz.mem_1490_sv2v_reg ;
  assign \nz.mem [1489] = \nz.mem_1489_sv2v_reg ;
  assign \nz.mem [1488] = \nz.mem_1488_sv2v_reg ;
  assign \nz.mem [1487] = \nz.mem_1487_sv2v_reg ;
  assign \nz.mem [1486] = \nz.mem_1486_sv2v_reg ;
  assign \nz.mem [1485] = \nz.mem_1485_sv2v_reg ;
  assign \nz.mem [1484] = \nz.mem_1484_sv2v_reg ;
  assign \nz.mem [1483] = \nz.mem_1483_sv2v_reg ;
  assign \nz.mem [1482] = \nz.mem_1482_sv2v_reg ;
  assign \nz.mem [1481] = \nz.mem_1481_sv2v_reg ;
  assign \nz.mem [1480] = \nz.mem_1480_sv2v_reg ;
  assign \nz.mem [1479] = \nz.mem_1479_sv2v_reg ;
  assign \nz.mem [1478] = \nz.mem_1478_sv2v_reg ;
  assign \nz.mem [1477] = \nz.mem_1477_sv2v_reg ;
  assign \nz.mem [1476] = \nz.mem_1476_sv2v_reg ;
  assign \nz.mem [1475] = \nz.mem_1475_sv2v_reg ;
  assign \nz.mem [1474] = \nz.mem_1474_sv2v_reg ;
  assign \nz.mem [1473] = \nz.mem_1473_sv2v_reg ;
  assign \nz.mem [1472] = \nz.mem_1472_sv2v_reg ;
  assign \nz.mem [1471] = \nz.mem_1471_sv2v_reg ;
  assign \nz.mem [1470] = \nz.mem_1470_sv2v_reg ;
  assign \nz.mem [1469] = \nz.mem_1469_sv2v_reg ;
  assign \nz.mem [1468] = \nz.mem_1468_sv2v_reg ;
  assign \nz.mem [1467] = \nz.mem_1467_sv2v_reg ;
  assign \nz.mem [1466] = \nz.mem_1466_sv2v_reg ;
  assign \nz.mem [1465] = \nz.mem_1465_sv2v_reg ;
  assign \nz.mem [1464] = \nz.mem_1464_sv2v_reg ;
  assign \nz.mem [1463] = \nz.mem_1463_sv2v_reg ;
  assign \nz.mem [1462] = \nz.mem_1462_sv2v_reg ;
  assign \nz.mem [1461] = \nz.mem_1461_sv2v_reg ;
  assign \nz.mem [1460] = \nz.mem_1460_sv2v_reg ;
  assign \nz.mem [1459] = \nz.mem_1459_sv2v_reg ;
  assign \nz.mem [1458] = \nz.mem_1458_sv2v_reg ;
  assign \nz.mem [1457] = \nz.mem_1457_sv2v_reg ;
  assign \nz.mem [1456] = \nz.mem_1456_sv2v_reg ;
  assign \nz.mem [1455] = \nz.mem_1455_sv2v_reg ;
  assign \nz.mem [1454] = \nz.mem_1454_sv2v_reg ;
  assign \nz.mem [1453] = \nz.mem_1453_sv2v_reg ;
  assign \nz.mem [1452] = \nz.mem_1452_sv2v_reg ;
  assign \nz.mem [1451] = \nz.mem_1451_sv2v_reg ;
  assign \nz.mem [1450] = \nz.mem_1450_sv2v_reg ;
  assign \nz.mem [1449] = \nz.mem_1449_sv2v_reg ;
  assign \nz.mem [1448] = \nz.mem_1448_sv2v_reg ;
  assign \nz.mem [1447] = \nz.mem_1447_sv2v_reg ;
  assign \nz.mem [1446] = \nz.mem_1446_sv2v_reg ;
  assign \nz.mem [1445] = \nz.mem_1445_sv2v_reg ;
  assign \nz.mem [1444] = \nz.mem_1444_sv2v_reg ;
  assign \nz.mem [1443] = \nz.mem_1443_sv2v_reg ;
  assign \nz.mem [1442] = \nz.mem_1442_sv2v_reg ;
  assign \nz.mem [1441] = \nz.mem_1441_sv2v_reg ;
  assign \nz.mem [1440] = \nz.mem_1440_sv2v_reg ;
  assign \nz.mem [1439] = \nz.mem_1439_sv2v_reg ;
  assign \nz.mem [1438] = \nz.mem_1438_sv2v_reg ;
  assign \nz.mem [1437] = \nz.mem_1437_sv2v_reg ;
  assign \nz.mem [1436] = \nz.mem_1436_sv2v_reg ;
  assign \nz.mem [1435] = \nz.mem_1435_sv2v_reg ;
  assign \nz.mem [1434] = \nz.mem_1434_sv2v_reg ;
  assign \nz.mem [1433] = \nz.mem_1433_sv2v_reg ;
  assign \nz.mem [1432] = \nz.mem_1432_sv2v_reg ;
  assign \nz.mem [1431] = \nz.mem_1431_sv2v_reg ;
  assign \nz.mem [1430] = \nz.mem_1430_sv2v_reg ;
  assign \nz.mem [1429] = \nz.mem_1429_sv2v_reg ;
  assign \nz.mem [1428] = \nz.mem_1428_sv2v_reg ;
  assign \nz.mem [1427] = \nz.mem_1427_sv2v_reg ;
  assign \nz.mem [1426] = \nz.mem_1426_sv2v_reg ;
  assign \nz.mem [1425] = \nz.mem_1425_sv2v_reg ;
  assign \nz.mem [1424] = \nz.mem_1424_sv2v_reg ;
  assign \nz.mem [1423] = \nz.mem_1423_sv2v_reg ;
  assign \nz.mem [1422] = \nz.mem_1422_sv2v_reg ;
  assign \nz.mem [1421] = \nz.mem_1421_sv2v_reg ;
  assign \nz.mem [1420] = \nz.mem_1420_sv2v_reg ;
  assign \nz.mem [1419] = \nz.mem_1419_sv2v_reg ;
  assign \nz.mem [1418] = \nz.mem_1418_sv2v_reg ;
  assign \nz.mem [1417] = \nz.mem_1417_sv2v_reg ;
  assign \nz.mem [1416] = \nz.mem_1416_sv2v_reg ;
  assign \nz.mem [1415] = \nz.mem_1415_sv2v_reg ;
  assign \nz.mem [1414] = \nz.mem_1414_sv2v_reg ;
  assign \nz.mem [1413] = \nz.mem_1413_sv2v_reg ;
  assign \nz.mem [1412] = \nz.mem_1412_sv2v_reg ;
  assign \nz.mem [1411] = \nz.mem_1411_sv2v_reg ;
  assign \nz.mem [1410] = \nz.mem_1410_sv2v_reg ;
  assign \nz.mem [1409] = \nz.mem_1409_sv2v_reg ;
  assign \nz.mem [1408] = \nz.mem_1408_sv2v_reg ;
  assign \nz.mem [1407] = \nz.mem_1407_sv2v_reg ;
  assign \nz.mem [1406] = \nz.mem_1406_sv2v_reg ;
  assign \nz.mem [1405] = \nz.mem_1405_sv2v_reg ;
  assign \nz.mem [1404] = \nz.mem_1404_sv2v_reg ;
  assign \nz.mem [1403] = \nz.mem_1403_sv2v_reg ;
  assign \nz.mem [1402] = \nz.mem_1402_sv2v_reg ;
  assign \nz.mem [1401] = \nz.mem_1401_sv2v_reg ;
  assign \nz.mem [1400] = \nz.mem_1400_sv2v_reg ;
  assign \nz.mem [1399] = \nz.mem_1399_sv2v_reg ;
  assign \nz.mem [1398] = \nz.mem_1398_sv2v_reg ;
  assign \nz.mem [1397] = \nz.mem_1397_sv2v_reg ;
  assign \nz.mem [1396] = \nz.mem_1396_sv2v_reg ;
  assign \nz.mem [1395] = \nz.mem_1395_sv2v_reg ;
  assign \nz.mem [1394] = \nz.mem_1394_sv2v_reg ;
  assign \nz.mem [1393] = \nz.mem_1393_sv2v_reg ;
  assign \nz.mem [1392] = \nz.mem_1392_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign N424 = ~w_addr_i[5];
  assign N425 = w_addr_i[3] & w_addr_i[4];
  assign N426 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N427 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N428 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N429 = w_addr_i[5] & N426;
  assign N430 = w_addr_i[5] & N427;
  assign N431 = w_addr_i[5] & N428;
  assign N432 = N424 & N425;
  assign N433 = N424 & N426;
  assign N434 = N424 & N427;
  assign N435 = N424 & N428;
  assign N436 = ~w_addr_i[2];
  assign N437 = w_addr_i[0] & w_addr_i[1];
  assign N438 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N439 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N440 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N441 = w_addr_i[2] & N437;
  assign N442 = w_addr_i[2] & N438;
  assign N443 = w_addr_i[2] & N439;
  assign N444 = w_addr_i[2] & N440;
  assign N445 = N436 & N437;
  assign N446 = N436 & N438;
  assign N447 = N436 & N439;
  assign N448 = N436 & N440;
  assign N373 = N429 & N447;
  assign N372 = N429 & N448;
  assign N371 = N430 & N441;
  assign N370 = N430 & N442;
  assign N369 = N430 & N443;
  assign N368 = N430 & N444;
  assign N367 = N430 & N445;
  assign N366 = N430 & N446;
  assign N365 = N430 & N447;
  assign N364 = N430 & N448;
  assign N363 = N431 & N441;
  assign N362 = N431 & N442;
  assign N361 = N431 & N443;
  assign N360 = N431 & N444;
  assign N359 = N431 & N445;
  assign N358 = N431 & N446;
  assign N357 = N431 & N447;
  assign N356 = N431 & N448;
  assign N355 = N432 & N441;
  assign N354 = N432 & N442;
  assign N353 = N432 & N443;
  assign N352 = N432 & N444;
  assign N351 = N432 & N445;
  assign N350 = N432 & N446;
  assign N349 = N432 & N447;
  assign N348 = N432 & N448;
  assign N347 = N433 & N441;
  assign N346 = N433 & N442;
  assign N345 = N433 & N443;
  assign N344 = N433 & N444;
  assign N343 = N433 & N445;
  assign N342 = N433 & N446;
  assign N341 = N433 & N447;
  assign N340 = N433 & N448;
  assign N339 = N434 & N441;
  assign N338 = N434 & N442;
  assign N337 = N434 & N443;
  assign N336 = N434 & N444;
  assign N335 = N434 & N445;
  assign N334 = N434 & N446;
  assign N333 = N434 & N447;
  assign N332 = N434 & N448;
  assign N331 = N435 & N441;
  assign N330 = N435 & N442;
  assign N329 = N435 & N443;
  assign N328 = N435 & N444;
  assign N327 = N435 & N445;
  assign N326 = N435 & N446;
  assign N325 = N435 & N447;
  assign N324 = N435 & N448;
  assign N8 = N12 & N13;
  assign N9 = N8 & N14;
  assign N10 = N9 & N15;
  assign N11 = N10 & N16;
  assign N273 = N11 & N17;
  assign N12 = ~r_addr_i[5];
  assign N13 = ~r_addr_i[4];
  assign N14 = ~r_addr_i[3];
  assign N15 = ~r_addr_i[2];
  assign N16 = ~r_addr_i[0];
  assign N17 = ~r_addr_i[1];
  assign N18 = r_addr_i[5] & N22;
  assign N19 = N18 & N23;
  assign N20 = N19 & N24;
  assign N21 = N20 & N25;
  assign N274 = N21 & N26;
  assign N22 = ~r_addr_i[4];
  assign N23 = ~r_addr_i[3];
  assign N24 = ~r_addr_i[2];
  assign N25 = ~r_addr_i[0];
  assign N26 = ~r_addr_i[1];
  assign N27 = N31 & N32;
  assign N28 = N27 & N33;
  assign N29 = N28 & N34;
  assign N30 = N29 & r_addr_i[0];
  assign N275 = N30 & N35;
  assign N31 = ~r_addr_i[5];
  assign N32 = ~r_addr_i[4];
  assign N33 = ~r_addr_i[3];
  assign N34 = ~r_addr_i[2];
  assign N35 = ~r_addr_i[1];
  assign N36 = N40 & N41;
  assign N37 = N36 & N42;
  assign N38 = N37 & N43;
  assign N39 = N38 & N44;
  assign N277 = N39 & r_addr_i[1];
  assign N40 = ~r_addr_i[5];
  assign N41 = ~r_addr_i[4];
  assign N42 = ~r_addr_i[3];
  assign N43 = ~r_addr_i[2];
  assign N44 = ~r_addr_i[0];
  assign N45 = N49 & N50;
  assign N46 = N45 & N51;
  assign N47 = N46 & N52;
  assign N48 = N47 & r_addr_i[0];
  assign N279 = N48 & r_addr_i[1];
  assign N49 = ~r_addr_i[5];
  assign N50 = ~r_addr_i[4];
  assign N51 = ~r_addr_i[3];
  assign N52 = ~r_addr_i[2];
  assign N53 = N57 & N58;
  assign N54 = N53 & N59;
  assign N55 = N54 & r_addr_i[2];
  assign N56 = N55 & N60;
  assign N281 = N56 & N61;
  assign N57 = ~r_addr_i[5];
  assign N58 = ~r_addr_i[4];
  assign N59 = ~r_addr_i[3];
  assign N60 = ~r_addr_i[0];
  assign N61 = ~r_addr_i[1];
  assign N62 = N66 & N67;
  assign N63 = N62 & N68;
  assign N64 = N63 & r_addr_i[2];
  assign N65 = N64 & r_addr_i[0];
  assign N283 = N65 & N69;
  assign N66 = ~r_addr_i[5];
  assign N67 = ~r_addr_i[4];
  assign N68 = ~r_addr_i[3];
  assign N69 = ~r_addr_i[1];
  assign N70 = N74 & N75;
  assign N71 = N70 & N76;
  assign N72 = N71 & r_addr_i[2];
  assign N73 = N72 & N77;
  assign N285 = N73 & r_addr_i[1];
  assign N74 = ~r_addr_i[5];
  assign N75 = ~r_addr_i[4];
  assign N76 = ~r_addr_i[3];
  assign N77 = ~r_addr_i[0];
  assign N78 = N82 & N83;
  assign N79 = N78 & N84;
  assign N80 = N79 & r_addr_i[2];
  assign N81 = N80 & r_addr_i[0];
  assign N287 = N81 & r_addr_i[1];
  assign N82 = ~r_addr_i[5];
  assign N83 = ~r_addr_i[4];
  assign N84 = ~r_addr_i[3];
  assign N85 = N89 & N90;
  assign N86 = N85 & r_addr_i[3];
  assign N87 = N86 & N91;
  assign N88 = N87 & N92;
  assign N289 = N88 & N93;
  assign N89 = ~r_addr_i[5];
  assign N90 = ~r_addr_i[4];
  assign N91 = ~r_addr_i[2];
  assign N92 = ~r_addr_i[0];
  assign N93 = ~r_addr_i[1];
  assign N94 = N98 & N99;
  assign N95 = N94 & r_addr_i[3];
  assign N96 = N95 & N100;
  assign N97 = N96 & r_addr_i[0];
  assign N291 = N97 & N101;
  assign N98 = ~r_addr_i[5];
  assign N99 = ~r_addr_i[4];
  assign N100 = ~r_addr_i[2];
  assign N101 = ~r_addr_i[1];
  assign N102 = N106 & N107;
  assign N103 = N102 & r_addr_i[3];
  assign N104 = N103 & N108;
  assign N105 = N104 & N109;
  assign N293 = N105 & r_addr_i[1];
  assign N106 = ~r_addr_i[5];
  assign N107 = ~r_addr_i[4];
  assign N108 = ~r_addr_i[2];
  assign N109 = ~r_addr_i[0];
  assign N110 = N114 & N115;
  assign N111 = N110 & r_addr_i[3];
  assign N112 = N111 & N116;
  assign N113 = N112 & r_addr_i[0];
  assign N295 = N113 & r_addr_i[1];
  assign N114 = ~r_addr_i[5];
  assign N115 = ~r_addr_i[4];
  assign N116 = ~r_addr_i[2];
  assign N117 = N121 & N122;
  assign N118 = N117 & r_addr_i[3];
  assign N119 = N118 & r_addr_i[2];
  assign N120 = N119 & N123;
  assign N297 = N120 & N124;
  assign N121 = ~r_addr_i[5];
  assign N122 = ~r_addr_i[4];
  assign N123 = ~r_addr_i[0];
  assign N124 = ~r_addr_i[1];
  assign N125 = N129 & N130;
  assign N126 = N125 & r_addr_i[3];
  assign N127 = N126 & r_addr_i[2];
  assign N128 = N127 & r_addr_i[0];
  assign N299 = N128 & N131;
  assign N129 = ~r_addr_i[5];
  assign N130 = ~r_addr_i[4];
  assign N131 = ~r_addr_i[1];
  assign N132 = N136 & N137;
  assign N133 = N132 & r_addr_i[3];
  assign N134 = N133 & r_addr_i[2];
  assign N135 = N134 & N138;
  assign N301 = N135 & r_addr_i[1];
  assign N136 = ~r_addr_i[5];
  assign N137 = ~r_addr_i[4];
  assign N138 = ~r_addr_i[0];
  assign N139 = N143 & N144;
  assign N140 = N139 & r_addr_i[3];
  assign N141 = N140 & r_addr_i[2];
  assign N142 = N141 & r_addr_i[0];
  assign N303 = N142 & r_addr_i[1];
  assign N143 = ~r_addr_i[5];
  assign N144 = ~r_addr_i[4];
  assign N145 = N149 & r_addr_i[4];
  assign N146 = N145 & N150;
  assign N147 = N146 & N151;
  assign N148 = N147 & N152;
  assign N305 = N148 & N153;
  assign N149 = ~r_addr_i[5];
  assign N150 = ~r_addr_i[3];
  assign N151 = ~r_addr_i[2];
  assign N152 = ~r_addr_i[0];
  assign N153 = ~r_addr_i[1];
  assign N154 = N158 & r_addr_i[4];
  assign N155 = N154 & N159;
  assign N156 = N155 & N160;
  assign N157 = N156 & r_addr_i[0];
  assign N307 = N157 & N161;
  assign N158 = ~r_addr_i[5];
  assign N159 = ~r_addr_i[3];
  assign N160 = ~r_addr_i[2];
  assign N161 = ~r_addr_i[1];
  assign N309 = r_addr_i[4] & N162 & (N163 & N164) & r_addr_i[1];
  assign N162 = ~r_addr_i[3];
  assign N163 = ~r_addr_i[2];
  assign N164 = ~r_addr_i[0];
  assign N310 = r_addr_i[4] & N165 & (N166 & r_addr_i[0]) & r_addr_i[1];
  assign N165 = ~r_addr_i[3];
  assign N166 = ~r_addr_i[2];
  assign N311 = r_addr_i[4] & N167 & (r_addr_i[2] & N168) & N169;
  assign N167 = ~r_addr_i[3];
  assign N168 = ~r_addr_i[0];
  assign N169 = ~r_addr_i[1];
  assign N312 = r_addr_i[4] & N170 & (r_addr_i[2] & r_addr_i[0]) & N171;
  assign N170 = ~r_addr_i[3];
  assign N171 = ~r_addr_i[1];
  assign N313 = r_addr_i[4] & N172 & (r_addr_i[2] & N173) & r_addr_i[1];
  assign N172 = ~r_addr_i[3];
  assign N173 = ~r_addr_i[0];
  assign N314 = r_addr_i[4] & N174 & (r_addr_i[2] & r_addr_i[0]) & r_addr_i[1];
  assign N174 = ~r_addr_i[3];
  assign N315 = r_addr_i[4] & r_addr_i[3] & (N175 & N176) & N177;
  assign N175 = ~r_addr_i[2];
  assign N176 = ~r_addr_i[0];
  assign N177 = ~r_addr_i[1];
  assign N316 = r_addr_i[4] & r_addr_i[3] & (N178 & r_addr_i[0]) & N179;
  assign N178 = ~r_addr_i[2];
  assign N179 = ~r_addr_i[1];
  assign N317 = r_addr_i[4] & r_addr_i[3] & (N180 & N181) & r_addr_i[1];
  assign N180 = ~r_addr_i[2];
  assign N181 = ~r_addr_i[0];
  assign N318 = r_addr_i[4] & r_addr_i[3] & (N182 & r_addr_i[0]) & r_addr_i[1];
  assign N182 = ~r_addr_i[2];
  assign N319 = r_addr_i[4] & r_addr_i[3] & (r_addr_i[2] & N183) & N184;
  assign N183 = ~r_addr_i[0];
  assign N184 = ~r_addr_i[1];
  assign N320 = r_addr_i[4] & r_addr_i[3] & (r_addr_i[2] & r_addr_i[0]) & N185;
  assign N185 = ~r_addr_i[1];
  assign N321 = r_addr_i[4] & r_addr_i[3] & (r_addr_i[2] & N186) & r_addr_i[1];
  assign N186 = ~r_addr_i[0];
  assign N322 = r_addr_i[4] & r_addr_i[3] & (r_addr_i[2] & r_addr_i[0]) & r_addr_i[1];
  assign N187 = r_addr_i[5] & N191;
  assign N188 = N187 & N192;
  assign N189 = N188 & N193;
  assign N190 = N189 & r_addr_i[0];
  assign N276 = N190 & N194;
  assign N191 = ~r_addr_i[4];
  assign N192 = ~r_addr_i[3];
  assign N193 = ~r_addr_i[2];
  assign N194 = ~r_addr_i[1];
  assign N278 = r_addr_i[5] & N195 & (N196 & N197) & r_addr_i[1];
  assign N195 = ~r_addr_i[3];
  assign N196 = ~r_addr_i[2];
  assign N197 = ~r_addr_i[0];
  assign N280 = r_addr_i[5] & N198 & (N199 & r_addr_i[0]) & r_addr_i[1];
  assign N198 = ~r_addr_i[3];
  assign N199 = ~r_addr_i[2];
  assign N282 = r_addr_i[5] & N200 & (r_addr_i[2] & N201) & N202;
  assign N200 = ~r_addr_i[3];
  assign N201 = ~r_addr_i[0];
  assign N202 = ~r_addr_i[1];
  assign N284 = r_addr_i[5] & N203 & (r_addr_i[2] & r_addr_i[0]) & N204;
  assign N203 = ~r_addr_i[3];
  assign N204 = ~r_addr_i[1];
  assign N286 = r_addr_i[5] & N205 & (r_addr_i[2] & N206) & r_addr_i[1];
  assign N205 = ~r_addr_i[3];
  assign N206 = ~r_addr_i[0];
  assign N288 = r_addr_i[5] & N207 & (r_addr_i[2] & r_addr_i[0]) & r_addr_i[1];
  assign N207 = ~r_addr_i[3];
  assign N290 = r_addr_i[5] & r_addr_i[3] & (N208 & N209) & N210;
  assign N208 = ~r_addr_i[2];
  assign N209 = ~r_addr_i[0];
  assign N210 = ~r_addr_i[1];
  assign N292 = r_addr_i[5] & r_addr_i[3] & (N211 & r_addr_i[0]) & N212;
  assign N211 = ~r_addr_i[2];
  assign N212 = ~r_addr_i[1];
  assign N294 = r_addr_i[5] & r_addr_i[3] & (N213 & N214) & r_addr_i[1];
  assign N213 = ~r_addr_i[2];
  assign N214 = ~r_addr_i[0];
  assign N296 = r_addr_i[5] & r_addr_i[3] & (N215 & r_addr_i[0]) & r_addr_i[1];
  assign N215 = ~r_addr_i[2];
  assign N298 = r_addr_i[5] & r_addr_i[3] & (r_addr_i[2] & N216) & N217;
  assign N216 = ~r_addr_i[0];
  assign N217 = ~r_addr_i[1];
  assign N300 = r_addr_i[5] & r_addr_i[3] & (r_addr_i[2] & r_addr_i[0]) & N218;
  assign N218 = ~r_addr_i[1];
  assign N302 = r_addr_i[5] & r_addr_i[3] & (r_addr_i[2] & N219) & r_addr_i[1];
  assign N219 = ~r_addr_i[0];
  assign N304 = r_addr_i[5] & r_addr_i[3] & (r_addr_i[2] & r_addr_i[0]) & r_addr_i[1];
  assign N306 = r_addr_i[5] & r_addr_i[4] & N220;
  assign N220 = ~r_addr_i[0];
  assign N308 = r_addr_i[5] & r_addr_i[4] & r_addr_i[0];
  assign { N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } = (N221)? { N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324 } : 
                                                                                                                                                                                                                                                                                                                          (N222)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N221 = w_v_i;
  assign N222 = N323;
  assign r_data_o[31] = (N223)? \nz.mem [31] : 
                        (N224)? \nz.mem [63] : 
                        (N225)? \nz.mem [95] : 
                        (N226)? \nz.mem [127] : 
                        (N227)? \nz.mem [159] : 
                        (N228)? \nz.mem [191] : 
                        (N229)? \nz.mem [223] : 
                        (N230)? \nz.mem [255] : 
                        (N231)? \nz.mem [287] : 
                        (N232)? \nz.mem [319] : 
                        (N233)? \nz.mem [351] : 
                        (N234)? \nz.mem [383] : 
                        (N235)? \nz.mem [415] : 
                        (N236)? \nz.mem [447] : 
                        (N237)? \nz.mem [479] : 
                        (N238)? \nz.mem [511] : 
                        (N239)? \nz.mem [543] : 
                        (N240)? \nz.mem [575] : 
                        (N241)? \nz.mem [607] : 
                        (N242)? \nz.mem [639] : 
                        (N243)? \nz.mem [671] : 
                        (N244)? \nz.mem [703] : 
                        (N245)? \nz.mem [735] : 
                        (N246)? \nz.mem [767] : 
                        (N247)? \nz.mem [799] : 
                        (N248)? \nz.mem [831] : 
                        (N249)? \nz.mem [863] : 
                        (N250)? \nz.mem [895] : 
                        (N251)? \nz.mem [927] : 
                        (N252)? \nz.mem [959] : 
                        (N253)? \nz.mem [991] : 
                        (N254)? \nz.mem [1023] : 
                        (N255)? \nz.mem [1055] : 
                        (N256)? \nz.mem [1087] : 
                        (N257)? \nz.mem [1119] : 
                        (N258)? \nz.mem [1151] : 
                        (N259)? \nz.mem [1183] : 
                        (N260)? \nz.mem [1215] : 
                        (N261)? \nz.mem [1247] : 
                        (N262)? \nz.mem [1279] : 
                        (N263)? \nz.mem [1311] : 
                        (N264)? \nz.mem [1343] : 
                        (N265)? \nz.mem [1375] : 
                        (N266)? \nz.mem [1407] : 
                        (N267)? \nz.mem [1439] : 
                        (N268)? \nz.mem [1471] : 
                        (N269)? \nz.mem [1503] : 
                        (N270)? \nz.mem [1535] : 
                        (N271)? \nz.mem [1567] : 
                        (N272)? \nz.mem [1599] : 1'b0;
  assign N223 = N273;
  assign N224 = N275;
  assign N225 = N277;
  assign N226 = N279;
  assign N227 = N281;
  assign N228 = N283;
  assign N229 = N285;
  assign N230 = N287;
  assign N231 = N289;
  assign N232 = N291;
  assign N233 = N293;
  assign N234 = N295;
  assign N235 = N297;
  assign N236 = N299;
  assign N237 = N301;
  assign N238 = N303;
  assign N239 = N305;
  assign N240 = N307;
  assign N241 = N309;
  assign N242 = N310;
  assign N243 = N311;
  assign N244 = N312;
  assign N245 = N313;
  assign N246 = N314;
  assign N247 = N315;
  assign N248 = N316;
  assign N249 = N317;
  assign N250 = N318;
  assign N251 = N319;
  assign N252 = N320;
  assign N253 = N321;
  assign N254 = N322;
  assign N255 = N274;
  assign N256 = N276;
  assign N257 = N278;
  assign N258 = N280;
  assign N259 = N282;
  assign N260 = N284;
  assign N261 = N286;
  assign N262 = N288;
  assign N263 = N290;
  assign N264 = N292;
  assign N265 = N294;
  assign N266 = N296;
  assign N267 = N298;
  assign N268 = N300;
  assign N269 = N302;
  assign N270 = N304;
  assign N271 = N306;
  assign N272 = N308;
  assign r_data_o[30] = (N223)? \nz.mem [30] : 
                        (N224)? \nz.mem [62] : 
                        (N225)? \nz.mem [94] : 
                        (N226)? \nz.mem [126] : 
                        (N227)? \nz.mem [158] : 
                        (N228)? \nz.mem [190] : 
                        (N229)? \nz.mem [222] : 
                        (N230)? \nz.mem [254] : 
                        (N231)? \nz.mem [286] : 
                        (N232)? \nz.mem [318] : 
                        (N233)? \nz.mem [350] : 
                        (N234)? \nz.mem [382] : 
                        (N235)? \nz.mem [414] : 
                        (N236)? \nz.mem [446] : 
                        (N237)? \nz.mem [478] : 
                        (N238)? \nz.mem [510] : 
                        (N239)? \nz.mem [542] : 
                        (N240)? \nz.mem [574] : 
                        (N241)? \nz.mem [606] : 
                        (N242)? \nz.mem [638] : 
                        (N243)? \nz.mem [670] : 
                        (N244)? \nz.mem [702] : 
                        (N245)? \nz.mem [734] : 
                        (N246)? \nz.mem [766] : 
                        (N247)? \nz.mem [798] : 
                        (N248)? \nz.mem [830] : 
                        (N249)? \nz.mem [862] : 
                        (N250)? \nz.mem [894] : 
                        (N251)? \nz.mem [926] : 
                        (N252)? \nz.mem [958] : 
                        (N253)? \nz.mem [990] : 
                        (N254)? \nz.mem [1022] : 
                        (N255)? \nz.mem [1054] : 
                        (N256)? \nz.mem [1086] : 
                        (N257)? \nz.mem [1118] : 
                        (N258)? \nz.mem [1150] : 
                        (N259)? \nz.mem [1182] : 
                        (N260)? \nz.mem [1214] : 
                        (N261)? \nz.mem [1246] : 
                        (N262)? \nz.mem [1278] : 
                        (N263)? \nz.mem [1310] : 
                        (N264)? \nz.mem [1342] : 
                        (N265)? \nz.mem [1374] : 
                        (N266)? \nz.mem [1406] : 
                        (N267)? \nz.mem [1438] : 
                        (N268)? \nz.mem [1470] : 
                        (N269)? \nz.mem [1502] : 
                        (N270)? \nz.mem [1534] : 
                        (N271)? \nz.mem [1566] : 
                        (N272)? \nz.mem [1598] : 1'b0;
  assign r_data_o[29] = (N223)? \nz.mem [29] : 
                        (N224)? \nz.mem [61] : 
                        (N225)? \nz.mem [93] : 
                        (N226)? \nz.mem [125] : 
                        (N227)? \nz.mem [157] : 
                        (N228)? \nz.mem [189] : 
                        (N229)? \nz.mem [221] : 
                        (N230)? \nz.mem [253] : 
                        (N231)? \nz.mem [285] : 
                        (N232)? \nz.mem [317] : 
                        (N233)? \nz.mem [349] : 
                        (N234)? \nz.mem [381] : 
                        (N235)? \nz.mem [413] : 
                        (N236)? \nz.mem [445] : 
                        (N237)? \nz.mem [477] : 
                        (N238)? \nz.mem [509] : 
                        (N239)? \nz.mem [541] : 
                        (N240)? \nz.mem [573] : 
                        (N241)? \nz.mem [605] : 
                        (N242)? \nz.mem [637] : 
                        (N243)? \nz.mem [669] : 
                        (N244)? \nz.mem [701] : 
                        (N245)? \nz.mem [733] : 
                        (N246)? \nz.mem [765] : 
                        (N247)? \nz.mem [797] : 
                        (N248)? \nz.mem [829] : 
                        (N249)? \nz.mem [861] : 
                        (N250)? \nz.mem [893] : 
                        (N251)? \nz.mem [925] : 
                        (N252)? \nz.mem [957] : 
                        (N253)? \nz.mem [989] : 
                        (N254)? \nz.mem [1021] : 
                        (N255)? \nz.mem [1053] : 
                        (N256)? \nz.mem [1085] : 
                        (N257)? \nz.mem [1117] : 
                        (N258)? \nz.mem [1149] : 
                        (N259)? \nz.mem [1181] : 
                        (N260)? \nz.mem [1213] : 
                        (N261)? \nz.mem [1245] : 
                        (N262)? \nz.mem [1277] : 
                        (N263)? \nz.mem [1309] : 
                        (N264)? \nz.mem [1341] : 
                        (N265)? \nz.mem [1373] : 
                        (N266)? \nz.mem [1405] : 
                        (N267)? \nz.mem [1437] : 
                        (N268)? \nz.mem [1469] : 
                        (N269)? \nz.mem [1501] : 
                        (N270)? \nz.mem [1533] : 
                        (N271)? \nz.mem [1565] : 
                        (N272)? \nz.mem [1597] : 1'b0;
  assign r_data_o[28] = (N223)? \nz.mem [28] : 
                        (N224)? \nz.mem [60] : 
                        (N225)? \nz.mem [92] : 
                        (N226)? \nz.mem [124] : 
                        (N227)? \nz.mem [156] : 
                        (N228)? \nz.mem [188] : 
                        (N229)? \nz.mem [220] : 
                        (N230)? \nz.mem [252] : 
                        (N231)? \nz.mem [284] : 
                        (N232)? \nz.mem [316] : 
                        (N233)? \nz.mem [348] : 
                        (N234)? \nz.mem [380] : 
                        (N235)? \nz.mem [412] : 
                        (N236)? \nz.mem [444] : 
                        (N237)? \nz.mem [476] : 
                        (N238)? \nz.mem [508] : 
                        (N239)? \nz.mem [540] : 
                        (N240)? \nz.mem [572] : 
                        (N241)? \nz.mem [604] : 
                        (N242)? \nz.mem [636] : 
                        (N243)? \nz.mem [668] : 
                        (N244)? \nz.mem [700] : 
                        (N245)? \nz.mem [732] : 
                        (N246)? \nz.mem [764] : 
                        (N247)? \nz.mem [796] : 
                        (N248)? \nz.mem [828] : 
                        (N249)? \nz.mem [860] : 
                        (N250)? \nz.mem [892] : 
                        (N251)? \nz.mem [924] : 
                        (N252)? \nz.mem [956] : 
                        (N253)? \nz.mem [988] : 
                        (N254)? \nz.mem [1020] : 
                        (N255)? \nz.mem [1052] : 
                        (N256)? \nz.mem [1084] : 
                        (N257)? \nz.mem [1116] : 
                        (N258)? \nz.mem [1148] : 
                        (N259)? \nz.mem [1180] : 
                        (N260)? \nz.mem [1212] : 
                        (N261)? \nz.mem [1244] : 
                        (N262)? \nz.mem [1276] : 
                        (N263)? \nz.mem [1308] : 
                        (N264)? \nz.mem [1340] : 
                        (N265)? \nz.mem [1372] : 
                        (N266)? \nz.mem [1404] : 
                        (N267)? \nz.mem [1436] : 
                        (N268)? \nz.mem [1468] : 
                        (N269)? \nz.mem [1500] : 
                        (N270)? \nz.mem [1532] : 
                        (N271)? \nz.mem [1564] : 
                        (N272)? \nz.mem [1596] : 1'b0;
  assign r_data_o[27] = (N223)? \nz.mem [27] : 
                        (N224)? \nz.mem [59] : 
                        (N225)? \nz.mem [91] : 
                        (N226)? \nz.mem [123] : 
                        (N227)? \nz.mem [155] : 
                        (N228)? \nz.mem [187] : 
                        (N229)? \nz.mem [219] : 
                        (N230)? \nz.mem [251] : 
                        (N231)? \nz.mem [283] : 
                        (N232)? \nz.mem [315] : 
                        (N233)? \nz.mem [347] : 
                        (N234)? \nz.mem [379] : 
                        (N235)? \nz.mem [411] : 
                        (N236)? \nz.mem [443] : 
                        (N237)? \nz.mem [475] : 
                        (N238)? \nz.mem [507] : 
                        (N239)? \nz.mem [539] : 
                        (N240)? \nz.mem [571] : 
                        (N241)? \nz.mem [603] : 
                        (N242)? \nz.mem [635] : 
                        (N243)? \nz.mem [667] : 
                        (N244)? \nz.mem [699] : 
                        (N245)? \nz.mem [731] : 
                        (N246)? \nz.mem [763] : 
                        (N247)? \nz.mem [795] : 
                        (N248)? \nz.mem [827] : 
                        (N249)? \nz.mem [859] : 
                        (N250)? \nz.mem [891] : 
                        (N251)? \nz.mem [923] : 
                        (N252)? \nz.mem [955] : 
                        (N253)? \nz.mem [987] : 
                        (N254)? \nz.mem [1019] : 
                        (N255)? \nz.mem [1051] : 
                        (N256)? \nz.mem [1083] : 
                        (N257)? \nz.mem [1115] : 
                        (N258)? \nz.mem [1147] : 
                        (N259)? \nz.mem [1179] : 
                        (N260)? \nz.mem [1211] : 
                        (N261)? \nz.mem [1243] : 
                        (N262)? \nz.mem [1275] : 
                        (N263)? \nz.mem [1307] : 
                        (N264)? \nz.mem [1339] : 
                        (N265)? \nz.mem [1371] : 
                        (N266)? \nz.mem [1403] : 
                        (N267)? \nz.mem [1435] : 
                        (N268)? \nz.mem [1467] : 
                        (N269)? \nz.mem [1499] : 
                        (N270)? \nz.mem [1531] : 
                        (N271)? \nz.mem [1563] : 
                        (N272)? \nz.mem [1595] : 1'b0;
  assign r_data_o[26] = (N223)? \nz.mem [26] : 
                        (N224)? \nz.mem [58] : 
                        (N225)? \nz.mem [90] : 
                        (N226)? \nz.mem [122] : 
                        (N227)? \nz.mem [154] : 
                        (N228)? \nz.mem [186] : 
                        (N229)? \nz.mem [218] : 
                        (N230)? \nz.mem [250] : 
                        (N231)? \nz.mem [282] : 
                        (N232)? \nz.mem [314] : 
                        (N233)? \nz.mem [346] : 
                        (N234)? \nz.mem [378] : 
                        (N235)? \nz.mem [410] : 
                        (N236)? \nz.mem [442] : 
                        (N237)? \nz.mem [474] : 
                        (N238)? \nz.mem [506] : 
                        (N239)? \nz.mem [538] : 
                        (N240)? \nz.mem [570] : 
                        (N241)? \nz.mem [602] : 
                        (N242)? \nz.mem [634] : 
                        (N243)? \nz.mem [666] : 
                        (N244)? \nz.mem [698] : 
                        (N245)? \nz.mem [730] : 
                        (N246)? \nz.mem [762] : 
                        (N247)? \nz.mem [794] : 
                        (N248)? \nz.mem [826] : 
                        (N249)? \nz.mem [858] : 
                        (N250)? \nz.mem [890] : 
                        (N251)? \nz.mem [922] : 
                        (N252)? \nz.mem [954] : 
                        (N253)? \nz.mem [986] : 
                        (N254)? \nz.mem [1018] : 
                        (N255)? \nz.mem [1050] : 
                        (N256)? \nz.mem [1082] : 
                        (N257)? \nz.mem [1114] : 
                        (N258)? \nz.mem [1146] : 
                        (N259)? \nz.mem [1178] : 
                        (N260)? \nz.mem [1210] : 
                        (N261)? \nz.mem [1242] : 
                        (N262)? \nz.mem [1274] : 
                        (N263)? \nz.mem [1306] : 
                        (N264)? \nz.mem [1338] : 
                        (N265)? \nz.mem [1370] : 
                        (N266)? \nz.mem [1402] : 
                        (N267)? \nz.mem [1434] : 
                        (N268)? \nz.mem [1466] : 
                        (N269)? \nz.mem [1498] : 
                        (N270)? \nz.mem [1530] : 
                        (N271)? \nz.mem [1562] : 
                        (N272)? \nz.mem [1594] : 1'b0;
  assign r_data_o[25] = (N223)? \nz.mem [25] : 
                        (N224)? \nz.mem [57] : 
                        (N225)? \nz.mem [89] : 
                        (N226)? \nz.mem [121] : 
                        (N227)? \nz.mem [153] : 
                        (N228)? \nz.mem [185] : 
                        (N229)? \nz.mem [217] : 
                        (N230)? \nz.mem [249] : 
                        (N231)? \nz.mem [281] : 
                        (N232)? \nz.mem [313] : 
                        (N233)? \nz.mem [345] : 
                        (N234)? \nz.mem [377] : 
                        (N235)? \nz.mem [409] : 
                        (N236)? \nz.mem [441] : 
                        (N237)? \nz.mem [473] : 
                        (N238)? \nz.mem [505] : 
                        (N239)? \nz.mem [537] : 
                        (N240)? \nz.mem [569] : 
                        (N241)? \nz.mem [601] : 
                        (N242)? \nz.mem [633] : 
                        (N243)? \nz.mem [665] : 
                        (N244)? \nz.mem [697] : 
                        (N245)? \nz.mem [729] : 
                        (N246)? \nz.mem [761] : 
                        (N247)? \nz.mem [793] : 
                        (N248)? \nz.mem [825] : 
                        (N249)? \nz.mem [857] : 
                        (N250)? \nz.mem [889] : 
                        (N251)? \nz.mem [921] : 
                        (N252)? \nz.mem [953] : 
                        (N253)? \nz.mem [985] : 
                        (N254)? \nz.mem [1017] : 
                        (N255)? \nz.mem [1049] : 
                        (N256)? \nz.mem [1081] : 
                        (N257)? \nz.mem [1113] : 
                        (N258)? \nz.mem [1145] : 
                        (N259)? \nz.mem [1177] : 
                        (N260)? \nz.mem [1209] : 
                        (N261)? \nz.mem [1241] : 
                        (N262)? \nz.mem [1273] : 
                        (N263)? \nz.mem [1305] : 
                        (N264)? \nz.mem [1337] : 
                        (N265)? \nz.mem [1369] : 
                        (N266)? \nz.mem [1401] : 
                        (N267)? \nz.mem [1433] : 
                        (N268)? \nz.mem [1465] : 
                        (N269)? \nz.mem [1497] : 
                        (N270)? \nz.mem [1529] : 
                        (N271)? \nz.mem [1561] : 
                        (N272)? \nz.mem [1593] : 1'b0;
  assign r_data_o[24] = (N223)? \nz.mem [24] : 
                        (N224)? \nz.mem [56] : 
                        (N225)? \nz.mem [88] : 
                        (N226)? \nz.mem [120] : 
                        (N227)? \nz.mem [152] : 
                        (N228)? \nz.mem [184] : 
                        (N229)? \nz.mem [216] : 
                        (N230)? \nz.mem [248] : 
                        (N231)? \nz.mem [280] : 
                        (N232)? \nz.mem [312] : 
                        (N233)? \nz.mem [344] : 
                        (N234)? \nz.mem [376] : 
                        (N235)? \nz.mem [408] : 
                        (N236)? \nz.mem [440] : 
                        (N237)? \nz.mem [472] : 
                        (N238)? \nz.mem [504] : 
                        (N239)? \nz.mem [536] : 
                        (N240)? \nz.mem [568] : 
                        (N241)? \nz.mem [600] : 
                        (N242)? \nz.mem [632] : 
                        (N243)? \nz.mem [664] : 
                        (N244)? \nz.mem [696] : 
                        (N245)? \nz.mem [728] : 
                        (N246)? \nz.mem [760] : 
                        (N247)? \nz.mem [792] : 
                        (N248)? \nz.mem [824] : 
                        (N249)? \nz.mem [856] : 
                        (N250)? \nz.mem [888] : 
                        (N251)? \nz.mem [920] : 
                        (N252)? \nz.mem [952] : 
                        (N253)? \nz.mem [984] : 
                        (N254)? \nz.mem [1016] : 
                        (N255)? \nz.mem [1048] : 
                        (N256)? \nz.mem [1080] : 
                        (N257)? \nz.mem [1112] : 
                        (N258)? \nz.mem [1144] : 
                        (N259)? \nz.mem [1176] : 
                        (N260)? \nz.mem [1208] : 
                        (N261)? \nz.mem [1240] : 
                        (N262)? \nz.mem [1272] : 
                        (N263)? \nz.mem [1304] : 
                        (N264)? \nz.mem [1336] : 
                        (N265)? \nz.mem [1368] : 
                        (N266)? \nz.mem [1400] : 
                        (N267)? \nz.mem [1432] : 
                        (N268)? \nz.mem [1464] : 
                        (N269)? \nz.mem [1496] : 
                        (N270)? \nz.mem [1528] : 
                        (N271)? \nz.mem [1560] : 
                        (N272)? \nz.mem [1592] : 1'b0;
  assign r_data_o[23] = (N223)? \nz.mem [23] : 
                        (N224)? \nz.mem [55] : 
                        (N225)? \nz.mem [87] : 
                        (N226)? \nz.mem [119] : 
                        (N227)? \nz.mem [151] : 
                        (N228)? \nz.mem [183] : 
                        (N229)? \nz.mem [215] : 
                        (N230)? \nz.mem [247] : 
                        (N231)? \nz.mem [279] : 
                        (N232)? \nz.mem [311] : 
                        (N233)? \nz.mem [343] : 
                        (N234)? \nz.mem [375] : 
                        (N235)? \nz.mem [407] : 
                        (N236)? \nz.mem [439] : 
                        (N237)? \nz.mem [471] : 
                        (N238)? \nz.mem [503] : 
                        (N239)? \nz.mem [535] : 
                        (N240)? \nz.mem [567] : 
                        (N241)? \nz.mem [599] : 
                        (N242)? \nz.mem [631] : 
                        (N243)? \nz.mem [663] : 
                        (N244)? \nz.mem [695] : 
                        (N245)? \nz.mem [727] : 
                        (N246)? \nz.mem [759] : 
                        (N247)? \nz.mem [791] : 
                        (N248)? \nz.mem [823] : 
                        (N249)? \nz.mem [855] : 
                        (N250)? \nz.mem [887] : 
                        (N251)? \nz.mem [919] : 
                        (N252)? \nz.mem [951] : 
                        (N253)? \nz.mem [983] : 
                        (N254)? \nz.mem [1015] : 
                        (N255)? \nz.mem [1047] : 
                        (N256)? \nz.mem [1079] : 
                        (N257)? \nz.mem [1111] : 
                        (N258)? \nz.mem [1143] : 
                        (N259)? \nz.mem [1175] : 
                        (N260)? \nz.mem [1207] : 
                        (N261)? \nz.mem [1239] : 
                        (N262)? \nz.mem [1271] : 
                        (N263)? \nz.mem [1303] : 
                        (N264)? \nz.mem [1335] : 
                        (N265)? \nz.mem [1367] : 
                        (N266)? \nz.mem [1399] : 
                        (N267)? \nz.mem [1431] : 
                        (N268)? \nz.mem [1463] : 
                        (N269)? \nz.mem [1495] : 
                        (N270)? \nz.mem [1527] : 
                        (N271)? \nz.mem [1559] : 
                        (N272)? \nz.mem [1591] : 1'b0;
  assign r_data_o[22] = (N223)? \nz.mem [22] : 
                        (N224)? \nz.mem [54] : 
                        (N225)? \nz.mem [86] : 
                        (N226)? \nz.mem [118] : 
                        (N227)? \nz.mem [150] : 
                        (N228)? \nz.mem [182] : 
                        (N229)? \nz.mem [214] : 
                        (N230)? \nz.mem [246] : 
                        (N231)? \nz.mem [278] : 
                        (N232)? \nz.mem [310] : 
                        (N233)? \nz.mem [342] : 
                        (N234)? \nz.mem [374] : 
                        (N235)? \nz.mem [406] : 
                        (N236)? \nz.mem [438] : 
                        (N237)? \nz.mem [470] : 
                        (N238)? \nz.mem [502] : 
                        (N239)? \nz.mem [534] : 
                        (N240)? \nz.mem [566] : 
                        (N241)? \nz.mem [598] : 
                        (N242)? \nz.mem [630] : 
                        (N243)? \nz.mem [662] : 
                        (N244)? \nz.mem [694] : 
                        (N245)? \nz.mem [726] : 
                        (N246)? \nz.mem [758] : 
                        (N247)? \nz.mem [790] : 
                        (N248)? \nz.mem [822] : 
                        (N249)? \nz.mem [854] : 
                        (N250)? \nz.mem [886] : 
                        (N251)? \nz.mem [918] : 
                        (N252)? \nz.mem [950] : 
                        (N253)? \nz.mem [982] : 
                        (N254)? \nz.mem [1014] : 
                        (N255)? \nz.mem [1046] : 
                        (N256)? \nz.mem [1078] : 
                        (N257)? \nz.mem [1110] : 
                        (N258)? \nz.mem [1142] : 
                        (N259)? \nz.mem [1174] : 
                        (N260)? \nz.mem [1206] : 
                        (N261)? \nz.mem [1238] : 
                        (N262)? \nz.mem [1270] : 
                        (N263)? \nz.mem [1302] : 
                        (N264)? \nz.mem [1334] : 
                        (N265)? \nz.mem [1366] : 
                        (N266)? \nz.mem [1398] : 
                        (N267)? \nz.mem [1430] : 
                        (N268)? \nz.mem [1462] : 
                        (N269)? \nz.mem [1494] : 
                        (N270)? \nz.mem [1526] : 
                        (N271)? \nz.mem [1558] : 
                        (N272)? \nz.mem [1590] : 1'b0;
  assign r_data_o[21] = (N223)? \nz.mem [21] : 
                        (N224)? \nz.mem [53] : 
                        (N225)? \nz.mem [85] : 
                        (N226)? \nz.mem [117] : 
                        (N227)? \nz.mem [149] : 
                        (N228)? \nz.mem [181] : 
                        (N229)? \nz.mem [213] : 
                        (N230)? \nz.mem [245] : 
                        (N231)? \nz.mem [277] : 
                        (N232)? \nz.mem [309] : 
                        (N233)? \nz.mem [341] : 
                        (N234)? \nz.mem [373] : 
                        (N235)? \nz.mem [405] : 
                        (N236)? \nz.mem [437] : 
                        (N237)? \nz.mem [469] : 
                        (N238)? \nz.mem [501] : 
                        (N239)? \nz.mem [533] : 
                        (N240)? \nz.mem [565] : 
                        (N241)? \nz.mem [597] : 
                        (N242)? \nz.mem [629] : 
                        (N243)? \nz.mem [661] : 
                        (N244)? \nz.mem [693] : 
                        (N245)? \nz.mem [725] : 
                        (N246)? \nz.mem [757] : 
                        (N247)? \nz.mem [789] : 
                        (N248)? \nz.mem [821] : 
                        (N249)? \nz.mem [853] : 
                        (N250)? \nz.mem [885] : 
                        (N251)? \nz.mem [917] : 
                        (N252)? \nz.mem [949] : 
                        (N253)? \nz.mem [981] : 
                        (N254)? \nz.mem [1013] : 
                        (N255)? \nz.mem [1045] : 
                        (N256)? \nz.mem [1077] : 
                        (N257)? \nz.mem [1109] : 
                        (N258)? \nz.mem [1141] : 
                        (N259)? \nz.mem [1173] : 
                        (N260)? \nz.mem [1205] : 
                        (N261)? \nz.mem [1237] : 
                        (N262)? \nz.mem [1269] : 
                        (N263)? \nz.mem [1301] : 
                        (N264)? \nz.mem [1333] : 
                        (N265)? \nz.mem [1365] : 
                        (N266)? \nz.mem [1397] : 
                        (N267)? \nz.mem [1429] : 
                        (N268)? \nz.mem [1461] : 
                        (N269)? \nz.mem [1493] : 
                        (N270)? \nz.mem [1525] : 
                        (N271)? \nz.mem [1557] : 
                        (N272)? \nz.mem [1589] : 1'b0;
  assign r_data_o[20] = (N223)? \nz.mem [20] : 
                        (N224)? \nz.mem [52] : 
                        (N225)? \nz.mem [84] : 
                        (N226)? \nz.mem [116] : 
                        (N227)? \nz.mem [148] : 
                        (N228)? \nz.mem [180] : 
                        (N229)? \nz.mem [212] : 
                        (N230)? \nz.mem [244] : 
                        (N231)? \nz.mem [276] : 
                        (N232)? \nz.mem [308] : 
                        (N233)? \nz.mem [340] : 
                        (N234)? \nz.mem [372] : 
                        (N235)? \nz.mem [404] : 
                        (N236)? \nz.mem [436] : 
                        (N237)? \nz.mem [468] : 
                        (N238)? \nz.mem [500] : 
                        (N239)? \nz.mem [532] : 
                        (N240)? \nz.mem [564] : 
                        (N241)? \nz.mem [596] : 
                        (N242)? \nz.mem [628] : 
                        (N243)? \nz.mem [660] : 
                        (N244)? \nz.mem [692] : 
                        (N245)? \nz.mem [724] : 
                        (N246)? \nz.mem [756] : 
                        (N247)? \nz.mem [788] : 
                        (N248)? \nz.mem [820] : 
                        (N249)? \nz.mem [852] : 
                        (N250)? \nz.mem [884] : 
                        (N251)? \nz.mem [916] : 
                        (N252)? \nz.mem [948] : 
                        (N253)? \nz.mem [980] : 
                        (N254)? \nz.mem [1012] : 
                        (N255)? \nz.mem [1044] : 
                        (N256)? \nz.mem [1076] : 
                        (N257)? \nz.mem [1108] : 
                        (N258)? \nz.mem [1140] : 
                        (N259)? \nz.mem [1172] : 
                        (N260)? \nz.mem [1204] : 
                        (N261)? \nz.mem [1236] : 
                        (N262)? \nz.mem [1268] : 
                        (N263)? \nz.mem [1300] : 
                        (N264)? \nz.mem [1332] : 
                        (N265)? \nz.mem [1364] : 
                        (N266)? \nz.mem [1396] : 
                        (N267)? \nz.mem [1428] : 
                        (N268)? \nz.mem [1460] : 
                        (N269)? \nz.mem [1492] : 
                        (N270)? \nz.mem [1524] : 
                        (N271)? \nz.mem [1556] : 
                        (N272)? \nz.mem [1588] : 1'b0;
  assign r_data_o[19] = (N223)? \nz.mem [19] : 
                        (N224)? \nz.mem [51] : 
                        (N225)? \nz.mem [83] : 
                        (N226)? \nz.mem [115] : 
                        (N227)? \nz.mem [147] : 
                        (N228)? \nz.mem [179] : 
                        (N229)? \nz.mem [211] : 
                        (N230)? \nz.mem [243] : 
                        (N231)? \nz.mem [275] : 
                        (N232)? \nz.mem [307] : 
                        (N233)? \nz.mem [339] : 
                        (N234)? \nz.mem [371] : 
                        (N235)? \nz.mem [403] : 
                        (N236)? \nz.mem [435] : 
                        (N237)? \nz.mem [467] : 
                        (N238)? \nz.mem [499] : 
                        (N239)? \nz.mem [531] : 
                        (N240)? \nz.mem [563] : 
                        (N241)? \nz.mem [595] : 
                        (N242)? \nz.mem [627] : 
                        (N243)? \nz.mem [659] : 
                        (N244)? \nz.mem [691] : 
                        (N245)? \nz.mem [723] : 
                        (N246)? \nz.mem [755] : 
                        (N247)? \nz.mem [787] : 
                        (N248)? \nz.mem [819] : 
                        (N249)? \nz.mem [851] : 
                        (N250)? \nz.mem [883] : 
                        (N251)? \nz.mem [915] : 
                        (N252)? \nz.mem [947] : 
                        (N253)? \nz.mem [979] : 
                        (N254)? \nz.mem [1011] : 
                        (N255)? \nz.mem [1043] : 
                        (N256)? \nz.mem [1075] : 
                        (N257)? \nz.mem [1107] : 
                        (N258)? \nz.mem [1139] : 
                        (N259)? \nz.mem [1171] : 
                        (N260)? \nz.mem [1203] : 
                        (N261)? \nz.mem [1235] : 
                        (N262)? \nz.mem [1267] : 
                        (N263)? \nz.mem [1299] : 
                        (N264)? \nz.mem [1331] : 
                        (N265)? \nz.mem [1363] : 
                        (N266)? \nz.mem [1395] : 
                        (N267)? \nz.mem [1427] : 
                        (N268)? \nz.mem [1459] : 
                        (N269)? \nz.mem [1491] : 
                        (N270)? \nz.mem [1523] : 
                        (N271)? \nz.mem [1555] : 
                        (N272)? \nz.mem [1587] : 1'b0;
  assign r_data_o[18] = (N223)? \nz.mem [18] : 
                        (N224)? \nz.mem [50] : 
                        (N225)? \nz.mem [82] : 
                        (N226)? \nz.mem [114] : 
                        (N227)? \nz.mem [146] : 
                        (N228)? \nz.mem [178] : 
                        (N229)? \nz.mem [210] : 
                        (N230)? \nz.mem [242] : 
                        (N231)? \nz.mem [274] : 
                        (N232)? \nz.mem [306] : 
                        (N233)? \nz.mem [338] : 
                        (N234)? \nz.mem [370] : 
                        (N235)? \nz.mem [402] : 
                        (N236)? \nz.mem [434] : 
                        (N237)? \nz.mem [466] : 
                        (N238)? \nz.mem [498] : 
                        (N239)? \nz.mem [530] : 
                        (N240)? \nz.mem [562] : 
                        (N241)? \nz.mem [594] : 
                        (N242)? \nz.mem [626] : 
                        (N243)? \nz.mem [658] : 
                        (N244)? \nz.mem [690] : 
                        (N245)? \nz.mem [722] : 
                        (N246)? \nz.mem [754] : 
                        (N247)? \nz.mem [786] : 
                        (N248)? \nz.mem [818] : 
                        (N249)? \nz.mem [850] : 
                        (N250)? \nz.mem [882] : 
                        (N251)? \nz.mem [914] : 
                        (N252)? \nz.mem [946] : 
                        (N253)? \nz.mem [978] : 
                        (N254)? \nz.mem [1010] : 
                        (N255)? \nz.mem [1042] : 
                        (N256)? \nz.mem [1074] : 
                        (N257)? \nz.mem [1106] : 
                        (N258)? \nz.mem [1138] : 
                        (N259)? \nz.mem [1170] : 
                        (N260)? \nz.mem [1202] : 
                        (N261)? \nz.mem [1234] : 
                        (N262)? \nz.mem [1266] : 
                        (N263)? \nz.mem [1298] : 
                        (N264)? \nz.mem [1330] : 
                        (N265)? \nz.mem [1362] : 
                        (N266)? \nz.mem [1394] : 
                        (N267)? \nz.mem [1426] : 
                        (N268)? \nz.mem [1458] : 
                        (N269)? \nz.mem [1490] : 
                        (N270)? \nz.mem [1522] : 
                        (N271)? \nz.mem [1554] : 
                        (N272)? \nz.mem [1586] : 1'b0;
  assign r_data_o[17] = (N223)? \nz.mem [17] : 
                        (N224)? \nz.mem [49] : 
                        (N225)? \nz.mem [81] : 
                        (N226)? \nz.mem [113] : 
                        (N227)? \nz.mem [145] : 
                        (N228)? \nz.mem [177] : 
                        (N229)? \nz.mem [209] : 
                        (N230)? \nz.mem [241] : 
                        (N231)? \nz.mem [273] : 
                        (N232)? \nz.mem [305] : 
                        (N233)? \nz.mem [337] : 
                        (N234)? \nz.mem [369] : 
                        (N235)? \nz.mem [401] : 
                        (N236)? \nz.mem [433] : 
                        (N237)? \nz.mem [465] : 
                        (N238)? \nz.mem [497] : 
                        (N239)? \nz.mem [529] : 
                        (N240)? \nz.mem [561] : 
                        (N241)? \nz.mem [593] : 
                        (N242)? \nz.mem [625] : 
                        (N243)? \nz.mem [657] : 
                        (N244)? \nz.mem [689] : 
                        (N245)? \nz.mem [721] : 
                        (N246)? \nz.mem [753] : 
                        (N247)? \nz.mem [785] : 
                        (N248)? \nz.mem [817] : 
                        (N249)? \nz.mem [849] : 
                        (N250)? \nz.mem [881] : 
                        (N251)? \nz.mem [913] : 
                        (N252)? \nz.mem [945] : 
                        (N253)? \nz.mem [977] : 
                        (N254)? \nz.mem [1009] : 
                        (N255)? \nz.mem [1041] : 
                        (N256)? \nz.mem [1073] : 
                        (N257)? \nz.mem [1105] : 
                        (N258)? \nz.mem [1137] : 
                        (N259)? \nz.mem [1169] : 
                        (N260)? \nz.mem [1201] : 
                        (N261)? \nz.mem [1233] : 
                        (N262)? \nz.mem [1265] : 
                        (N263)? \nz.mem [1297] : 
                        (N264)? \nz.mem [1329] : 
                        (N265)? \nz.mem [1361] : 
                        (N266)? \nz.mem [1393] : 
                        (N267)? \nz.mem [1425] : 
                        (N268)? \nz.mem [1457] : 
                        (N269)? \nz.mem [1489] : 
                        (N270)? \nz.mem [1521] : 
                        (N271)? \nz.mem [1553] : 
                        (N272)? \nz.mem [1585] : 1'b0;
  assign r_data_o[16] = (N223)? \nz.mem [16] : 
                        (N224)? \nz.mem [48] : 
                        (N225)? \nz.mem [80] : 
                        (N226)? \nz.mem [112] : 
                        (N227)? \nz.mem [144] : 
                        (N228)? \nz.mem [176] : 
                        (N229)? \nz.mem [208] : 
                        (N230)? \nz.mem [240] : 
                        (N231)? \nz.mem [272] : 
                        (N232)? \nz.mem [304] : 
                        (N233)? \nz.mem [336] : 
                        (N234)? \nz.mem [368] : 
                        (N235)? \nz.mem [400] : 
                        (N236)? \nz.mem [432] : 
                        (N237)? \nz.mem [464] : 
                        (N238)? \nz.mem [496] : 
                        (N239)? \nz.mem [528] : 
                        (N240)? \nz.mem [560] : 
                        (N241)? \nz.mem [592] : 
                        (N242)? \nz.mem [624] : 
                        (N243)? \nz.mem [656] : 
                        (N244)? \nz.mem [688] : 
                        (N245)? \nz.mem [720] : 
                        (N246)? \nz.mem [752] : 
                        (N247)? \nz.mem [784] : 
                        (N248)? \nz.mem [816] : 
                        (N249)? \nz.mem [848] : 
                        (N250)? \nz.mem [880] : 
                        (N251)? \nz.mem [912] : 
                        (N252)? \nz.mem [944] : 
                        (N253)? \nz.mem [976] : 
                        (N254)? \nz.mem [1008] : 
                        (N255)? \nz.mem [1040] : 
                        (N256)? \nz.mem [1072] : 
                        (N257)? \nz.mem [1104] : 
                        (N258)? \nz.mem [1136] : 
                        (N259)? \nz.mem [1168] : 
                        (N260)? \nz.mem [1200] : 
                        (N261)? \nz.mem [1232] : 
                        (N262)? \nz.mem [1264] : 
                        (N263)? \nz.mem [1296] : 
                        (N264)? \nz.mem [1328] : 
                        (N265)? \nz.mem [1360] : 
                        (N266)? \nz.mem [1392] : 
                        (N267)? \nz.mem [1424] : 
                        (N268)? \nz.mem [1456] : 
                        (N269)? \nz.mem [1488] : 
                        (N270)? \nz.mem [1520] : 
                        (N271)? \nz.mem [1552] : 
                        (N272)? \nz.mem [1584] : 1'b0;
  assign r_data_o[15] = (N223)? \nz.mem [15] : 
                        (N224)? \nz.mem [47] : 
                        (N225)? \nz.mem [79] : 
                        (N226)? \nz.mem [111] : 
                        (N227)? \nz.mem [143] : 
                        (N228)? \nz.mem [175] : 
                        (N229)? \nz.mem [207] : 
                        (N230)? \nz.mem [239] : 
                        (N231)? \nz.mem [271] : 
                        (N232)? \nz.mem [303] : 
                        (N233)? \nz.mem [335] : 
                        (N234)? \nz.mem [367] : 
                        (N235)? \nz.mem [399] : 
                        (N236)? \nz.mem [431] : 
                        (N237)? \nz.mem [463] : 
                        (N238)? \nz.mem [495] : 
                        (N239)? \nz.mem [527] : 
                        (N240)? \nz.mem [559] : 
                        (N241)? \nz.mem [591] : 
                        (N242)? \nz.mem [623] : 
                        (N243)? \nz.mem [655] : 
                        (N244)? \nz.mem [687] : 
                        (N245)? \nz.mem [719] : 
                        (N246)? \nz.mem [751] : 
                        (N247)? \nz.mem [783] : 
                        (N248)? \nz.mem [815] : 
                        (N249)? \nz.mem [847] : 
                        (N250)? \nz.mem [879] : 
                        (N251)? \nz.mem [911] : 
                        (N252)? \nz.mem [943] : 
                        (N253)? \nz.mem [975] : 
                        (N254)? \nz.mem [1007] : 
                        (N255)? \nz.mem [1039] : 
                        (N256)? \nz.mem [1071] : 
                        (N257)? \nz.mem [1103] : 
                        (N258)? \nz.mem [1135] : 
                        (N259)? \nz.mem [1167] : 
                        (N260)? \nz.mem [1199] : 
                        (N261)? \nz.mem [1231] : 
                        (N262)? \nz.mem [1263] : 
                        (N263)? \nz.mem [1295] : 
                        (N264)? \nz.mem [1327] : 
                        (N265)? \nz.mem [1359] : 
                        (N266)? \nz.mem [1391] : 
                        (N267)? \nz.mem [1423] : 
                        (N268)? \nz.mem [1455] : 
                        (N269)? \nz.mem [1487] : 
                        (N270)? \nz.mem [1519] : 
                        (N271)? \nz.mem [1551] : 
                        (N272)? \nz.mem [1583] : 1'b0;
  assign r_data_o[14] = (N223)? \nz.mem [14] : 
                        (N224)? \nz.mem [46] : 
                        (N225)? \nz.mem [78] : 
                        (N226)? \nz.mem [110] : 
                        (N227)? \nz.mem [142] : 
                        (N228)? \nz.mem [174] : 
                        (N229)? \nz.mem [206] : 
                        (N230)? \nz.mem [238] : 
                        (N231)? \nz.mem [270] : 
                        (N232)? \nz.mem [302] : 
                        (N233)? \nz.mem [334] : 
                        (N234)? \nz.mem [366] : 
                        (N235)? \nz.mem [398] : 
                        (N236)? \nz.mem [430] : 
                        (N237)? \nz.mem [462] : 
                        (N238)? \nz.mem [494] : 
                        (N239)? \nz.mem [526] : 
                        (N240)? \nz.mem [558] : 
                        (N241)? \nz.mem [590] : 
                        (N242)? \nz.mem [622] : 
                        (N243)? \nz.mem [654] : 
                        (N244)? \nz.mem [686] : 
                        (N245)? \nz.mem [718] : 
                        (N246)? \nz.mem [750] : 
                        (N247)? \nz.mem [782] : 
                        (N248)? \nz.mem [814] : 
                        (N249)? \nz.mem [846] : 
                        (N250)? \nz.mem [878] : 
                        (N251)? \nz.mem [910] : 
                        (N252)? \nz.mem [942] : 
                        (N253)? \nz.mem [974] : 
                        (N254)? \nz.mem [1006] : 
                        (N255)? \nz.mem [1038] : 
                        (N256)? \nz.mem [1070] : 
                        (N257)? \nz.mem [1102] : 
                        (N258)? \nz.mem [1134] : 
                        (N259)? \nz.mem [1166] : 
                        (N260)? \nz.mem [1198] : 
                        (N261)? \nz.mem [1230] : 
                        (N262)? \nz.mem [1262] : 
                        (N263)? \nz.mem [1294] : 
                        (N264)? \nz.mem [1326] : 
                        (N265)? \nz.mem [1358] : 
                        (N266)? \nz.mem [1390] : 
                        (N267)? \nz.mem [1422] : 
                        (N268)? \nz.mem [1454] : 
                        (N269)? \nz.mem [1486] : 
                        (N270)? \nz.mem [1518] : 
                        (N271)? \nz.mem [1550] : 
                        (N272)? \nz.mem [1582] : 1'b0;
  assign r_data_o[13] = (N223)? \nz.mem [13] : 
                        (N224)? \nz.mem [45] : 
                        (N225)? \nz.mem [77] : 
                        (N226)? \nz.mem [109] : 
                        (N227)? \nz.mem [141] : 
                        (N228)? \nz.mem [173] : 
                        (N229)? \nz.mem [205] : 
                        (N230)? \nz.mem [237] : 
                        (N231)? \nz.mem [269] : 
                        (N232)? \nz.mem [301] : 
                        (N233)? \nz.mem [333] : 
                        (N234)? \nz.mem [365] : 
                        (N235)? \nz.mem [397] : 
                        (N236)? \nz.mem [429] : 
                        (N237)? \nz.mem [461] : 
                        (N238)? \nz.mem [493] : 
                        (N239)? \nz.mem [525] : 
                        (N240)? \nz.mem [557] : 
                        (N241)? \nz.mem [589] : 
                        (N242)? \nz.mem [621] : 
                        (N243)? \nz.mem [653] : 
                        (N244)? \nz.mem [685] : 
                        (N245)? \nz.mem [717] : 
                        (N246)? \nz.mem [749] : 
                        (N247)? \nz.mem [781] : 
                        (N248)? \nz.mem [813] : 
                        (N249)? \nz.mem [845] : 
                        (N250)? \nz.mem [877] : 
                        (N251)? \nz.mem [909] : 
                        (N252)? \nz.mem [941] : 
                        (N253)? \nz.mem [973] : 
                        (N254)? \nz.mem [1005] : 
                        (N255)? \nz.mem [1037] : 
                        (N256)? \nz.mem [1069] : 
                        (N257)? \nz.mem [1101] : 
                        (N258)? \nz.mem [1133] : 
                        (N259)? \nz.mem [1165] : 
                        (N260)? \nz.mem [1197] : 
                        (N261)? \nz.mem [1229] : 
                        (N262)? \nz.mem [1261] : 
                        (N263)? \nz.mem [1293] : 
                        (N264)? \nz.mem [1325] : 
                        (N265)? \nz.mem [1357] : 
                        (N266)? \nz.mem [1389] : 
                        (N267)? \nz.mem [1421] : 
                        (N268)? \nz.mem [1453] : 
                        (N269)? \nz.mem [1485] : 
                        (N270)? \nz.mem [1517] : 
                        (N271)? \nz.mem [1549] : 
                        (N272)? \nz.mem [1581] : 1'b0;
  assign r_data_o[12] = (N223)? \nz.mem [12] : 
                        (N224)? \nz.mem [44] : 
                        (N225)? \nz.mem [76] : 
                        (N226)? \nz.mem [108] : 
                        (N227)? \nz.mem [140] : 
                        (N228)? \nz.mem [172] : 
                        (N229)? \nz.mem [204] : 
                        (N230)? \nz.mem [236] : 
                        (N231)? \nz.mem [268] : 
                        (N232)? \nz.mem [300] : 
                        (N233)? \nz.mem [332] : 
                        (N234)? \nz.mem [364] : 
                        (N235)? \nz.mem [396] : 
                        (N236)? \nz.mem [428] : 
                        (N237)? \nz.mem [460] : 
                        (N238)? \nz.mem [492] : 
                        (N239)? \nz.mem [524] : 
                        (N240)? \nz.mem [556] : 
                        (N241)? \nz.mem [588] : 
                        (N242)? \nz.mem [620] : 
                        (N243)? \nz.mem [652] : 
                        (N244)? \nz.mem [684] : 
                        (N245)? \nz.mem [716] : 
                        (N246)? \nz.mem [748] : 
                        (N247)? \nz.mem [780] : 
                        (N248)? \nz.mem [812] : 
                        (N249)? \nz.mem [844] : 
                        (N250)? \nz.mem [876] : 
                        (N251)? \nz.mem [908] : 
                        (N252)? \nz.mem [940] : 
                        (N253)? \nz.mem [972] : 
                        (N254)? \nz.mem [1004] : 
                        (N255)? \nz.mem [1036] : 
                        (N256)? \nz.mem [1068] : 
                        (N257)? \nz.mem [1100] : 
                        (N258)? \nz.mem [1132] : 
                        (N259)? \nz.mem [1164] : 
                        (N260)? \nz.mem [1196] : 
                        (N261)? \nz.mem [1228] : 
                        (N262)? \nz.mem [1260] : 
                        (N263)? \nz.mem [1292] : 
                        (N264)? \nz.mem [1324] : 
                        (N265)? \nz.mem [1356] : 
                        (N266)? \nz.mem [1388] : 
                        (N267)? \nz.mem [1420] : 
                        (N268)? \nz.mem [1452] : 
                        (N269)? \nz.mem [1484] : 
                        (N270)? \nz.mem [1516] : 
                        (N271)? \nz.mem [1548] : 
                        (N272)? \nz.mem [1580] : 1'b0;
  assign r_data_o[11] = (N223)? \nz.mem [11] : 
                        (N224)? \nz.mem [43] : 
                        (N225)? \nz.mem [75] : 
                        (N226)? \nz.mem [107] : 
                        (N227)? \nz.mem [139] : 
                        (N228)? \nz.mem [171] : 
                        (N229)? \nz.mem [203] : 
                        (N230)? \nz.mem [235] : 
                        (N231)? \nz.mem [267] : 
                        (N232)? \nz.mem [299] : 
                        (N233)? \nz.mem [331] : 
                        (N234)? \nz.mem [363] : 
                        (N235)? \nz.mem [395] : 
                        (N236)? \nz.mem [427] : 
                        (N237)? \nz.mem [459] : 
                        (N238)? \nz.mem [491] : 
                        (N239)? \nz.mem [523] : 
                        (N240)? \nz.mem [555] : 
                        (N241)? \nz.mem [587] : 
                        (N242)? \nz.mem [619] : 
                        (N243)? \nz.mem [651] : 
                        (N244)? \nz.mem [683] : 
                        (N245)? \nz.mem [715] : 
                        (N246)? \nz.mem [747] : 
                        (N247)? \nz.mem [779] : 
                        (N248)? \nz.mem [811] : 
                        (N249)? \nz.mem [843] : 
                        (N250)? \nz.mem [875] : 
                        (N251)? \nz.mem [907] : 
                        (N252)? \nz.mem [939] : 
                        (N253)? \nz.mem [971] : 
                        (N254)? \nz.mem [1003] : 
                        (N255)? \nz.mem [1035] : 
                        (N256)? \nz.mem [1067] : 
                        (N257)? \nz.mem [1099] : 
                        (N258)? \nz.mem [1131] : 
                        (N259)? \nz.mem [1163] : 
                        (N260)? \nz.mem [1195] : 
                        (N261)? \nz.mem [1227] : 
                        (N262)? \nz.mem [1259] : 
                        (N263)? \nz.mem [1291] : 
                        (N264)? \nz.mem [1323] : 
                        (N265)? \nz.mem [1355] : 
                        (N266)? \nz.mem [1387] : 
                        (N267)? \nz.mem [1419] : 
                        (N268)? \nz.mem [1451] : 
                        (N269)? \nz.mem [1483] : 
                        (N270)? \nz.mem [1515] : 
                        (N271)? \nz.mem [1547] : 
                        (N272)? \nz.mem [1579] : 1'b0;
  assign r_data_o[10] = (N223)? \nz.mem [10] : 
                        (N224)? \nz.mem [42] : 
                        (N225)? \nz.mem [74] : 
                        (N226)? \nz.mem [106] : 
                        (N227)? \nz.mem [138] : 
                        (N228)? \nz.mem [170] : 
                        (N229)? \nz.mem [202] : 
                        (N230)? \nz.mem [234] : 
                        (N231)? \nz.mem [266] : 
                        (N232)? \nz.mem [298] : 
                        (N233)? \nz.mem [330] : 
                        (N234)? \nz.mem [362] : 
                        (N235)? \nz.mem [394] : 
                        (N236)? \nz.mem [426] : 
                        (N237)? \nz.mem [458] : 
                        (N238)? \nz.mem [490] : 
                        (N239)? \nz.mem [522] : 
                        (N240)? \nz.mem [554] : 
                        (N241)? \nz.mem [586] : 
                        (N242)? \nz.mem [618] : 
                        (N243)? \nz.mem [650] : 
                        (N244)? \nz.mem [682] : 
                        (N245)? \nz.mem [714] : 
                        (N246)? \nz.mem [746] : 
                        (N247)? \nz.mem [778] : 
                        (N248)? \nz.mem [810] : 
                        (N249)? \nz.mem [842] : 
                        (N250)? \nz.mem [874] : 
                        (N251)? \nz.mem [906] : 
                        (N252)? \nz.mem [938] : 
                        (N253)? \nz.mem [970] : 
                        (N254)? \nz.mem [1002] : 
                        (N255)? \nz.mem [1034] : 
                        (N256)? \nz.mem [1066] : 
                        (N257)? \nz.mem [1098] : 
                        (N258)? \nz.mem [1130] : 
                        (N259)? \nz.mem [1162] : 
                        (N260)? \nz.mem [1194] : 
                        (N261)? \nz.mem [1226] : 
                        (N262)? \nz.mem [1258] : 
                        (N263)? \nz.mem [1290] : 
                        (N264)? \nz.mem [1322] : 
                        (N265)? \nz.mem [1354] : 
                        (N266)? \nz.mem [1386] : 
                        (N267)? \nz.mem [1418] : 
                        (N268)? \nz.mem [1450] : 
                        (N269)? \nz.mem [1482] : 
                        (N270)? \nz.mem [1514] : 
                        (N271)? \nz.mem [1546] : 
                        (N272)? \nz.mem [1578] : 1'b0;
  assign r_data_o[9] = (N223)? \nz.mem [9] : 
                       (N224)? \nz.mem [41] : 
                       (N225)? \nz.mem [73] : 
                       (N226)? \nz.mem [105] : 
                       (N227)? \nz.mem [137] : 
                       (N228)? \nz.mem [169] : 
                       (N229)? \nz.mem [201] : 
                       (N230)? \nz.mem [233] : 
                       (N231)? \nz.mem [265] : 
                       (N232)? \nz.mem [297] : 
                       (N233)? \nz.mem [329] : 
                       (N234)? \nz.mem [361] : 
                       (N235)? \nz.mem [393] : 
                       (N236)? \nz.mem [425] : 
                       (N237)? \nz.mem [457] : 
                       (N238)? \nz.mem [489] : 
                       (N239)? \nz.mem [521] : 
                       (N240)? \nz.mem [553] : 
                       (N241)? \nz.mem [585] : 
                       (N242)? \nz.mem [617] : 
                       (N243)? \nz.mem [649] : 
                       (N244)? \nz.mem [681] : 
                       (N245)? \nz.mem [713] : 
                       (N246)? \nz.mem [745] : 
                       (N247)? \nz.mem [777] : 
                       (N248)? \nz.mem [809] : 
                       (N249)? \nz.mem [841] : 
                       (N250)? \nz.mem [873] : 
                       (N251)? \nz.mem [905] : 
                       (N252)? \nz.mem [937] : 
                       (N253)? \nz.mem [969] : 
                       (N254)? \nz.mem [1001] : 
                       (N255)? \nz.mem [1033] : 
                       (N256)? \nz.mem [1065] : 
                       (N257)? \nz.mem [1097] : 
                       (N258)? \nz.mem [1129] : 
                       (N259)? \nz.mem [1161] : 
                       (N260)? \nz.mem [1193] : 
                       (N261)? \nz.mem [1225] : 
                       (N262)? \nz.mem [1257] : 
                       (N263)? \nz.mem [1289] : 
                       (N264)? \nz.mem [1321] : 
                       (N265)? \nz.mem [1353] : 
                       (N266)? \nz.mem [1385] : 
                       (N267)? \nz.mem [1417] : 
                       (N268)? \nz.mem [1449] : 
                       (N269)? \nz.mem [1481] : 
                       (N270)? \nz.mem [1513] : 
                       (N271)? \nz.mem [1545] : 
                       (N272)? \nz.mem [1577] : 1'b0;
  assign r_data_o[8] = (N223)? \nz.mem [8] : 
                       (N224)? \nz.mem [40] : 
                       (N225)? \nz.mem [72] : 
                       (N226)? \nz.mem [104] : 
                       (N227)? \nz.mem [136] : 
                       (N228)? \nz.mem [168] : 
                       (N229)? \nz.mem [200] : 
                       (N230)? \nz.mem [232] : 
                       (N231)? \nz.mem [264] : 
                       (N232)? \nz.mem [296] : 
                       (N233)? \nz.mem [328] : 
                       (N234)? \nz.mem [360] : 
                       (N235)? \nz.mem [392] : 
                       (N236)? \nz.mem [424] : 
                       (N237)? \nz.mem [456] : 
                       (N238)? \nz.mem [488] : 
                       (N239)? \nz.mem [520] : 
                       (N240)? \nz.mem [552] : 
                       (N241)? \nz.mem [584] : 
                       (N242)? \nz.mem [616] : 
                       (N243)? \nz.mem [648] : 
                       (N244)? \nz.mem [680] : 
                       (N245)? \nz.mem [712] : 
                       (N246)? \nz.mem [744] : 
                       (N247)? \nz.mem [776] : 
                       (N248)? \nz.mem [808] : 
                       (N249)? \nz.mem [840] : 
                       (N250)? \nz.mem [872] : 
                       (N251)? \nz.mem [904] : 
                       (N252)? \nz.mem [936] : 
                       (N253)? \nz.mem [968] : 
                       (N254)? \nz.mem [1000] : 
                       (N255)? \nz.mem [1032] : 
                       (N256)? \nz.mem [1064] : 
                       (N257)? \nz.mem [1096] : 
                       (N258)? \nz.mem [1128] : 
                       (N259)? \nz.mem [1160] : 
                       (N260)? \nz.mem [1192] : 
                       (N261)? \nz.mem [1224] : 
                       (N262)? \nz.mem [1256] : 
                       (N263)? \nz.mem [1288] : 
                       (N264)? \nz.mem [1320] : 
                       (N265)? \nz.mem [1352] : 
                       (N266)? \nz.mem [1384] : 
                       (N267)? \nz.mem [1416] : 
                       (N268)? \nz.mem [1448] : 
                       (N269)? \nz.mem [1480] : 
                       (N270)? \nz.mem [1512] : 
                       (N271)? \nz.mem [1544] : 
                       (N272)? \nz.mem [1576] : 1'b0;
  assign r_data_o[7] = (N223)? \nz.mem [7] : 
                       (N224)? \nz.mem [39] : 
                       (N225)? \nz.mem [71] : 
                       (N226)? \nz.mem [103] : 
                       (N227)? \nz.mem [135] : 
                       (N228)? \nz.mem [167] : 
                       (N229)? \nz.mem [199] : 
                       (N230)? \nz.mem [231] : 
                       (N231)? \nz.mem [263] : 
                       (N232)? \nz.mem [295] : 
                       (N233)? \nz.mem [327] : 
                       (N234)? \nz.mem [359] : 
                       (N235)? \nz.mem [391] : 
                       (N236)? \nz.mem [423] : 
                       (N237)? \nz.mem [455] : 
                       (N238)? \nz.mem [487] : 
                       (N239)? \nz.mem [519] : 
                       (N240)? \nz.mem [551] : 
                       (N241)? \nz.mem [583] : 
                       (N242)? \nz.mem [615] : 
                       (N243)? \nz.mem [647] : 
                       (N244)? \nz.mem [679] : 
                       (N245)? \nz.mem [711] : 
                       (N246)? \nz.mem [743] : 
                       (N247)? \nz.mem [775] : 
                       (N248)? \nz.mem [807] : 
                       (N249)? \nz.mem [839] : 
                       (N250)? \nz.mem [871] : 
                       (N251)? \nz.mem [903] : 
                       (N252)? \nz.mem [935] : 
                       (N253)? \nz.mem [967] : 
                       (N254)? \nz.mem [999] : 
                       (N255)? \nz.mem [1031] : 
                       (N256)? \nz.mem [1063] : 
                       (N257)? \nz.mem [1095] : 
                       (N258)? \nz.mem [1127] : 
                       (N259)? \nz.mem [1159] : 
                       (N260)? \nz.mem [1191] : 
                       (N261)? \nz.mem [1223] : 
                       (N262)? \nz.mem [1255] : 
                       (N263)? \nz.mem [1287] : 
                       (N264)? \nz.mem [1319] : 
                       (N265)? \nz.mem [1351] : 
                       (N266)? \nz.mem [1383] : 
                       (N267)? \nz.mem [1415] : 
                       (N268)? \nz.mem [1447] : 
                       (N269)? \nz.mem [1479] : 
                       (N270)? \nz.mem [1511] : 
                       (N271)? \nz.mem [1543] : 
                       (N272)? \nz.mem [1575] : 1'b0;
  assign r_data_o[6] = (N223)? \nz.mem [6] : 
                       (N224)? \nz.mem [38] : 
                       (N225)? \nz.mem [70] : 
                       (N226)? \nz.mem [102] : 
                       (N227)? \nz.mem [134] : 
                       (N228)? \nz.mem [166] : 
                       (N229)? \nz.mem [198] : 
                       (N230)? \nz.mem [230] : 
                       (N231)? \nz.mem [262] : 
                       (N232)? \nz.mem [294] : 
                       (N233)? \nz.mem [326] : 
                       (N234)? \nz.mem [358] : 
                       (N235)? \nz.mem [390] : 
                       (N236)? \nz.mem [422] : 
                       (N237)? \nz.mem [454] : 
                       (N238)? \nz.mem [486] : 
                       (N239)? \nz.mem [518] : 
                       (N240)? \nz.mem [550] : 
                       (N241)? \nz.mem [582] : 
                       (N242)? \nz.mem [614] : 
                       (N243)? \nz.mem [646] : 
                       (N244)? \nz.mem [678] : 
                       (N245)? \nz.mem [710] : 
                       (N246)? \nz.mem [742] : 
                       (N247)? \nz.mem [774] : 
                       (N248)? \nz.mem [806] : 
                       (N249)? \nz.mem [838] : 
                       (N250)? \nz.mem [870] : 
                       (N251)? \nz.mem [902] : 
                       (N252)? \nz.mem [934] : 
                       (N253)? \nz.mem [966] : 
                       (N254)? \nz.mem [998] : 
                       (N255)? \nz.mem [1030] : 
                       (N256)? \nz.mem [1062] : 
                       (N257)? \nz.mem [1094] : 
                       (N258)? \nz.mem [1126] : 
                       (N259)? \nz.mem [1158] : 
                       (N260)? \nz.mem [1190] : 
                       (N261)? \nz.mem [1222] : 
                       (N262)? \nz.mem [1254] : 
                       (N263)? \nz.mem [1286] : 
                       (N264)? \nz.mem [1318] : 
                       (N265)? \nz.mem [1350] : 
                       (N266)? \nz.mem [1382] : 
                       (N267)? \nz.mem [1414] : 
                       (N268)? \nz.mem [1446] : 
                       (N269)? \nz.mem [1478] : 
                       (N270)? \nz.mem [1510] : 
                       (N271)? \nz.mem [1542] : 
                       (N272)? \nz.mem [1574] : 1'b0;
  assign r_data_o[5] = (N223)? \nz.mem [5] : 
                       (N224)? \nz.mem [37] : 
                       (N225)? \nz.mem [69] : 
                       (N226)? \nz.mem [101] : 
                       (N227)? \nz.mem [133] : 
                       (N228)? \nz.mem [165] : 
                       (N229)? \nz.mem [197] : 
                       (N230)? \nz.mem [229] : 
                       (N231)? \nz.mem [261] : 
                       (N232)? \nz.mem [293] : 
                       (N233)? \nz.mem [325] : 
                       (N234)? \nz.mem [357] : 
                       (N235)? \nz.mem [389] : 
                       (N236)? \nz.mem [421] : 
                       (N237)? \nz.mem [453] : 
                       (N238)? \nz.mem [485] : 
                       (N239)? \nz.mem [517] : 
                       (N240)? \nz.mem [549] : 
                       (N241)? \nz.mem [581] : 
                       (N242)? \nz.mem [613] : 
                       (N243)? \nz.mem [645] : 
                       (N244)? \nz.mem [677] : 
                       (N245)? \nz.mem [709] : 
                       (N246)? \nz.mem [741] : 
                       (N247)? \nz.mem [773] : 
                       (N248)? \nz.mem [805] : 
                       (N249)? \nz.mem [837] : 
                       (N250)? \nz.mem [869] : 
                       (N251)? \nz.mem [901] : 
                       (N252)? \nz.mem [933] : 
                       (N253)? \nz.mem [965] : 
                       (N254)? \nz.mem [997] : 
                       (N255)? \nz.mem [1029] : 
                       (N256)? \nz.mem [1061] : 
                       (N257)? \nz.mem [1093] : 
                       (N258)? \nz.mem [1125] : 
                       (N259)? \nz.mem [1157] : 
                       (N260)? \nz.mem [1189] : 
                       (N261)? \nz.mem [1221] : 
                       (N262)? \nz.mem [1253] : 
                       (N263)? \nz.mem [1285] : 
                       (N264)? \nz.mem [1317] : 
                       (N265)? \nz.mem [1349] : 
                       (N266)? \nz.mem [1381] : 
                       (N267)? \nz.mem [1413] : 
                       (N268)? \nz.mem [1445] : 
                       (N269)? \nz.mem [1477] : 
                       (N270)? \nz.mem [1509] : 
                       (N271)? \nz.mem [1541] : 
                       (N272)? \nz.mem [1573] : 1'b0;
  assign r_data_o[4] = (N223)? \nz.mem [4] : 
                       (N224)? \nz.mem [36] : 
                       (N225)? \nz.mem [68] : 
                       (N226)? \nz.mem [100] : 
                       (N227)? \nz.mem [132] : 
                       (N228)? \nz.mem [164] : 
                       (N229)? \nz.mem [196] : 
                       (N230)? \nz.mem [228] : 
                       (N231)? \nz.mem [260] : 
                       (N232)? \nz.mem [292] : 
                       (N233)? \nz.mem [324] : 
                       (N234)? \nz.mem [356] : 
                       (N235)? \nz.mem [388] : 
                       (N236)? \nz.mem [420] : 
                       (N237)? \nz.mem [452] : 
                       (N238)? \nz.mem [484] : 
                       (N239)? \nz.mem [516] : 
                       (N240)? \nz.mem [548] : 
                       (N241)? \nz.mem [580] : 
                       (N242)? \nz.mem [612] : 
                       (N243)? \nz.mem [644] : 
                       (N244)? \nz.mem [676] : 
                       (N245)? \nz.mem [708] : 
                       (N246)? \nz.mem [740] : 
                       (N247)? \nz.mem [772] : 
                       (N248)? \nz.mem [804] : 
                       (N249)? \nz.mem [836] : 
                       (N250)? \nz.mem [868] : 
                       (N251)? \nz.mem [900] : 
                       (N252)? \nz.mem [932] : 
                       (N253)? \nz.mem [964] : 
                       (N254)? \nz.mem [996] : 
                       (N255)? \nz.mem [1028] : 
                       (N256)? \nz.mem [1060] : 
                       (N257)? \nz.mem [1092] : 
                       (N258)? \nz.mem [1124] : 
                       (N259)? \nz.mem [1156] : 
                       (N260)? \nz.mem [1188] : 
                       (N261)? \nz.mem [1220] : 
                       (N262)? \nz.mem [1252] : 
                       (N263)? \nz.mem [1284] : 
                       (N264)? \nz.mem [1316] : 
                       (N265)? \nz.mem [1348] : 
                       (N266)? \nz.mem [1380] : 
                       (N267)? \nz.mem [1412] : 
                       (N268)? \nz.mem [1444] : 
                       (N269)? \nz.mem [1476] : 
                       (N270)? \nz.mem [1508] : 
                       (N271)? \nz.mem [1540] : 
                       (N272)? \nz.mem [1572] : 1'b0;
  assign r_data_o[3] = (N223)? \nz.mem [3] : 
                       (N224)? \nz.mem [35] : 
                       (N225)? \nz.mem [67] : 
                       (N226)? \nz.mem [99] : 
                       (N227)? \nz.mem [131] : 
                       (N228)? \nz.mem [163] : 
                       (N229)? \nz.mem [195] : 
                       (N230)? \nz.mem [227] : 
                       (N231)? \nz.mem [259] : 
                       (N232)? \nz.mem [291] : 
                       (N233)? \nz.mem [323] : 
                       (N234)? \nz.mem [355] : 
                       (N235)? \nz.mem [387] : 
                       (N236)? \nz.mem [419] : 
                       (N237)? \nz.mem [451] : 
                       (N238)? \nz.mem [483] : 
                       (N239)? \nz.mem [515] : 
                       (N240)? \nz.mem [547] : 
                       (N241)? \nz.mem [579] : 
                       (N242)? \nz.mem [611] : 
                       (N243)? \nz.mem [643] : 
                       (N244)? \nz.mem [675] : 
                       (N245)? \nz.mem [707] : 
                       (N246)? \nz.mem [739] : 
                       (N247)? \nz.mem [771] : 
                       (N248)? \nz.mem [803] : 
                       (N249)? \nz.mem [835] : 
                       (N250)? \nz.mem [867] : 
                       (N251)? \nz.mem [899] : 
                       (N252)? \nz.mem [931] : 
                       (N253)? \nz.mem [963] : 
                       (N254)? \nz.mem [995] : 
                       (N255)? \nz.mem [1027] : 
                       (N256)? \nz.mem [1059] : 
                       (N257)? \nz.mem [1091] : 
                       (N258)? \nz.mem [1123] : 
                       (N259)? \nz.mem [1155] : 
                       (N260)? \nz.mem [1187] : 
                       (N261)? \nz.mem [1219] : 
                       (N262)? \nz.mem [1251] : 
                       (N263)? \nz.mem [1283] : 
                       (N264)? \nz.mem [1315] : 
                       (N265)? \nz.mem [1347] : 
                       (N266)? \nz.mem [1379] : 
                       (N267)? \nz.mem [1411] : 
                       (N268)? \nz.mem [1443] : 
                       (N269)? \nz.mem [1475] : 
                       (N270)? \nz.mem [1507] : 
                       (N271)? \nz.mem [1539] : 
                       (N272)? \nz.mem [1571] : 1'b0;
  assign r_data_o[2] = (N223)? \nz.mem [2] : 
                       (N224)? \nz.mem [34] : 
                       (N225)? \nz.mem [66] : 
                       (N226)? \nz.mem [98] : 
                       (N227)? \nz.mem [130] : 
                       (N228)? \nz.mem [162] : 
                       (N229)? \nz.mem [194] : 
                       (N230)? \nz.mem [226] : 
                       (N231)? \nz.mem [258] : 
                       (N232)? \nz.mem [290] : 
                       (N233)? \nz.mem [322] : 
                       (N234)? \nz.mem [354] : 
                       (N235)? \nz.mem [386] : 
                       (N236)? \nz.mem [418] : 
                       (N237)? \nz.mem [450] : 
                       (N238)? \nz.mem [482] : 
                       (N239)? \nz.mem [514] : 
                       (N240)? \nz.mem [546] : 
                       (N241)? \nz.mem [578] : 
                       (N242)? \nz.mem [610] : 
                       (N243)? \nz.mem [642] : 
                       (N244)? \nz.mem [674] : 
                       (N245)? \nz.mem [706] : 
                       (N246)? \nz.mem [738] : 
                       (N247)? \nz.mem [770] : 
                       (N248)? \nz.mem [802] : 
                       (N249)? \nz.mem [834] : 
                       (N250)? \nz.mem [866] : 
                       (N251)? \nz.mem [898] : 
                       (N252)? \nz.mem [930] : 
                       (N253)? \nz.mem [962] : 
                       (N254)? \nz.mem [994] : 
                       (N255)? \nz.mem [1026] : 
                       (N256)? \nz.mem [1058] : 
                       (N257)? \nz.mem [1090] : 
                       (N258)? \nz.mem [1122] : 
                       (N259)? \nz.mem [1154] : 
                       (N260)? \nz.mem [1186] : 
                       (N261)? \nz.mem [1218] : 
                       (N262)? \nz.mem [1250] : 
                       (N263)? \nz.mem [1282] : 
                       (N264)? \nz.mem [1314] : 
                       (N265)? \nz.mem [1346] : 
                       (N266)? \nz.mem [1378] : 
                       (N267)? \nz.mem [1410] : 
                       (N268)? \nz.mem [1442] : 
                       (N269)? \nz.mem [1474] : 
                       (N270)? \nz.mem [1506] : 
                       (N271)? \nz.mem [1538] : 
                       (N272)? \nz.mem [1570] : 1'b0;
  assign r_data_o[1] = (N223)? \nz.mem [1] : 
                       (N224)? \nz.mem [33] : 
                       (N225)? \nz.mem [65] : 
                       (N226)? \nz.mem [97] : 
                       (N227)? \nz.mem [129] : 
                       (N228)? \nz.mem [161] : 
                       (N229)? \nz.mem [193] : 
                       (N230)? \nz.mem [225] : 
                       (N231)? \nz.mem [257] : 
                       (N232)? \nz.mem [289] : 
                       (N233)? \nz.mem [321] : 
                       (N234)? \nz.mem [353] : 
                       (N235)? \nz.mem [385] : 
                       (N236)? \nz.mem [417] : 
                       (N237)? \nz.mem [449] : 
                       (N238)? \nz.mem [481] : 
                       (N239)? \nz.mem [513] : 
                       (N240)? \nz.mem [545] : 
                       (N241)? \nz.mem [577] : 
                       (N242)? \nz.mem [609] : 
                       (N243)? \nz.mem [641] : 
                       (N244)? \nz.mem [673] : 
                       (N245)? \nz.mem [705] : 
                       (N246)? \nz.mem [737] : 
                       (N247)? \nz.mem [769] : 
                       (N248)? \nz.mem [801] : 
                       (N249)? \nz.mem [833] : 
                       (N250)? \nz.mem [865] : 
                       (N251)? \nz.mem [897] : 
                       (N252)? \nz.mem [929] : 
                       (N253)? \nz.mem [961] : 
                       (N254)? \nz.mem [993] : 
                       (N255)? \nz.mem [1025] : 
                       (N256)? \nz.mem [1057] : 
                       (N257)? \nz.mem [1089] : 
                       (N258)? \nz.mem [1121] : 
                       (N259)? \nz.mem [1153] : 
                       (N260)? \nz.mem [1185] : 
                       (N261)? \nz.mem [1217] : 
                       (N262)? \nz.mem [1249] : 
                       (N263)? \nz.mem [1281] : 
                       (N264)? \nz.mem [1313] : 
                       (N265)? \nz.mem [1345] : 
                       (N266)? \nz.mem [1377] : 
                       (N267)? \nz.mem [1409] : 
                       (N268)? \nz.mem [1441] : 
                       (N269)? \nz.mem [1473] : 
                       (N270)? \nz.mem [1505] : 
                       (N271)? \nz.mem [1537] : 
                       (N272)? \nz.mem [1569] : 1'b0;
  assign r_data_o[0] = (N223)? \nz.mem [0] : 
                       (N224)? \nz.mem [32] : 
                       (N225)? \nz.mem [64] : 
                       (N226)? \nz.mem [96] : 
                       (N227)? \nz.mem [128] : 
                       (N228)? \nz.mem [160] : 
                       (N229)? \nz.mem [192] : 
                       (N230)? \nz.mem [224] : 
                       (N231)? \nz.mem [256] : 
                       (N232)? \nz.mem [288] : 
                       (N233)? \nz.mem [320] : 
                       (N234)? \nz.mem [352] : 
                       (N235)? \nz.mem [384] : 
                       (N236)? \nz.mem [416] : 
                       (N237)? \nz.mem [448] : 
                       (N238)? \nz.mem [480] : 
                       (N239)? \nz.mem [512] : 
                       (N240)? \nz.mem [544] : 
                       (N241)? \nz.mem [576] : 
                       (N242)? \nz.mem [608] : 
                       (N243)? \nz.mem [640] : 
                       (N244)? \nz.mem [672] : 
                       (N245)? \nz.mem [704] : 
                       (N246)? \nz.mem [736] : 
                       (N247)? \nz.mem [768] : 
                       (N248)? \nz.mem [800] : 
                       (N249)? \nz.mem [832] : 
                       (N250)? \nz.mem [864] : 
                       (N251)? \nz.mem [896] : 
                       (N252)? \nz.mem [928] : 
                       (N253)? \nz.mem [960] : 
                       (N254)? \nz.mem [992] : 
                       (N255)? \nz.mem [1024] : 
                       (N256)? \nz.mem [1056] : 
                       (N257)? \nz.mem [1088] : 
                       (N258)? \nz.mem [1120] : 
                       (N259)? \nz.mem [1152] : 
                       (N260)? \nz.mem [1184] : 
                       (N261)? \nz.mem [1216] : 
                       (N262)? \nz.mem [1248] : 
                       (N263)? \nz.mem [1280] : 
                       (N264)? \nz.mem [1312] : 
                       (N265)? \nz.mem [1344] : 
                       (N266)? \nz.mem [1376] : 
                       (N267)? \nz.mem [1408] : 
                       (N268)? \nz.mem [1440] : 
                       (N269)? \nz.mem [1472] : 
                       (N270)? \nz.mem [1504] : 
                       (N271)? \nz.mem [1536] : 
                       (N272)? \nz.mem [1568] : 1'b0;
  assign N323 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N423) begin
      \nz.mem_1599_sv2v_reg  <= w_data_i[31];
      \nz.mem_1598_sv2v_reg  <= w_data_i[30];
      \nz.mem_1597_sv2v_reg  <= w_data_i[29];
      \nz.mem_1596_sv2v_reg  <= w_data_i[28];
      \nz.mem_1595_sv2v_reg  <= w_data_i[27];
      \nz.mem_1594_sv2v_reg  <= w_data_i[26];
      \nz.mem_1593_sv2v_reg  <= w_data_i[25];
      \nz.mem_1592_sv2v_reg  <= w_data_i[24];
      \nz.mem_1591_sv2v_reg  <= w_data_i[23];
      \nz.mem_1590_sv2v_reg  <= w_data_i[22];
      \nz.mem_1589_sv2v_reg  <= w_data_i[21];
      \nz.mem_1588_sv2v_reg  <= w_data_i[20];
      \nz.mem_1587_sv2v_reg  <= w_data_i[19];
      \nz.mem_1586_sv2v_reg  <= w_data_i[18];
      \nz.mem_1585_sv2v_reg  <= w_data_i[17];
      \nz.mem_1584_sv2v_reg  <= w_data_i[16];
      \nz.mem_1583_sv2v_reg  <= w_data_i[15];
      \nz.mem_1582_sv2v_reg  <= w_data_i[14];
      \nz.mem_1581_sv2v_reg  <= w_data_i[13];
      \nz.mem_1580_sv2v_reg  <= w_data_i[12];
      \nz.mem_1579_sv2v_reg  <= w_data_i[11];
      \nz.mem_1578_sv2v_reg  <= w_data_i[10];
      \nz.mem_1577_sv2v_reg  <= w_data_i[9];
      \nz.mem_1576_sv2v_reg  <= w_data_i[8];
      \nz.mem_1575_sv2v_reg  <= w_data_i[7];
      \nz.mem_1574_sv2v_reg  <= w_data_i[6];
      \nz.mem_1573_sv2v_reg  <= w_data_i[5];
      \nz.mem_1572_sv2v_reg  <= w_data_i[4];
      \nz.mem_1571_sv2v_reg  <= w_data_i[3];
      \nz.mem_1570_sv2v_reg  <= w_data_i[2];
      \nz.mem_1569_sv2v_reg  <= w_data_i[1];
      \nz.mem_1568_sv2v_reg  <= w_data_i[0];
    end 
    if(N422) begin
      \nz.mem_1567_sv2v_reg  <= w_data_i[31];
      \nz.mem_1566_sv2v_reg  <= w_data_i[30];
      \nz.mem_1565_sv2v_reg  <= w_data_i[29];
      \nz.mem_1564_sv2v_reg  <= w_data_i[28];
      \nz.mem_1563_sv2v_reg  <= w_data_i[27];
      \nz.mem_1562_sv2v_reg  <= w_data_i[26];
      \nz.mem_1561_sv2v_reg  <= w_data_i[25];
      \nz.mem_1560_sv2v_reg  <= w_data_i[24];
      \nz.mem_1559_sv2v_reg  <= w_data_i[23];
      \nz.mem_1558_sv2v_reg  <= w_data_i[22];
      \nz.mem_1557_sv2v_reg  <= w_data_i[21];
      \nz.mem_1556_sv2v_reg  <= w_data_i[20];
      \nz.mem_1555_sv2v_reg  <= w_data_i[19];
      \nz.mem_1554_sv2v_reg  <= w_data_i[18];
      \nz.mem_1553_sv2v_reg  <= w_data_i[17];
      \nz.mem_1552_sv2v_reg  <= w_data_i[16];
      \nz.mem_1551_sv2v_reg  <= w_data_i[15];
      \nz.mem_1550_sv2v_reg  <= w_data_i[14];
      \nz.mem_1549_sv2v_reg  <= w_data_i[13];
      \nz.mem_1548_sv2v_reg  <= w_data_i[12];
      \nz.mem_1547_sv2v_reg  <= w_data_i[11];
      \nz.mem_1546_sv2v_reg  <= w_data_i[10];
      \nz.mem_1545_sv2v_reg  <= w_data_i[9];
      \nz.mem_1544_sv2v_reg  <= w_data_i[8];
      \nz.mem_1543_sv2v_reg  <= w_data_i[7];
      \nz.mem_1542_sv2v_reg  <= w_data_i[6];
      \nz.mem_1541_sv2v_reg  <= w_data_i[5];
      \nz.mem_1540_sv2v_reg  <= w_data_i[4];
      \nz.mem_1539_sv2v_reg  <= w_data_i[3];
      \nz.mem_1538_sv2v_reg  <= w_data_i[2];
      \nz.mem_1537_sv2v_reg  <= w_data_i[1];
      \nz.mem_1536_sv2v_reg  <= w_data_i[0];
    end 
    if(N421) begin
      \nz.mem_1535_sv2v_reg  <= w_data_i[31];
      \nz.mem_1534_sv2v_reg  <= w_data_i[30];
      \nz.mem_1533_sv2v_reg  <= w_data_i[29];
      \nz.mem_1532_sv2v_reg  <= w_data_i[28];
      \nz.mem_1531_sv2v_reg  <= w_data_i[27];
      \nz.mem_1530_sv2v_reg  <= w_data_i[26];
      \nz.mem_1529_sv2v_reg  <= w_data_i[25];
      \nz.mem_1528_sv2v_reg  <= w_data_i[24];
      \nz.mem_1527_sv2v_reg  <= w_data_i[23];
      \nz.mem_1526_sv2v_reg  <= w_data_i[22];
      \nz.mem_1525_sv2v_reg  <= w_data_i[21];
      \nz.mem_1524_sv2v_reg  <= w_data_i[20];
      \nz.mem_1523_sv2v_reg  <= w_data_i[19];
      \nz.mem_1522_sv2v_reg  <= w_data_i[18];
      \nz.mem_1521_sv2v_reg  <= w_data_i[17];
      \nz.mem_1520_sv2v_reg  <= w_data_i[16];
      \nz.mem_1519_sv2v_reg  <= w_data_i[15];
      \nz.mem_1518_sv2v_reg  <= w_data_i[14];
      \nz.mem_1517_sv2v_reg  <= w_data_i[13];
      \nz.mem_1516_sv2v_reg  <= w_data_i[12];
      \nz.mem_1515_sv2v_reg  <= w_data_i[11];
      \nz.mem_1514_sv2v_reg  <= w_data_i[10];
      \nz.mem_1513_sv2v_reg  <= w_data_i[9];
      \nz.mem_1512_sv2v_reg  <= w_data_i[8];
      \nz.mem_1511_sv2v_reg  <= w_data_i[7];
      \nz.mem_1510_sv2v_reg  <= w_data_i[6];
      \nz.mem_1509_sv2v_reg  <= w_data_i[5];
      \nz.mem_1508_sv2v_reg  <= w_data_i[4];
      \nz.mem_1507_sv2v_reg  <= w_data_i[3];
      \nz.mem_1506_sv2v_reg  <= w_data_i[2];
      \nz.mem_1505_sv2v_reg  <= w_data_i[1];
      \nz.mem_1504_sv2v_reg  <= w_data_i[0];
    end 
    if(N420) begin
      \nz.mem_1503_sv2v_reg  <= w_data_i[31];
      \nz.mem_1502_sv2v_reg  <= w_data_i[30];
      \nz.mem_1501_sv2v_reg  <= w_data_i[29];
      \nz.mem_1500_sv2v_reg  <= w_data_i[28];
      \nz.mem_1499_sv2v_reg  <= w_data_i[27];
      \nz.mem_1498_sv2v_reg  <= w_data_i[26];
      \nz.mem_1497_sv2v_reg  <= w_data_i[25];
      \nz.mem_1496_sv2v_reg  <= w_data_i[24];
      \nz.mem_1495_sv2v_reg  <= w_data_i[23];
      \nz.mem_1494_sv2v_reg  <= w_data_i[22];
      \nz.mem_1493_sv2v_reg  <= w_data_i[21];
      \nz.mem_1492_sv2v_reg  <= w_data_i[20];
      \nz.mem_1491_sv2v_reg  <= w_data_i[19];
      \nz.mem_1490_sv2v_reg  <= w_data_i[18];
      \nz.mem_1489_sv2v_reg  <= w_data_i[17];
      \nz.mem_1488_sv2v_reg  <= w_data_i[16];
      \nz.mem_1487_sv2v_reg  <= w_data_i[15];
      \nz.mem_1486_sv2v_reg  <= w_data_i[14];
      \nz.mem_1485_sv2v_reg  <= w_data_i[13];
      \nz.mem_1484_sv2v_reg  <= w_data_i[12];
      \nz.mem_1483_sv2v_reg  <= w_data_i[11];
      \nz.mem_1482_sv2v_reg  <= w_data_i[10];
      \nz.mem_1481_sv2v_reg  <= w_data_i[9];
      \nz.mem_1480_sv2v_reg  <= w_data_i[8];
      \nz.mem_1479_sv2v_reg  <= w_data_i[7];
      \nz.mem_1478_sv2v_reg  <= w_data_i[6];
      \nz.mem_1477_sv2v_reg  <= w_data_i[5];
      \nz.mem_1476_sv2v_reg  <= w_data_i[4];
      \nz.mem_1475_sv2v_reg  <= w_data_i[3];
      \nz.mem_1474_sv2v_reg  <= w_data_i[2];
      \nz.mem_1473_sv2v_reg  <= w_data_i[1];
      \nz.mem_1472_sv2v_reg  <= w_data_i[0];
    end 
    if(N419) begin
      \nz.mem_1471_sv2v_reg  <= w_data_i[31];
      \nz.mem_1470_sv2v_reg  <= w_data_i[30];
      \nz.mem_1469_sv2v_reg  <= w_data_i[29];
      \nz.mem_1468_sv2v_reg  <= w_data_i[28];
      \nz.mem_1467_sv2v_reg  <= w_data_i[27];
      \nz.mem_1466_sv2v_reg  <= w_data_i[26];
      \nz.mem_1465_sv2v_reg  <= w_data_i[25];
      \nz.mem_1464_sv2v_reg  <= w_data_i[24];
      \nz.mem_1463_sv2v_reg  <= w_data_i[23];
      \nz.mem_1462_sv2v_reg  <= w_data_i[22];
      \nz.mem_1461_sv2v_reg  <= w_data_i[21];
      \nz.mem_1460_sv2v_reg  <= w_data_i[20];
      \nz.mem_1459_sv2v_reg  <= w_data_i[19];
      \nz.mem_1458_sv2v_reg  <= w_data_i[18];
      \nz.mem_1457_sv2v_reg  <= w_data_i[17];
      \nz.mem_1456_sv2v_reg  <= w_data_i[16];
      \nz.mem_1455_sv2v_reg  <= w_data_i[15];
      \nz.mem_1454_sv2v_reg  <= w_data_i[14];
      \nz.mem_1453_sv2v_reg  <= w_data_i[13];
      \nz.mem_1452_sv2v_reg  <= w_data_i[12];
      \nz.mem_1451_sv2v_reg  <= w_data_i[11];
      \nz.mem_1450_sv2v_reg  <= w_data_i[10];
      \nz.mem_1449_sv2v_reg  <= w_data_i[9];
      \nz.mem_1448_sv2v_reg  <= w_data_i[8];
      \nz.mem_1447_sv2v_reg  <= w_data_i[7];
      \nz.mem_1446_sv2v_reg  <= w_data_i[6];
      \nz.mem_1445_sv2v_reg  <= w_data_i[5];
      \nz.mem_1444_sv2v_reg  <= w_data_i[4];
      \nz.mem_1443_sv2v_reg  <= w_data_i[3];
      \nz.mem_1442_sv2v_reg  <= w_data_i[2];
      \nz.mem_1441_sv2v_reg  <= w_data_i[1];
      \nz.mem_1440_sv2v_reg  <= w_data_i[0];
    end 
    if(N418) begin
      \nz.mem_1439_sv2v_reg  <= w_data_i[31];
      \nz.mem_1438_sv2v_reg  <= w_data_i[30];
      \nz.mem_1437_sv2v_reg  <= w_data_i[29];
      \nz.mem_1436_sv2v_reg  <= w_data_i[28];
      \nz.mem_1435_sv2v_reg  <= w_data_i[27];
      \nz.mem_1434_sv2v_reg  <= w_data_i[26];
      \nz.mem_1433_sv2v_reg  <= w_data_i[25];
      \nz.mem_1432_sv2v_reg  <= w_data_i[24];
      \nz.mem_1431_sv2v_reg  <= w_data_i[23];
      \nz.mem_1430_sv2v_reg  <= w_data_i[22];
      \nz.mem_1429_sv2v_reg  <= w_data_i[21];
      \nz.mem_1428_sv2v_reg  <= w_data_i[20];
      \nz.mem_1427_sv2v_reg  <= w_data_i[19];
      \nz.mem_1426_sv2v_reg  <= w_data_i[18];
      \nz.mem_1425_sv2v_reg  <= w_data_i[17];
      \nz.mem_1424_sv2v_reg  <= w_data_i[16];
      \nz.mem_1423_sv2v_reg  <= w_data_i[15];
      \nz.mem_1422_sv2v_reg  <= w_data_i[14];
      \nz.mem_1421_sv2v_reg  <= w_data_i[13];
      \nz.mem_1420_sv2v_reg  <= w_data_i[12];
      \nz.mem_1419_sv2v_reg  <= w_data_i[11];
      \nz.mem_1418_sv2v_reg  <= w_data_i[10];
      \nz.mem_1417_sv2v_reg  <= w_data_i[9];
      \nz.mem_1416_sv2v_reg  <= w_data_i[8];
      \nz.mem_1415_sv2v_reg  <= w_data_i[7];
      \nz.mem_1414_sv2v_reg  <= w_data_i[6];
      \nz.mem_1413_sv2v_reg  <= w_data_i[5];
      \nz.mem_1412_sv2v_reg  <= w_data_i[4];
      \nz.mem_1411_sv2v_reg  <= w_data_i[3];
      \nz.mem_1410_sv2v_reg  <= w_data_i[2];
      \nz.mem_1409_sv2v_reg  <= w_data_i[1];
      \nz.mem_1408_sv2v_reg  <= w_data_i[0];
    end 
    if(N417) begin
      \nz.mem_1407_sv2v_reg  <= w_data_i[31];
      \nz.mem_1406_sv2v_reg  <= w_data_i[30];
      \nz.mem_1405_sv2v_reg  <= w_data_i[29];
      \nz.mem_1404_sv2v_reg  <= w_data_i[28];
      \nz.mem_1403_sv2v_reg  <= w_data_i[27];
      \nz.mem_1402_sv2v_reg  <= w_data_i[26];
      \nz.mem_1401_sv2v_reg  <= w_data_i[25];
      \nz.mem_1400_sv2v_reg  <= w_data_i[24];
      \nz.mem_1399_sv2v_reg  <= w_data_i[23];
      \nz.mem_1398_sv2v_reg  <= w_data_i[22];
      \nz.mem_1397_sv2v_reg  <= w_data_i[21];
      \nz.mem_1396_sv2v_reg  <= w_data_i[20];
      \nz.mem_1395_sv2v_reg  <= w_data_i[19];
      \nz.mem_1394_sv2v_reg  <= w_data_i[18];
      \nz.mem_1393_sv2v_reg  <= w_data_i[17];
      \nz.mem_1392_sv2v_reg  <= w_data_i[16];
      \nz.mem_1391_sv2v_reg  <= w_data_i[15];
      \nz.mem_1390_sv2v_reg  <= w_data_i[14];
      \nz.mem_1389_sv2v_reg  <= w_data_i[13];
      \nz.mem_1388_sv2v_reg  <= w_data_i[12];
      \nz.mem_1387_sv2v_reg  <= w_data_i[11];
      \nz.mem_1386_sv2v_reg  <= w_data_i[10];
      \nz.mem_1385_sv2v_reg  <= w_data_i[9];
      \nz.mem_1384_sv2v_reg  <= w_data_i[8];
      \nz.mem_1383_sv2v_reg  <= w_data_i[7];
      \nz.mem_1382_sv2v_reg  <= w_data_i[6];
      \nz.mem_1381_sv2v_reg  <= w_data_i[5];
      \nz.mem_1380_sv2v_reg  <= w_data_i[4];
      \nz.mem_1379_sv2v_reg  <= w_data_i[3];
      \nz.mem_1378_sv2v_reg  <= w_data_i[2];
      \nz.mem_1377_sv2v_reg  <= w_data_i[1];
      \nz.mem_1376_sv2v_reg  <= w_data_i[0];
    end 
    if(N416) begin
      \nz.mem_1375_sv2v_reg  <= w_data_i[31];
      \nz.mem_1374_sv2v_reg  <= w_data_i[30];
      \nz.mem_1373_sv2v_reg  <= w_data_i[29];
      \nz.mem_1372_sv2v_reg  <= w_data_i[28];
      \nz.mem_1371_sv2v_reg  <= w_data_i[27];
      \nz.mem_1370_sv2v_reg  <= w_data_i[26];
      \nz.mem_1369_sv2v_reg  <= w_data_i[25];
      \nz.mem_1368_sv2v_reg  <= w_data_i[24];
      \nz.mem_1367_sv2v_reg  <= w_data_i[23];
      \nz.mem_1366_sv2v_reg  <= w_data_i[22];
      \nz.mem_1365_sv2v_reg  <= w_data_i[21];
      \nz.mem_1364_sv2v_reg  <= w_data_i[20];
      \nz.mem_1363_sv2v_reg  <= w_data_i[19];
      \nz.mem_1362_sv2v_reg  <= w_data_i[18];
      \nz.mem_1361_sv2v_reg  <= w_data_i[17];
      \nz.mem_1360_sv2v_reg  <= w_data_i[16];
      \nz.mem_1359_sv2v_reg  <= w_data_i[15];
      \nz.mem_1358_sv2v_reg  <= w_data_i[14];
      \nz.mem_1357_sv2v_reg  <= w_data_i[13];
      \nz.mem_1356_sv2v_reg  <= w_data_i[12];
      \nz.mem_1355_sv2v_reg  <= w_data_i[11];
      \nz.mem_1354_sv2v_reg  <= w_data_i[10];
      \nz.mem_1353_sv2v_reg  <= w_data_i[9];
      \nz.mem_1352_sv2v_reg  <= w_data_i[8];
      \nz.mem_1351_sv2v_reg  <= w_data_i[7];
      \nz.mem_1350_sv2v_reg  <= w_data_i[6];
      \nz.mem_1349_sv2v_reg  <= w_data_i[5];
      \nz.mem_1348_sv2v_reg  <= w_data_i[4];
      \nz.mem_1347_sv2v_reg  <= w_data_i[3];
      \nz.mem_1346_sv2v_reg  <= w_data_i[2];
      \nz.mem_1345_sv2v_reg  <= w_data_i[1];
      \nz.mem_1344_sv2v_reg  <= w_data_i[0];
    end 
    if(N415) begin
      \nz.mem_1343_sv2v_reg  <= w_data_i[31];
      \nz.mem_1342_sv2v_reg  <= w_data_i[30];
      \nz.mem_1341_sv2v_reg  <= w_data_i[29];
      \nz.mem_1340_sv2v_reg  <= w_data_i[28];
      \nz.mem_1339_sv2v_reg  <= w_data_i[27];
      \nz.mem_1338_sv2v_reg  <= w_data_i[26];
      \nz.mem_1337_sv2v_reg  <= w_data_i[25];
      \nz.mem_1336_sv2v_reg  <= w_data_i[24];
      \nz.mem_1335_sv2v_reg  <= w_data_i[23];
      \nz.mem_1334_sv2v_reg  <= w_data_i[22];
      \nz.mem_1333_sv2v_reg  <= w_data_i[21];
      \nz.mem_1332_sv2v_reg  <= w_data_i[20];
      \nz.mem_1331_sv2v_reg  <= w_data_i[19];
      \nz.mem_1330_sv2v_reg  <= w_data_i[18];
      \nz.mem_1329_sv2v_reg  <= w_data_i[17];
      \nz.mem_1328_sv2v_reg  <= w_data_i[16];
      \nz.mem_1327_sv2v_reg  <= w_data_i[15];
      \nz.mem_1326_sv2v_reg  <= w_data_i[14];
      \nz.mem_1325_sv2v_reg  <= w_data_i[13];
      \nz.mem_1324_sv2v_reg  <= w_data_i[12];
      \nz.mem_1323_sv2v_reg  <= w_data_i[11];
      \nz.mem_1322_sv2v_reg  <= w_data_i[10];
      \nz.mem_1321_sv2v_reg  <= w_data_i[9];
      \nz.mem_1320_sv2v_reg  <= w_data_i[8];
      \nz.mem_1319_sv2v_reg  <= w_data_i[7];
      \nz.mem_1318_sv2v_reg  <= w_data_i[6];
      \nz.mem_1317_sv2v_reg  <= w_data_i[5];
      \nz.mem_1316_sv2v_reg  <= w_data_i[4];
      \nz.mem_1315_sv2v_reg  <= w_data_i[3];
      \nz.mem_1314_sv2v_reg  <= w_data_i[2];
      \nz.mem_1313_sv2v_reg  <= w_data_i[1];
      \nz.mem_1312_sv2v_reg  <= w_data_i[0];
    end 
    if(N414) begin
      \nz.mem_1311_sv2v_reg  <= w_data_i[31];
      \nz.mem_1310_sv2v_reg  <= w_data_i[30];
      \nz.mem_1309_sv2v_reg  <= w_data_i[29];
      \nz.mem_1308_sv2v_reg  <= w_data_i[28];
      \nz.mem_1307_sv2v_reg  <= w_data_i[27];
      \nz.mem_1306_sv2v_reg  <= w_data_i[26];
      \nz.mem_1305_sv2v_reg  <= w_data_i[25];
      \nz.mem_1304_sv2v_reg  <= w_data_i[24];
      \nz.mem_1303_sv2v_reg  <= w_data_i[23];
      \nz.mem_1302_sv2v_reg  <= w_data_i[22];
      \nz.mem_1301_sv2v_reg  <= w_data_i[21];
      \nz.mem_1300_sv2v_reg  <= w_data_i[20];
      \nz.mem_1299_sv2v_reg  <= w_data_i[19];
      \nz.mem_1298_sv2v_reg  <= w_data_i[18];
      \nz.mem_1297_sv2v_reg  <= w_data_i[17];
      \nz.mem_1296_sv2v_reg  <= w_data_i[16];
      \nz.mem_1295_sv2v_reg  <= w_data_i[15];
      \nz.mem_1294_sv2v_reg  <= w_data_i[14];
      \nz.mem_1293_sv2v_reg  <= w_data_i[13];
      \nz.mem_1292_sv2v_reg  <= w_data_i[12];
      \nz.mem_1291_sv2v_reg  <= w_data_i[11];
      \nz.mem_1290_sv2v_reg  <= w_data_i[10];
      \nz.mem_1289_sv2v_reg  <= w_data_i[9];
      \nz.mem_1288_sv2v_reg  <= w_data_i[8];
      \nz.mem_1287_sv2v_reg  <= w_data_i[7];
      \nz.mem_1286_sv2v_reg  <= w_data_i[6];
      \nz.mem_1285_sv2v_reg  <= w_data_i[5];
      \nz.mem_1284_sv2v_reg  <= w_data_i[4];
      \nz.mem_1283_sv2v_reg  <= w_data_i[3];
      \nz.mem_1282_sv2v_reg  <= w_data_i[2];
      \nz.mem_1281_sv2v_reg  <= w_data_i[1];
      \nz.mem_1280_sv2v_reg  <= w_data_i[0];
    end 
    if(N413) begin
      \nz.mem_1279_sv2v_reg  <= w_data_i[31];
      \nz.mem_1278_sv2v_reg  <= w_data_i[30];
      \nz.mem_1277_sv2v_reg  <= w_data_i[29];
      \nz.mem_1276_sv2v_reg  <= w_data_i[28];
      \nz.mem_1275_sv2v_reg  <= w_data_i[27];
      \nz.mem_1274_sv2v_reg  <= w_data_i[26];
      \nz.mem_1273_sv2v_reg  <= w_data_i[25];
      \nz.mem_1272_sv2v_reg  <= w_data_i[24];
      \nz.mem_1271_sv2v_reg  <= w_data_i[23];
      \nz.mem_1270_sv2v_reg  <= w_data_i[22];
      \nz.mem_1269_sv2v_reg  <= w_data_i[21];
      \nz.mem_1268_sv2v_reg  <= w_data_i[20];
      \nz.mem_1267_sv2v_reg  <= w_data_i[19];
      \nz.mem_1266_sv2v_reg  <= w_data_i[18];
      \nz.mem_1265_sv2v_reg  <= w_data_i[17];
      \nz.mem_1264_sv2v_reg  <= w_data_i[16];
      \nz.mem_1263_sv2v_reg  <= w_data_i[15];
      \nz.mem_1262_sv2v_reg  <= w_data_i[14];
      \nz.mem_1261_sv2v_reg  <= w_data_i[13];
      \nz.mem_1260_sv2v_reg  <= w_data_i[12];
      \nz.mem_1259_sv2v_reg  <= w_data_i[11];
      \nz.mem_1258_sv2v_reg  <= w_data_i[10];
      \nz.mem_1257_sv2v_reg  <= w_data_i[9];
      \nz.mem_1256_sv2v_reg  <= w_data_i[8];
      \nz.mem_1255_sv2v_reg  <= w_data_i[7];
      \nz.mem_1254_sv2v_reg  <= w_data_i[6];
      \nz.mem_1253_sv2v_reg  <= w_data_i[5];
      \nz.mem_1252_sv2v_reg  <= w_data_i[4];
      \nz.mem_1251_sv2v_reg  <= w_data_i[3];
      \nz.mem_1250_sv2v_reg  <= w_data_i[2];
      \nz.mem_1249_sv2v_reg  <= w_data_i[1];
      \nz.mem_1248_sv2v_reg  <= w_data_i[0];
    end 
    if(N412) begin
      \nz.mem_1247_sv2v_reg  <= w_data_i[31];
      \nz.mem_1246_sv2v_reg  <= w_data_i[30];
      \nz.mem_1245_sv2v_reg  <= w_data_i[29];
      \nz.mem_1244_sv2v_reg  <= w_data_i[28];
      \nz.mem_1243_sv2v_reg  <= w_data_i[27];
      \nz.mem_1242_sv2v_reg  <= w_data_i[26];
      \nz.mem_1241_sv2v_reg  <= w_data_i[25];
      \nz.mem_1240_sv2v_reg  <= w_data_i[24];
      \nz.mem_1239_sv2v_reg  <= w_data_i[23];
      \nz.mem_1238_sv2v_reg  <= w_data_i[22];
      \nz.mem_1237_sv2v_reg  <= w_data_i[21];
      \nz.mem_1236_sv2v_reg  <= w_data_i[20];
      \nz.mem_1235_sv2v_reg  <= w_data_i[19];
      \nz.mem_1234_sv2v_reg  <= w_data_i[18];
      \nz.mem_1233_sv2v_reg  <= w_data_i[17];
      \nz.mem_1232_sv2v_reg  <= w_data_i[16];
      \nz.mem_1231_sv2v_reg  <= w_data_i[15];
      \nz.mem_1230_sv2v_reg  <= w_data_i[14];
      \nz.mem_1229_sv2v_reg  <= w_data_i[13];
      \nz.mem_1228_sv2v_reg  <= w_data_i[12];
      \nz.mem_1227_sv2v_reg  <= w_data_i[11];
      \nz.mem_1226_sv2v_reg  <= w_data_i[10];
      \nz.mem_1225_sv2v_reg  <= w_data_i[9];
      \nz.mem_1224_sv2v_reg  <= w_data_i[8];
      \nz.mem_1223_sv2v_reg  <= w_data_i[7];
      \nz.mem_1222_sv2v_reg  <= w_data_i[6];
      \nz.mem_1221_sv2v_reg  <= w_data_i[5];
      \nz.mem_1220_sv2v_reg  <= w_data_i[4];
      \nz.mem_1219_sv2v_reg  <= w_data_i[3];
      \nz.mem_1218_sv2v_reg  <= w_data_i[2];
      \nz.mem_1217_sv2v_reg  <= w_data_i[1];
      \nz.mem_1216_sv2v_reg  <= w_data_i[0];
    end 
    if(N411) begin
      \nz.mem_1215_sv2v_reg  <= w_data_i[31];
      \nz.mem_1214_sv2v_reg  <= w_data_i[30];
      \nz.mem_1213_sv2v_reg  <= w_data_i[29];
      \nz.mem_1212_sv2v_reg  <= w_data_i[28];
      \nz.mem_1211_sv2v_reg  <= w_data_i[27];
      \nz.mem_1210_sv2v_reg  <= w_data_i[26];
      \nz.mem_1209_sv2v_reg  <= w_data_i[25];
      \nz.mem_1208_sv2v_reg  <= w_data_i[24];
      \nz.mem_1207_sv2v_reg  <= w_data_i[23];
      \nz.mem_1206_sv2v_reg  <= w_data_i[22];
      \nz.mem_1205_sv2v_reg  <= w_data_i[21];
      \nz.mem_1204_sv2v_reg  <= w_data_i[20];
      \nz.mem_1203_sv2v_reg  <= w_data_i[19];
      \nz.mem_1202_sv2v_reg  <= w_data_i[18];
      \nz.mem_1201_sv2v_reg  <= w_data_i[17];
      \nz.mem_1200_sv2v_reg  <= w_data_i[16];
      \nz.mem_1199_sv2v_reg  <= w_data_i[15];
      \nz.mem_1198_sv2v_reg  <= w_data_i[14];
      \nz.mem_1197_sv2v_reg  <= w_data_i[13];
      \nz.mem_1196_sv2v_reg  <= w_data_i[12];
      \nz.mem_1195_sv2v_reg  <= w_data_i[11];
      \nz.mem_1194_sv2v_reg  <= w_data_i[10];
      \nz.mem_1193_sv2v_reg  <= w_data_i[9];
      \nz.mem_1192_sv2v_reg  <= w_data_i[8];
      \nz.mem_1191_sv2v_reg  <= w_data_i[7];
      \nz.mem_1190_sv2v_reg  <= w_data_i[6];
      \nz.mem_1189_sv2v_reg  <= w_data_i[5];
      \nz.mem_1188_sv2v_reg  <= w_data_i[4];
      \nz.mem_1187_sv2v_reg  <= w_data_i[3];
      \nz.mem_1186_sv2v_reg  <= w_data_i[2];
      \nz.mem_1185_sv2v_reg  <= w_data_i[1];
      \nz.mem_1184_sv2v_reg  <= w_data_i[0];
    end 
    if(N410) begin
      \nz.mem_1183_sv2v_reg  <= w_data_i[31];
      \nz.mem_1182_sv2v_reg  <= w_data_i[30];
      \nz.mem_1181_sv2v_reg  <= w_data_i[29];
      \nz.mem_1180_sv2v_reg  <= w_data_i[28];
      \nz.mem_1179_sv2v_reg  <= w_data_i[27];
      \nz.mem_1178_sv2v_reg  <= w_data_i[26];
      \nz.mem_1177_sv2v_reg  <= w_data_i[25];
      \nz.mem_1176_sv2v_reg  <= w_data_i[24];
      \nz.mem_1175_sv2v_reg  <= w_data_i[23];
      \nz.mem_1174_sv2v_reg  <= w_data_i[22];
      \nz.mem_1173_sv2v_reg  <= w_data_i[21];
      \nz.mem_1172_sv2v_reg  <= w_data_i[20];
      \nz.mem_1171_sv2v_reg  <= w_data_i[19];
      \nz.mem_1170_sv2v_reg  <= w_data_i[18];
      \nz.mem_1169_sv2v_reg  <= w_data_i[17];
      \nz.mem_1168_sv2v_reg  <= w_data_i[16];
      \nz.mem_1167_sv2v_reg  <= w_data_i[15];
      \nz.mem_1166_sv2v_reg  <= w_data_i[14];
      \nz.mem_1165_sv2v_reg  <= w_data_i[13];
      \nz.mem_1164_sv2v_reg  <= w_data_i[12];
      \nz.mem_1163_sv2v_reg  <= w_data_i[11];
      \nz.mem_1162_sv2v_reg  <= w_data_i[10];
      \nz.mem_1161_sv2v_reg  <= w_data_i[9];
      \nz.mem_1160_sv2v_reg  <= w_data_i[8];
      \nz.mem_1159_sv2v_reg  <= w_data_i[7];
      \nz.mem_1158_sv2v_reg  <= w_data_i[6];
      \nz.mem_1157_sv2v_reg  <= w_data_i[5];
      \nz.mem_1156_sv2v_reg  <= w_data_i[4];
      \nz.mem_1155_sv2v_reg  <= w_data_i[3];
      \nz.mem_1154_sv2v_reg  <= w_data_i[2];
      \nz.mem_1153_sv2v_reg  <= w_data_i[1];
      \nz.mem_1152_sv2v_reg  <= w_data_i[0];
    end 
    if(N409) begin
      \nz.mem_1151_sv2v_reg  <= w_data_i[31];
      \nz.mem_1150_sv2v_reg  <= w_data_i[30];
      \nz.mem_1149_sv2v_reg  <= w_data_i[29];
      \nz.mem_1148_sv2v_reg  <= w_data_i[28];
      \nz.mem_1147_sv2v_reg  <= w_data_i[27];
      \nz.mem_1146_sv2v_reg  <= w_data_i[26];
      \nz.mem_1145_sv2v_reg  <= w_data_i[25];
      \nz.mem_1144_sv2v_reg  <= w_data_i[24];
      \nz.mem_1143_sv2v_reg  <= w_data_i[23];
      \nz.mem_1142_sv2v_reg  <= w_data_i[22];
      \nz.mem_1141_sv2v_reg  <= w_data_i[21];
      \nz.mem_1140_sv2v_reg  <= w_data_i[20];
      \nz.mem_1139_sv2v_reg  <= w_data_i[19];
      \nz.mem_1138_sv2v_reg  <= w_data_i[18];
      \nz.mem_1137_sv2v_reg  <= w_data_i[17];
      \nz.mem_1136_sv2v_reg  <= w_data_i[16];
      \nz.mem_1135_sv2v_reg  <= w_data_i[15];
      \nz.mem_1134_sv2v_reg  <= w_data_i[14];
      \nz.mem_1133_sv2v_reg  <= w_data_i[13];
      \nz.mem_1132_sv2v_reg  <= w_data_i[12];
      \nz.mem_1131_sv2v_reg  <= w_data_i[11];
      \nz.mem_1130_sv2v_reg  <= w_data_i[10];
      \nz.mem_1129_sv2v_reg  <= w_data_i[9];
      \nz.mem_1128_sv2v_reg  <= w_data_i[8];
      \nz.mem_1127_sv2v_reg  <= w_data_i[7];
      \nz.mem_1126_sv2v_reg  <= w_data_i[6];
      \nz.mem_1125_sv2v_reg  <= w_data_i[5];
      \nz.mem_1124_sv2v_reg  <= w_data_i[4];
      \nz.mem_1123_sv2v_reg  <= w_data_i[3];
      \nz.mem_1122_sv2v_reg  <= w_data_i[2];
      \nz.mem_1121_sv2v_reg  <= w_data_i[1];
      \nz.mem_1120_sv2v_reg  <= w_data_i[0];
    end 
    if(N408) begin
      \nz.mem_1119_sv2v_reg  <= w_data_i[31];
      \nz.mem_1118_sv2v_reg  <= w_data_i[30];
      \nz.mem_1117_sv2v_reg  <= w_data_i[29];
      \nz.mem_1116_sv2v_reg  <= w_data_i[28];
      \nz.mem_1115_sv2v_reg  <= w_data_i[27];
      \nz.mem_1114_sv2v_reg  <= w_data_i[26];
      \nz.mem_1113_sv2v_reg  <= w_data_i[25];
      \nz.mem_1112_sv2v_reg  <= w_data_i[24];
      \nz.mem_1111_sv2v_reg  <= w_data_i[23];
      \nz.mem_1110_sv2v_reg  <= w_data_i[22];
      \nz.mem_1109_sv2v_reg  <= w_data_i[21];
      \nz.mem_1108_sv2v_reg  <= w_data_i[20];
      \nz.mem_1107_sv2v_reg  <= w_data_i[19];
      \nz.mem_1106_sv2v_reg  <= w_data_i[18];
      \nz.mem_1105_sv2v_reg  <= w_data_i[17];
      \nz.mem_1104_sv2v_reg  <= w_data_i[16];
      \nz.mem_1103_sv2v_reg  <= w_data_i[15];
      \nz.mem_1102_sv2v_reg  <= w_data_i[14];
      \nz.mem_1101_sv2v_reg  <= w_data_i[13];
      \nz.mem_1100_sv2v_reg  <= w_data_i[12];
      \nz.mem_1099_sv2v_reg  <= w_data_i[11];
      \nz.mem_1098_sv2v_reg  <= w_data_i[10];
      \nz.mem_1097_sv2v_reg  <= w_data_i[9];
      \nz.mem_1096_sv2v_reg  <= w_data_i[8];
      \nz.mem_1095_sv2v_reg  <= w_data_i[7];
      \nz.mem_1094_sv2v_reg  <= w_data_i[6];
      \nz.mem_1093_sv2v_reg  <= w_data_i[5];
      \nz.mem_1092_sv2v_reg  <= w_data_i[4];
      \nz.mem_1091_sv2v_reg  <= w_data_i[3];
      \nz.mem_1090_sv2v_reg  <= w_data_i[2];
      \nz.mem_1089_sv2v_reg  <= w_data_i[1];
      \nz.mem_1088_sv2v_reg  <= w_data_i[0];
    end 
    if(N407) begin
      \nz.mem_1087_sv2v_reg  <= w_data_i[31];
      \nz.mem_1086_sv2v_reg  <= w_data_i[30];
      \nz.mem_1085_sv2v_reg  <= w_data_i[29];
      \nz.mem_1084_sv2v_reg  <= w_data_i[28];
      \nz.mem_1083_sv2v_reg  <= w_data_i[27];
      \nz.mem_1082_sv2v_reg  <= w_data_i[26];
      \nz.mem_1081_sv2v_reg  <= w_data_i[25];
      \nz.mem_1080_sv2v_reg  <= w_data_i[24];
      \nz.mem_1079_sv2v_reg  <= w_data_i[23];
      \nz.mem_1078_sv2v_reg  <= w_data_i[22];
      \nz.mem_1077_sv2v_reg  <= w_data_i[21];
      \nz.mem_1076_sv2v_reg  <= w_data_i[20];
      \nz.mem_1075_sv2v_reg  <= w_data_i[19];
      \nz.mem_1074_sv2v_reg  <= w_data_i[18];
      \nz.mem_1073_sv2v_reg  <= w_data_i[17];
      \nz.mem_1072_sv2v_reg  <= w_data_i[16];
      \nz.mem_1071_sv2v_reg  <= w_data_i[15];
      \nz.mem_1070_sv2v_reg  <= w_data_i[14];
      \nz.mem_1069_sv2v_reg  <= w_data_i[13];
      \nz.mem_1068_sv2v_reg  <= w_data_i[12];
      \nz.mem_1067_sv2v_reg  <= w_data_i[11];
      \nz.mem_1066_sv2v_reg  <= w_data_i[10];
      \nz.mem_1065_sv2v_reg  <= w_data_i[9];
      \nz.mem_1064_sv2v_reg  <= w_data_i[8];
      \nz.mem_1063_sv2v_reg  <= w_data_i[7];
      \nz.mem_1062_sv2v_reg  <= w_data_i[6];
      \nz.mem_1061_sv2v_reg  <= w_data_i[5];
      \nz.mem_1060_sv2v_reg  <= w_data_i[4];
      \nz.mem_1059_sv2v_reg  <= w_data_i[3];
      \nz.mem_1058_sv2v_reg  <= w_data_i[2];
      \nz.mem_1057_sv2v_reg  <= w_data_i[1];
      \nz.mem_1056_sv2v_reg  <= w_data_i[0];
    end 
    if(N406) begin
      \nz.mem_1055_sv2v_reg  <= w_data_i[31];
      \nz.mem_1054_sv2v_reg  <= w_data_i[30];
      \nz.mem_1053_sv2v_reg  <= w_data_i[29];
      \nz.mem_1052_sv2v_reg  <= w_data_i[28];
      \nz.mem_1051_sv2v_reg  <= w_data_i[27];
      \nz.mem_1050_sv2v_reg  <= w_data_i[26];
      \nz.mem_1049_sv2v_reg  <= w_data_i[25];
      \nz.mem_1048_sv2v_reg  <= w_data_i[24];
      \nz.mem_1047_sv2v_reg  <= w_data_i[23];
      \nz.mem_1046_sv2v_reg  <= w_data_i[22];
      \nz.mem_1045_sv2v_reg  <= w_data_i[21];
      \nz.mem_1044_sv2v_reg  <= w_data_i[20];
      \nz.mem_1043_sv2v_reg  <= w_data_i[19];
      \nz.mem_1042_sv2v_reg  <= w_data_i[18];
      \nz.mem_1041_sv2v_reg  <= w_data_i[17];
      \nz.mem_1040_sv2v_reg  <= w_data_i[16];
      \nz.mem_1039_sv2v_reg  <= w_data_i[15];
      \nz.mem_1038_sv2v_reg  <= w_data_i[14];
      \nz.mem_1037_sv2v_reg  <= w_data_i[13];
      \nz.mem_1036_sv2v_reg  <= w_data_i[12];
      \nz.mem_1035_sv2v_reg  <= w_data_i[11];
      \nz.mem_1034_sv2v_reg  <= w_data_i[10];
      \nz.mem_1033_sv2v_reg  <= w_data_i[9];
      \nz.mem_1032_sv2v_reg  <= w_data_i[8];
      \nz.mem_1031_sv2v_reg  <= w_data_i[7];
      \nz.mem_1030_sv2v_reg  <= w_data_i[6];
      \nz.mem_1029_sv2v_reg  <= w_data_i[5];
      \nz.mem_1028_sv2v_reg  <= w_data_i[4];
      \nz.mem_1027_sv2v_reg  <= w_data_i[3];
      \nz.mem_1026_sv2v_reg  <= w_data_i[2];
      \nz.mem_1025_sv2v_reg  <= w_data_i[1];
      \nz.mem_1024_sv2v_reg  <= w_data_i[0];
    end 
    if(N405) begin
      \nz.mem_1023_sv2v_reg  <= w_data_i[31];
      \nz.mem_1022_sv2v_reg  <= w_data_i[30];
      \nz.mem_1021_sv2v_reg  <= w_data_i[29];
      \nz.mem_1020_sv2v_reg  <= w_data_i[28];
      \nz.mem_1019_sv2v_reg  <= w_data_i[27];
      \nz.mem_1018_sv2v_reg  <= w_data_i[26];
      \nz.mem_1017_sv2v_reg  <= w_data_i[25];
      \nz.mem_1016_sv2v_reg  <= w_data_i[24];
      \nz.mem_1015_sv2v_reg  <= w_data_i[23];
      \nz.mem_1014_sv2v_reg  <= w_data_i[22];
      \nz.mem_1013_sv2v_reg  <= w_data_i[21];
      \nz.mem_1012_sv2v_reg  <= w_data_i[20];
      \nz.mem_1011_sv2v_reg  <= w_data_i[19];
      \nz.mem_1010_sv2v_reg  <= w_data_i[18];
      \nz.mem_1009_sv2v_reg  <= w_data_i[17];
      \nz.mem_1008_sv2v_reg  <= w_data_i[16];
      \nz.mem_1007_sv2v_reg  <= w_data_i[15];
      \nz.mem_1006_sv2v_reg  <= w_data_i[14];
      \nz.mem_1005_sv2v_reg  <= w_data_i[13];
      \nz.mem_1004_sv2v_reg  <= w_data_i[12];
      \nz.mem_1003_sv2v_reg  <= w_data_i[11];
      \nz.mem_1002_sv2v_reg  <= w_data_i[10];
      \nz.mem_1001_sv2v_reg  <= w_data_i[9];
      \nz.mem_1000_sv2v_reg  <= w_data_i[8];
      \nz.mem_999_sv2v_reg  <= w_data_i[7];
      \nz.mem_998_sv2v_reg  <= w_data_i[6];
      \nz.mem_997_sv2v_reg  <= w_data_i[5];
      \nz.mem_996_sv2v_reg  <= w_data_i[4];
      \nz.mem_995_sv2v_reg  <= w_data_i[3];
      \nz.mem_994_sv2v_reg  <= w_data_i[2];
      \nz.mem_993_sv2v_reg  <= w_data_i[1];
      \nz.mem_992_sv2v_reg  <= w_data_i[0];
    end 
    if(N404) begin
      \nz.mem_991_sv2v_reg  <= w_data_i[31];
      \nz.mem_990_sv2v_reg  <= w_data_i[30];
      \nz.mem_989_sv2v_reg  <= w_data_i[29];
      \nz.mem_988_sv2v_reg  <= w_data_i[28];
      \nz.mem_987_sv2v_reg  <= w_data_i[27];
      \nz.mem_986_sv2v_reg  <= w_data_i[26];
      \nz.mem_985_sv2v_reg  <= w_data_i[25];
      \nz.mem_984_sv2v_reg  <= w_data_i[24];
      \nz.mem_983_sv2v_reg  <= w_data_i[23];
      \nz.mem_982_sv2v_reg  <= w_data_i[22];
      \nz.mem_981_sv2v_reg  <= w_data_i[21];
      \nz.mem_980_sv2v_reg  <= w_data_i[20];
      \nz.mem_979_sv2v_reg  <= w_data_i[19];
      \nz.mem_978_sv2v_reg  <= w_data_i[18];
      \nz.mem_977_sv2v_reg  <= w_data_i[17];
      \nz.mem_976_sv2v_reg  <= w_data_i[16];
      \nz.mem_975_sv2v_reg  <= w_data_i[15];
      \nz.mem_974_sv2v_reg  <= w_data_i[14];
      \nz.mem_973_sv2v_reg  <= w_data_i[13];
      \nz.mem_972_sv2v_reg  <= w_data_i[12];
      \nz.mem_971_sv2v_reg  <= w_data_i[11];
      \nz.mem_970_sv2v_reg  <= w_data_i[10];
      \nz.mem_969_sv2v_reg  <= w_data_i[9];
      \nz.mem_968_sv2v_reg  <= w_data_i[8];
      \nz.mem_967_sv2v_reg  <= w_data_i[7];
      \nz.mem_966_sv2v_reg  <= w_data_i[6];
      \nz.mem_965_sv2v_reg  <= w_data_i[5];
      \nz.mem_964_sv2v_reg  <= w_data_i[4];
      \nz.mem_963_sv2v_reg  <= w_data_i[3];
      \nz.mem_962_sv2v_reg  <= w_data_i[2];
      \nz.mem_961_sv2v_reg  <= w_data_i[1];
      \nz.mem_960_sv2v_reg  <= w_data_i[0];
    end 
    if(N403) begin
      \nz.mem_959_sv2v_reg  <= w_data_i[31];
      \nz.mem_958_sv2v_reg  <= w_data_i[30];
      \nz.mem_957_sv2v_reg  <= w_data_i[29];
      \nz.mem_956_sv2v_reg  <= w_data_i[28];
      \nz.mem_955_sv2v_reg  <= w_data_i[27];
      \nz.mem_954_sv2v_reg  <= w_data_i[26];
      \nz.mem_953_sv2v_reg  <= w_data_i[25];
      \nz.mem_952_sv2v_reg  <= w_data_i[24];
      \nz.mem_951_sv2v_reg  <= w_data_i[23];
      \nz.mem_950_sv2v_reg  <= w_data_i[22];
      \nz.mem_949_sv2v_reg  <= w_data_i[21];
      \nz.mem_948_sv2v_reg  <= w_data_i[20];
      \nz.mem_947_sv2v_reg  <= w_data_i[19];
      \nz.mem_946_sv2v_reg  <= w_data_i[18];
      \nz.mem_945_sv2v_reg  <= w_data_i[17];
      \nz.mem_944_sv2v_reg  <= w_data_i[16];
      \nz.mem_943_sv2v_reg  <= w_data_i[15];
      \nz.mem_942_sv2v_reg  <= w_data_i[14];
      \nz.mem_941_sv2v_reg  <= w_data_i[13];
      \nz.mem_940_sv2v_reg  <= w_data_i[12];
      \nz.mem_939_sv2v_reg  <= w_data_i[11];
      \nz.mem_938_sv2v_reg  <= w_data_i[10];
      \nz.mem_937_sv2v_reg  <= w_data_i[9];
      \nz.mem_936_sv2v_reg  <= w_data_i[8];
      \nz.mem_935_sv2v_reg  <= w_data_i[7];
      \nz.mem_934_sv2v_reg  <= w_data_i[6];
      \nz.mem_933_sv2v_reg  <= w_data_i[5];
      \nz.mem_932_sv2v_reg  <= w_data_i[4];
      \nz.mem_931_sv2v_reg  <= w_data_i[3];
      \nz.mem_930_sv2v_reg  <= w_data_i[2];
      \nz.mem_929_sv2v_reg  <= w_data_i[1];
      \nz.mem_928_sv2v_reg  <= w_data_i[0];
    end 
    if(N402) begin
      \nz.mem_927_sv2v_reg  <= w_data_i[31];
      \nz.mem_926_sv2v_reg  <= w_data_i[30];
      \nz.mem_925_sv2v_reg  <= w_data_i[29];
      \nz.mem_924_sv2v_reg  <= w_data_i[28];
      \nz.mem_923_sv2v_reg  <= w_data_i[27];
      \nz.mem_922_sv2v_reg  <= w_data_i[26];
      \nz.mem_921_sv2v_reg  <= w_data_i[25];
      \nz.mem_920_sv2v_reg  <= w_data_i[24];
      \nz.mem_919_sv2v_reg  <= w_data_i[23];
      \nz.mem_918_sv2v_reg  <= w_data_i[22];
      \nz.mem_917_sv2v_reg  <= w_data_i[21];
      \nz.mem_916_sv2v_reg  <= w_data_i[20];
      \nz.mem_915_sv2v_reg  <= w_data_i[19];
      \nz.mem_914_sv2v_reg  <= w_data_i[18];
      \nz.mem_913_sv2v_reg  <= w_data_i[17];
      \nz.mem_912_sv2v_reg  <= w_data_i[16];
      \nz.mem_911_sv2v_reg  <= w_data_i[15];
      \nz.mem_910_sv2v_reg  <= w_data_i[14];
      \nz.mem_909_sv2v_reg  <= w_data_i[13];
      \nz.mem_908_sv2v_reg  <= w_data_i[12];
      \nz.mem_907_sv2v_reg  <= w_data_i[11];
      \nz.mem_906_sv2v_reg  <= w_data_i[10];
      \nz.mem_905_sv2v_reg  <= w_data_i[9];
      \nz.mem_904_sv2v_reg  <= w_data_i[8];
      \nz.mem_903_sv2v_reg  <= w_data_i[7];
      \nz.mem_902_sv2v_reg  <= w_data_i[6];
      \nz.mem_901_sv2v_reg  <= w_data_i[5];
      \nz.mem_900_sv2v_reg  <= w_data_i[4];
      \nz.mem_899_sv2v_reg  <= w_data_i[3];
      \nz.mem_898_sv2v_reg  <= w_data_i[2];
      \nz.mem_897_sv2v_reg  <= w_data_i[1];
      \nz.mem_896_sv2v_reg  <= w_data_i[0];
    end 
    if(N401) begin
      \nz.mem_895_sv2v_reg  <= w_data_i[31];
      \nz.mem_894_sv2v_reg  <= w_data_i[30];
      \nz.mem_893_sv2v_reg  <= w_data_i[29];
      \nz.mem_892_sv2v_reg  <= w_data_i[28];
      \nz.mem_891_sv2v_reg  <= w_data_i[27];
      \nz.mem_890_sv2v_reg  <= w_data_i[26];
      \nz.mem_889_sv2v_reg  <= w_data_i[25];
      \nz.mem_888_sv2v_reg  <= w_data_i[24];
      \nz.mem_887_sv2v_reg  <= w_data_i[23];
      \nz.mem_886_sv2v_reg  <= w_data_i[22];
      \nz.mem_885_sv2v_reg  <= w_data_i[21];
      \nz.mem_884_sv2v_reg  <= w_data_i[20];
      \nz.mem_883_sv2v_reg  <= w_data_i[19];
      \nz.mem_882_sv2v_reg  <= w_data_i[18];
      \nz.mem_881_sv2v_reg  <= w_data_i[17];
      \nz.mem_880_sv2v_reg  <= w_data_i[16];
      \nz.mem_879_sv2v_reg  <= w_data_i[15];
      \nz.mem_878_sv2v_reg  <= w_data_i[14];
      \nz.mem_877_sv2v_reg  <= w_data_i[13];
      \nz.mem_876_sv2v_reg  <= w_data_i[12];
      \nz.mem_875_sv2v_reg  <= w_data_i[11];
      \nz.mem_874_sv2v_reg  <= w_data_i[10];
      \nz.mem_873_sv2v_reg  <= w_data_i[9];
      \nz.mem_872_sv2v_reg  <= w_data_i[8];
      \nz.mem_871_sv2v_reg  <= w_data_i[7];
      \nz.mem_870_sv2v_reg  <= w_data_i[6];
      \nz.mem_869_sv2v_reg  <= w_data_i[5];
      \nz.mem_868_sv2v_reg  <= w_data_i[4];
      \nz.mem_867_sv2v_reg  <= w_data_i[3];
      \nz.mem_866_sv2v_reg  <= w_data_i[2];
      \nz.mem_865_sv2v_reg  <= w_data_i[1];
      \nz.mem_864_sv2v_reg  <= w_data_i[0];
    end 
    if(N400) begin
      \nz.mem_863_sv2v_reg  <= w_data_i[31];
      \nz.mem_862_sv2v_reg  <= w_data_i[30];
      \nz.mem_861_sv2v_reg  <= w_data_i[29];
      \nz.mem_860_sv2v_reg  <= w_data_i[28];
      \nz.mem_859_sv2v_reg  <= w_data_i[27];
      \nz.mem_858_sv2v_reg  <= w_data_i[26];
      \nz.mem_857_sv2v_reg  <= w_data_i[25];
      \nz.mem_856_sv2v_reg  <= w_data_i[24];
      \nz.mem_855_sv2v_reg  <= w_data_i[23];
      \nz.mem_854_sv2v_reg  <= w_data_i[22];
      \nz.mem_853_sv2v_reg  <= w_data_i[21];
      \nz.mem_852_sv2v_reg  <= w_data_i[20];
      \nz.mem_851_sv2v_reg  <= w_data_i[19];
      \nz.mem_850_sv2v_reg  <= w_data_i[18];
      \nz.mem_849_sv2v_reg  <= w_data_i[17];
      \nz.mem_848_sv2v_reg  <= w_data_i[16];
      \nz.mem_847_sv2v_reg  <= w_data_i[15];
      \nz.mem_846_sv2v_reg  <= w_data_i[14];
      \nz.mem_845_sv2v_reg  <= w_data_i[13];
      \nz.mem_844_sv2v_reg  <= w_data_i[12];
      \nz.mem_843_sv2v_reg  <= w_data_i[11];
      \nz.mem_842_sv2v_reg  <= w_data_i[10];
      \nz.mem_841_sv2v_reg  <= w_data_i[9];
      \nz.mem_840_sv2v_reg  <= w_data_i[8];
      \nz.mem_839_sv2v_reg  <= w_data_i[7];
      \nz.mem_838_sv2v_reg  <= w_data_i[6];
      \nz.mem_837_sv2v_reg  <= w_data_i[5];
      \nz.mem_836_sv2v_reg  <= w_data_i[4];
      \nz.mem_835_sv2v_reg  <= w_data_i[3];
      \nz.mem_834_sv2v_reg  <= w_data_i[2];
      \nz.mem_833_sv2v_reg  <= w_data_i[1];
      \nz.mem_832_sv2v_reg  <= w_data_i[0];
    end 
    if(N399) begin
      \nz.mem_831_sv2v_reg  <= w_data_i[31];
      \nz.mem_830_sv2v_reg  <= w_data_i[30];
      \nz.mem_829_sv2v_reg  <= w_data_i[29];
      \nz.mem_828_sv2v_reg  <= w_data_i[28];
      \nz.mem_827_sv2v_reg  <= w_data_i[27];
      \nz.mem_826_sv2v_reg  <= w_data_i[26];
      \nz.mem_825_sv2v_reg  <= w_data_i[25];
      \nz.mem_824_sv2v_reg  <= w_data_i[24];
      \nz.mem_823_sv2v_reg  <= w_data_i[23];
      \nz.mem_822_sv2v_reg  <= w_data_i[22];
      \nz.mem_821_sv2v_reg  <= w_data_i[21];
      \nz.mem_820_sv2v_reg  <= w_data_i[20];
      \nz.mem_819_sv2v_reg  <= w_data_i[19];
      \nz.mem_818_sv2v_reg  <= w_data_i[18];
      \nz.mem_817_sv2v_reg  <= w_data_i[17];
      \nz.mem_816_sv2v_reg  <= w_data_i[16];
      \nz.mem_815_sv2v_reg  <= w_data_i[15];
      \nz.mem_814_sv2v_reg  <= w_data_i[14];
      \nz.mem_813_sv2v_reg  <= w_data_i[13];
      \nz.mem_812_sv2v_reg  <= w_data_i[12];
      \nz.mem_811_sv2v_reg  <= w_data_i[11];
      \nz.mem_810_sv2v_reg  <= w_data_i[10];
      \nz.mem_809_sv2v_reg  <= w_data_i[9];
      \nz.mem_808_sv2v_reg  <= w_data_i[8];
      \nz.mem_807_sv2v_reg  <= w_data_i[7];
      \nz.mem_806_sv2v_reg  <= w_data_i[6];
      \nz.mem_805_sv2v_reg  <= w_data_i[5];
      \nz.mem_804_sv2v_reg  <= w_data_i[4];
      \nz.mem_803_sv2v_reg  <= w_data_i[3];
      \nz.mem_802_sv2v_reg  <= w_data_i[2];
      \nz.mem_801_sv2v_reg  <= w_data_i[1];
      \nz.mem_800_sv2v_reg  <= w_data_i[0];
    end 
    if(N398) begin
      \nz.mem_799_sv2v_reg  <= w_data_i[31];
      \nz.mem_798_sv2v_reg  <= w_data_i[30];
      \nz.mem_797_sv2v_reg  <= w_data_i[29];
      \nz.mem_796_sv2v_reg  <= w_data_i[28];
      \nz.mem_795_sv2v_reg  <= w_data_i[27];
      \nz.mem_794_sv2v_reg  <= w_data_i[26];
      \nz.mem_793_sv2v_reg  <= w_data_i[25];
      \nz.mem_792_sv2v_reg  <= w_data_i[24];
      \nz.mem_791_sv2v_reg  <= w_data_i[23];
      \nz.mem_790_sv2v_reg  <= w_data_i[22];
      \nz.mem_789_sv2v_reg  <= w_data_i[21];
      \nz.mem_788_sv2v_reg  <= w_data_i[20];
      \nz.mem_787_sv2v_reg  <= w_data_i[19];
      \nz.mem_786_sv2v_reg  <= w_data_i[18];
      \nz.mem_785_sv2v_reg  <= w_data_i[17];
      \nz.mem_784_sv2v_reg  <= w_data_i[16];
      \nz.mem_783_sv2v_reg  <= w_data_i[15];
      \nz.mem_782_sv2v_reg  <= w_data_i[14];
      \nz.mem_781_sv2v_reg  <= w_data_i[13];
      \nz.mem_780_sv2v_reg  <= w_data_i[12];
      \nz.mem_779_sv2v_reg  <= w_data_i[11];
      \nz.mem_778_sv2v_reg  <= w_data_i[10];
      \nz.mem_777_sv2v_reg  <= w_data_i[9];
      \nz.mem_776_sv2v_reg  <= w_data_i[8];
      \nz.mem_775_sv2v_reg  <= w_data_i[7];
      \nz.mem_774_sv2v_reg  <= w_data_i[6];
      \nz.mem_773_sv2v_reg  <= w_data_i[5];
      \nz.mem_772_sv2v_reg  <= w_data_i[4];
      \nz.mem_771_sv2v_reg  <= w_data_i[3];
      \nz.mem_770_sv2v_reg  <= w_data_i[2];
      \nz.mem_769_sv2v_reg  <= w_data_i[1];
      \nz.mem_768_sv2v_reg  <= w_data_i[0];
    end 
    if(N397) begin
      \nz.mem_767_sv2v_reg  <= w_data_i[31];
      \nz.mem_766_sv2v_reg  <= w_data_i[30];
      \nz.mem_765_sv2v_reg  <= w_data_i[29];
      \nz.mem_764_sv2v_reg  <= w_data_i[28];
      \nz.mem_763_sv2v_reg  <= w_data_i[27];
      \nz.mem_762_sv2v_reg  <= w_data_i[26];
      \nz.mem_761_sv2v_reg  <= w_data_i[25];
      \nz.mem_760_sv2v_reg  <= w_data_i[24];
      \nz.mem_759_sv2v_reg  <= w_data_i[23];
      \nz.mem_758_sv2v_reg  <= w_data_i[22];
      \nz.mem_757_sv2v_reg  <= w_data_i[21];
      \nz.mem_756_sv2v_reg  <= w_data_i[20];
      \nz.mem_755_sv2v_reg  <= w_data_i[19];
      \nz.mem_754_sv2v_reg  <= w_data_i[18];
      \nz.mem_753_sv2v_reg  <= w_data_i[17];
      \nz.mem_752_sv2v_reg  <= w_data_i[16];
      \nz.mem_751_sv2v_reg  <= w_data_i[15];
      \nz.mem_750_sv2v_reg  <= w_data_i[14];
      \nz.mem_749_sv2v_reg  <= w_data_i[13];
      \nz.mem_748_sv2v_reg  <= w_data_i[12];
      \nz.mem_747_sv2v_reg  <= w_data_i[11];
      \nz.mem_746_sv2v_reg  <= w_data_i[10];
      \nz.mem_745_sv2v_reg  <= w_data_i[9];
      \nz.mem_744_sv2v_reg  <= w_data_i[8];
      \nz.mem_743_sv2v_reg  <= w_data_i[7];
      \nz.mem_742_sv2v_reg  <= w_data_i[6];
      \nz.mem_741_sv2v_reg  <= w_data_i[5];
      \nz.mem_740_sv2v_reg  <= w_data_i[4];
      \nz.mem_739_sv2v_reg  <= w_data_i[3];
      \nz.mem_738_sv2v_reg  <= w_data_i[2];
      \nz.mem_737_sv2v_reg  <= w_data_i[1];
      \nz.mem_736_sv2v_reg  <= w_data_i[0];
    end 
    if(N396) begin
      \nz.mem_735_sv2v_reg  <= w_data_i[31];
      \nz.mem_734_sv2v_reg  <= w_data_i[30];
      \nz.mem_733_sv2v_reg  <= w_data_i[29];
      \nz.mem_732_sv2v_reg  <= w_data_i[28];
      \nz.mem_731_sv2v_reg  <= w_data_i[27];
      \nz.mem_730_sv2v_reg  <= w_data_i[26];
      \nz.mem_729_sv2v_reg  <= w_data_i[25];
      \nz.mem_728_sv2v_reg  <= w_data_i[24];
      \nz.mem_727_sv2v_reg  <= w_data_i[23];
      \nz.mem_726_sv2v_reg  <= w_data_i[22];
      \nz.mem_725_sv2v_reg  <= w_data_i[21];
      \nz.mem_724_sv2v_reg  <= w_data_i[20];
      \nz.mem_723_sv2v_reg  <= w_data_i[19];
      \nz.mem_722_sv2v_reg  <= w_data_i[18];
      \nz.mem_721_sv2v_reg  <= w_data_i[17];
      \nz.mem_720_sv2v_reg  <= w_data_i[16];
      \nz.mem_719_sv2v_reg  <= w_data_i[15];
      \nz.mem_718_sv2v_reg  <= w_data_i[14];
      \nz.mem_717_sv2v_reg  <= w_data_i[13];
      \nz.mem_716_sv2v_reg  <= w_data_i[12];
      \nz.mem_715_sv2v_reg  <= w_data_i[11];
      \nz.mem_714_sv2v_reg  <= w_data_i[10];
      \nz.mem_713_sv2v_reg  <= w_data_i[9];
      \nz.mem_712_sv2v_reg  <= w_data_i[8];
      \nz.mem_711_sv2v_reg  <= w_data_i[7];
      \nz.mem_710_sv2v_reg  <= w_data_i[6];
      \nz.mem_709_sv2v_reg  <= w_data_i[5];
      \nz.mem_708_sv2v_reg  <= w_data_i[4];
      \nz.mem_707_sv2v_reg  <= w_data_i[3];
      \nz.mem_706_sv2v_reg  <= w_data_i[2];
      \nz.mem_705_sv2v_reg  <= w_data_i[1];
      \nz.mem_704_sv2v_reg  <= w_data_i[0];
    end 
    if(N395) begin
      \nz.mem_703_sv2v_reg  <= w_data_i[31];
      \nz.mem_702_sv2v_reg  <= w_data_i[30];
      \nz.mem_701_sv2v_reg  <= w_data_i[29];
      \nz.mem_700_sv2v_reg  <= w_data_i[28];
      \nz.mem_699_sv2v_reg  <= w_data_i[27];
      \nz.mem_698_sv2v_reg  <= w_data_i[26];
      \nz.mem_697_sv2v_reg  <= w_data_i[25];
      \nz.mem_696_sv2v_reg  <= w_data_i[24];
      \nz.mem_695_sv2v_reg  <= w_data_i[23];
      \nz.mem_694_sv2v_reg  <= w_data_i[22];
      \nz.mem_693_sv2v_reg  <= w_data_i[21];
      \nz.mem_692_sv2v_reg  <= w_data_i[20];
      \nz.mem_691_sv2v_reg  <= w_data_i[19];
      \nz.mem_690_sv2v_reg  <= w_data_i[18];
      \nz.mem_689_sv2v_reg  <= w_data_i[17];
      \nz.mem_688_sv2v_reg  <= w_data_i[16];
      \nz.mem_687_sv2v_reg  <= w_data_i[15];
      \nz.mem_686_sv2v_reg  <= w_data_i[14];
      \nz.mem_685_sv2v_reg  <= w_data_i[13];
      \nz.mem_684_sv2v_reg  <= w_data_i[12];
      \nz.mem_683_sv2v_reg  <= w_data_i[11];
      \nz.mem_682_sv2v_reg  <= w_data_i[10];
      \nz.mem_681_sv2v_reg  <= w_data_i[9];
      \nz.mem_680_sv2v_reg  <= w_data_i[8];
      \nz.mem_679_sv2v_reg  <= w_data_i[7];
      \nz.mem_678_sv2v_reg  <= w_data_i[6];
      \nz.mem_677_sv2v_reg  <= w_data_i[5];
      \nz.mem_676_sv2v_reg  <= w_data_i[4];
      \nz.mem_675_sv2v_reg  <= w_data_i[3];
      \nz.mem_674_sv2v_reg  <= w_data_i[2];
      \nz.mem_673_sv2v_reg  <= w_data_i[1];
      \nz.mem_672_sv2v_reg  <= w_data_i[0];
    end 
    if(N394) begin
      \nz.mem_671_sv2v_reg  <= w_data_i[31];
      \nz.mem_670_sv2v_reg  <= w_data_i[30];
      \nz.mem_669_sv2v_reg  <= w_data_i[29];
      \nz.mem_668_sv2v_reg  <= w_data_i[28];
      \nz.mem_667_sv2v_reg  <= w_data_i[27];
      \nz.mem_666_sv2v_reg  <= w_data_i[26];
      \nz.mem_665_sv2v_reg  <= w_data_i[25];
      \nz.mem_664_sv2v_reg  <= w_data_i[24];
      \nz.mem_663_sv2v_reg  <= w_data_i[23];
      \nz.mem_662_sv2v_reg  <= w_data_i[22];
      \nz.mem_661_sv2v_reg  <= w_data_i[21];
      \nz.mem_660_sv2v_reg  <= w_data_i[20];
      \nz.mem_659_sv2v_reg  <= w_data_i[19];
      \nz.mem_658_sv2v_reg  <= w_data_i[18];
      \nz.mem_657_sv2v_reg  <= w_data_i[17];
      \nz.mem_656_sv2v_reg  <= w_data_i[16];
      \nz.mem_655_sv2v_reg  <= w_data_i[15];
      \nz.mem_654_sv2v_reg  <= w_data_i[14];
      \nz.mem_653_sv2v_reg  <= w_data_i[13];
      \nz.mem_652_sv2v_reg  <= w_data_i[12];
      \nz.mem_651_sv2v_reg  <= w_data_i[11];
      \nz.mem_650_sv2v_reg  <= w_data_i[10];
      \nz.mem_649_sv2v_reg  <= w_data_i[9];
      \nz.mem_648_sv2v_reg  <= w_data_i[8];
      \nz.mem_647_sv2v_reg  <= w_data_i[7];
      \nz.mem_646_sv2v_reg  <= w_data_i[6];
      \nz.mem_645_sv2v_reg  <= w_data_i[5];
      \nz.mem_644_sv2v_reg  <= w_data_i[4];
      \nz.mem_643_sv2v_reg  <= w_data_i[3];
      \nz.mem_642_sv2v_reg  <= w_data_i[2];
      \nz.mem_641_sv2v_reg  <= w_data_i[1];
      \nz.mem_640_sv2v_reg  <= w_data_i[0];
    end 
    if(N393) begin
      \nz.mem_639_sv2v_reg  <= w_data_i[31];
      \nz.mem_638_sv2v_reg  <= w_data_i[30];
      \nz.mem_637_sv2v_reg  <= w_data_i[29];
      \nz.mem_636_sv2v_reg  <= w_data_i[28];
      \nz.mem_635_sv2v_reg  <= w_data_i[27];
      \nz.mem_634_sv2v_reg  <= w_data_i[26];
      \nz.mem_633_sv2v_reg  <= w_data_i[25];
      \nz.mem_632_sv2v_reg  <= w_data_i[24];
      \nz.mem_631_sv2v_reg  <= w_data_i[23];
      \nz.mem_630_sv2v_reg  <= w_data_i[22];
      \nz.mem_629_sv2v_reg  <= w_data_i[21];
      \nz.mem_628_sv2v_reg  <= w_data_i[20];
      \nz.mem_627_sv2v_reg  <= w_data_i[19];
      \nz.mem_626_sv2v_reg  <= w_data_i[18];
      \nz.mem_625_sv2v_reg  <= w_data_i[17];
      \nz.mem_624_sv2v_reg  <= w_data_i[16];
      \nz.mem_623_sv2v_reg  <= w_data_i[15];
      \nz.mem_622_sv2v_reg  <= w_data_i[14];
      \nz.mem_621_sv2v_reg  <= w_data_i[13];
      \nz.mem_620_sv2v_reg  <= w_data_i[12];
      \nz.mem_619_sv2v_reg  <= w_data_i[11];
      \nz.mem_618_sv2v_reg  <= w_data_i[10];
      \nz.mem_617_sv2v_reg  <= w_data_i[9];
      \nz.mem_616_sv2v_reg  <= w_data_i[8];
      \nz.mem_615_sv2v_reg  <= w_data_i[7];
      \nz.mem_614_sv2v_reg  <= w_data_i[6];
      \nz.mem_613_sv2v_reg  <= w_data_i[5];
      \nz.mem_612_sv2v_reg  <= w_data_i[4];
      \nz.mem_611_sv2v_reg  <= w_data_i[3];
      \nz.mem_610_sv2v_reg  <= w_data_i[2];
      \nz.mem_609_sv2v_reg  <= w_data_i[1];
      \nz.mem_608_sv2v_reg  <= w_data_i[0];
    end 
    if(N392) begin
      \nz.mem_607_sv2v_reg  <= w_data_i[31];
      \nz.mem_606_sv2v_reg  <= w_data_i[30];
      \nz.mem_605_sv2v_reg  <= w_data_i[29];
      \nz.mem_604_sv2v_reg  <= w_data_i[28];
      \nz.mem_603_sv2v_reg  <= w_data_i[27];
      \nz.mem_602_sv2v_reg  <= w_data_i[26];
      \nz.mem_601_sv2v_reg  <= w_data_i[25];
      \nz.mem_600_sv2v_reg  <= w_data_i[24];
      \nz.mem_599_sv2v_reg  <= w_data_i[23];
      \nz.mem_598_sv2v_reg  <= w_data_i[22];
      \nz.mem_597_sv2v_reg  <= w_data_i[21];
      \nz.mem_596_sv2v_reg  <= w_data_i[20];
      \nz.mem_595_sv2v_reg  <= w_data_i[19];
      \nz.mem_594_sv2v_reg  <= w_data_i[18];
      \nz.mem_593_sv2v_reg  <= w_data_i[17];
      \nz.mem_592_sv2v_reg  <= w_data_i[16];
      \nz.mem_591_sv2v_reg  <= w_data_i[15];
      \nz.mem_590_sv2v_reg  <= w_data_i[14];
      \nz.mem_589_sv2v_reg  <= w_data_i[13];
      \nz.mem_588_sv2v_reg  <= w_data_i[12];
      \nz.mem_587_sv2v_reg  <= w_data_i[11];
      \nz.mem_586_sv2v_reg  <= w_data_i[10];
      \nz.mem_585_sv2v_reg  <= w_data_i[9];
      \nz.mem_584_sv2v_reg  <= w_data_i[8];
      \nz.mem_583_sv2v_reg  <= w_data_i[7];
      \nz.mem_582_sv2v_reg  <= w_data_i[6];
      \nz.mem_581_sv2v_reg  <= w_data_i[5];
      \nz.mem_580_sv2v_reg  <= w_data_i[4];
      \nz.mem_579_sv2v_reg  <= w_data_i[3];
      \nz.mem_578_sv2v_reg  <= w_data_i[2];
      \nz.mem_577_sv2v_reg  <= w_data_i[1];
      \nz.mem_576_sv2v_reg  <= w_data_i[0];
    end 
    if(N391) begin
      \nz.mem_575_sv2v_reg  <= w_data_i[31];
      \nz.mem_574_sv2v_reg  <= w_data_i[30];
      \nz.mem_573_sv2v_reg  <= w_data_i[29];
      \nz.mem_572_sv2v_reg  <= w_data_i[28];
      \nz.mem_571_sv2v_reg  <= w_data_i[27];
      \nz.mem_570_sv2v_reg  <= w_data_i[26];
      \nz.mem_569_sv2v_reg  <= w_data_i[25];
      \nz.mem_568_sv2v_reg  <= w_data_i[24];
      \nz.mem_567_sv2v_reg  <= w_data_i[23];
      \nz.mem_566_sv2v_reg  <= w_data_i[22];
      \nz.mem_565_sv2v_reg  <= w_data_i[21];
      \nz.mem_564_sv2v_reg  <= w_data_i[20];
      \nz.mem_563_sv2v_reg  <= w_data_i[19];
      \nz.mem_562_sv2v_reg  <= w_data_i[18];
      \nz.mem_561_sv2v_reg  <= w_data_i[17];
      \nz.mem_560_sv2v_reg  <= w_data_i[16];
      \nz.mem_559_sv2v_reg  <= w_data_i[15];
      \nz.mem_558_sv2v_reg  <= w_data_i[14];
      \nz.mem_557_sv2v_reg  <= w_data_i[13];
      \nz.mem_556_sv2v_reg  <= w_data_i[12];
      \nz.mem_555_sv2v_reg  <= w_data_i[11];
      \nz.mem_554_sv2v_reg  <= w_data_i[10];
      \nz.mem_553_sv2v_reg  <= w_data_i[9];
      \nz.mem_552_sv2v_reg  <= w_data_i[8];
      \nz.mem_551_sv2v_reg  <= w_data_i[7];
      \nz.mem_550_sv2v_reg  <= w_data_i[6];
      \nz.mem_549_sv2v_reg  <= w_data_i[5];
      \nz.mem_548_sv2v_reg  <= w_data_i[4];
      \nz.mem_547_sv2v_reg  <= w_data_i[3];
      \nz.mem_546_sv2v_reg  <= w_data_i[2];
      \nz.mem_545_sv2v_reg  <= w_data_i[1];
      \nz.mem_544_sv2v_reg  <= w_data_i[0];
    end 
    if(N390) begin
      \nz.mem_543_sv2v_reg  <= w_data_i[31];
      \nz.mem_542_sv2v_reg  <= w_data_i[30];
      \nz.mem_541_sv2v_reg  <= w_data_i[29];
      \nz.mem_540_sv2v_reg  <= w_data_i[28];
      \nz.mem_539_sv2v_reg  <= w_data_i[27];
      \nz.mem_538_sv2v_reg  <= w_data_i[26];
      \nz.mem_537_sv2v_reg  <= w_data_i[25];
      \nz.mem_536_sv2v_reg  <= w_data_i[24];
      \nz.mem_535_sv2v_reg  <= w_data_i[23];
      \nz.mem_534_sv2v_reg  <= w_data_i[22];
      \nz.mem_533_sv2v_reg  <= w_data_i[21];
      \nz.mem_532_sv2v_reg  <= w_data_i[20];
      \nz.mem_531_sv2v_reg  <= w_data_i[19];
      \nz.mem_530_sv2v_reg  <= w_data_i[18];
      \nz.mem_529_sv2v_reg  <= w_data_i[17];
      \nz.mem_528_sv2v_reg  <= w_data_i[16];
      \nz.mem_527_sv2v_reg  <= w_data_i[15];
      \nz.mem_526_sv2v_reg  <= w_data_i[14];
      \nz.mem_525_sv2v_reg  <= w_data_i[13];
      \nz.mem_524_sv2v_reg  <= w_data_i[12];
      \nz.mem_523_sv2v_reg  <= w_data_i[11];
      \nz.mem_522_sv2v_reg  <= w_data_i[10];
      \nz.mem_521_sv2v_reg  <= w_data_i[9];
      \nz.mem_520_sv2v_reg  <= w_data_i[8];
      \nz.mem_519_sv2v_reg  <= w_data_i[7];
      \nz.mem_518_sv2v_reg  <= w_data_i[6];
      \nz.mem_517_sv2v_reg  <= w_data_i[5];
      \nz.mem_516_sv2v_reg  <= w_data_i[4];
      \nz.mem_515_sv2v_reg  <= w_data_i[3];
      \nz.mem_514_sv2v_reg  <= w_data_i[2];
      \nz.mem_513_sv2v_reg  <= w_data_i[1];
      \nz.mem_512_sv2v_reg  <= w_data_i[0];
    end 
    if(N389) begin
      \nz.mem_511_sv2v_reg  <= w_data_i[31];
      \nz.mem_510_sv2v_reg  <= w_data_i[30];
      \nz.mem_509_sv2v_reg  <= w_data_i[29];
      \nz.mem_508_sv2v_reg  <= w_data_i[28];
      \nz.mem_507_sv2v_reg  <= w_data_i[27];
      \nz.mem_506_sv2v_reg  <= w_data_i[26];
      \nz.mem_505_sv2v_reg  <= w_data_i[25];
      \nz.mem_504_sv2v_reg  <= w_data_i[24];
      \nz.mem_503_sv2v_reg  <= w_data_i[23];
      \nz.mem_502_sv2v_reg  <= w_data_i[22];
      \nz.mem_501_sv2v_reg  <= w_data_i[21];
      \nz.mem_500_sv2v_reg  <= w_data_i[20];
      \nz.mem_499_sv2v_reg  <= w_data_i[19];
      \nz.mem_498_sv2v_reg  <= w_data_i[18];
      \nz.mem_497_sv2v_reg  <= w_data_i[17];
      \nz.mem_496_sv2v_reg  <= w_data_i[16];
      \nz.mem_495_sv2v_reg  <= w_data_i[15];
      \nz.mem_494_sv2v_reg  <= w_data_i[14];
      \nz.mem_493_sv2v_reg  <= w_data_i[13];
      \nz.mem_492_sv2v_reg  <= w_data_i[12];
      \nz.mem_491_sv2v_reg  <= w_data_i[11];
      \nz.mem_490_sv2v_reg  <= w_data_i[10];
      \nz.mem_489_sv2v_reg  <= w_data_i[9];
      \nz.mem_488_sv2v_reg  <= w_data_i[8];
      \nz.mem_487_sv2v_reg  <= w_data_i[7];
      \nz.mem_486_sv2v_reg  <= w_data_i[6];
      \nz.mem_485_sv2v_reg  <= w_data_i[5];
      \nz.mem_484_sv2v_reg  <= w_data_i[4];
      \nz.mem_483_sv2v_reg  <= w_data_i[3];
      \nz.mem_482_sv2v_reg  <= w_data_i[2];
      \nz.mem_481_sv2v_reg  <= w_data_i[1];
      \nz.mem_480_sv2v_reg  <= w_data_i[0];
    end 
    if(N388) begin
      \nz.mem_479_sv2v_reg  <= w_data_i[31];
      \nz.mem_478_sv2v_reg  <= w_data_i[30];
      \nz.mem_477_sv2v_reg  <= w_data_i[29];
      \nz.mem_476_sv2v_reg  <= w_data_i[28];
      \nz.mem_475_sv2v_reg  <= w_data_i[27];
      \nz.mem_474_sv2v_reg  <= w_data_i[26];
      \nz.mem_473_sv2v_reg  <= w_data_i[25];
      \nz.mem_472_sv2v_reg  <= w_data_i[24];
      \nz.mem_471_sv2v_reg  <= w_data_i[23];
      \nz.mem_470_sv2v_reg  <= w_data_i[22];
      \nz.mem_469_sv2v_reg  <= w_data_i[21];
      \nz.mem_468_sv2v_reg  <= w_data_i[20];
      \nz.mem_467_sv2v_reg  <= w_data_i[19];
      \nz.mem_466_sv2v_reg  <= w_data_i[18];
      \nz.mem_465_sv2v_reg  <= w_data_i[17];
      \nz.mem_464_sv2v_reg  <= w_data_i[16];
      \nz.mem_463_sv2v_reg  <= w_data_i[15];
      \nz.mem_462_sv2v_reg  <= w_data_i[14];
      \nz.mem_461_sv2v_reg  <= w_data_i[13];
      \nz.mem_460_sv2v_reg  <= w_data_i[12];
      \nz.mem_459_sv2v_reg  <= w_data_i[11];
      \nz.mem_458_sv2v_reg  <= w_data_i[10];
      \nz.mem_457_sv2v_reg  <= w_data_i[9];
      \nz.mem_456_sv2v_reg  <= w_data_i[8];
      \nz.mem_455_sv2v_reg  <= w_data_i[7];
      \nz.mem_454_sv2v_reg  <= w_data_i[6];
      \nz.mem_453_sv2v_reg  <= w_data_i[5];
      \nz.mem_452_sv2v_reg  <= w_data_i[4];
      \nz.mem_451_sv2v_reg  <= w_data_i[3];
      \nz.mem_450_sv2v_reg  <= w_data_i[2];
      \nz.mem_449_sv2v_reg  <= w_data_i[1];
      \nz.mem_448_sv2v_reg  <= w_data_i[0];
    end 
    if(N387) begin
      \nz.mem_447_sv2v_reg  <= w_data_i[31];
      \nz.mem_446_sv2v_reg  <= w_data_i[30];
      \nz.mem_445_sv2v_reg  <= w_data_i[29];
      \nz.mem_444_sv2v_reg  <= w_data_i[28];
      \nz.mem_443_sv2v_reg  <= w_data_i[27];
      \nz.mem_442_sv2v_reg  <= w_data_i[26];
      \nz.mem_441_sv2v_reg  <= w_data_i[25];
      \nz.mem_440_sv2v_reg  <= w_data_i[24];
      \nz.mem_439_sv2v_reg  <= w_data_i[23];
      \nz.mem_438_sv2v_reg  <= w_data_i[22];
      \nz.mem_437_sv2v_reg  <= w_data_i[21];
      \nz.mem_436_sv2v_reg  <= w_data_i[20];
      \nz.mem_435_sv2v_reg  <= w_data_i[19];
      \nz.mem_434_sv2v_reg  <= w_data_i[18];
      \nz.mem_433_sv2v_reg  <= w_data_i[17];
      \nz.mem_432_sv2v_reg  <= w_data_i[16];
      \nz.mem_431_sv2v_reg  <= w_data_i[15];
      \nz.mem_430_sv2v_reg  <= w_data_i[14];
      \nz.mem_429_sv2v_reg  <= w_data_i[13];
      \nz.mem_428_sv2v_reg  <= w_data_i[12];
      \nz.mem_427_sv2v_reg  <= w_data_i[11];
      \nz.mem_426_sv2v_reg  <= w_data_i[10];
      \nz.mem_425_sv2v_reg  <= w_data_i[9];
      \nz.mem_424_sv2v_reg  <= w_data_i[8];
      \nz.mem_423_sv2v_reg  <= w_data_i[7];
      \nz.mem_422_sv2v_reg  <= w_data_i[6];
      \nz.mem_421_sv2v_reg  <= w_data_i[5];
      \nz.mem_420_sv2v_reg  <= w_data_i[4];
      \nz.mem_419_sv2v_reg  <= w_data_i[3];
      \nz.mem_418_sv2v_reg  <= w_data_i[2];
      \nz.mem_417_sv2v_reg  <= w_data_i[1];
      \nz.mem_416_sv2v_reg  <= w_data_i[0];
    end 
    if(N386) begin
      \nz.mem_415_sv2v_reg  <= w_data_i[31];
      \nz.mem_414_sv2v_reg  <= w_data_i[30];
      \nz.mem_413_sv2v_reg  <= w_data_i[29];
      \nz.mem_412_sv2v_reg  <= w_data_i[28];
      \nz.mem_411_sv2v_reg  <= w_data_i[27];
      \nz.mem_410_sv2v_reg  <= w_data_i[26];
      \nz.mem_409_sv2v_reg  <= w_data_i[25];
      \nz.mem_408_sv2v_reg  <= w_data_i[24];
      \nz.mem_407_sv2v_reg  <= w_data_i[23];
      \nz.mem_406_sv2v_reg  <= w_data_i[22];
      \nz.mem_405_sv2v_reg  <= w_data_i[21];
      \nz.mem_404_sv2v_reg  <= w_data_i[20];
      \nz.mem_403_sv2v_reg  <= w_data_i[19];
      \nz.mem_402_sv2v_reg  <= w_data_i[18];
      \nz.mem_401_sv2v_reg  <= w_data_i[17];
      \nz.mem_400_sv2v_reg  <= w_data_i[16];
      \nz.mem_399_sv2v_reg  <= w_data_i[15];
      \nz.mem_398_sv2v_reg  <= w_data_i[14];
      \nz.mem_397_sv2v_reg  <= w_data_i[13];
      \nz.mem_396_sv2v_reg  <= w_data_i[12];
      \nz.mem_395_sv2v_reg  <= w_data_i[11];
      \nz.mem_394_sv2v_reg  <= w_data_i[10];
      \nz.mem_393_sv2v_reg  <= w_data_i[9];
      \nz.mem_392_sv2v_reg  <= w_data_i[8];
      \nz.mem_391_sv2v_reg  <= w_data_i[7];
      \nz.mem_390_sv2v_reg  <= w_data_i[6];
      \nz.mem_389_sv2v_reg  <= w_data_i[5];
      \nz.mem_388_sv2v_reg  <= w_data_i[4];
      \nz.mem_387_sv2v_reg  <= w_data_i[3];
      \nz.mem_386_sv2v_reg  <= w_data_i[2];
      \nz.mem_385_sv2v_reg  <= w_data_i[1];
      \nz.mem_384_sv2v_reg  <= w_data_i[0];
    end 
    if(N385) begin
      \nz.mem_383_sv2v_reg  <= w_data_i[31];
      \nz.mem_382_sv2v_reg  <= w_data_i[30];
      \nz.mem_381_sv2v_reg  <= w_data_i[29];
      \nz.mem_380_sv2v_reg  <= w_data_i[28];
      \nz.mem_379_sv2v_reg  <= w_data_i[27];
      \nz.mem_378_sv2v_reg  <= w_data_i[26];
      \nz.mem_377_sv2v_reg  <= w_data_i[25];
      \nz.mem_376_sv2v_reg  <= w_data_i[24];
      \nz.mem_375_sv2v_reg  <= w_data_i[23];
      \nz.mem_374_sv2v_reg  <= w_data_i[22];
      \nz.mem_373_sv2v_reg  <= w_data_i[21];
      \nz.mem_372_sv2v_reg  <= w_data_i[20];
      \nz.mem_371_sv2v_reg  <= w_data_i[19];
      \nz.mem_370_sv2v_reg  <= w_data_i[18];
      \nz.mem_369_sv2v_reg  <= w_data_i[17];
      \nz.mem_368_sv2v_reg  <= w_data_i[16];
      \nz.mem_367_sv2v_reg  <= w_data_i[15];
      \nz.mem_366_sv2v_reg  <= w_data_i[14];
      \nz.mem_365_sv2v_reg  <= w_data_i[13];
      \nz.mem_364_sv2v_reg  <= w_data_i[12];
      \nz.mem_363_sv2v_reg  <= w_data_i[11];
      \nz.mem_362_sv2v_reg  <= w_data_i[10];
      \nz.mem_361_sv2v_reg  <= w_data_i[9];
      \nz.mem_360_sv2v_reg  <= w_data_i[8];
      \nz.mem_359_sv2v_reg  <= w_data_i[7];
      \nz.mem_358_sv2v_reg  <= w_data_i[6];
      \nz.mem_357_sv2v_reg  <= w_data_i[5];
      \nz.mem_356_sv2v_reg  <= w_data_i[4];
      \nz.mem_355_sv2v_reg  <= w_data_i[3];
      \nz.mem_354_sv2v_reg  <= w_data_i[2];
      \nz.mem_353_sv2v_reg  <= w_data_i[1];
      \nz.mem_352_sv2v_reg  <= w_data_i[0];
    end 
    if(N384) begin
      \nz.mem_351_sv2v_reg  <= w_data_i[31];
      \nz.mem_350_sv2v_reg  <= w_data_i[30];
      \nz.mem_349_sv2v_reg  <= w_data_i[29];
      \nz.mem_348_sv2v_reg  <= w_data_i[28];
      \nz.mem_347_sv2v_reg  <= w_data_i[27];
      \nz.mem_346_sv2v_reg  <= w_data_i[26];
      \nz.mem_345_sv2v_reg  <= w_data_i[25];
      \nz.mem_344_sv2v_reg  <= w_data_i[24];
      \nz.mem_343_sv2v_reg  <= w_data_i[23];
      \nz.mem_342_sv2v_reg  <= w_data_i[22];
      \nz.mem_341_sv2v_reg  <= w_data_i[21];
      \nz.mem_340_sv2v_reg  <= w_data_i[20];
      \nz.mem_339_sv2v_reg  <= w_data_i[19];
      \nz.mem_338_sv2v_reg  <= w_data_i[18];
      \nz.mem_337_sv2v_reg  <= w_data_i[17];
      \nz.mem_336_sv2v_reg  <= w_data_i[16];
      \nz.mem_335_sv2v_reg  <= w_data_i[15];
      \nz.mem_334_sv2v_reg  <= w_data_i[14];
      \nz.mem_333_sv2v_reg  <= w_data_i[13];
      \nz.mem_332_sv2v_reg  <= w_data_i[12];
      \nz.mem_331_sv2v_reg  <= w_data_i[11];
      \nz.mem_330_sv2v_reg  <= w_data_i[10];
      \nz.mem_329_sv2v_reg  <= w_data_i[9];
      \nz.mem_328_sv2v_reg  <= w_data_i[8];
      \nz.mem_327_sv2v_reg  <= w_data_i[7];
      \nz.mem_326_sv2v_reg  <= w_data_i[6];
      \nz.mem_325_sv2v_reg  <= w_data_i[5];
      \nz.mem_324_sv2v_reg  <= w_data_i[4];
      \nz.mem_323_sv2v_reg  <= w_data_i[3];
      \nz.mem_322_sv2v_reg  <= w_data_i[2];
      \nz.mem_321_sv2v_reg  <= w_data_i[1];
      \nz.mem_320_sv2v_reg  <= w_data_i[0];
    end 
    if(N383) begin
      \nz.mem_319_sv2v_reg  <= w_data_i[31];
      \nz.mem_318_sv2v_reg  <= w_data_i[30];
      \nz.mem_317_sv2v_reg  <= w_data_i[29];
      \nz.mem_316_sv2v_reg  <= w_data_i[28];
      \nz.mem_315_sv2v_reg  <= w_data_i[27];
      \nz.mem_314_sv2v_reg  <= w_data_i[26];
      \nz.mem_313_sv2v_reg  <= w_data_i[25];
      \nz.mem_312_sv2v_reg  <= w_data_i[24];
      \nz.mem_311_sv2v_reg  <= w_data_i[23];
      \nz.mem_310_sv2v_reg  <= w_data_i[22];
      \nz.mem_309_sv2v_reg  <= w_data_i[21];
      \nz.mem_308_sv2v_reg  <= w_data_i[20];
      \nz.mem_307_sv2v_reg  <= w_data_i[19];
      \nz.mem_306_sv2v_reg  <= w_data_i[18];
      \nz.mem_305_sv2v_reg  <= w_data_i[17];
      \nz.mem_304_sv2v_reg  <= w_data_i[16];
      \nz.mem_303_sv2v_reg  <= w_data_i[15];
      \nz.mem_302_sv2v_reg  <= w_data_i[14];
      \nz.mem_301_sv2v_reg  <= w_data_i[13];
      \nz.mem_300_sv2v_reg  <= w_data_i[12];
      \nz.mem_299_sv2v_reg  <= w_data_i[11];
      \nz.mem_298_sv2v_reg  <= w_data_i[10];
      \nz.mem_297_sv2v_reg  <= w_data_i[9];
      \nz.mem_296_sv2v_reg  <= w_data_i[8];
      \nz.mem_295_sv2v_reg  <= w_data_i[7];
      \nz.mem_294_sv2v_reg  <= w_data_i[6];
      \nz.mem_293_sv2v_reg  <= w_data_i[5];
      \nz.mem_292_sv2v_reg  <= w_data_i[4];
      \nz.mem_291_sv2v_reg  <= w_data_i[3];
      \nz.mem_290_sv2v_reg  <= w_data_i[2];
      \nz.mem_289_sv2v_reg  <= w_data_i[1];
      \nz.mem_288_sv2v_reg  <= w_data_i[0];
    end 
    if(N382) begin
      \nz.mem_287_sv2v_reg  <= w_data_i[31];
      \nz.mem_286_sv2v_reg  <= w_data_i[30];
      \nz.mem_285_sv2v_reg  <= w_data_i[29];
      \nz.mem_284_sv2v_reg  <= w_data_i[28];
      \nz.mem_283_sv2v_reg  <= w_data_i[27];
      \nz.mem_282_sv2v_reg  <= w_data_i[26];
      \nz.mem_281_sv2v_reg  <= w_data_i[25];
      \nz.mem_280_sv2v_reg  <= w_data_i[24];
      \nz.mem_279_sv2v_reg  <= w_data_i[23];
      \nz.mem_278_sv2v_reg  <= w_data_i[22];
      \nz.mem_277_sv2v_reg  <= w_data_i[21];
      \nz.mem_276_sv2v_reg  <= w_data_i[20];
      \nz.mem_275_sv2v_reg  <= w_data_i[19];
      \nz.mem_274_sv2v_reg  <= w_data_i[18];
      \nz.mem_273_sv2v_reg  <= w_data_i[17];
      \nz.mem_272_sv2v_reg  <= w_data_i[16];
      \nz.mem_271_sv2v_reg  <= w_data_i[15];
      \nz.mem_270_sv2v_reg  <= w_data_i[14];
      \nz.mem_269_sv2v_reg  <= w_data_i[13];
      \nz.mem_268_sv2v_reg  <= w_data_i[12];
      \nz.mem_267_sv2v_reg  <= w_data_i[11];
      \nz.mem_266_sv2v_reg  <= w_data_i[10];
      \nz.mem_265_sv2v_reg  <= w_data_i[9];
      \nz.mem_264_sv2v_reg  <= w_data_i[8];
      \nz.mem_263_sv2v_reg  <= w_data_i[7];
      \nz.mem_262_sv2v_reg  <= w_data_i[6];
      \nz.mem_261_sv2v_reg  <= w_data_i[5];
      \nz.mem_260_sv2v_reg  <= w_data_i[4];
      \nz.mem_259_sv2v_reg  <= w_data_i[3];
      \nz.mem_258_sv2v_reg  <= w_data_i[2];
      \nz.mem_257_sv2v_reg  <= w_data_i[1];
      \nz.mem_256_sv2v_reg  <= w_data_i[0];
    end 
    if(N381) begin
      \nz.mem_255_sv2v_reg  <= w_data_i[31];
      \nz.mem_254_sv2v_reg  <= w_data_i[30];
      \nz.mem_253_sv2v_reg  <= w_data_i[29];
      \nz.mem_252_sv2v_reg  <= w_data_i[28];
      \nz.mem_251_sv2v_reg  <= w_data_i[27];
      \nz.mem_250_sv2v_reg  <= w_data_i[26];
      \nz.mem_249_sv2v_reg  <= w_data_i[25];
      \nz.mem_248_sv2v_reg  <= w_data_i[24];
      \nz.mem_247_sv2v_reg  <= w_data_i[23];
      \nz.mem_246_sv2v_reg  <= w_data_i[22];
      \nz.mem_245_sv2v_reg  <= w_data_i[21];
      \nz.mem_244_sv2v_reg  <= w_data_i[20];
      \nz.mem_243_sv2v_reg  <= w_data_i[19];
      \nz.mem_242_sv2v_reg  <= w_data_i[18];
      \nz.mem_241_sv2v_reg  <= w_data_i[17];
      \nz.mem_240_sv2v_reg  <= w_data_i[16];
      \nz.mem_239_sv2v_reg  <= w_data_i[15];
      \nz.mem_238_sv2v_reg  <= w_data_i[14];
      \nz.mem_237_sv2v_reg  <= w_data_i[13];
      \nz.mem_236_sv2v_reg  <= w_data_i[12];
      \nz.mem_235_sv2v_reg  <= w_data_i[11];
      \nz.mem_234_sv2v_reg  <= w_data_i[10];
      \nz.mem_233_sv2v_reg  <= w_data_i[9];
      \nz.mem_232_sv2v_reg  <= w_data_i[8];
      \nz.mem_231_sv2v_reg  <= w_data_i[7];
      \nz.mem_230_sv2v_reg  <= w_data_i[6];
      \nz.mem_229_sv2v_reg  <= w_data_i[5];
      \nz.mem_228_sv2v_reg  <= w_data_i[4];
      \nz.mem_227_sv2v_reg  <= w_data_i[3];
      \nz.mem_226_sv2v_reg  <= w_data_i[2];
      \nz.mem_225_sv2v_reg  <= w_data_i[1];
      \nz.mem_224_sv2v_reg  <= w_data_i[0];
    end 
    if(N380) begin
      \nz.mem_223_sv2v_reg  <= w_data_i[31];
      \nz.mem_222_sv2v_reg  <= w_data_i[30];
      \nz.mem_221_sv2v_reg  <= w_data_i[29];
      \nz.mem_220_sv2v_reg  <= w_data_i[28];
      \nz.mem_219_sv2v_reg  <= w_data_i[27];
      \nz.mem_218_sv2v_reg  <= w_data_i[26];
      \nz.mem_217_sv2v_reg  <= w_data_i[25];
      \nz.mem_216_sv2v_reg  <= w_data_i[24];
      \nz.mem_215_sv2v_reg  <= w_data_i[23];
      \nz.mem_214_sv2v_reg  <= w_data_i[22];
      \nz.mem_213_sv2v_reg  <= w_data_i[21];
      \nz.mem_212_sv2v_reg  <= w_data_i[20];
      \nz.mem_211_sv2v_reg  <= w_data_i[19];
      \nz.mem_210_sv2v_reg  <= w_data_i[18];
      \nz.mem_209_sv2v_reg  <= w_data_i[17];
      \nz.mem_208_sv2v_reg  <= w_data_i[16];
      \nz.mem_207_sv2v_reg  <= w_data_i[15];
      \nz.mem_206_sv2v_reg  <= w_data_i[14];
      \nz.mem_205_sv2v_reg  <= w_data_i[13];
      \nz.mem_204_sv2v_reg  <= w_data_i[12];
      \nz.mem_203_sv2v_reg  <= w_data_i[11];
      \nz.mem_202_sv2v_reg  <= w_data_i[10];
      \nz.mem_201_sv2v_reg  <= w_data_i[9];
      \nz.mem_200_sv2v_reg  <= w_data_i[8];
      \nz.mem_199_sv2v_reg  <= w_data_i[7];
      \nz.mem_198_sv2v_reg  <= w_data_i[6];
      \nz.mem_197_sv2v_reg  <= w_data_i[5];
      \nz.mem_196_sv2v_reg  <= w_data_i[4];
      \nz.mem_195_sv2v_reg  <= w_data_i[3];
      \nz.mem_194_sv2v_reg  <= w_data_i[2];
      \nz.mem_193_sv2v_reg  <= w_data_i[1];
      \nz.mem_192_sv2v_reg  <= w_data_i[0];
    end 
    if(N379) begin
      \nz.mem_191_sv2v_reg  <= w_data_i[31];
      \nz.mem_190_sv2v_reg  <= w_data_i[30];
      \nz.mem_189_sv2v_reg  <= w_data_i[29];
      \nz.mem_188_sv2v_reg  <= w_data_i[28];
      \nz.mem_187_sv2v_reg  <= w_data_i[27];
      \nz.mem_186_sv2v_reg  <= w_data_i[26];
      \nz.mem_185_sv2v_reg  <= w_data_i[25];
      \nz.mem_184_sv2v_reg  <= w_data_i[24];
      \nz.mem_183_sv2v_reg  <= w_data_i[23];
      \nz.mem_182_sv2v_reg  <= w_data_i[22];
      \nz.mem_181_sv2v_reg  <= w_data_i[21];
      \nz.mem_180_sv2v_reg  <= w_data_i[20];
      \nz.mem_179_sv2v_reg  <= w_data_i[19];
      \nz.mem_178_sv2v_reg  <= w_data_i[18];
      \nz.mem_177_sv2v_reg  <= w_data_i[17];
      \nz.mem_176_sv2v_reg  <= w_data_i[16];
      \nz.mem_175_sv2v_reg  <= w_data_i[15];
      \nz.mem_174_sv2v_reg  <= w_data_i[14];
      \nz.mem_173_sv2v_reg  <= w_data_i[13];
      \nz.mem_172_sv2v_reg  <= w_data_i[12];
      \nz.mem_171_sv2v_reg  <= w_data_i[11];
      \nz.mem_170_sv2v_reg  <= w_data_i[10];
      \nz.mem_169_sv2v_reg  <= w_data_i[9];
      \nz.mem_168_sv2v_reg  <= w_data_i[8];
      \nz.mem_167_sv2v_reg  <= w_data_i[7];
      \nz.mem_166_sv2v_reg  <= w_data_i[6];
      \nz.mem_165_sv2v_reg  <= w_data_i[5];
      \nz.mem_164_sv2v_reg  <= w_data_i[4];
      \nz.mem_163_sv2v_reg  <= w_data_i[3];
      \nz.mem_162_sv2v_reg  <= w_data_i[2];
      \nz.mem_161_sv2v_reg  <= w_data_i[1];
      \nz.mem_160_sv2v_reg  <= w_data_i[0];
    end 
    if(N378) begin
      \nz.mem_159_sv2v_reg  <= w_data_i[31];
      \nz.mem_158_sv2v_reg  <= w_data_i[30];
      \nz.mem_157_sv2v_reg  <= w_data_i[29];
      \nz.mem_156_sv2v_reg  <= w_data_i[28];
      \nz.mem_155_sv2v_reg  <= w_data_i[27];
      \nz.mem_154_sv2v_reg  <= w_data_i[26];
      \nz.mem_153_sv2v_reg  <= w_data_i[25];
      \nz.mem_152_sv2v_reg  <= w_data_i[24];
      \nz.mem_151_sv2v_reg  <= w_data_i[23];
      \nz.mem_150_sv2v_reg  <= w_data_i[22];
      \nz.mem_149_sv2v_reg  <= w_data_i[21];
      \nz.mem_148_sv2v_reg  <= w_data_i[20];
      \nz.mem_147_sv2v_reg  <= w_data_i[19];
      \nz.mem_146_sv2v_reg  <= w_data_i[18];
      \nz.mem_145_sv2v_reg  <= w_data_i[17];
      \nz.mem_144_sv2v_reg  <= w_data_i[16];
      \nz.mem_143_sv2v_reg  <= w_data_i[15];
      \nz.mem_142_sv2v_reg  <= w_data_i[14];
      \nz.mem_141_sv2v_reg  <= w_data_i[13];
      \nz.mem_140_sv2v_reg  <= w_data_i[12];
      \nz.mem_139_sv2v_reg  <= w_data_i[11];
      \nz.mem_138_sv2v_reg  <= w_data_i[10];
      \nz.mem_137_sv2v_reg  <= w_data_i[9];
      \nz.mem_136_sv2v_reg  <= w_data_i[8];
      \nz.mem_135_sv2v_reg  <= w_data_i[7];
      \nz.mem_134_sv2v_reg  <= w_data_i[6];
      \nz.mem_133_sv2v_reg  <= w_data_i[5];
      \nz.mem_132_sv2v_reg  <= w_data_i[4];
      \nz.mem_131_sv2v_reg  <= w_data_i[3];
      \nz.mem_130_sv2v_reg  <= w_data_i[2];
      \nz.mem_129_sv2v_reg  <= w_data_i[1];
      \nz.mem_128_sv2v_reg  <= w_data_i[0];
    end 
    if(N377) begin
      \nz.mem_127_sv2v_reg  <= w_data_i[31];
      \nz.mem_126_sv2v_reg  <= w_data_i[30];
      \nz.mem_125_sv2v_reg  <= w_data_i[29];
      \nz.mem_124_sv2v_reg  <= w_data_i[28];
      \nz.mem_123_sv2v_reg  <= w_data_i[27];
      \nz.mem_122_sv2v_reg  <= w_data_i[26];
      \nz.mem_121_sv2v_reg  <= w_data_i[25];
      \nz.mem_120_sv2v_reg  <= w_data_i[24];
      \nz.mem_119_sv2v_reg  <= w_data_i[23];
      \nz.mem_118_sv2v_reg  <= w_data_i[22];
      \nz.mem_117_sv2v_reg  <= w_data_i[21];
      \nz.mem_116_sv2v_reg  <= w_data_i[20];
      \nz.mem_115_sv2v_reg  <= w_data_i[19];
      \nz.mem_114_sv2v_reg  <= w_data_i[18];
      \nz.mem_113_sv2v_reg  <= w_data_i[17];
      \nz.mem_112_sv2v_reg  <= w_data_i[16];
      \nz.mem_111_sv2v_reg  <= w_data_i[15];
      \nz.mem_110_sv2v_reg  <= w_data_i[14];
      \nz.mem_109_sv2v_reg  <= w_data_i[13];
      \nz.mem_108_sv2v_reg  <= w_data_i[12];
      \nz.mem_107_sv2v_reg  <= w_data_i[11];
      \nz.mem_106_sv2v_reg  <= w_data_i[10];
      \nz.mem_105_sv2v_reg  <= w_data_i[9];
      \nz.mem_104_sv2v_reg  <= w_data_i[8];
      \nz.mem_103_sv2v_reg  <= w_data_i[7];
      \nz.mem_102_sv2v_reg  <= w_data_i[6];
      \nz.mem_101_sv2v_reg  <= w_data_i[5];
      \nz.mem_100_sv2v_reg  <= w_data_i[4];
      \nz.mem_99_sv2v_reg  <= w_data_i[3];
      \nz.mem_98_sv2v_reg  <= w_data_i[2];
      \nz.mem_97_sv2v_reg  <= w_data_i[1];
      \nz.mem_96_sv2v_reg  <= w_data_i[0];
    end 
    if(N376) begin
      \nz.mem_95_sv2v_reg  <= w_data_i[31];
      \nz.mem_94_sv2v_reg  <= w_data_i[30];
      \nz.mem_93_sv2v_reg  <= w_data_i[29];
      \nz.mem_92_sv2v_reg  <= w_data_i[28];
      \nz.mem_91_sv2v_reg  <= w_data_i[27];
      \nz.mem_90_sv2v_reg  <= w_data_i[26];
      \nz.mem_89_sv2v_reg  <= w_data_i[25];
      \nz.mem_88_sv2v_reg  <= w_data_i[24];
      \nz.mem_87_sv2v_reg  <= w_data_i[23];
      \nz.mem_86_sv2v_reg  <= w_data_i[22];
      \nz.mem_85_sv2v_reg  <= w_data_i[21];
      \nz.mem_84_sv2v_reg  <= w_data_i[20];
      \nz.mem_83_sv2v_reg  <= w_data_i[19];
      \nz.mem_82_sv2v_reg  <= w_data_i[18];
      \nz.mem_81_sv2v_reg  <= w_data_i[17];
      \nz.mem_80_sv2v_reg  <= w_data_i[16];
      \nz.mem_79_sv2v_reg  <= w_data_i[15];
      \nz.mem_78_sv2v_reg  <= w_data_i[14];
      \nz.mem_77_sv2v_reg  <= w_data_i[13];
      \nz.mem_76_sv2v_reg  <= w_data_i[12];
      \nz.mem_75_sv2v_reg  <= w_data_i[11];
      \nz.mem_74_sv2v_reg  <= w_data_i[10];
      \nz.mem_73_sv2v_reg  <= w_data_i[9];
      \nz.mem_72_sv2v_reg  <= w_data_i[8];
      \nz.mem_71_sv2v_reg  <= w_data_i[7];
      \nz.mem_70_sv2v_reg  <= w_data_i[6];
      \nz.mem_69_sv2v_reg  <= w_data_i[5];
      \nz.mem_68_sv2v_reg  <= w_data_i[4];
      \nz.mem_67_sv2v_reg  <= w_data_i[3];
      \nz.mem_66_sv2v_reg  <= w_data_i[2];
      \nz.mem_65_sv2v_reg  <= w_data_i[1];
      \nz.mem_64_sv2v_reg  <= w_data_i[0];
    end 
    if(N375) begin
      \nz.mem_63_sv2v_reg  <= w_data_i[31];
      \nz.mem_62_sv2v_reg  <= w_data_i[30];
      \nz.mem_61_sv2v_reg  <= w_data_i[29];
      \nz.mem_60_sv2v_reg  <= w_data_i[28];
      \nz.mem_59_sv2v_reg  <= w_data_i[27];
      \nz.mem_58_sv2v_reg  <= w_data_i[26];
      \nz.mem_57_sv2v_reg  <= w_data_i[25];
      \nz.mem_56_sv2v_reg  <= w_data_i[24];
      \nz.mem_55_sv2v_reg  <= w_data_i[23];
      \nz.mem_54_sv2v_reg  <= w_data_i[22];
      \nz.mem_53_sv2v_reg  <= w_data_i[21];
      \nz.mem_52_sv2v_reg  <= w_data_i[20];
      \nz.mem_51_sv2v_reg  <= w_data_i[19];
      \nz.mem_50_sv2v_reg  <= w_data_i[18];
      \nz.mem_49_sv2v_reg  <= w_data_i[17];
      \nz.mem_48_sv2v_reg  <= w_data_i[16];
      \nz.mem_47_sv2v_reg  <= w_data_i[15];
      \nz.mem_46_sv2v_reg  <= w_data_i[14];
      \nz.mem_45_sv2v_reg  <= w_data_i[13];
      \nz.mem_44_sv2v_reg  <= w_data_i[12];
      \nz.mem_43_sv2v_reg  <= w_data_i[11];
      \nz.mem_42_sv2v_reg  <= w_data_i[10];
      \nz.mem_41_sv2v_reg  <= w_data_i[9];
      \nz.mem_40_sv2v_reg  <= w_data_i[8];
      \nz.mem_39_sv2v_reg  <= w_data_i[7];
      \nz.mem_38_sv2v_reg  <= w_data_i[6];
      \nz.mem_37_sv2v_reg  <= w_data_i[5];
      \nz.mem_36_sv2v_reg  <= w_data_i[4];
      \nz.mem_35_sv2v_reg  <= w_data_i[3];
      \nz.mem_34_sv2v_reg  <= w_data_i[2];
      \nz.mem_33_sv2v_reg  <= w_data_i[1];
      \nz.mem_32_sv2v_reg  <= w_data_i[0];
    end 
    if(N374) begin
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p50_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [31:0] w_data_i;
  input [5:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p50_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p32_els_p50_ready_THEN_valid_p1
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,full,empty,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,
  sv2v_dc_6;
  wire [5:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p50
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(v_i),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p32_els_p50_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(v_i),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p32_els_p50_harden_p0_ready_THEN_valid_p1
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p32_els_p50_ready_THEN_valid_p1
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_fifo_1r1w_small_credit_on_input
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  credit_o,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output credit_o;
  output v_o;
  wire [31:0] data_o;
  wire credit_o,v_o,ready;
  reg credit_o_sv2v_reg;
  assign credit_o = credit_o_sv2v_reg;

  bsg_fifo_1r1w_small_width_p32_els_p50_harden_p0_ready_THEN_valid_p1
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


  always @(posedge clk_i) begin
    if(reset_i) begin
      credit_o_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      credit_o_sv2v_reg <= yumi_i;
    end 
  end


endmodule

