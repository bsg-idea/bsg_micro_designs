

module top
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [68:0] cache_pkt_i;
  output [31:0] data_o;
  output [28:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output ready_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output v_we_o;

  bsg_cache
  wrapper
  (
    .cache_pkt_i(cache_pkt_i),
    .data_o(data_o),
    .dma_pkt_o(dma_pkt_o),
    .dma_data_i(dma_data_i),
    .dma_data_o(dma_data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_yumi_i(dma_data_yumi_i),
    .ready_o(ready_o),
    .v_o(v_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_data_ready_o(dma_data_ready_o),
    .dma_data_v_o(dma_data_v_o),
    .v_we_o(v_we_o)
  );


endmodule



module bsg_cache_pkt_decode_data_width_p32_addr_width_p28
(
  cache_pkt_i,
  decode_o
);

  input [68:0] cache_pkt_i;
  output [15:0] decode_o;
  wire [15:0] decode_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N42,
  N43,N44,N46,N48,N49,N50,N51,N52,N54,N56,N57,N59,N61,N62,N63,N64,N66,N67,N68,N69,
  N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,
  N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,
  N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,
  N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135;
  assign N7 = cache_pkt_i[67] | cache_pkt_i[66];
  assign N8 = N42 | N36;
  assign N9 = N7 | N8;
  assign N10 = N48 | cache_pkt_i[66];
  assign N11 = N10 | N8;
  assign N12 = cache_pkt_i[67] | N61;
  assign N13 = N12 | N8;
  assign N15 = N42 | cache_pkt_i[64];
  assign N16 = N7 | N15;
  assign N17 = N10 | N15;
  assign N18 = N12 | N15;
  assign N20 = cache_pkt_i[65] | N36;
  assign N21 = N7 | N20;
  assign N22 = N10 | N20;
  assign N23 = N12 | N20;
  assign N25 = N48 & N61;
  assign N26 = N42 & N36;
  assign N27 = N25 & N26;
  assign N28 = cache_pkt_i[65] | cache_pkt_i[64];
  assign N29 = N10 | N28;
  assign N30 = N12 | N28;
  assign N32 = cache_pkt_i[67] & cache_pkt_i[66];
  assign N35 = ~cache_pkt_i[68];
  assign N36 = ~cache_pkt_i[64];
  assign N37 = cache_pkt_i[67] | N35;
  assign N38 = cache_pkt_i[66] | N37;
  assign N39 = cache_pkt_i[65] | N38;
  assign N40 = N36 | N39;
  assign decode_o[8] = ~N40;
  assign N42 = ~cache_pkt_i[65];
  assign N43 = N42 | N38;
  assign N44 = cache_pkt_i[64] | N43;
  assign decode_o[7] = ~N44;
  assign N46 = N36 | N43;
  assign decode_o[6] = ~N46;
  assign N48 = ~cache_pkt_i[67];
  assign N49 = N48 | N35;
  assign N50 = cache_pkt_i[66] | N49;
  assign N51 = cache_pkt_i[65] | N50;
  assign N52 = cache_pkt_i[64] | N51;
  assign decode_o[5] = ~N52;
  assign N54 = N36 | N51;
  assign decode_o[4] = ~N54;
  assign N56 = N42 | N50;
  assign N57 = cache_pkt_i[64] | N56;
  assign decode_o[3] = ~N57;
  assign N59 = N36 | N56;
  assign decode_o[2] = ~N59;
  assign N61 = ~cache_pkt_i[66];
  assign N62 = N61 | N49;
  assign N63 = cache_pkt_i[65] | N62;
  assign N64 = cache_pkt_i[64] | N63;
  assign decode_o[1] = ~N64;
  assign N66 = cache_pkt_i[67] | cache_pkt_i[68];
  assign N67 = cache_pkt_i[66] | N66;
  assign N68 = cache_pkt_i[65] | N67;
  assign N69 = cache_pkt_i[64] | N68;
  assign N70 = ~N69;
  assign N71 = N36 | N68;
  assign N72 = ~N71;
  assign N73 = N42 | N67;
  assign N74 = cache_pkt_i[64] | N73;
  assign N75 = ~N74;
  assign N76 = N36 | N73;
  assign N77 = ~N76;
  assign N78 = N48 | cache_pkt_i[68];
  assign N79 = N61 | N78;
  assign N80 = cache_pkt_i[65] | N79;
  assign N81 = cache_pkt_i[64] | N80;
  assign N82 = ~N81;
  assign N83 = N36 | N80;
  assign N84 = ~N83;
  assign N85 = N61 | N66;
  assign N86 = cache_pkt_i[65] | N85;
  assign N87 = cache_pkt_i[64] | N86;
  assign N88 = ~N87;
  assign N89 = N36 | N86;
  assign N90 = ~N89;
  assign N91 = N42 | N85;
  assign N92 = cache_pkt_i[64] | N91;
  assign N93 = ~N92;
  assign N94 = N36 | N91;
  assign N95 = ~N94;
  assign N96 = cache_pkt_i[66] | N78;
  assign N97 = cache_pkt_i[65] | N96;
  assign N98 = cache_pkt_i[64] | N97;
  assign N99 = ~N98;
  assign N100 = N36 | N97;
  assign N101 = ~N100;
  assign N102 = N42 | N96;
  assign N103 = cache_pkt_i[64] | N102;
  assign N104 = ~N103;
  assign N105 = N36 | N102;
  assign N106 = ~N105;
  assign N107 = cache_pkt_i[64] | N39;
  assign decode_o[9] = ~N107;
  assign { N34, N33 } = (N0)? { 1'b1, 1'b1 } : 
                        (N1)? { 1'b1, 1'b0 } : 
                        (N2)? { 1'b0, 1'b1 } : 
                        (N3)? { 1'b0, 1'b0 } : 
                        (N4)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = N14;
  assign N1 = N19;
  assign N2 = N24;
  assign N3 = N31;
  assign N4 = N32;
  assign decode_o[15:14] = (N5)? { N34, N33 } : 
                           (N6)? { 1'b0, 1'b0 } : 1'b0;
  assign N5 = N35;
  assign N6 = cache_pkt_i[68];
  assign N14 = N111 | N112;
  assign N111 = N109 | N110;
  assign N109 = ~N9;
  assign N110 = ~N11;
  assign N112 = ~N13;
  assign N19 = N115 | N116;
  assign N115 = N113 | N114;
  assign N113 = ~N16;
  assign N114 = ~N17;
  assign N116 = ~N18;
  assign N24 = N119 | N120;
  assign N119 = N117 | N118;
  assign N117 = ~N21;
  assign N118 = ~N22;
  assign N120 = ~N23;
  assign N31 = N122 | N123;
  assign N122 = N27 | N121;
  assign N121 = ~N29;
  assign N123 = ~N30;
  assign decode_o[12] = N82 | N84;
  assign decode_o[13] = N125 | N77;
  assign N125 = N124 | N75;
  assign N124 = N70 | N72;
  assign decode_o[11] = N132 | N82;
  assign N132 = N131 | N95;
  assign N131 = N130 | N93;
  assign N130 = N129 | N90;
  assign N129 = N128 | N88;
  assign N128 = N127 | N77;
  assign N127 = N126 | N75;
  assign N126 = N70 | N72;
  assign decode_o[10] = N135 | N84;
  assign N135 = N134 | N106;
  assign N134 = N133 | N104;
  assign N133 = N99 | N101;
  assign decode_o[0] = ~decode_o[9];

endmodule



module bsg_dff_width_p1
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  reg [0:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[0:0] } <= { data_i[0:0] };
    end 
  end


endmodule



module bsg_dff_en_width_p40_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [39:0] data_i;
  output [39:0] data_o;
  input clk_i;
  input en_i;
  reg [39:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[39:0] } <= { data_i[39:0] };
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p40
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [39:0] data_i;
  output [39:0] data_o;
  input clk_i;
  input en_i;
  wire [39:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p40_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p40_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [39:0] data_i;
  input [5:0] addr_i;
  input [39:0] w_mask_i;
  output [39:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [39:0] data_o,data_out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,read_en,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  llr_read_en_r,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,
  N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,
  N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,
  N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,
  N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,
  N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,
  N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,
  N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,
  N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,
  N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,
  N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,
  N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,
  N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,
  N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,
  N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,
  N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,
  N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,
  N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,
  N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,
  N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,
  N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,
  N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,
  N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,
  N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,
  N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,
  N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,
  N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,
  N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,
  N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,
  N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,
  N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,
  N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,
  N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,
  N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,
  N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,
  N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,
  N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,
  N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,
  N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,
  N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,
  N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,
  N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,
  N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,
  N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,
  N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,
  N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,
  N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,
  N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,
  N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,
  N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,
  N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,
  N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,
  N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,
  N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,
  N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,
  N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,
  N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,
  N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,
  N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,
  N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,
  N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,
  N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,
  N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,
  N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,
  N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,
  N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,
  N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,
  N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,
  N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,
  N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,
  N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,
  N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,
  N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,
  N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,
  N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,
  N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,
  N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,
  N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,
  N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
  N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,
  N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,
  N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,
  N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,
  N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,
  N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,
  N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,
  N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,
  N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,
  N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,
  N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,
  N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,
  N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,
  N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,
  N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,
  N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,
  N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,
  N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,
  N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,
  N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,
  N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,
  N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,
  N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,
  N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,
  N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,
  N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,
  N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,
  N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,
  N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,
  N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,
  N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,
  N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,
  N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,
  N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,
  N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,
  N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,
  N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,
  N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,
  N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,
  N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,
  N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,
  N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,
  N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,
  N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,
  N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,
  N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,
  N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,
  N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,
  N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,
  N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,
  N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,
  N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,
  N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,
  N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,
  N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,
  N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,
  N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,
  N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,
  N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,
  N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,
  N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,
  N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,
  N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,
  N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,
  N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
  N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,
  N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,
  N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,
  N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,
  N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,
  N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,
  N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,
  N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,
  N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,
  N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,
  N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,
  N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,
  N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,
  N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,
  N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,
  N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,
  N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,
  N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,
  N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,
  N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,
  N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,
  N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,
  N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,
  N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,
  N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,
  N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,
  N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,
  N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,
  N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,
  N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,
  N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,
  N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,
  N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,
  N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,
  N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,
  N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,
  N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,
  N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,
  N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,
  N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,
  N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,
  N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,
  N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,
  N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,
  N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,
  N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,
  N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,
  N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,
  N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,
  N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,
  N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,
  N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,
  N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,
  N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,
  N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,
  N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,
  N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,
  N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,
  N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,
  N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,
  N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,
  N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,
  N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,
  N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,
  N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,
  N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,
  N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,
  N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,
  N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,
  N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,
  N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,
  N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,
  N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,
  N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,
  N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,
  N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,
  N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,
  N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,
  N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,
  N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,
  N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,
  N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,
  N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,
  N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,
  N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,
  N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,
  N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,
  N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,
  N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,
  N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,
  N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,
  N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,
  N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,
  N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,
  N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,
  N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,
  N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,
  N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,
  N4208,N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,
  N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,
  N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,
  N4248,N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,
  N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,
  N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,
  N4288,N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,
  N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,
  N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,
  N4328,N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,
  N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,
  N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,
  N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,
  N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,
  N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,
  N4408,N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,
  N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,
  N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,
  N4448,N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,
  N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,
  N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,
  N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,
  N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,
  N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,
  N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,
  N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,
  N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,
  N4568,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,
  N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,
  N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,
  N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,
  N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,
  N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,
  N4648,N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,
  N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,
  N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,
  N4688,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,
  N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,
  N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,
  N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,
  N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,
  N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,
  N4768,N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,
  N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,
  N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,
  N4808,N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,
  N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,
  N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,
  N4848,N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,
  N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,
  N4874,N4875,N4876,N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,
  N4888,N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,N4900,
  N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,
  N4914,N4915,N4916,N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,
  N4928,N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,
  N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,
  N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,
  N4968,N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,
  N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,
  N4994,N4995,N4996,N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,
  N5008,N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,
  N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,
  N5034,N5035,N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,
  N5048,N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,
  N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,
  N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,
  N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,
  N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,
  N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,
  N5128,N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,
  N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,
  N5154,N5155,N5156,N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,
  N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,
  N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,
  N5194,N5195,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,
  N5208,N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,
  N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,
  N5234,N5235,N5236,N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,
  N5248,N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,
  N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,
  N5274,N5275,N5276,N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,
  N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,
  N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,
  N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,
  N5328,N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,
  N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,
  N5354,N5355,N5356,N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,
  N5368,N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,
  N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,
  N5394,N5395,N5396,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,
  N5408,N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,
  N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,
  N5434,N5435,N5436,N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,
  N5448,N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,
  N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,
  N5474,N5475,N5476,N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,
  N5488,N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,
  N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,
  N5514,N5515,N5516,N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,
  N5528,N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,
  N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,
  N5554,N5555,N5556,N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,
  N5568,N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,
  N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,
  N5594,N5595,N5596,N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,
  N5608,N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,
  N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,
  N5634,N5635,N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,
  N5648,N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,
  N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,
  N5674,N5675,N5676,N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,
  N5688,N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,
  N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,
  N5714,N5715,N5716,N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,
  N5728,N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,
  N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,
  N5754,N5755,N5756,N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,
  N5768,N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,N5780,
  N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,
  N5794,N5795,N5796,N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,
  N5808,N5809,N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,N5820,
  N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,
  N5834,N5835,N5836,N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,
  N5848,N5849,N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860,
  N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,
  N5874,N5875,N5876,N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,
  N5888,N5889,N5890,N5891,N5892,N5893;
  reg [5:0] addr_r;
  reg [2559:0] mem;
  assign data_out[39] = (N115)? mem[39] : 
                        (N117)? mem[79] : 
                        (N119)? mem[119] : 
                        (N121)? mem[159] : 
                        (N123)? mem[199] : 
                        (N125)? mem[239] : 
                        (N127)? mem[279] : 
                        (N129)? mem[319] : 
                        (N131)? mem[359] : 
                        (N133)? mem[399] : 
                        (N135)? mem[439] : 
                        (N137)? mem[479] : 
                        (N139)? mem[519] : 
                        (N141)? mem[559] : 
                        (N143)? mem[599] : 
                        (N145)? mem[639] : 
                        (N147)? mem[679] : 
                        (N149)? mem[719] : 
                        (N151)? mem[759] : 
                        (N153)? mem[799] : 
                        (N155)? mem[839] : 
                        (N157)? mem[879] : 
                        (N159)? mem[919] : 
                        (N161)? mem[959] : 
                        (N163)? mem[999] : 
                        (N165)? mem[1039] : 
                        (N167)? mem[1079] : 
                        (N169)? mem[1119] : 
                        (N171)? mem[1159] : 
                        (N173)? mem[1199] : 
                        (N175)? mem[1239] : 
                        (N177)? mem[1279] : 
                        (N116)? mem[1319] : 
                        (N118)? mem[1359] : 
                        (N120)? mem[1399] : 
                        (N122)? mem[1439] : 
                        (N124)? mem[1479] : 
                        (N126)? mem[1519] : 
                        (N128)? mem[1559] : 
                        (N130)? mem[1599] : 
                        (N132)? mem[1639] : 
                        (N134)? mem[1679] : 
                        (N136)? mem[1719] : 
                        (N138)? mem[1759] : 
                        (N140)? mem[1799] : 
                        (N142)? mem[1839] : 
                        (N144)? mem[1879] : 
                        (N146)? mem[1919] : 
                        (N148)? mem[1959] : 
                        (N150)? mem[1999] : 
                        (N152)? mem[2039] : 
                        (N154)? mem[2079] : 
                        (N156)? mem[2119] : 
                        (N158)? mem[2159] : 
                        (N160)? mem[2199] : 
                        (N162)? mem[2239] : 
                        (N164)? mem[2279] : 
                        (N166)? mem[2319] : 
                        (N168)? mem[2359] : 
                        (N170)? mem[2399] : 
                        (N172)? mem[2439] : 
                        (N174)? mem[2479] : 
                        (N176)? mem[2519] : 
                        (N178)? mem[2559] : 1'b0;
  assign data_out[38] = (N115)? mem[38] : 
                        (N117)? mem[78] : 
                        (N119)? mem[118] : 
                        (N121)? mem[158] : 
                        (N123)? mem[198] : 
                        (N125)? mem[238] : 
                        (N127)? mem[278] : 
                        (N129)? mem[318] : 
                        (N131)? mem[358] : 
                        (N133)? mem[398] : 
                        (N135)? mem[438] : 
                        (N137)? mem[478] : 
                        (N139)? mem[518] : 
                        (N141)? mem[558] : 
                        (N143)? mem[598] : 
                        (N145)? mem[638] : 
                        (N147)? mem[678] : 
                        (N149)? mem[718] : 
                        (N151)? mem[758] : 
                        (N153)? mem[798] : 
                        (N155)? mem[838] : 
                        (N157)? mem[878] : 
                        (N159)? mem[918] : 
                        (N161)? mem[958] : 
                        (N163)? mem[998] : 
                        (N165)? mem[1038] : 
                        (N167)? mem[1078] : 
                        (N169)? mem[1118] : 
                        (N171)? mem[1158] : 
                        (N173)? mem[1198] : 
                        (N175)? mem[1238] : 
                        (N177)? mem[1278] : 
                        (N116)? mem[1318] : 
                        (N118)? mem[1358] : 
                        (N120)? mem[1398] : 
                        (N122)? mem[1438] : 
                        (N124)? mem[1478] : 
                        (N126)? mem[1518] : 
                        (N128)? mem[1558] : 
                        (N130)? mem[1598] : 
                        (N132)? mem[1638] : 
                        (N134)? mem[1678] : 
                        (N136)? mem[1718] : 
                        (N138)? mem[1758] : 
                        (N140)? mem[1798] : 
                        (N142)? mem[1838] : 
                        (N144)? mem[1878] : 
                        (N146)? mem[1918] : 
                        (N148)? mem[1958] : 
                        (N150)? mem[1998] : 
                        (N152)? mem[2038] : 
                        (N154)? mem[2078] : 
                        (N156)? mem[2118] : 
                        (N158)? mem[2158] : 
                        (N160)? mem[2198] : 
                        (N162)? mem[2238] : 
                        (N164)? mem[2278] : 
                        (N166)? mem[2318] : 
                        (N168)? mem[2358] : 
                        (N170)? mem[2398] : 
                        (N172)? mem[2438] : 
                        (N174)? mem[2478] : 
                        (N176)? mem[2518] : 
                        (N178)? mem[2558] : 1'b0;
  assign data_out[37] = (N115)? mem[37] : 
                        (N117)? mem[77] : 
                        (N119)? mem[117] : 
                        (N121)? mem[157] : 
                        (N123)? mem[197] : 
                        (N125)? mem[237] : 
                        (N127)? mem[277] : 
                        (N129)? mem[317] : 
                        (N131)? mem[357] : 
                        (N133)? mem[397] : 
                        (N135)? mem[437] : 
                        (N137)? mem[477] : 
                        (N139)? mem[517] : 
                        (N141)? mem[557] : 
                        (N143)? mem[597] : 
                        (N145)? mem[637] : 
                        (N147)? mem[677] : 
                        (N149)? mem[717] : 
                        (N151)? mem[757] : 
                        (N153)? mem[797] : 
                        (N155)? mem[837] : 
                        (N157)? mem[877] : 
                        (N159)? mem[917] : 
                        (N161)? mem[957] : 
                        (N163)? mem[997] : 
                        (N165)? mem[1037] : 
                        (N167)? mem[1077] : 
                        (N169)? mem[1117] : 
                        (N171)? mem[1157] : 
                        (N173)? mem[1197] : 
                        (N175)? mem[1237] : 
                        (N177)? mem[1277] : 
                        (N116)? mem[1317] : 
                        (N118)? mem[1357] : 
                        (N120)? mem[1397] : 
                        (N122)? mem[1437] : 
                        (N124)? mem[1477] : 
                        (N126)? mem[1517] : 
                        (N128)? mem[1557] : 
                        (N130)? mem[1597] : 
                        (N132)? mem[1637] : 
                        (N134)? mem[1677] : 
                        (N136)? mem[1717] : 
                        (N138)? mem[1757] : 
                        (N140)? mem[1797] : 
                        (N142)? mem[1837] : 
                        (N144)? mem[1877] : 
                        (N146)? mem[1917] : 
                        (N148)? mem[1957] : 
                        (N150)? mem[1997] : 
                        (N152)? mem[2037] : 
                        (N154)? mem[2077] : 
                        (N156)? mem[2117] : 
                        (N158)? mem[2157] : 
                        (N160)? mem[2197] : 
                        (N162)? mem[2237] : 
                        (N164)? mem[2277] : 
                        (N166)? mem[2317] : 
                        (N168)? mem[2357] : 
                        (N170)? mem[2397] : 
                        (N172)? mem[2437] : 
                        (N174)? mem[2477] : 
                        (N176)? mem[2517] : 
                        (N178)? mem[2557] : 1'b0;
  assign data_out[36] = (N115)? mem[36] : 
                        (N117)? mem[76] : 
                        (N119)? mem[116] : 
                        (N121)? mem[156] : 
                        (N123)? mem[196] : 
                        (N125)? mem[236] : 
                        (N127)? mem[276] : 
                        (N129)? mem[316] : 
                        (N131)? mem[356] : 
                        (N133)? mem[396] : 
                        (N135)? mem[436] : 
                        (N137)? mem[476] : 
                        (N139)? mem[516] : 
                        (N141)? mem[556] : 
                        (N143)? mem[596] : 
                        (N145)? mem[636] : 
                        (N147)? mem[676] : 
                        (N149)? mem[716] : 
                        (N151)? mem[756] : 
                        (N153)? mem[796] : 
                        (N155)? mem[836] : 
                        (N157)? mem[876] : 
                        (N159)? mem[916] : 
                        (N161)? mem[956] : 
                        (N163)? mem[996] : 
                        (N165)? mem[1036] : 
                        (N167)? mem[1076] : 
                        (N169)? mem[1116] : 
                        (N171)? mem[1156] : 
                        (N173)? mem[1196] : 
                        (N175)? mem[1236] : 
                        (N177)? mem[1276] : 
                        (N116)? mem[1316] : 
                        (N118)? mem[1356] : 
                        (N120)? mem[1396] : 
                        (N122)? mem[1436] : 
                        (N124)? mem[1476] : 
                        (N126)? mem[1516] : 
                        (N128)? mem[1556] : 
                        (N130)? mem[1596] : 
                        (N132)? mem[1636] : 
                        (N134)? mem[1676] : 
                        (N136)? mem[1716] : 
                        (N138)? mem[1756] : 
                        (N140)? mem[1796] : 
                        (N142)? mem[1836] : 
                        (N144)? mem[1876] : 
                        (N146)? mem[1916] : 
                        (N148)? mem[1956] : 
                        (N150)? mem[1996] : 
                        (N152)? mem[2036] : 
                        (N154)? mem[2076] : 
                        (N156)? mem[2116] : 
                        (N158)? mem[2156] : 
                        (N160)? mem[2196] : 
                        (N162)? mem[2236] : 
                        (N164)? mem[2276] : 
                        (N166)? mem[2316] : 
                        (N168)? mem[2356] : 
                        (N170)? mem[2396] : 
                        (N172)? mem[2436] : 
                        (N174)? mem[2476] : 
                        (N176)? mem[2516] : 
                        (N178)? mem[2556] : 1'b0;
  assign data_out[35] = (N115)? mem[35] : 
                        (N117)? mem[75] : 
                        (N119)? mem[115] : 
                        (N121)? mem[155] : 
                        (N123)? mem[195] : 
                        (N125)? mem[235] : 
                        (N127)? mem[275] : 
                        (N129)? mem[315] : 
                        (N131)? mem[355] : 
                        (N133)? mem[395] : 
                        (N135)? mem[435] : 
                        (N137)? mem[475] : 
                        (N139)? mem[515] : 
                        (N141)? mem[555] : 
                        (N143)? mem[595] : 
                        (N145)? mem[635] : 
                        (N147)? mem[675] : 
                        (N149)? mem[715] : 
                        (N151)? mem[755] : 
                        (N153)? mem[795] : 
                        (N155)? mem[835] : 
                        (N157)? mem[875] : 
                        (N159)? mem[915] : 
                        (N161)? mem[955] : 
                        (N163)? mem[995] : 
                        (N165)? mem[1035] : 
                        (N167)? mem[1075] : 
                        (N169)? mem[1115] : 
                        (N171)? mem[1155] : 
                        (N173)? mem[1195] : 
                        (N175)? mem[1235] : 
                        (N177)? mem[1275] : 
                        (N116)? mem[1315] : 
                        (N118)? mem[1355] : 
                        (N120)? mem[1395] : 
                        (N122)? mem[1435] : 
                        (N124)? mem[1475] : 
                        (N126)? mem[1515] : 
                        (N128)? mem[1555] : 
                        (N130)? mem[1595] : 
                        (N132)? mem[1635] : 
                        (N134)? mem[1675] : 
                        (N136)? mem[1715] : 
                        (N138)? mem[1755] : 
                        (N140)? mem[1795] : 
                        (N142)? mem[1835] : 
                        (N144)? mem[1875] : 
                        (N146)? mem[1915] : 
                        (N148)? mem[1955] : 
                        (N150)? mem[1995] : 
                        (N152)? mem[2035] : 
                        (N154)? mem[2075] : 
                        (N156)? mem[2115] : 
                        (N158)? mem[2155] : 
                        (N160)? mem[2195] : 
                        (N162)? mem[2235] : 
                        (N164)? mem[2275] : 
                        (N166)? mem[2315] : 
                        (N168)? mem[2355] : 
                        (N170)? mem[2395] : 
                        (N172)? mem[2435] : 
                        (N174)? mem[2475] : 
                        (N176)? mem[2515] : 
                        (N178)? mem[2555] : 1'b0;
  assign data_out[34] = (N115)? mem[34] : 
                        (N117)? mem[74] : 
                        (N119)? mem[114] : 
                        (N121)? mem[154] : 
                        (N123)? mem[194] : 
                        (N125)? mem[234] : 
                        (N127)? mem[274] : 
                        (N129)? mem[314] : 
                        (N131)? mem[354] : 
                        (N133)? mem[394] : 
                        (N135)? mem[434] : 
                        (N137)? mem[474] : 
                        (N139)? mem[514] : 
                        (N141)? mem[554] : 
                        (N143)? mem[594] : 
                        (N145)? mem[634] : 
                        (N147)? mem[674] : 
                        (N149)? mem[714] : 
                        (N151)? mem[754] : 
                        (N153)? mem[794] : 
                        (N155)? mem[834] : 
                        (N157)? mem[874] : 
                        (N159)? mem[914] : 
                        (N161)? mem[954] : 
                        (N163)? mem[994] : 
                        (N165)? mem[1034] : 
                        (N167)? mem[1074] : 
                        (N169)? mem[1114] : 
                        (N171)? mem[1154] : 
                        (N173)? mem[1194] : 
                        (N175)? mem[1234] : 
                        (N177)? mem[1274] : 
                        (N116)? mem[1314] : 
                        (N118)? mem[1354] : 
                        (N120)? mem[1394] : 
                        (N122)? mem[1434] : 
                        (N124)? mem[1474] : 
                        (N126)? mem[1514] : 
                        (N128)? mem[1554] : 
                        (N130)? mem[1594] : 
                        (N132)? mem[1634] : 
                        (N134)? mem[1674] : 
                        (N136)? mem[1714] : 
                        (N138)? mem[1754] : 
                        (N140)? mem[1794] : 
                        (N142)? mem[1834] : 
                        (N144)? mem[1874] : 
                        (N146)? mem[1914] : 
                        (N148)? mem[1954] : 
                        (N150)? mem[1994] : 
                        (N152)? mem[2034] : 
                        (N154)? mem[2074] : 
                        (N156)? mem[2114] : 
                        (N158)? mem[2154] : 
                        (N160)? mem[2194] : 
                        (N162)? mem[2234] : 
                        (N164)? mem[2274] : 
                        (N166)? mem[2314] : 
                        (N168)? mem[2354] : 
                        (N170)? mem[2394] : 
                        (N172)? mem[2434] : 
                        (N174)? mem[2474] : 
                        (N176)? mem[2514] : 
                        (N178)? mem[2554] : 1'b0;
  assign data_out[33] = (N115)? mem[33] : 
                        (N117)? mem[73] : 
                        (N119)? mem[113] : 
                        (N121)? mem[153] : 
                        (N123)? mem[193] : 
                        (N125)? mem[233] : 
                        (N127)? mem[273] : 
                        (N129)? mem[313] : 
                        (N131)? mem[353] : 
                        (N133)? mem[393] : 
                        (N135)? mem[433] : 
                        (N137)? mem[473] : 
                        (N139)? mem[513] : 
                        (N141)? mem[553] : 
                        (N143)? mem[593] : 
                        (N145)? mem[633] : 
                        (N147)? mem[673] : 
                        (N149)? mem[713] : 
                        (N151)? mem[753] : 
                        (N153)? mem[793] : 
                        (N155)? mem[833] : 
                        (N157)? mem[873] : 
                        (N159)? mem[913] : 
                        (N161)? mem[953] : 
                        (N163)? mem[993] : 
                        (N165)? mem[1033] : 
                        (N167)? mem[1073] : 
                        (N169)? mem[1113] : 
                        (N171)? mem[1153] : 
                        (N173)? mem[1193] : 
                        (N175)? mem[1233] : 
                        (N177)? mem[1273] : 
                        (N116)? mem[1313] : 
                        (N118)? mem[1353] : 
                        (N120)? mem[1393] : 
                        (N122)? mem[1433] : 
                        (N124)? mem[1473] : 
                        (N126)? mem[1513] : 
                        (N128)? mem[1553] : 
                        (N130)? mem[1593] : 
                        (N132)? mem[1633] : 
                        (N134)? mem[1673] : 
                        (N136)? mem[1713] : 
                        (N138)? mem[1753] : 
                        (N140)? mem[1793] : 
                        (N142)? mem[1833] : 
                        (N144)? mem[1873] : 
                        (N146)? mem[1913] : 
                        (N148)? mem[1953] : 
                        (N150)? mem[1993] : 
                        (N152)? mem[2033] : 
                        (N154)? mem[2073] : 
                        (N156)? mem[2113] : 
                        (N158)? mem[2153] : 
                        (N160)? mem[2193] : 
                        (N162)? mem[2233] : 
                        (N164)? mem[2273] : 
                        (N166)? mem[2313] : 
                        (N168)? mem[2353] : 
                        (N170)? mem[2393] : 
                        (N172)? mem[2433] : 
                        (N174)? mem[2473] : 
                        (N176)? mem[2513] : 
                        (N178)? mem[2553] : 1'b0;
  assign data_out[32] = (N115)? mem[32] : 
                        (N117)? mem[72] : 
                        (N119)? mem[112] : 
                        (N121)? mem[152] : 
                        (N123)? mem[192] : 
                        (N125)? mem[232] : 
                        (N127)? mem[272] : 
                        (N129)? mem[312] : 
                        (N131)? mem[352] : 
                        (N133)? mem[392] : 
                        (N135)? mem[432] : 
                        (N137)? mem[472] : 
                        (N139)? mem[512] : 
                        (N141)? mem[552] : 
                        (N143)? mem[592] : 
                        (N145)? mem[632] : 
                        (N147)? mem[672] : 
                        (N149)? mem[712] : 
                        (N151)? mem[752] : 
                        (N153)? mem[792] : 
                        (N155)? mem[832] : 
                        (N157)? mem[872] : 
                        (N159)? mem[912] : 
                        (N161)? mem[952] : 
                        (N163)? mem[992] : 
                        (N165)? mem[1032] : 
                        (N167)? mem[1072] : 
                        (N169)? mem[1112] : 
                        (N171)? mem[1152] : 
                        (N173)? mem[1192] : 
                        (N175)? mem[1232] : 
                        (N177)? mem[1272] : 
                        (N116)? mem[1312] : 
                        (N118)? mem[1352] : 
                        (N120)? mem[1392] : 
                        (N122)? mem[1432] : 
                        (N124)? mem[1472] : 
                        (N126)? mem[1512] : 
                        (N128)? mem[1552] : 
                        (N130)? mem[1592] : 
                        (N132)? mem[1632] : 
                        (N134)? mem[1672] : 
                        (N136)? mem[1712] : 
                        (N138)? mem[1752] : 
                        (N140)? mem[1792] : 
                        (N142)? mem[1832] : 
                        (N144)? mem[1872] : 
                        (N146)? mem[1912] : 
                        (N148)? mem[1952] : 
                        (N150)? mem[1992] : 
                        (N152)? mem[2032] : 
                        (N154)? mem[2072] : 
                        (N156)? mem[2112] : 
                        (N158)? mem[2152] : 
                        (N160)? mem[2192] : 
                        (N162)? mem[2232] : 
                        (N164)? mem[2272] : 
                        (N166)? mem[2312] : 
                        (N168)? mem[2352] : 
                        (N170)? mem[2392] : 
                        (N172)? mem[2432] : 
                        (N174)? mem[2472] : 
                        (N176)? mem[2512] : 
                        (N178)? mem[2552] : 1'b0;
  assign data_out[31] = (N115)? mem[31] : 
                        (N117)? mem[71] : 
                        (N119)? mem[111] : 
                        (N121)? mem[151] : 
                        (N123)? mem[191] : 
                        (N125)? mem[231] : 
                        (N127)? mem[271] : 
                        (N129)? mem[311] : 
                        (N131)? mem[351] : 
                        (N133)? mem[391] : 
                        (N135)? mem[431] : 
                        (N137)? mem[471] : 
                        (N139)? mem[511] : 
                        (N141)? mem[551] : 
                        (N143)? mem[591] : 
                        (N145)? mem[631] : 
                        (N147)? mem[671] : 
                        (N149)? mem[711] : 
                        (N151)? mem[751] : 
                        (N153)? mem[791] : 
                        (N155)? mem[831] : 
                        (N157)? mem[871] : 
                        (N159)? mem[911] : 
                        (N161)? mem[951] : 
                        (N163)? mem[991] : 
                        (N165)? mem[1031] : 
                        (N167)? mem[1071] : 
                        (N169)? mem[1111] : 
                        (N171)? mem[1151] : 
                        (N173)? mem[1191] : 
                        (N175)? mem[1231] : 
                        (N177)? mem[1271] : 
                        (N116)? mem[1311] : 
                        (N118)? mem[1351] : 
                        (N120)? mem[1391] : 
                        (N122)? mem[1431] : 
                        (N124)? mem[1471] : 
                        (N126)? mem[1511] : 
                        (N128)? mem[1551] : 
                        (N130)? mem[1591] : 
                        (N132)? mem[1631] : 
                        (N134)? mem[1671] : 
                        (N136)? mem[1711] : 
                        (N138)? mem[1751] : 
                        (N140)? mem[1791] : 
                        (N142)? mem[1831] : 
                        (N144)? mem[1871] : 
                        (N146)? mem[1911] : 
                        (N148)? mem[1951] : 
                        (N150)? mem[1991] : 
                        (N152)? mem[2031] : 
                        (N154)? mem[2071] : 
                        (N156)? mem[2111] : 
                        (N158)? mem[2151] : 
                        (N160)? mem[2191] : 
                        (N162)? mem[2231] : 
                        (N164)? mem[2271] : 
                        (N166)? mem[2311] : 
                        (N168)? mem[2351] : 
                        (N170)? mem[2391] : 
                        (N172)? mem[2431] : 
                        (N174)? mem[2471] : 
                        (N176)? mem[2511] : 
                        (N178)? mem[2551] : 1'b0;
  assign data_out[30] = (N115)? mem[30] : 
                        (N117)? mem[70] : 
                        (N119)? mem[110] : 
                        (N121)? mem[150] : 
                        (N123)? mem[190] : 
                        (N125)? mem[230] : 
                        (N127)? mem[270] : 
                        (N129)? mem[310] : 
                        (N131)? mem[350] : 
                        (N133)? mem[390] : 
                        (N135)? mem[430] : 
                        (N137)? mem[470] : 
                        (N139)? mem[510] : 
                        (N141)? mem[550] : 
                        (N143)? mem[590] : 
                        (N145)? mem[630] : 
                        (N147)? mem[670] : 
                        (N149)? mem[710] : 
                        (N151)? mem[750] : 
                        (N153)? mem[790] : 
                        (N155)? mem[830] : 
                        (N157)? mem[870] : 
                        (N159)? mem[910] : 
                        (N161)? mem[950] : 
                        (N163)? mem[990] : 
                        (N165)? mem[1030] : 
                        (N167)? mem[1070] : 
                        (N169)? mem[1110] : 
                        (N171)? mem[1150] : 
                        (N173)? mem[1190] : 
                        (N175)? mem[1230] : 
                        (N177)? mem[1270] : 
                        (N116)? mem[1310] : 
                        (N118)? mem[1350] : 
                        (N120)? mem[1390] : 
                        (N122)? mem[1430] : 
                        (N124)? mem[1470] : 
                        (N126)? mem[1510] : 
                        (N128)? mem[1550] : 
                        (N130)? mem[1590] : 
                        (N132)? mem[1630] : 
                        (N134)? mem[1670] : 
                        (N136)? mem[1710] : 
                        (N138)? mem[1750] : 
                        (N140)? mem[1790] : 
                        (N142)? mem[1830] : 
                        (N144)? mem[1870] : 
                        (N146)? mem[1910] : 
                        (N148)? mem[1950] : 
                        (N150)? mem[1990] : 
                        (N152)? mem[2030] : 
                        (N154)? mem[2070] : 
                        (N156)? mem[2110] : 
                        (N158)? mem[2150] : 
                        (N160)? mem[2190] : 
                        (N162)? mem[2230] : 
                        (N164)? mem[2270] : 
                        (N166)? mem[2310] : 
                        (N168)? mem[2350] : 
                        (N170)? mem[2390] : 
                        (N172)? mem[2430] : 
                        (N174)? mem[2470] : 
                        (N176)? mem[2510] : 
                        (N178)? mem[2550] : 1'b0;
  assign data_out[29] = (N115)? mem[29] : 
                        (N117)? mem[69] : 
                        (N119)? mem[109] : 
                        (N121)? mem[149] : 
                        (N123)? mem[189] : 
                        (N125)? mem[229] : 
                        (N127)? mem[269] : 
                        (N129)? mem[309] : 
                        (N131)? mem[349] : 
                        (N133)? mem[389] : 
                        (N135)? mem[429] : 
                        (N137)? mem[469] : 
                        (N139)? mem[509] : 
                        (N141)? mem[549] : 
                        (N143)? mem[589] : 
                        (N145)? mem[629] : 
                        (N147)? mem[669] : 
                        (N149)? mem[709] : 
                        (N151)? mem[749] : 
                        (N153)? mem[789] : 
                        (N155)? mem[829] : 
                        (N157)? mem[869] : 
                        (N159)? mem[909] : 
                        (N161)? mem[949] : 
                        (N163)? mem[989] : 
                        (N165)? mem[1029] : 
                        (N167)? mem[1069] : 
                        (N169)? mem[1109] : 
                        (N171)? mem[1149] : 
                        (N173)? mem[1189] : 
                        (N175)? mem[1229] : 
                        (N177)? mem[1269] : 
                        (N116)? mem[1309] : 
                        (N118)? mem[1349] : 
                        (N120)? mem[1389] : 
                        (N122)? mem[1429] : 
                        (N124)? mem[1469] : 
                        (N126)? mem[1509] : 
                        (N128)? mem[1549] : 
                        (N130)? mem[1589] : 
                        (N132)? mem[1629] : 
                        (N134)? mem[1669] : 
                        (N136)? mem[1709] : 
                        (N138)? mem[1749] : 
                        (N140)? mem[1789] : 
                        (N142)? mem[1829] : 
                        (N144)? mem[1869] : 
                        (N146)? mem[1909] : 
                        (N148)? mem[1949] : 
                        (N150)? mem[1989] : 
                        (N152)? mem[2029] : 
                        (N154)? mem[2069] : 
                        (N156)? mem[2109] : 
                        (N158)? mem[2149] : 
                        (N160)? mem[2189] : 
                        (N162)? mem[2229] : 
                        (N164)? mem[2269] : 
                        (N166)? mem[2309] : 
                        (N168)? mem[2349] : 
                        (N170)? mem[2389] : 
                        (N172)? mem[2429] : 
                        (N174)? mem[2469] : 
                        (N176)? mem[2509] : 
                        (N178)? mem[2549] : 1'b0;
  assign data_out[28] = (N115)? mem[28] : 
                        (N117)? mem[68] : 
                        (N119)? mem[108] : 
                        (N121)? mem[148] : 
                        (N123)? mem[188] : 
                        (N125)? mem[228] : 
                        (N127)? mem[268] : 
                        (N129)? mem[308] : 
                        (N131)? mem[348] : 
                        (N133)? mem[388] : 
                        (N135)? mem[428] : 
                        (N137)? mem[468] : 
                        (N139)? mem[508] : 
                        (N141)? mem[548] : 
                        (N143)? mem[588] : 
                        (N145)? mem[628] : 
                        (N147)? mem[668] : 
                        (N149)? mem[708] : 
                        (N151)? mem[748] : 
                        (N153)? mem[788] : 
                        (N155)? mem[828] : 
                        (N157)? mem[868] : 
                        (N159)? mem[908] : 
                        (N161)? mem[948] : 
                        (N163)? mem[988] : 
                        (N165)? mem[1028] : 
                        (N167)? mem[1068] : 
                        (N169)? mem[1108] : 
                        (N171)? mem[1148] : 
                        (N173)? mem[1188] : 
                        (N175)? mem[1228] : 
                        (N177)? mem[1268] : 
                        (N116)? mem[1308] : 
                        (N118)? mem[1348] : 
                        (N120)? mem[1388] : 
                        (N122)? mem[1428] : 
                        (N124)? mem[1468] : 
                        (N126)? mem[1508] : 
                        (N128)? mem[1548] : 
                        (N130)? mem[1588] : 
                        (N132)? mem[1628] : 
                        (N134)? mem[1668] : 
                        (N136)? mem[1708] : 
                        (N138)? mem[1748] : 
                        (N140)? mem[1788] : 
                        (N142)? mem[1828] : 
                        (N144)? mem[1868] : 
                        (N146)? mem[1908] : 
                        (N148)? mem[1948] : 
                        (N150)? mem[1988] : 
                        (N152)? mem[2028] : 
                        (N154)? mem[2068] : 
                        (N156)? mem[2108] : 
                        (N158)? mem[2148] : 
                        (N160)? mem[2188] : 
                        (N162)? mem[2228] : 
                        (N164)? mem[2268] : 
                        (N166)? mem[2308] : 
                        (N168)? mem[2348] : 
                        (N170)? mem[2388] : 
                        (N172)? mem[2428] : 
                        (N174)? mem[2468] : 
                        (N176)? mem[2508] : 
                        (N178)? mem[2548] : 1'b0;
  assign data_out[27] = (N115)? mem[27] : 
                        (N117)? mem[67] : 
                        (N119)? mem[107] : 
                        (N121)? mem[147] : 
                        (N123)? mem[187] : 
                        (N125)? mem[227] : 
                        (N127)? mem[267] : 
                        (N129)? mem[307] : 
                        (N131)? mem[347] : 
                        (N133)? mem[387] : 
                        (N135)? mem[427] : 
                        (N137)? mem[467] : 
                        (N139)? mem[507] : 
                        (N141)? mem[547] : 
                        (N143)? mem[587] : 
                        (N145)? mem[627] : 
                        (N147)? mem[667] : 
                        (N149)? mem[707] : 
                        (N151)? mem[747] : 
                        (N153)? mem[787] : 
                        (N155)? mem[827] : 
                        (N157)? mem[867] : 
                        (N159)? mem[907] : 
                        (N161)? mem[947] : 
                        (N163)? mem[987] : 
                        (N165)? mem[1027] : 
                        (N167)? mem[1067] : 
                        (N169)? mem[1107] : 
                        (N171)? mem[1147] : 
                        (N173)? mem[1187] : 
                        (N175)? mem[1227] : 
                        (N177)? mem[1267] : 
                        (N116)? mem[1307] : 
                        (N118)? mem[1347] : 
                        (N120)? mem[1387] : 
                        (N122)? mem[1427] : 
                        (N124)? mem[1467] : 
                        (N126)? mem[1507] : 
                        (N128)? mem[1547] : 
                        (N130)? mem[1587] : 
                        (N132)? mem[1627] : 
                        (N134)? mem[1667] : 
                        (N136)? mem[1707] : 
                        (N138)? mem[1747] : 
                        (N140)? mem[1787] : 
                        (N142)? mem[1827] : 
                        (N144)? mem[1867] : 
                        (N146)? mem[1907] : 
                        (N148)? mem[1947] : 
                        (N150)? mem[1987] : 
                        (N152)? mem[2027] : 
                        (N154)? mem[2067] : 
                        (N156)? mem[2107] : 
                        (N158)? mem[2147] : 
                        (N160)? mem[2187] : 
                        (N162)? mem[2227] : 
                        (N164)? mem[2267] : 
                        (N166)? mem[2307] : 
                        (N168)? mem[2347] : 
                        (N170)? mem[2387] : 
                        (N172)? mem[2427] : 
                        (N174)? mem[2467] : 
                        (N176)? mem[2507] : 
                        (N178)? mem[2547] : 1'b0;
  assign data_out[26] = (N115)? mem[26] : 
                        (N117)? mem[66] : 
                        (N119)? mem[106] : 
                        (N121)? mem[146] : 
                        (N123)? mem[186] : 
                        (N125)? mem[226] : 
                        (N127)? mem[266] : 
                        (N129)? mem[306] : 
                        (N131)? mem[346] : 
                        (N133)? mem[386] : 
                        (N135)? mem[426] : 
                        (N137)? mem[466] : 
                        (N139)? mem[506] : 
                        (N141)? mem[546] : 
                        (N143)? mem[586] : 
                        (N145)? mem[626] : 
                        (N147)? mem[666] : 
                        (N149)? mem[706] : 
                        (N151)? mem[746] : 
                        (N153)? mem[786] : 
                        (N155)? mem[826] : 
                        (N157)? mem[866] : 
                        (N159)? mem[906] : 
                        (N161)? mem[946] : 
                        (N163)? mem[986] : 
                        (N165)? mem[1026] : 
                        (N167)? mem[1066] : 
                        (N169)? mem[1106] : 
                        (N171)? mem[1146] : 
                        (N173)? mem[1186] : 
                        (N175)? mem[1226] : 
                        (N177)? mem[1266] : 
                        (N116)? mem[1306] : 
                        (N118)? mem[1346] : 
                        (N120)? mem[1386] : 
                        (N122)? mem[1426] : 
                        (N124)? mem[1466] : 
                        (N126)? mem[1506] : 
                        (N128)? mem[1546] : 
                        (N130)? mem[1586] : 
                        (N132)? mem[1626] : 
                        (N134)? mem[1666] : 
                        (N136)? mem[1706] : 
                        (N138)? mem[1746] : 
                        (N140)? mem[1786] : 
                        (N142)? mem[1826] : 
                        (N144)? mem[1866] : 
                        (N146)? mem[1906] : 
                        (N148)? mem[1946] : 
                        (N150)? mem[1986] : 
                        (N152)? mem[2026] : 
                        (N154)? mem[2066] : 
                        (N156)? mem[2106] : 
                        (N158)? mem[2146] : 
                        (N160)? mem[2186] : 
                        (N162)? mem[2226] : 
                        (N164)? mem[2266] : 
                        (N166)? mem[2306] : 
                        (N168)? mem[2346] : 
                        (N170)? mem[2386] : 
                        (N172)? mem[2426] : 
                        (N174)? mem[2466] : 
                        (N176)? mem[2506] : 
                        (N178)? mem[2546] : 1'b0;
  assign data_out[25] = (N115)? mem[25] : 
                        (N117)? mem[65] : 
                        (N119)? mem[105] : 
                        (N121)? mem[145] : 
                        (N123)? mem[185] : 
                        (N125)? mem[225] : 
                        (N127)? mem[265] : 
                        (N129)? mem[305] : 
                        (N131)? mem[345] : 
                        (N133)? mem[385] : 
                        (N135)? mem[425] : 
                        (N137)? mem[465] : 
                        (N139)? mem[505] : 
                        (N141)? mem[545] : 
                        (N143)? mem[585] : 
                        (N145)? mem[625] : 
                        (N147)? mem[665] : 
                        (N149)? mem[705] : 
                        (N151)? mem[745] : 
                        (N153)? mem[785] : 
                        (N155)? mem[825] : 
                        (N157)? mem[865] : 
                        (N159)? mem[905] : 
                        (N161)? mem[945] : 
                        (N163)? mem[985] : 
                        (N165)? mem[1025] : 
                        (N167)? mem[1065] : 
                        (N169)? mem[1105] : 
                        (N171)? mem[1145] : 
                        (N173)? mem[1185] : 
                        (N175)? mem[1225] : 
                        (N177)? mem[1265] : 
                        (N116)? mem[1305] : 
                        (N118)? mem[1345] : 
                        (N120)? mem[1385] : 
                        (N122)? mem[1425] : 
                        (N124)? mem[1465] : 
                        (N126)? mem[1505] : 
                        (N128)? mem[1545] : 
                        (N130)? mem[1585] : 
                        (N132)? mem[1625] : 
                        (N134)? mem[1665] : 
                        (N136)? mem[1705] : 
                        (N138)? mem[1745] : 
                        (N140)? mem[1785] : 
                        (N142)? mem[1825] : 
                        (N144)? mem[1865] : 
                        (N146)? mem[1905] : 
                        (N148)? mem[1945] : 
                        (N150)? mem[1985] : 
                        (N152)? mem[2025] : 
                        (N154)? mem[2065] : 
                        (N156)? mem[2105] : 
                        (N158)? mem[2145] : 
                        (N160)? mem[2185] : 
                        (N162)? mem[2225] : 
                        (N164)? mem[2265] : 
                        (N166)? mem[2305] : 
                        (N168)? mem[2345] : 
                        (N170)? mem[2385] : 
                        (N172)? mem[2425] : 
                        (N174)? mem[2465] : 
                        (N176)? mem[2505] : 
                        (N178)? mem[2545] : 1'b0;
  assign data_out[24] = (N115)? mem[24] : 
                        (N117)? mem[64] : 
                        (N119)? mem[104] : 
                        (N121)? mem[144] : 
                        (N123)? mem[184] : 
                        (N125)? mem[224] : 
                        (N127)? mem[264] : 
                        (N129)? mem[304] : 
                        (N131)? mem[344] : 
                        (N133)? mem[384] : 
                        (N135)? mem[424] : 
                        (N137)? mem[464] : 
                        (N139)? mem[504] : 
                        (N141)? mem[544] : 
                        (N143)? mem[584] : 
                        (N145)? mem[624] : 
                        (N147)? mem[664] : 
                        (N149)? mem[704] : 
                        (N151)? mem[744] : 
                        (N153)? mem[784] : 
                        (N155)? mem[824] : 
                        (N157)? mem[864] : 
                        (N159)? mem[904] : 
                        (N161)? mem[944] : 
                        (N163)? mem[984] : 
                        (N165)? mem[1024] : 
                        (N167)? mem[1064] : 
                        (N169)? mem[1104] : 
                        (N171)? mem[1144] : 
                        (N173)? mem[1184] : 
                        (N175)? mem[1224] : 
                        (N177)? mem[1264] : 
                        (N116)? mem[1304] : 
                        (N118)? mem[1344] : 
                        (N120)? mem[1384] : 
                        (N122)? mem[1424] : 
                        (N124)? mem[1464] : 
                        (N126)? mem[1504] : 
                        (N128)? mem[1544] : 
                        (N130)? mem[1584] : 
                        (N132)? mem[1624] : 
                        (N134)? mem[1664] : 
                        (N136)? mem[1704] : 
                        (N138)? mem[1744] : 
                        (N140)? mem[1784] : 
                        (N142)? mem[1824] : 
                        (N144)? mem[1864] : 
                        (N146)? mem[1904] : 
                        (N148)? mem[1944] : 
                        (N150)? mem[1984] : 
                        (N152)? mem[2024] : 
                        (N154)? mem[2064] : 
                        (N156)? mem[2104] : 
                        (N158)? mem[2144] : 
                        (N160)? mem[2184] : 
                        (N162)? mem[2224] : 
                        (N164)? mem[2264] : 
                        (N166)? mem[2304] : 
                        (N168)? mem[2344] : 
                        (N170)? mem[2384] : 
                        (N172)? mem[2424] : 
                        (N174)? mem[2464] : 
                        (N176)? mem[2504] : 
                        (N178)? mem[2544] : 1'b0;
  assign data_out[23] = (N115)? mem[23] : 
                        (N117)? mem[63] : 
                        (N119)? mem[103] : 
                        (N121)? mem[143] : 
                        (N123)? mem[183] : 
                        (N125)? mem[223] : 
                        (N127)? mem[263] : 
                        (N129)? mem[303] : 
                        (N131)? mem[343] : 
                        (N133)? mem[383] : 
                        (N135)? mem[423] : 
                        (N137)? mem[463] : 
                        (N139)? mem[503] : 
                        (N141)? mem[543] : 
                        (N143)? mem[583] : 
                        (N145)? mem[623] : 
                        (N147)? mem[663] : 
                        (N149)? mem[703] : 
                        (N151)? mem[743] : 
                        (N153)? mem[783] : 
                        (N155)? mem[823] : 
                        (N157)? mem[863] : 
                        (N159)? mem[903] : 
                        (N161)? mem[943] : 
                        (N163)? mem[983] : 
                        (N165)? mem[1023] : 
                        (N167)? mem[1063] : 
                        (N169)? mem[1103] : 
                        (N171)? mem[1143] : 
                        (N173)? mem[1183] : 
                        (N175)? mem[1223] : 
                        (N177)? mem[1263] : 
                        (N116)? mem[1303] : 
                        (N118)? mem[1343] : 
                        (N120)? mem[1383] : 
                        (N122)? mem[1423] : 
                        (N124)? mem[1463] : 
                        (N126)? mem[1503] : 
                        (N128)? mem[1543] : 
                        (N130)? mem[1583] : 
                        (N132)? mem[1623] : 
                        (N134)? mem[1663] : 
                        (N136)? mem[1703] : 
                        (N138)? mem[1743] : 
                        (N140)? mem[1783] : 
                        (N142)? mem[1823] : 
                        (N144)? mem[1863] : 
                        (N146)? mem[1903] : 
                        (N148)? mem[1943] : 
                        (N150)? mem[1983] : 
                        (N152)? mem[2023] : 
                        (N154)? mem[2063] : 
                        (N156)? mem[2103] : 
                        (N158)? mem[2143] : 
                        (N160)? mem[2183] : 
                        (N162)? mem[2223] : 
                        (N164)? mem[2263] : 
                        (N166)? mem[2303] : 
                        (N168)? mem[2343] : 
                        (N170)? mem[2383] : 
                        (N172)? mem[2423] : 
                        (N174)? mem[2463] : 
                        (N176)? mem[2503] : 
                        (N178)? mem[2543] : 1'b0;
  assign data_out[22] = (N115)? mem[22] : 
                        (N117)? mem[62] : 
                        (N119)? mem[102] : 
                        (N121)? mem[142] : 
                        (N123)? mem[182] : 
                        (N125)? mem[222] : 
                        (N127)? mem[262] : 
                        (N129)? mem[302] : 
                        (N131)? mem[342] : 
                        (N133)? mem[382] : 
                        (N135)? mem[422] : 
                        (N137)? mem[462] : 
                        (N139)? mem[502] : 
                        (N141)? mem[542] : 
                        (N143)? mem[582] : 
                        (N145)? mem[622] : 
                        (N147)? mem[662] : 
                        (N149)? mem[702] : 
                        (N151)? mem[742] : 
                        (N153)? mem[782] : 
                        (N155)? mem[822] : 
                        (N157)? mem[862] : 
                        (N159)? mem[902] : 
                        (N161)? mem[942] : 
                        (N163)? mem[982] : 
                        (N165)? mem[1022] : 
                        (N167)? mem[1062] : 
                        (N169)? mem[1102] : 
                        (N171)? mem[1142] : 
                        (N173)? mem[1182] : 
                        (N175)? mem[1222] : 
                        (N177)? mem[1262] : 
                        (N116)? mem[1302] : 
                        (N118)? mem[1342] : 
                        (N120)? mem[1382] : 
                        (N122)? mem[1422] : 
                        (N124)? mem[1462] : 
                        (N126)? mem[1502] : 
                        (N128)? mem[1542] : 
                        (N130)? mem[1582] : 
                        (N132)? mem[1622] : 
                        (N134)? mem[1662] : 
                        (N136)? mem[1702] : 
                        (N138)? mem[1742] : 
                        (N140)? mem[1782] : 
                        (N142)? mem[1822] : 
                        (N144)? mem[1862] : 
                        (N146)? mem[1902] : 
                        (N148)? mem[1942] : 
                        (N150)? mem[1982] : 
                        (N152)? mem[2022] : 
                        (N154)? mem[2062] : 
                        (N156)? mem[2102] : 
                        (N158)? mem[2142] : 
                        (N160)? mem[2182] : 
                        (N162)? mem[2222] : 
                        (N164)? mem[2262] : 
                        (N166)? mem[2302] : 
                        (N168)? mem[2342] : 
                        (N170)? mem[2382] : 
                        (N172)? mem[2422] : 
                        (N174)? mem[2462] : 
                        (N176)? mem[2502] : 
                        (N178)? mem[2542] : 1'b0;
  assign data_out[21] = (N115)? mem[21] : 
                        (N117)? mem[61] : 
                        (N119)? mem[101] : 
                        (N121)? mem[141] : 
                        (N123)? mem[181] : 
                        (N125)? mem[221] : 
                        (N127)? mem[261] : 
                        (N129)? mem[301] : 
                        (N131)? mem[341] : 
                        (N133)? mem[381] : 
                        (N135)? mem[421] : 
                        (N137)? mem[461] : 
                        (N139)? mem[501] : 
                        (N141)? mem[541] : 
                        (N143)? mem[581] : 
                        (N145)? mem[621] : 
                        (N147)? mem[661] : 
                        (N149)? mem[701] : 
                        (N151)? mem[741] : 
                        (N153)? mem[781] : 
                        (N155)? mem[821] : 
                        (N157)? mem[861] : 
                        (N159)? mem[901] : 
                        (N161)? mem[941] : 
                        (N163)? mem[981] : 
                        (N165)? mem[1021] : 
                        (N167)? mem[1061] : 
                        (N169)? mem[1101] : 
                        (N171)? mem[1141] : 
                        (N173)? mem[1181] : 
                        (N175)? mem[1221] : 
                        (N177)? mem[1261] : 
                        (N116)? mem[1301] : 
                        (N118)? mem[1341] : 
                        (N120)? mem[1381] : 
                        (N122)? mem[1421] : 
                        (N124)? mem[1461] : 
                        (N126)? mem[1501] : 
                        (N128)? mem[1541] : 
                        (N130)? mem[1581] : 
                        (N132)? mem[1621] : 
                        (N134)? mem[1661] : 
                        (N136)? mem[1701] : 
                        (N138)? mem[1741] : 
                        (N140)? mem[1781] : 
                        (N142)? mem[1821] : 
                        (N144)? mem[1861] : 
                        (N146)? mem[1901] : 
                        (N148)? mem[1941] : 
                        (N150)? mem[1981] : 
                        (N152)? mem[2021] : 
                        (N154)? mem[2061] : 
                        (N156)? mem[2101] : 
                        (N158)? mem[2141] : 
                        (N160)? mem[2181] : 
                        (N162)? mem[2221] : 
                        (N164)? mem[2261] : 
                        (N166)? mem[2301] : 
                        (N168)? mem[2341] : 
                        (N170)? mem[2381] : 
                        (N172)? mem[2421] : 
                        (N174)? mem[2461] : 
                        (N176)? mem[2501] : 
                        (N178)? mem[2541] : 1'b0;
  assign data_out[20] = (N115)? mem[20] : 
                        (N117)? mem[60] : 
                        (N119)? mem[100] : 
                        (N121)? mem[140] : 
                        (N123)? mem[180] : 
                        (N125)? mem[220] : 
                        (N127)? mem[260] : 
                        (N129)? mem[300] : 
                        (N131)? mem[340] : 
                        (N133)? mem[380] : 
                        (N135)? mem[420] : 
                        (N137)? mem[460] : 
                        (N139)? mem[500] : 
                        (N141)? mem[540] : 
                        (N143)? mem[580] : 
                        (N145)? mem[620] : 
                        (N147)? mem[660] : 
                        (N149)? mem[700] : 
                        (N151)? mem[740] : 
                        (N153)? mem[780] : 
                        (N155)? mem[820] : 
                        (N157)? mem[860] : 
                        (N159)? mem[900] : 
                        (N161)? mem[940] : 
                        (N163)? mem[980] : 
                        (N165)? mem[1020] : 
                        (N167)? mem[1060] : 
                        (N169)? mem[1100] : 
                        (N171)? mem[1140] : 
                        (N173)? mem[1180] : 
                        (N175)? mem[1220] : 
                        (N177)? mem[1260] : 
                        (N116)? mem[1300] : 
                        (N118)? mem[1340] : 
                        (N120)? mem[1380] : 
                        (N122)? mem[1420] : 
                        (N124)? mem[1460] : 
                        (N126)? mem[1500] : 
                        (N128)? mem[1540] : 
                        (N130)? mem[1580] : 
                        (N132)? mem[1620] : 
                        (N134)? mem[1660] : 
                        (N136)? mem[1700] : 
                        (N138)? mem[1740] : 
                        (N140)? mem[1780] : 
                        (N142)? mem[1820] : 
                        (N144)? mem[1860] : 
                        (N146)? mem[1900] : 
                        (N148)? mem[1940] : 
                        (N150)? mem[1980] : 
                        (N152)? mem[2020] : 
                        (N154)? mem[2060] : 
                        (N156)? mem[2100] : 
                        (N158)? mem[2140] : 
                        (N160)? mem[2180] : 
                        (N162)? mem[2220] : 
                        (N164)? mem[2260] : 
                        (N166)? mem[2300] : 
                        (N168)? mem[2340] : 
                        (N170)? mem[2380] : 
                        (N172)? mem[2420] : 
                        (N174)? mem[2460] : 
                        (N176)? mem[2500] : 
                        (N178)? mem[2540] : 1'b0;
  assign data_out[19] = (N115)? mem[19] : 
                        (N117)? mem[59] : 
                        (N119)? mem[99] : 
                        (N121)? mem[139] : 
                        (N123)? mem[179] : 
                        (N125)? mem[219] : 
                        (N127)? mem[259] : 
                        (N129)? mem[299] : 
                        (N131)? mem[339] : 
                        (N133)? mem[379] : 
                        (N135)? mem[419] : 
                        (N137)? mem[459] : 
                        (N139)? mem[499] : 
                        (N141)? mem[539] : 
                        (N143)? mem[579] : 
                        (N145)? mem[619] : 
                        (N147)? mem[659] : 
                        (N149)? mem[699] : 
                        (N151)? mem[739] : 
                        (N153)? mem[779] : 
                        (N155)? mem[819] : 
                        (N157)? mem[859] : 
                        (N159)? mem[899] : 
                        (N161)? mem[939] : 
                        (N163)? mem[979] : 
                        (N165)? mem[1019] : 
                        (N167)? mem[1059] : 
                        (N169)? mem[1099] : 
                        (N171)? mem[1139] : 
                        (N173)? mem[1179] : 
                        (N175)? mem[1219] : 
                        (N177)? mem[1259] : 
                        (N116)? mem[1299] : 
                        (N118)? mem[1339] : 
                        (N120)? mem[1379] : 
                        (N122)? mem[1419] : 
                        (N124)? mem[1459] : 
                        (N126)? mem[1499] : 
                        (N128)? mem[1539] : 
                        (N130)? mem[1579] : 
                        (N132)? mem[1619] : 
                        (N134)? mem[1659] : 
                        (N136)? mem[1699] : 
                        (N138)? mem[1739] : 
                        (N140)? mem[1779] : 
                        (N142)? mem[1819] : 
                        (N144)? mem[1859] : 
                        (N146)? mem[1899] : 
                        (N148)? mem[1939] : 
                        (N150)? mem[1979] : 
                        (N152)? mem[2019] : 
                        (N154)? mem[2059] : 
                        (N156)? mem[2099] : 
                        (N158)? mem[2139] : 
                        (N160)? mem[2179] : 
                        (N162)? mem[2219] : 
                        (N164)? mem[2259] : 
                        (N166)? mem[2299] : 
                        (N168)? mem[2339] : 
                        (N170)? mem[2379] : 
                        (N172)? mem[2419] : 
                        (N174)? mem[2459] : 
                        (N176)? mem[2499] : 
                        (N178)? mem[2539] : 1'b0;
  assign data_out[18] = (N115)? mem[18] : 
                        (N117)? mem[58] : 
                        (N119)? mem[98] : 
                        (N121)? mem[138] : 
                        (N123)? mem[178] : 
                        (N125)? mem[218] : 
                        (N127)? mem[258] : 
                        (N129)? mem[298] : 
                        (N131)? mem[338] : 
                        (N133)? mem[378] : 
                        (N135)? mem[418] : 
                        (N137)? mem[458] : 
                        (N139)? mem[498] : 
                        (N141)? mem[538] : 
                        (N143)? mem[578] : 
                        (N145)? mem[618] : 
                        (N147)? mem[658] : 
                        (N149)? mem[698] : 
                        (N151)? mem[738] : 
                        (N153)? mem[778] : 
                        (N155)? mem[818] : 
                        (N157)? mem[858] : 
                        (N159)? mem[898] : 
                        (N161)? mem[938] : 
                        (N163)? mem[978] : 
                        (N165)? mem[1018] : 
                        (N167)? mem[1058] : 
                        (N169)? mem[1098] : 
                        (N171)? mem[1138] : 
                        (N173)? mem[1178] : 
                        (N175)? mem[1218] : 
                        (N177)? mem[1258] : 
                        (N116)? mem[1298] : 
                        (N118)? mem[1338] : 
                        (N120)? mem[1378] : 
                        (N122)? mem[1418] : 
                        (N124)? mem[1458] : 
                        (N126)? mem[1498] : 
                        (N128)? mem[1538] : 
                        (N130)? mem[1578] : 
                        (N132)? mem[1618] : 
                        (N134)? mem[1658] : 
                        (N136)? mem[1698] : 
                        (N138)? mem[1738] : 
                        (N140)? mem[1778] : 
                        (N142)? mem[1818] : 
                        (N144)? mem[1858] : 
                        (N146)? mem[1898] : 
                        (N148)? mem[1938] : 
                        (N150)? mem[1978] : 
                        (N152)? mem[2018] : 
                        (N154)? mem[2058] : 
                        (N156)? mem[2098] : 
                        (N158)? mem[2138] : 
                        (N160)? mem[2178] : 
                        (N162)? mem[2218] : 
                        (N164)? mem[2258] : 
                        (N166)? mem[2298] : 
                        (N168)? mem[2338] : 
                        (N170)? mem[2378] : 
                        (N172)? mem[2418] : 
                        (N174)? mem[2458] : 
                        (N176)? mem[2498] : 
                        (N178)? mem[2538] : 1'b0;
  assign data_out[17] = (N115)? mem[17] : 
                        (N117)? mem[57] : 
                        (N119)? mem[97] : 
                        (N121)? mem[137] : 
                        (N123)? mem[177] : 
                        (N125)? mem[217] : 
                        (N127)? mem[257] : 
                        (N129)? mem[297] : 
                        (N131)? mem[337] : 
                        (N133)? mem[377] : 
                        (N135)? mem[417] : 
                        (N137)? mem[457] : 
                        (N139)? mem[497] : 
                        (N141)? mem[537] : 
                        (N143)? mem[577] : 
                        (N145)? mem[617] : 
                        (N147)? mem[657] : 
                        (N149)? mem[697] : 
                        (N151)? mem[737] : 
                        (N153)? mem[777] : 
                        (N155)? mem[817] : 
                        (N157)? mem[857] : 
                        (N159)? mem[897] : 
                        (N161)? mem[937] : 
                        (N163)? mem[977] : 
                        (N165)? mem[1017] : 
                        (N167)? mem[1057] : 
                        (N169)? mem[1097] : 
                        (N171)? mem[1137] : 
                        (N173)? mem[1177] : 
                        (N175)? mem[1217] : 
                        (N177)? mem[1257] : 
                        (N116)? mem[1297] : 
                        (N118)? mem[1337] : 
                        (N120)? mem[1377] : 
                        (N122)? mem[1417] : 
                        (N124)? mem[1457] : 
                        (N126)? mem[1497] : 
                        (N128)? mem[1537] : 
                        (N130)? mem[1577] : 
                        (N132)? mem[1617] : 
                        (N134)? mem[1657] : 
                        (N136)? mem[1697] : 
                        (N138)? mem[1737] : 
                        (N140)? mem[1777] : 
                        (N142)? mem[1817] : 
                        (N144)? mem[1857] : 
                        (N146)? mem[1897] : 
                        (N148)? mem[1937] : 
                        (N150)? mem[1977] : 
                        (N152)? mem[2017] : 
                        (N154)? mem[2057] : 
                        (N156)? mem[2097] : 
                        (N158)? mem[2137] : 
                        (N160)? mem[2177] : 
                        (N162)? mem[2217] : 
                        (N164)? mem[2257] : 
                        (N166)? mem[2297] : 
                        (N168)? mem[2337] : 
                        (N170)? mem[2377] : 
                        (N172)? mem[2417] : 
                        (N174)? mem[2457] : 
                        (N176)? mem[2497] : 
                        (N178)? mem[2537] : 1'b0;
  assign data_out[16] = (N115)? mem[16] : 
                        (N117)? mem[56] : 
                        (N119)? mem[96] : 
                        (N121)? mem[136] : 
                        (N123)? mem[176] : 
                        (N125)? mem[216] : 
                        (N127)? mem[256] : 
                        (N129)? mem[296] : 
                        (N131)? mem[336] : 
                        (N133)? mem[376] : 
                        (N135)? mem[416] : 
                        (N137)? mem[456] : 
                        (N139)? mem[496] : 
                        (N141)? mem[536] : 
                        (N143)? mem[576] : 
                        (N145)? mem[616] : 
                        (N147)? mem[656] : 
                        (N149)? mem[696] : 
                        (N151)? mem[736] : 
                        (N153)? mem[776] : 
                        (N155)? mem[816] : 
                        (N157)? mem[856] : 
                        (N159)? mem[896] : 
                        (N161)? mem[936] : 
                        (N163)? mem[976] : 
                        (N165)? mem[1016] : 
                        (N167)? mem[1056] : 
                        (N169)? mem[1096] : 
                        (N171)? mem[1136] : 
                        (N173)? mem[1176] : 
                        (N175)? mem[1216] : 
                        (N177)? mem[1256] : 
                        (N116)? mem[1296] : 
                        (N118)? mem[1336] : 
                        (N120)? mem[1376] : 
                        (N122)? mem[1416] : 
                        (N124)? mem[1456] : 
                        (N126)? mem[1496] : 
                        (N128)? mem[1536] : 
                        (N130)? mem[1576] : 
                        (N132)? mem[1616] : 
                        (N134)? mem[1656] : 
                        (N136)? mem[1696] : 
                        (N138)? mem[1736] : 
                        (N140)? mem[1776] : 
                        (N142)? mem[1816] : 
                        (N144)? mem[1856] : 
                        (N146)? mem[1896] : 
                        (N148)? mem[1936] : 
                        (N150)? mem[1976] : 
                        (N152)? mem[2016] : 
                        (N154)? mem[2056] : 
                        (N156)? mem[2096] : 
                        (N158)? mem[2136] : 
                        (N160)? mem[2176] : 
                        (N162)? mem[2216] : 
                        (N164)? mem[2256] : 
                        (N166)? mem[2296] : 
                        (N168)? mem[2336] : 
                        (N170)? mem[2376] : 
                        (N172)? mem[2416] : 
                        (N174)? mem[2456] : 
                        (N176)? mem[2496] : 
                        (N178)? mem[2536] : 1'b0;
  assign data_out[15] = (N115)? mem[15] : 
                        (N117)? mem[55] : 
                        (N119)? mem[95] : 
                        (N121)? mem[135] : 
                        (N123)? mem[175] : 
                        (N125)? mem[215] : 
                        (N127)? mem[255] : 
                        (N129)? mem[295] : 
                        (N131)? mem[335] : 
                        (N133)? mem[375] : 
                        (N135)? mem[415] : 
                        (N137)? mem[455] : 
                        (N139)? mem[495] : 
                        (N141)? mem[535] : 
                        (N143)? mem[575] : 
                        (N145)? mem[615] : 
                        (N147)? mem[655] : 
                        (N149)? mem[695] : 
                        (N151)? mem[735] : 
                        (N153)? mem[775] : 
                        (N155)? mem[815] : 
                        (N157)? mem[855] : 
                        (N159)? mem[895] : 
                        (N161)? mem[935] : 
                        (N163)? mem[975] : 
                        (N165)? mem[1015] : 
                        (N167)? mem[1055] : 
                        (N169)? mem[1095] : 
                        (N171)? mem[1135] : 
                        (N173)? mem[1175] : 
                        (N175)? mem[1215] : 
                        (N177)? mem[1255] : 
                        (N116)? mem[1295] : 
                        (N118)? mem[1335] : 
                        (N120)? mem[1375] : 
                        (N122)? mem[1415] : 
                        (N124)? mem[1455] : 
                        (N126)? mem[1495] : 
                        (N128)? mem[1535] : 
                        (N130)? mem[1575] : 
                        (N132)? mem[1615] : 
                        (N134)? mem[1655] : 
                        (N136)? mem[1695] : 
                        (N138)? mem[1735] : 
                        (N140)? mem[1775] : 
                        (N142)? mem[1815] : 
                        (N144)? mem[1855] : 
                        (N146)? mem[1895] : 
                        (N148)? mem[1935] : 
                        (N150)? mem[1975] : 
                        (N152)? mem[2015] : 
                        (N154)? mem[2055] : 
                        (N156)? mem[2095] : 
                        (N158)? mem[2135] : 
                        (N160)? mem[2175] : 
                        (N162)? mem[2215] : 
                        (N164)? mem[2255] : 
                        (N166)? mem[2295] : 
                        (N168)? mem[2335] : 
                        (N170)? mem[2375] : 
                        (N172)? mem[2415] : 
                        (N174)? mem[2455] : 
                        (N176)? mem[2495] : 
                        (N178)? mem[2535] : 1'b0;
  assign data_out[14] = (N115)? mem[14] : 
                        (N117)? mem[54] : 
                        (N119)? mem[94] : 
                        (N121)? mem[134] : 
                        (N123)? mem[174] : 
                        (N125)? mem[214] : 
                        (N127)? mem[254] : 
                        (N129)? mem[294] : 
                        (N131)? mem[334] : 
                        (N133)? mem[374] : 
                        (N135)? mem[414] : 
                        (N137)? mem[454] : 
                        (N139)? mem[494] : 
                        (N141)? mem[534] : 
                        (N143)? mem[574] : 
                        (N145)? mem[614] : 
                        (N147)? mem[654] : 
                        (N149)? mem[694] : 
                        (N151)? mem[734] : 
                        (N153)? mem[774] : 
                        (N155)? mem[814] : 
                        (N157)? mem[854] : 
                        (N159)? mem[894] : 
                        (N161)? mem[934] : 
                        (N163)? mem[974] : 
                        (N165)? mem[1014] : 
                        (N167)? mem[1054] : 
                        (N169)? mem[1094] : 
                        (N171)? mem[1134] : 
                        (N173)? mem[1174] : 
                        (N175)? mem[1214] : 
                        (N177)? mem[1254] : 
                        (N116)? mem[1294] : 
                        (N118)? mem[1334] : 
                        (N120)? mem[1374] : 
                        (N122)? mem[1414] : 
                        (N124)? mem[1454] : 
                        (N126)? mem[1494] : 
                        (N128)? mem[1534] : 
                        (N130)? mem[1574] : 
                        (N132)? mem[1614] : 
                        (N134)? mem[1654] : 
                        (N136)? mem[1694] : 
                        (N138)? mem[1734] : 
                        (N140)? mem[1774] : 
                        (N142)? mem[1814] : 
                        (N144)? mem[1854] : 
                        (N146)? mem[1894] : 
                        (N148)? mem[1934] : 
                        (N150)? mem[1974] : 
                        (N152)? mem[2014] : 
                        (N154)? mem[2054] : 
                        (N156)? mem[2094] : 
                        (N158)? mem[2134] : 
                        (N160)? mem[2174] : 
                        (N162)? mem[2214] : 
                        (N164)? mem[2254] : 
                        (N166)? mem[2294] : 
                        (N168)? mem[2334] : 
                        (N170)? mem[2374] : 
                        (N172)? mem[2414] : 
                        (N174)? mem[2454] : 
                        (N176)? mem[2494] : 
                        (N178)? mem[2534] : 1'b0;
  assign data_out[13] = (N115)? mem[13] : 
                        (N117)? mem[53] : 
                        (N119)? mem[93] : 
                        (N121)? mem[133] : 
                        (N123)? mem[173] : 
                        (N125)? mem[213] : 
                        (N127)? mem[253] : 
                        (N129)? mem[293] : 
                        (N131)? mem[333] : 
                        (N133)? mem[373] : 
                        (N135)? mem[413] : 
                        (N137)? mem[453] : 
                        (N139)? mem[493] : 
                        (N141)? mem[533] : 
                        (N143)? mem[573] : 
                        (N145)? mem[613] : 
                        (N147)? mem[653] : 
                        (N149)? mem[693] : 
                        (N151)? mem[733] : 
                        (N153)? mem[773] : 
                        (N155)? mem[813] : 
                        (N157)? mem[853] : 
                        (N159)? mem[893] : 
                        (N161)? mem[933] : 
                        (N163)? mem[973] : 
                        (N165)? mem[1013] : 
                        (N167)? mem[1053] : 
                        (N169)? mem[1093] : 
                        (N171)? mem[1133] : 
                        (N173)? mem[1173] : 
                        (N175)? mem[1213] : 
                        (N177)? mem[1253] : 
                        (N116)? mem[1293] : 
                        (N118)? mem[1333] : 
                        (N120)? mem[1373] : 
                        (N122)? mem[1413] : 
                        (N124)? mem[1453] : 
                        (N126)? mem[1493] : 
                        (N128)? mem[1533] : 
                        (N130)? mem[1573] : 
                        (N132)? mem[1613] : 
                        (N134)? mem[1653] : 
                        (N136)? mem[1693] : 
                        (N138)? mem[1733] : 
                        (N140)? mem[1773] : 
                        (N142)? mem[1813] : 
                        (N144)? mem[1853] : 
                        (N146)? mem[1893] : 
                        (N148)? mem[1933] : 
                        (N150)? mem[1973] : 
                        (N152)? mem[2013] : 
                        (N154)? mem[2053] : 
                        (N156)? mem[2093] : 
                        (N158)? mem[2133] : 
                        (N160)? mem[2173] : 
                        (N162)? mem[2213] : 
                        (N164)? mem[2253] : 
                        (N166)? mem[2293] : 
                        (N168)? mem[2333] : 
                        (N170)? mem[2373] : 
                        (N172)? mem[2413] : 
                        (N174)? mem[2453] : 
                        (N176)? mem[2493] : 
                        (N178)? mem[2533] : 1'b0;
  assign data_out[12] = (N115)? mem[12] : 
                        (N117)? mem[52] : 
                        (N119)? mem[92] : 
                        (N121)? mem[132] : 
                        (N123)? mem[172] : 
                        (N125)? mem[212] : 
                        (N127)? mem[252] : 
                        (N129)? mem[292] : 
                        (N131)? mem[332] : 
                        (N133)? mem[372] : 
                        (N135)? mem[412] : 
                        (N137)? mem[452] : 
                        (N139)? mem[492] : 
                        (N141)? mem[532] : 
                        (N143)? mem[572] : 
                        (N145)? mem[612] : 
                        (N147)? mem[652] : 
                        (N149)? mem[692] : 
                        (N151)? mem[732] : 
                        (N153)? mem[772] : 
                        (N155)? mem[812] : 
                        (N157)? mem[852] : 
                        (N159)? mem[892] : 
                        (N161)? mem[932] : 
                        (N163)? mem[972] : 
                        (N165)? mem[1012] : 
                        (N167)? mem[1052] : 
                        (N169)? mem[1092] : 
                        (N171)? mem[1132] : 
                        (N173)? mem[1172] : 
                        (N175)? mem[1212] : 
                        (N177)? mem[1252] : 
                        (N116)? mem[1292] : 
                        (N118)? mem[1332] : 
                        (N120)? mem[1372] : 
                        (N122)? mem[1412] : 
                        (N124)? mem[1452] : 
                        (N126)? mem[1492] : 
                        (N128)? mem[1532] : 
                        (N130)? mem[1572] : 
                        (N132)? mem[1612] : 
                        (N134)? mem[1652] : 
                        (N136)? mem[1692] : 
                        (N138)? mem[1732] : 
                        (N140)? mem[1772] : 
                        (N142)? mem[1812] : 
                        (N144)? mem[1852] : 
                        (N146)? mem[1892] : 
                        (N148)? mem[1932] : 
                        (N150)? mem[1972] : 
                        (N152)? mem[2012] : 
                        (N154)? mem[2052] : 
                        (N156)? mem[2092] : 
                        (N158)? mem[2132] : 
                        (N160)? mem[2172] : 
                        (N162)? mem[2212] : 
                        (N164)? mem[2252] : 
                        (N166)? mem[2292] : 
                        (N168)? mem[2332] : 
                        (N170)? mem[2372] : 
                        (N172)? mem[2412] : 
                        (N174)? mem[2452] : 
                        (N176)? mem[2492] : 
                        (N178)? mem[2532] : 1'b0;
  assign data_out[11] = (N115)? mem[11] : 
                        (N117)? mem[51] : 
                        (N119)? mem[91] : 
                        (N121)? mem[131] : 
                        (N123)? mem[171] : 
                        (N125)? mem[211] : 
                        (N127)? mem[251] : 
                        (N129)? mem[291] : 
                        (N131)? mem[331] : 
                        (N133)? mem[371] : 
                        (N135)? mem[411] : 
                        (N137)? mem[451] : 
                        (N139)? mem[491] : 
                        (N141)? mem[531] : 
                        (N143)? mem[571] : 
                        (N145)? mem[611] : 
                        (N147)? mem[651] : 
                        (N149)? mem[691] : 
                        (N151)? mem[731] : 
                        (N153)? mem[771] : 
                        (N155)? mem[811] : 
                        (N157)? mem[851] : 
                        (N159)? mem[891] : 
                        (N161)? mem[931] : 
                        (N163)? mem[971] : 
                        (N165)? mem[1011] : 
                        (N167)? mem[1051] : 
                        (N169)? mem[1091] : 
                        (N171)? mem[1131] : 
                        (N173)? mem[1171] : 
                        (N175)? mem[1211] : 
                        (N177)? mem[1251] : 
                        (N116)? mem[1291] : 
                        (N118)? mem[1331] : 
                        (N120)? mem[1371] : 
                        (N122)? mem[1411] : 
                        (N124)? mem[1451] : 
                        (N126)? mem[1491] : 
                        (N128)? mem[1531] : 
                        (N130)? mem[1571] : 
                        (N132)? mem[1611] : 
                        (N134)? mem[1651] : 
                        (N136)? mem[1691] : 
                        (N138)? mem[1731] : 
                        (N140)? mem[1771] : 
                        (N142)? mem[1811] : 
                        (N144)? mem[1851] : 
                        (N146)? mem[1891] : 
                        (N148)? mem[1931] : 
                        (N150)? mem[1971] : 
                        (N152)? mem[2011] : 
                        (N154)? mem[2051] : 
                        (N156)? mem[2091] : 
                        (N158)? mem[2131] : 
                        (N160)? mem[2171] : 
                        (N162)? mem[2211] : 
                        (N164)? mem[2251] : 
                        (N166)? mem[2291] : 
                        (N168)? mem[2331] : 
                        (N170)? mem[2371] : 
                        (N172)? mem[2411] : 
                        (N174)? mem[2451] : 
                        (N176)? mem[2491] : 
                        (N178)? mem[2531] : 1'b0;
  assign data_out[10] = (N115)? mem[10] : 
                        (N117)? mem[50] : 
                        (N119)? mem[90] : 
                        (N121)? mem[130] : 
                        (N123)? mem[170] : 
                        (N125)? mem[210] : 
                        (N127)? mem[250] : 
                        (N129)? mem[290] : 
                        (N131)? mem[330] : 
                        (N133)? mem[370] : 
                        (N135)? mem[410] : 
                        (N137)? mem[450] : 
                        (N139)? mem[490] : 
                        (N141)? mem[530] : 
                        (N143)? mem[570] : 
                        (N145)? mem[610] : 
                        (N147)? mem[650] : 
                        (N149)? mem[690] : 
                        (N151)? mem[730] : 
                        (N153)? mem[770] : 
                        (N155)? mem[810] : 
                        (N157)? mem[850] : 
                        (N159)? mem[890] : 
                        (N161)? mem[930] : 
                        (N163)? mem[970] : 
                        (N165)? mem[1010] : 
                        (N167)? mem[1050] : 
                        (N169)? mem[1090] : 
                        (N171)? mem[1130] : 
                        (N173)? mem[1170] : 
                        (N175)? mem[1210] : 
                        (N177)? mem[1250] : 
                        (N116)? mem[1290] : 
                        (N118)? mem[1330] : 
                        (N120)? mem[1370] : 
                        (N122)? mem[1410] : 
                        (N124)? mem[1450] : 
                        (N126)? mem[1490] : 
                        (N128)? mem[1530] : 
                        (N130)? mem[1570] : 
                        (N132)? mem[1610] : 
                        (N134)? mem[1650] : 
                        (N136)? mem[1690] : 
                        (N138)? mem[1730] : 
                        (N140)? mem[1770] : 
                        (N142)? mem[1810] : 
                        (N144)? mem[1850] : 
                        (N146)? mem[1890] : 
                        (N148)? mem[1930] : 
                        (N150)? mem[1970] : 
                        (N152)? mem[2010] : 
                        (N154)? mem[2050] : 
                        (N156)? mem[2090] : 
                        (N158)? mem[2130] : 
                        (N160)? mem[2170] : 
                        (N162)? mem[2210] : 
                        (N164)? mem[2250] : 
                        (N166)? mem[2290] : 
                        (N168)? mem[2330] : 
                        (N170)? mem[2370] : 
                        (N172)? mem[2410] : 
                        (N174)? mem[2450] : 
                        (N176)? mem[2490] : 
                        (N178)? mem[2530] : 1'b0;
  assign data_out[9] = (N115)? mem[9] : 
                       (N117)? mem[49] : 
                       (N119)? mem[89] : 
                       (N121)? mem[129] : 
                       (N123)? mem[169] : 
                       (N125)? mem[209] : 
                       (N127)? mem[249] : 
                       (N129)? mem[289] : 
                       (N131)? mem[329] : 
                       (N133)? mem[369] : 
                       (N135)? mem[409] : 
                       (N137)? mem[449] : 
                       (N139)? mem[489] : 
                       (N141)? mem[529] : 
                       (N143)? mem[569] : 
                       (N145)? mem[609] : 
                       (N147)? mem[649] : 
                       (N149)? mem[689] : 
                       (N151)? mem[729] : 
                       (N153)? mem[769] : 
                       (N155)? mem[809] : 
                       (N157)? mem[849] : 
                       (N159)? mem[889] : 
                       (N161)? mem[929] : 
                       (N163)? mem[969] : 
                       (N165)? mem[1009] : 
                       (N167)? mem[1049] : 
                       (N169)? mem[1089] : 
                       (N171)? mem[1129] : 
                       (N173)? mem[1169] : 
                       (N175)? mem[1209] : 
                       (N177)? mem[1249] : 
                       (N116)? mem[1289] : 
                       (N118)? mem[1329] : 
                       (N120)? mem[1369] : 
                       (N122)? mem[1409] : 
                       (N124)? mem[1449] : 
                       (N126)? mem[1489] : 
                       (N128)? mem[1529] : 
                       (N130)? mem[1569] : 
                       (N132)? mem[1609] : 
                       (N134)? mem[1649] : 
                       (N136)? mem[1689] : 
                       (N138)? mem[1729] : 
                       (N140)? mem[1769] : 
                       (N142)? mem[1809] : 
                       (N144)? mem[1849] : 
                       (N146)? mem[1889] : 
                       (N148)? mem[1929] : 
                       (N150)? mem[1969] : 
                       (N152)? mem[2009] : 
                       (N154)? mem[2049] : 
                       (N156)? mem[2089] : 
                       (N158)? mem[2129] : 
                       (N160)? mem[2169] : 
                       (N162)? mem[2209] : 
                       (N164)? mem[2249] : 
                       (N166)? mem[2289] : 
                       (N168)? mem[2329] : 
                       (N170)? mem[2369] : 
                       (N172)? mem[2409] : 
                       (N174)? mem[2449] : 
                       (N176)? mem[2489] : 
                       (N178)? mem[2529] : 1'b0;
  assign data_out[8] = (N115)? mem[8] : 
                       (N117)? mem[48] : 
                       (N119)? mem[88] : 
                       (N121)? mem[128] : 
                       (N123)? mem[168] : 
                       (N125)? mem[208] : 
                       (N127)? mem[248] : 
                       (N129)? mem[288] : 
                       (N131)? mem[328] : 
                       (N133)? mem[368] : 
                       (N135)? mem[408] : 
                       (N137)? mem[448] : 
                       (N139)? mem[488] : 
                       (N141)? mem[528] : 
                       (N143)? mem[568] : 
                       (N145)? mem[608] : 
                       (N147)? mem[648] : 
                       (N149)? mem[688] : 
                       (N151)? mem[728] : 
                       (N153)? mem[768] : 
                       (N155)? mem[808] : 
                       (N157)? mem[848] : 
                       (N159)? mem[888] : 
                       (N161)? mem[928] : 
                       (N163)? mem[968] : 
                       (N165)? mem[1008] : 
                       (N167)? mem[1048] : 
                       (N169)? mem[1088] : 
                       (N171)? mem[1128] : 
                       (N173)? mem[1168] : 
                       (N175)? mem[1208] : 
                       (N177)? mem[1248] : 
                       (N116)? mem[1288] : 
                       (N118)? mem[1328] : 
                       (N120)? mem[1368] : 
                       (N122)? mem[1408] : 
                       (N124)? mem[1448] : 
                       (N126)? mem[1488] : 
                       (N128)? mem[1528] : 
                       (N130)? mem[1568] : 
                       (N132)? mem[1608] : 
                       (N134)? mem[1648] : 
                       (N136)? mem[1688] : 
                       (N138)? mem[1728] : 
                       (N140)? mem[1768] : 
                       (N142)? mem[1808] : 
                       (N144)? mem[1848] : 
                       (N146)? mem[1888] : 
                       (N148)? mem[1928] : 
                       (N150)? mem[1968] : 
                       (N152)? mem[2008] : 
                       (N154)? mem[2048] : 
                       (N156)? mem[2088] : 
                       (N158)? mem[2128] : 
                       (N160)? mem[2168] : 
                       (N162)? mem[2208] : 
                       (N164)? mem[2248] : 
                       (N166)? mem[2288] : 
                       (N168)? mem[2328] : 
                       (N170)? mem[2368] : 
                       (N172)? mem[2408] : 
                       (N174)? mem[2448] : 
                       (N176)? mem[2488] : 
                       (N178)? mem[2528] : 1'b0;
  assign data_out[7] = (N115)? mem[7] : 
                       (N117)? mem[47] : 
                       (N119)? mem[87] : 
                       (N121)? mem[127] : 
                       (N123)? mem[167] : 
                       (N125)? mem[207] : 
                       (N127)? mem[247] : 
                       (N129)? mem[287] : 
                       (N131)? mem[327] : 
                       (N133)? mem[367] : 
                       (N135)? mem[407] : 
                       (N137)? mem[447] : 
                       (N139)? mem[487] : 
                       (N141)? mem[527] : 
                       (N143)? mem[567] : 
                       (N145)? mem[607] : 
                       (N147)? mem[647] : 
                       (N149)? mem[687] : 
                       (N151)? mem[727] : 
                       (N153)? mem[767] : 
                       (N155)? mem[807] : 
                       (N157)? mem[847] : 
                       (N159)? mem[887] : 
                       (N161)? mem[927] : 
                       (N163)? mem[967] : 
                       (N165)? mem[1007] : 
                       (N167)? mem[1047] : 
                       (N169)? mem[1087] : 
                       (N171)? mem[1127] : 
                       (N173)? mem[1167] : 
                       (N175)? mem[1207] : 
                       (N177)? mem[1247] : 
                       (N116)? mem[1287] : 
                       (N118)? mem[1327] : 
                       (N120)? mem[1367] : 
                       (N122)? mem[1407] : 
                       (N124)? mem[1447] : 
                       (N126)? mem[1487] : 
                       (N128)? mem[1527] : 
                       (N130)? mem[1567] : 
                       (N132)? mem[1607] : 
                       (N134)? mem[1647] : 
                       (N136)? mem[1687] : 
                       (N138)? mem[1727] : 
                       (N140)? mem[1767] : 
                       (N142)? mem[1807] : 
                       (N144)? mem[1847] : 
                       (N146)? mem[1887] : 
                       (N148)? mem[1927] : 
                       (N150)? mem[1967] : 
                       (N152)? mem[2007] : 
                       (N154)? mem[2047] : 
                       (N156)? mem[2087] : 
                       (N158)? mem[2127] : 
                       (N160)? mem[2167] : 
                       (N162)? mem[2207] : 
                       (N164)? mem[2247] : 
                       (N166)? mem[2287] : 
                       (N168)? mem[2327] : 
                       (N170)? mem[2367] : 
                       (N172)? mem[2407] : 
                       (N174)? mem[2447] : 
                       (N176)? mem[2487] : 
                       (N178)? mem[2527] : 1'b0;
  assign data_out[6] = (N115)? mem[6] : 
                       (N117)? mem[46] : 
                       (N119)? mem[86] : 
                       (N121)? mem[126] : 
                       (N123)? mem[166] : 
                       (N125)? mem[206] : 
                       (N127)? mem[246] : 
                       (N129)? mem[286] : 
                       (N131)? mem[326] : 
                       (N133)? mem[366] : 
                       (N135)? mem[406] : 
                       (N137)? mem[446] : 
                       (N139)? mem[486] : 
                       (N141)? mem[526] : 
                       (N143)? mem[566] : 
                       (N145)? mem[606] : 
                       (N147)? mem[646] : 
                       (N149)? mem[686] : 
                       (N151)? mem[726] : 
                       (N153)? mem[766] : 
                       (N155)? mem[806] : 
                       (N157)? mem[846] : 
                       (N159)? mem[886] : 
                       (N161)? mem[926] : 
                       (N163)? mem[966] : 
                       (N165)? mem[1006] : 
                       (N167)? mem[1046] : 
                       (N169)? mem[1086] : 
                       (N171)? mem[1126] : 
                       (N173)? mem[1166] : 
                       (N175)? mem[1206] : 
                       (N177)? mem[1246] : 
                       (N116)? mem[1286] : 
                       (N118)? mem[1326] : 
                       (N120)? mem[1366] : 
                       (N122)? mem[1406] : 
                       (N124)? mem[1446] : 
                       (N126)? mem[1486] : 
                       (N128)? mem[1526] : 
                       (N130)? mem[1566] : 
                       (N132)? mem[1606] : 
                       (N134)? mem[1646] : 
                       (N136)? mem[1686] : 
                       (N138)? mem[1726] : 
                       (N140)? mem[1766] : 
                       (N142)? mem[1806] : 
                       (N144)? mem[1846] : 
                       (N146)? mem[1886] : 
                       (N148)? mem[1926] : 
                       (N150)? mem[1966] : 
                       (N152)? mem[2006] : 
                       (N154)? mem[2046] : 
                       (N156)? mem[2086] : 
                       (N158)? mem[2126] : 
                       (N160)? mem[2166] : 
                       (N162)? mem[2206] : 
                       (N164)? mem[2246] : 
                       (N166)? mem[2286] : 
                       (N168)? mem[2326] : 
                       (N170)? mem[2366] : 
                       (N172)? mem[2406] : 
                       (N174)? mem[2446] : 
                       (N176)? mem[2486] : 
                       (N178)? mem[2526] : 1'b0;
  assign data_out[5] = (N115)? mem[5] : 
                       (N117)? mem[45] : 
                       (N119)? mem[85] : 
                       (N121)? mem[125] : 
                       (N123)? mem[165] : 
                       (N125)? mem[205] : 
                       (N127)? mem[245] : 
                       (N129)? mem[285] : 
                       (N131)? mem[325] : 
                       (N133)? mem[365] : 
                       (N135)? mem[405] : 
                       (N137)? mem[445] : 
                       (N139)? mem[485] : 
                       (N141)? mem[525] : 
                       (N143)? mem[565] : 
                       (N145)? mem[605] : 
                       (N147)? mem[645] : 
                       (N149)? mem[685] : 
                       (N151)? mem[725] : 
                       (N153)? mem[765] : 
                       (N155)? mem[805] : 
                       (N157)? mem[845] : 
                       (N159)? mem[885] : 
                       (N161)? mem[925] : 
                       (N163)? mem[965] : 
                       (N165)? mem[1005] : 
                       (N167)? mem[1045] : 
                       (N169)? mem[1085] : 
                       (N171)? mem[1125] : 
                       (N173)? mem[1165] : 
                       (N175)? mem[1205] : 
                       (N177)? mem[1245] : 
                       (N116)? mem[1285] : 
                       (N118)? mem[1325] : 
                       (N120)? mem[1365] : 
                       (N122)? mem[1405] : 
                       (N124)? mem[1445] : 
                       (N126)? mem[1485] : 
                       (N128)? mem[1525] : 
                       (N130)? mem[1565] : 
                       (N132)? mem[1605] : 
                       (N134)? mem[1645] : 
                       (N136)? mem[1685] : 
                       (N138)? mem[1725] : 
                       (N140)? mem[1765] : 
                       (N142)? mem[1805] : 
                       (N144)? mem[1845] : 
                       (N146)? mem[1885] : 
                       (N148)? mem[1925] : 
                       (N150)? mem[1965] : 
                       (N152)? mem[2005] : 
                       (N154)? mem[2045] : 
                       (N156)? mem[2085] : 
                       (N158)? mem[2125] : 
                       (N160)? mem[2165] : 
                       (N162)? mem[2205] : 
                       (N164)? mem[2245] : 
                       (N166)? mem[2285] : 
                       (N168)? mem[2325] : 
                       (N170)? mem[2365] : 
                       (N172)? mem[2405] : 
                       (N174)? mem[2445] : 
                       (N176)? mem[2485] : 
                       (N178)? mem[2525] : 1'b0;
  assign data_out[4] = (N115)? mem[4] : 
                       (N117)? mem[44] : 
                       (N119)? mem[84] : 
                       (N121)? mem[124] : 
                       (N123)? mem[164] : 
                       (N125)? mem[204] : 
                       (N127)? mem[244] : 
                       (N129)? mem[284] : 
                       (N131)? mem[324] : 
                       (N133)? mem[364] : 
                       (N135)? mem[404] : 
                       (N137)? mem[444] : 
                       (N139)? mem[484] : 
                       (N141)? mem[524] : 
                       (N143)? mem[564] : 
                       (N145)? mem[604] : 
                       (N147)? mem[644] : 
                       (N149)? mem[684] : 
                       (N151)? mem[724] : 
                       (N153)? mem[764] : 
                       (N155)? mem[804] : 
                       (N157)? mem[844] : 
                       (N159)? mem[884] : 
                       (N161)? mem[924] : 
                       (N163)? mem[964] : 
                       (N165)? mem[1004] : 
                       (N167)? mem[1044] : 
                       (N169)? mem[1084] : 
                       (N171)? mem[1124] : 
                       (N173)? mem[1164] : 
                       (N175)? mem[1204] : 
                       (N177)? mem[1244] : 
                       (N116)? mem[1284] : 
                       (N118)? mem[1324] : 
                       (N120)? mem[1364] : 
                       (N122)? mem[1404] : 
                       (N124)? mem[1444] : 
                       (N126)? mem[1484] : 
                       (N128)? mem[1524] : 
                       (N130)? mem[1564] : 
                       (N132)? mem[1604] : 
                       (N134)? mem[1644] : 
                       (N136)? mem[1684] : 
                       (N138)? mem[1724] : 
                       (N140)? mem[1764] : 
                       (N142)? mem[1804] : 
                       (N144)? mem[1844] : 
                       (N146)? mem[1884] : 
                       (N148)? mem[1924] : 
                       (N150)? mem[1964] : 
                       (N152)? mem[2004] : 
                       (N154)? mem[2044] : 
                       (N156)? mem[2084] : 
                       (N158)? mem[2124] : 
                       (N160)? mem[2164] : 
                       (N162)? mem[2204] : 
                       (N164)? mem[2244] : 
                       (N166)? mem[2284] : 
                       (N168)? mem[2324] : 
                       (N170)? mem[2364] : 
                       (N172)? mem[2404] : 
                       (N174)? mem[2444] : 
                       (N176)? mem[2484] : 
                       (N178)? mem[2524] : 1'b0;
  assign data_out[3] = (N115)? mem[3] : 
                       (N117)? mem[43] : 
                       (N119)? mem[83] : 
                       (N121)? mem[123] : 
                       (N123)? mem[163] : 
                       (N125)? mem[203] : 
                       (N127)? mem[243] : 
                       (N129)? mem[283] : 
                       (N131)? mem[323] : 
                       (N133)? mem[363] : 
                       (N135)? mem[403] : 
                       (N137)? mem[443] : 
                       (N139)? mem[483] : 
                       (N141)? mem[523] : 
                       (N143)? mem[563] : 
                       (N145)? mem[603] : 
                       (N147)? mem[643] : 
                       (N149)? mem[683] : 
                       (N151)? mem[723] : 
                       (N153)? mem[763] : 
                       (N155)? mem[803] : 
                       (N157)? mem[843] : 
                       (N159)? mem[883] : 
                       (N161)? mem[923] : 
                       (N163)? mem[963] : 
                       (N165)? mem[1003] : 
                       (N167)? mem[1043] : 
                       (N169)? mem[1083] : 
                       (N171)? mem[1123] : 
                       (N173)? mem[1163] : 
                       (N175)? mem[1203] : 
                       (N177)? mem[1243] : 
                       (N116)? mem[1283] : 
                       (N118)? mem[1323] : 
                       (N120)? mem[1363] : 
                       (N122)? mem[1403] : 
                       (N124)? mem[1443] : 
                       (N126)? mem[1483] : 
                       (N128)? mem[1523] : 
                       (N130)? mem[1563] : 
                       (N132)? mem[1603] : 
                       (N134)? mem[1643] : 
                       (N136)? mem[1683] : 
                       (N138)? mem[1723] : 
                       (N140)? mem[1763] : 
                       (N142)? mem[1803] : 
                       (N144)? mem[1843] : 
                       (N146)? mem[1883] : 
                       (N148)? mem[1923] : 
                       (N150)? mem[1963] : 
                       (N152)? mem[2003] : 
                       (N154)? mem[2043] : 
                       (N156)? mem[2083] : 
                       (N158)? mem[2123] : 
                       (N160)? mem[2163] : 
                       (N162)? mem[2203] : 
                       (N164)? mem[2243] : 
                       (N166)? mem[2283] : 
                       (N168)? mem[2323] : 
                       (N170)? mem[2363] : 
                       (N172)? mem[2403] : 
                       (N174)? mem[2443] : 
                       (N176)? mem[2483] : 
                       (N178)? mem[2523] : 1'b0;
  assign data_out[2] = (N115)? mem[2] : 
                       (N117)? mem[42] : 
                       (N119)? mem[82] : 
                       (N121)? mem[122] : 
                       (N123)? mem[162] : 
                       (N125)? mem[202] : 
                       (N127)? mem[242] : 
                       (N129)? mem[282] : 
                       (N131)? mem[322] : 
                       (N133)? mem[362] : 
                       (N135)? mem[402] : 
                       (N137)? mem[442] : 
                       (N139)? mem[482] : 
                       (N141)? mem[522] : 
                       (N143)? mem[562] : 
                       (N145)? mem[602] : 
                       (N147)? mem[642] : 
                       (N149)? mem[682] : 
                       (N151)? mem[722] : 
                       (N153)? mem[762] : 
                       (N155)? mem[802] : 
                       (N157)? mem[842] : 
                       (N159)? mem[882] : 
                       (N161)? mem[922] : 
                       (N163)? mem[962] : 
                       (N165)? mem[1002] : 
                       (N167)? mem[1042] : 
                       (N169)? mem[1082] : 
                       (N171)? mem[1122] : 
                       (N173)? mem[1162] : 
                       (N175)? mem[1202] : 
                       (N177)? mem[1242] : 
                       (N116)? mem[1282] : 
                       (N118)? mem[1322] : 
                       (N120)? mem[1362] : 
                       (N122)? mem[1402] : 
                       (N124)? mem[1442] : 
                       (N126)? mem[1482] : 
                       (N128)? mem[1522] : 
                       (N130)? mem[1562] : 
                       (N132)? mem[1602] : 
                       (N134)? mem[1642] : 
                       (N136)? mem[1682] : 
                       (N138)? mem[1722] : 
                       (N140)? mem[1762] : 
                       (N142)? mem[1802] : 
                       (N144)? mem[1842] : 
                       (N146)? mem[1882] : 
                       (N148)? mem[1922] : 
                       (N150)? mem[1962] : 
                       (N152)? mem[2002] : 
                       (N154)? mem[2042] : 
                       (N156)? mem[2082] : 
                       (N158)? mem[2122] : 
                       (N160)? mem[2162] : 
                       (N162)? mem[2202] : 
                       (N164)? mem[2242] : 
                       (N166)? mem[2282] : 
                       (N168)? mem[2322] : 
                       (N170)? mem[2362] : 
                       (N172)? mem[2402] : 
                       (N174)? mem[2442] : 
                       (N176)? mem[2482] : 
                       (N178)? mem[2522] : 1'b0;
  assign data_out[1] = (N115)? mem[1] : 
                       (N117)? mem[41] : 
                       (N119)? mem[81] : 
                       (N121)? mem[121] : 
                       (N123)? mem[161] : 
                       (N125)? mem[201] : 
                       (N127)? mem[241] : 
                       (N129)? mem[281] : 
                       (N131)? mem[321] : 
                       (N133)? mem[361] : 
                       (N135)? mem[401] : 
                       (N137)? mem[441] : 
                       (N139)? mem[481] : 
                       (N141)? mem[521] : 
                       (N143)? mem[561] : 
                       (N145)? mem[601] : 
                       (N147)? mem[641] : 
                       (N149)? mem[681] : 
                       (N151)? mem[721] : 
                       (N153)? mem[761] : 
                       (N155)? mem[801] : 
                       (N157)? mem[841] : 
                       (N159)? mem[881] : 
                       (N161)? mem[921] : 
                       (N163)? mem[961] : 
                       (N165)? mem[1001] : 
                       (N167)? mem[1041] : 
                       (N169)? mem[1081] : 
                       (N171)? mem[1121] : 
                       (N173)? mem[1161] : 
                       (N175)? mem[1201] : 
                       (N177)? mem[1241] : 
                       (N116)? mem[1281] : 
                       (N118)? mem[1321] : 
                       (N120)? mem[1361] : 
                       (N122)? mem[1401] : 
                       (N124)? mem[1441] : 
                       (N126)? mem[1481] : 
                       (N128)? mem[1521] : 
                       (N130)? mem[1561] : 
                       (N132)? mem[1601] : 
                       (N134)? mem[1641] : 
                       (N136)? mem[1681] : 
                       (N138)? mem[1721] : 
                       (N140)? mem[1761] : 
                       (N142)? mem[1801] : 
                       (N144)? mem[1841] : 
                       (N146)? mem[1881] : 
                       (N148)? mem[1921] : 
                       (N150)? mem[1961] : 
                       (N152)? mem[2001] : 
                       (N154)? mem[2041] : 
                       (N156)? mem[2081] : 
                       (N158)? mem[2121] : 
                       (N160)? mem[2161] : 
                       (N162)? mem[2201] : 
                       (N164)? mem[2241] : 
                       (N166)? mem[2281] : 
                       (N168)? mem[2321] : 
                       (N170)? mem[2361] : 
                       (N172)? mem[2401] : 
                       (N174)? mem[2441] : 
                       (N176)? mem[2481] : 
                       (N178)? mem[2521] : 1'b0;
  assign data_out[0] = (N115)? mem[0] : 
                       (N117)? mem[40] : 
                       (N119)? mem[80] : 
                       (N121)? mem[120] : 
                       (N123)? mem[160] : 
                       (N125)? mem[200] : 
                       (N127)? mem[240] : 
                       (N129)? mem[280] : 
                       (N131)? mem[320] : 
                       (N133)? mem[360] : 
                       (N135)? mem[400] : 
                       (N137)? mem[440] : 
                       (N139)? mem[480] : 
                       (N141)? mem[520] : 
                       (N143)? mem[560] : 
                       (N145)? mem[600] : 
                       (N147)? mem[640] : 
                       (N149)? mem[680] : 
                       (N151)? mem[720] : 
                       (N153)? mem[760] : 
                       (N155)? mem[800] : 
                       (N157)? mem[840] : 
                       (N159)? mem[880] : 
                       (N161)? mem[920] : 
                       (N163)? mem[960] : 
                       (N165)? mem[1000] : 
                       (N167)? mem[1040] : 
                       (N169)? mem[1080] : 
                       (N171)? mem[1120] : 
                       (N173)? mem[1160] : 
                       (N175)? mem[1200] : 
                       (N177)? mem[1240] : 
                       (N116)? mem[1280] : 
                       (N118)? mem[1320] : 
                       (N120)? mem[1360] : 
                       (N122)? mem[1400] : 
                       (N124)? mem[1440] : 
                       (N126)? mem[1480] : 
                       (N128)? mem[1520] : 
                       (N130)? mem[1560] : 
                       (N132)? mem[1600] : 
                       (N134)? mem[1640] : 
                       (N136)? mem[1680] : 
                       (N138)? mem[1720] : 
                       (N140)? mem[1760] : 
                       (N142)? mem[1800] : 
                       (N144)? mem[1840] : 
                       (N146)? mem[1880] : 
                       (N148)? mem[1920] : 
                       (N150)? mem[1960] : 
                       (N152)? mem[2000] : 
                       (N154)? mem[2040] : 
                       (N156)? mem[2080] : 
                       (N158)? mem[2120] : 
                       (N160)? mem[2160] : 
                       (N162)? mem[2200] : 
                       (N164)? mem[2240] : 
                       (N166)? mem[2280] : 
                       (N168)? mem[2320] : 
                       (N170)? mem[2360] : 
                       (N172)? mem[2400] : 
                       (N174)? mem[2440] : 
                       (N176)? mem[2480] : 
                       (N178)? mem[2520] : 1'b0;

  bsg_dff_width_p1
  llr_read_en_dff
  (
    .clk_i(clk_i),
    .data_i(read_en),
    .data_o(llr_read_en_r)
  );


  bsg_dff_en_bypass_width_p40
  llr_dff_bypass
  (
    .clk_i(clk_i),
    .en_i(llr_read_en_r),
    .data_i(data_out),
    .data_o(data_o)
  );

  assign N5811 = addr_i[5] & N5869;
  assign N5812 = addr_i[5] & N5870;
  assign N5813 = addr_i[5] & N5871;
  assign N5814 = addr_i[2] & N5881;
  assign N5815 = addr_i[2] & N5882;
  assign N5816 = addr_i[2] & N5883;
  assign N415 = N5811 & N5814;
  assign N414 = N5811 & N5815;
  assign N413 = N5811 & N5816;
  assign N412 = N5811 & N5888;
  assign N411 = N5811 & N5831;
  assign N410 = N5811 & N5832;
  assign N409 = N5811 & N5833;
  assign N408 = N5811 & N5834;
  assign N407 = N5812 & N5814;
  assign N406 = N5812 & N5815;
  assign N405 = N5812 & N5816;
  assign N404 = N5812 & N5888;
  assign N403 = N5812 & N5831;
  assign N402 = N5812 & N5832;
  assign N401 = N5812 & N5833;
  assign N400 = N5812 & N5834;
  assign N399 = N5813 & N5814;
  assign N398 = N5813 & N5815;
  assign N397 = N5813 & N5816;
  assign N396 = N5813 & N5888;
  assign N395 = N5813 & N5831;
  assign N394 = N5813 & N5832;
  assign N393 = N5813 & N5833;
  assign N392 = N5813 & N5834;
  assign N391 = N5876 & N5814;
  assign N390 = N5876 & N5815;
  assign N389 = N5876 & N5816;
  assign N388 = N5826 & N5814;
  assign N387 = N5826 & N5815;
  assign N386 = N5826 & N5816;
  assign N385 = N5827 & N5814;
  assign N384 = N5827 & N5815;
  assign N383 = N5827 & N5816;
  assign N382 = N5828 & N5814;
  assign N381 = N5828 & N5815;
  assign N380 = N5828 & N5816;
  assign N379 = N5829 & N5814;
  assign N378 = N5829 & N5815;
  assign N377 = N5829 & N5816;
  assign N884 = N5835 & N5888;
  assign N883 = N5836 & N5888;
  assign N882 = N5837 & N5888;
  assign N881 = N5876 & N5838;
  assign N880 = N5876 & N5839;
  assign N879 = N5876 & N5840;
  assign N878 = N5876 & N5831;
  assign N877 = N5876 & N5832;
  assign N876 = N5876 & N5833;
  assign N875 = N5876 & N5834;
  assign N874 = N5826 & N5888;
  assign N873 = N5827 & N5888;
  assign N872 = N5828 & N5888;
  assign N871 = N5829 & N5888;
  assign N5817 = N5825 & N5869;
  assign N5818 = N5825 & N5870;
  assign N5819 = N5825 & N5871;
  assign N5820 = N5825 & N5872;
  assign N5821 = N5830 & N5881;
  assign N5822 = N5830 & N5882;
  assign N5823 = N5830 & N5883;
  assign N5824 = N5830 & N5884;
  assign N1127 = N5835 & N5821;
  assign N1126 = N5835 & N5822;
  assign N1125 = N5835 & N5823;
  assign N1124 = N5835 & N5824;
  assign N1123 = N5836 & N5821;
  assign N1122 = N5836 & N5822;
  assign N1121 = N5836 & N5823;
  assign N1120 = N5836 & N5824;
  assign N1119 = N5837 & N5821;
  assign N1118 = N5837 & N5822;
  assign N1117 = N5837 & N5823;
  assign N1116 = N5837 & N5824;
  assign N1115 = N5859 & N5821;
  assign N1114 = N5859 & N5822;
  assign N1113 = N5859 & N5823;
  assign N1112 = N5859 & N5824;
  assign N1111 = N5817 & N5838;
  assign N1110 = N5817 & N5839;
  assign N1109 = N5817 & N5840;
  assign N1108 = N5817 & N5864;
  assign N1107 = N5817 & N5821;
  assign N1106 = N5817 & N5822;
  assign N1105 = N5817 & N5823;
  assign N1104 = N5817 & N5824;
  assign N1103 = N5818 & N5838;
  assign N1102 = N5818 & N5839;
  assign N1101 = N5818 & N5840;
  assign N1100 = N5818 & N5864;
  assign N1099 = N5818 & N5821;
  assign N1098 = N5818 & N5822;
  assign N1097 = N5818 & N5823;
  assign N1096 = N5818 & N5824;
  assign N1095 = N5819 & N5838;
  assign N1094 = N5819 & N5839;
  assign N1093 = N5819 & N5840;
  assign N1092 = N5819 & N5864;
  assign N1091 = N5819 & N5821;
  assign N1090 = N5819 & N5822;
  assign N1089 = N5819 & N5823;
  assign N1088 = N5819 & N5824;
  assign N1087 = N5820 & N5838;
  assign N1086 = N5820 & N5839;
  assign N1085 = N5820 & N5840;
  assign N1084 = N5820 & N5864;
  assign N1083 = N5820 & N5821;
  assign N1082 = N5820 & N5822;
  assign N1081 = N5820 & N5823;
  assign N1080 = N5820 & N5824;
  assign N5825 = ~addr_i[5];
  assign N5826 = N5825 & N5869;
  assign N5827 = N5825 & N5870;
  assign N5828 = N5825 & N5871;
  assign N5829 = N5825 & N5872;
  assign N5830 = ~addr_i[2];
  assign N5831 = N5830 & N5881;
  assign N5832 = N5830 & N5882;
  assign N5833 = N5830 & N5883;
  assign N5834 = N5830 & N5884;
  assign N1240 = N5835 & N5831;
  assign N1239 = N5835 & N5832;
  assign N1238 = N5835 & N5833;
  assign N1237 = N5835 & N5834;
  assign N1236 = N5836 & N5831;
  assign N1235 = N5836 & N5832;
  assign N1234 = N5836 & N5833;
  assign N1233 = N5836 & N5834;
  assign N1232 = N5837 & N5831;
  assign N1231 = N5837 & N5832;
  assign N1230 = N5837 & N5833;
  assign N1229 = N5837 & N5834;
  assign N1228 = N5859 & N5831;
  assign N1227 = N5859 & N5832;
  assign N1226 = N5859 & N5833;
  assign N1225 = N5859 & N5834;
  assign N1224 = N5826 & N5838;
  assign N1223 = N5826 & N5839;
  assign N1222 = N5826 & N5840;
  assign N1221 = N5826 & N5864;
  assign N1220 = N5826 & N5831;
  assign N1219 = N5826 & N5832;
  assign N1218 = N5826 & N5833;
  assign N1217 = N5826 & N5834;
  assign N1216 = N5827 & N5838;
  assign N1215 = N5827 & N5839;
  assign N1214 = N5827 & N5840;
  assign N1213 = N5827 & N5864;
  assign N1212 = N5827 & N5831;
  assign N1211 = N5827 & N5832;
  assign N1210 = N5827 & N5833;
  assign N1209 = N5827 & N5834;
  assign N1208 = N5828 & N5838;
  assign N1207 = N5828 & N5839;
  assign N1206 = N5828 & N5840;
  assign N1205 = N5828 & N5864;
  assign N1204 = N5828 & N5831;
  assign N1203 = N5828 & N5832;
  assign N1202 = N5828 & N5833;
  assign N1201 = N5828 & N5834;
  assign N1200 = N5829 & N5838;
  assign N1199 = N5829 & N5839;
  assign N1198 = N5829 & N5840;
  assign N1197 = N5829 & N5864;
  assign N1196 = N5829 & N5831;
  assign N1195 = N5829 & N5832;
  assign N1194 = N5829 & N5833;
  assign N1193 = N5829 & N5834;
  assign N5835 = addr_i[5] & N5869;
  assign N5836 = addr_i[5] & N5870;
  assign N5837 = addr_i[5] & N5871;
  assign N5838 = addr_i[2] & N5881;
  assign N5839 = addr_i[2] & N5882;
  assign N5840 = addr_i[2] & N5883;
  assign N1344 = N5835 & N5838;
  assign N1343 = N5835 & N5839;
  assign N1342 = N5835 & N5840;
  assign N1341 = N5835 & N5864;
  assign N1340 = N5835 & N5889;
  assign N1339 = N5835 & N5890;
  assign N1338 = N5835 & N5891;
  assign N1337 = N5835 & N5892;
  assign N1336 = N5836 & N5838;
  assign N1335 = N5836 & N5839;
  assign N1334 = N5836 & N5840;
  assign N1333 = N5836 & N5864;
  assign N1332 = N5836 & N5889;
  assign N1331 = N5836 & N5890;
  assign N1330 = N5836 & N5891;
  assign N1329 = N5836 & N5892;
  assign N1328 = N5837 & N5838;
  assign N1327 = N5837 & N5839;
  assign N1326 = N5837 & N5840;
  assign N1325 = N5837 & N5864;
  assign N1324 = N5837 & N5889;
  assign N1323 = N5837 & N5890;
  assign N1322 = N5837 & N5891;
  assign N1321 = N5837 & N5892;
  assign N1320 = N5859 & N5838;
  assign N1319 = N5859 & N5839;
  assign N1318 = N5859 & N5840;
  assign N1317 = N5877 & N5838;
  assign N1316 = N5877 & N5839;
  assign N1315 = N5877 & N5840;
  assign N1314 = N5878 & N5838;
  assign N1313 = N5878 & N5839;
  assign N1312 = N5878 & N5840;
  assign N1311 = N5879 & N5838;
  assign N1310 = N5879 & N5839;
  assign N1309 = N5879 & N5840;
  assign N1308 = N5880 & N5838;
  assign N1307 = N5880 & N5839;
  assign N1306 = N5880 & N5840;
  assign N1748 = N5841 & N5864;
  assign N1747 = N5842 & N5864;
  assign N1746 = N5843 & N5864;
  assign N1745 = N5859 & N5844;
  assign N1744 = N5859 & N5845;
  assign N1743 = N5859 & N5846;
  assign N1742 = N5859 & N5889;
  assign N1741 = N5859 & N5890;
  assign N1740 = N5859 & N5891;
  assign N1739 = N5859 & N5892;
  assign N1738 = N5877 & N5864;
  assign N1737 = N5878 & N5864;
  assign N1736 = N5879 & N5864;
  assign N1735 = N5880 & N5864;
  assign N2040 = N5841 & N5889;
  assign N2039 = N5841 & N5890;
  assign N2038 = N5841 & N5891;
  assign N2037 = N5841 & N5892;
  assign N2036 = N5842 & N5889;
  assign N2035 = N5842 & N5890;
  assign N2034 = N5842 & N5891;
  assign N2033 = N5842 & N5892;
  assign N2032 = N5843 & N5889;
  assign N2031 = N5843 & N5890;
  assign N2030 = N5843 & N5891;
  assign N2029 = N5843 & N5892;
  assign N2028 = N5849 & N5889;
  assign N2027 = N5849 & N5890;
  assign N2026 = N5849 & N5891;
  assign N2025 = N5849 & N5892;
  assign N2024 = N5877 & N5844;
  assign N2023 = N5877 & N5845;
  assign N2022 = N5877 & N5846;
  assign N2021 = N5877 & N5854;
  assign N2020 = N5878 & N5844;
  assign N2019 = N5878 & N5845;
  assign N2018 = N5878 & N5846;
  assign N2017 = N5878 & N5854;
  assign N2016 = N5879 & N5844;
  assign N2015 = N5879 & N5845;
  assign N2014 = N5879 & N5846;
  assign N2013 = N5879 & N5854;
  assign N2012 = N5880 & N5844;
  assign N2011 = N5880 & N5845;
  assign N2010 = N5880 & N5846;
  assign N2009 = N5880 & N5854;
  assign N5841 = addr_i[5] & N5869;
  assign N5842 = addr_i[5] & N5870;
  assign N5843 = addr_i[5] & N5871;
  assign N5844 = addr_i[2] & N5881;
  assign N5845 = addr_i[2] & N5882;
  assign N5846 = addr_i[2] & N5883;
  assign N2209 = N5841 & N5844;
  assign N2208 = N5841 & N5845;
  assign N2207 = N5841 & N5846;
  assign N2206 = N5841 & N5854;
  assign N2205 = N5841 & N5865;
  assign N2204 = N5841 & N5866;
  assign N2203 = N5841 & N5867;
  assign N2202 = N5841 & N5868;
  assign N2201 = N5842 & N5844;
  assign N2200 = N5842 & N5845;
  assign N2199 = N5842 & N5846;
  assign N2198 = N5842 & N5854;
  assign N2197 = N5842 & N5865;
  assign N2196 = N5842 & N5866;
  assign N2195 = N5842 & N5867;
  assign N2194 = N5842 & N5868;
  assign N2193 = N5843 & N5844;
  assign N2192 = N5843 & N5845;
  assign N2191 = N5843 & N5846;
  assign N2190 = N5843 & N5854;
  assign N2189 = N5843 & N5865;
  assign N2188 = N5843 & N5866;
  assign N2187 = N5843 & N5867;
  assign N2186 = N5843 & N5868;
  assign N2185 = N5849 & N5844;
  assign N2184 = N5849 & N5845;
  assign N2183 = N5849 & N5846;
  assign N2182 = N5860 & N5844;
  assign N2181 = N5860 & N5845;
  assign N2180 = N5860 & N5846;
  assign N2179 = N5861 & N5844;
  assign N2178 = N5861 & N5845;
  assign N2177 = N5861 & N5846;
  assign N2176 = N5862 & N5844;
  assign N2175 = N5862 & N5845;
  assign N2174 = N5862 & N5846;
  assign N2173 = N5863 & N5844;
  assign N2172 = N5863 & N5845;
  assign N2171 = N5863 & N5846;
  assign N2542 = N5849 & N5865;
  assign N2541 = N5849 & N5866;
  assign N2540 = N5849 & N5867;
  assign N2539 = N5849 & N5868;
  assign N2538 = N5860 & N5854;
  assign N2537 = N5861 & N5854;
  assign N2536 = N5862 & N5854;
  assign N2535 = N5863 & N5854;
  assign N5847 = addr_i[5] & N5872;
  assign N5848 = addr_i[2] & N5884;
  assign N2817 = N5873 & N5848;
  assign N2816 = N5874 & N5848;
  assign N2815 = N5875 & N5848;
  assign N2814 = N5847 & N5885;
  assign N2813 = N5847 & N5886;
  assign N2812 = N5847 & N5887;
  assign N2811 = N5847 & N5848;
  assign N2810 = N5847 & N5865;
  assign N2809 = N5847 & N5866;
  assign N2808 = N5847 & N5867;
  assign N2807 = N5847 & N5868;
  assign N2806 = N5860 & N5848;
  assign N2805 = N5861 & N5848;
  assign N2804 = N5862 & N5848;
  assign N2803 = N5863 & N5848;
  assign N5849 = addr_i[5] & N5872;
  assign N5850 = N5825 & N5869;
  assign N5851 = N5825 & N5870;
  assign N5852 = N5825 & N5871;
  assign N5853 = N5825 & N5872;
  assign N5854 = addr_i[2] & N5884;
  assign N5855 = N5830 & N5881;
  assign N5856 = N5830 & N5882;
  assign N5857 = N5830 & N5883;
  assign N5858 = N5830 & N5884;
  assign N2937 = N5873 & N5854;
  assign N2936 = N5873 & N5855;
  assign N2935 = N5873 & N5856;
  assign N2934 = N5873 & N5857;
  assign N2933 = N5873 & N5858;
  assign N2932 = N5874 & N5854;
  assign N2931 = N5874 & N5855;
  assign N2930 = N5874 & N5856;
  assign N2929 = N5874 & N5857;
  assign N2928 = N5874 & N5858;
  assign N2927 = N5875 & N5854;
  assign N2926 = N5875 & N5855;
  assign N2925 = N5875 & N5856;
  assign N2924 = N5875 & N5857;
  assign N2923 = N5875 & N5858;
  assign N2922 = N5849 & N5885;
  assign N2921 = N5849 & N5886;
  assign N2920 = N5849 & N5887;
  assign N2919 = N5849 & N5854;
  assign N2918 = N5849 & N5855;
  assign N2917 = N5849 & N5856;
  assign N2916 = N5849 & N5857;
  assign N2915 = N5849 & N5858;
  assign N2914 = N5850 & N5885;
  assign N2913 = N5850 & N5886;
  assign N2912 = N5850 & N5887;
  assign N2911 = N5850 & N5854;
  assign N2910 = N5850 & N5855;
  assign N2909 = N5850 & N5856;
  assign N2908 = N5850 & N5857;
  assign N2907 = N5850 & N5858;
  assign N2906 = N5851 & N5885;
  assign N2905 = N5851 & N5886;
  assign N2904 = N5851 & N5887;
  assign N2903 = N5851 & N5854;
  assign N2902 = N5851 & N5855;
  assign N2901 = N5851 & N5856;
  assign N2900 = N5851 & N5857;
  assign N2899 = N5851 & N5858;
  assign N2898 = N5852 & N5885;
  assign N2897 = N5852 & N5886;
  assign N2896 = N5852 & N5887;
  assign N2895 = N5852 & N5854;
  assign N2894 = N5852 & N5855;
  assign N2893 = N5852 & N5856;
  assign N2892 = N5852 & N5857;
  assign N2891 = N5852 & N5858;
  assign N2890 = N5853 & N5885;
  assign N2889 = N5853 & N5886;
  assign N2888 = N5853 & N5887;
  assign N2887 = N5853 & N5854;
  assign N2886 = N5853 & N5855;
  assign N2885 = N5853 & N5856;
  assign N2884 = N5853 & N5857;
  assign N2883 = N5853 & N5858;
  assign N5859 = addr_i[5] & N5872;
  assign N5860 = N5825 & N5869;
  assign N5861 = N5825 & N5870;
  assign N5862 = N5825 & N5871;
  assign N5863 = N5825 & N5872;
  assign N5864 = addr_i[2] & N5884;
  assign N5865 = N5830 & N5881;
  assign N5866 = N5830 & N5882;
  assign N5867 = N5830 & N5883;
  assign N5868 = N5830 & N5884;
  assign N3057 = N5873 & N5864;
  assign N3056 = N5873 & N5865;
  assign N3055 = N5873 & N5866;
  assign N3054 = N5873 & N5867;
  assign N3053 = N5873 & N5868;
  assign N3052 = N5874 & N5864;
  assign N3051 = N5874 & N5865;
  assign N3050 = N5874 & N5866;
  assign N3049 = N5874 & N5867;
  assign N3048 = N5874 & N5868;
  assign N3047 = N5875 & N5864;
  assign N3046 = N5875 & N5865;
  assign N3045 = N5875 & N5866;
  assign N3044 = N5875 & N5867;
  assign N3043 = N5875 & N5868;
  assign N3042 = N5859 & N5885;
  assign N3041 = N5859 & N5886;
  assign N3040 = N5859 & N5887;
  assign N3039 = N5859 & N5864;
  assign N3038 = N5859 & N5865;
  assign N3037 = N5859 & N5866;
  assign N3036 = N5859 & N5867;
  assign N3035 = N5859 & N5868;
  assign N3034 = N5860 & N5885;
  assign N3033 = N5860 & N5886;
  assign N3032 = N5860 & N5887;
  assign N3031 = N5860 & N5864;
  assign N3030 = N5860 & N5865;
  assign N3029 = N5860 & N5866;
  assign N3028 = N5860 & N5867;
  assign N3027 = N5860 & N5868;
  assign N3026 = N5861 & N5885;
  assign N3025 = N5861 & N5886;
  assign N3024 = N5861 & N5887;
  assign N3023 = N5861 & N5864;
  assign N3022 = N5861 & N5865;
  assign N3021 = N5861 & N5866;
  assign N3020 = N5861 & N5867;
  assign N3019 = N5861 & N5868;
  assign N3018 = N5862 & N5885;
  assign N3017 = N5862 & N5886;
  assign N3016 = N5862 & N5887;
  assign N3015 = N5862 & N5864;
  assign N3014 = N5862 & N5865;
  assign N3013 = N5862 & N5866;
  assign N3012 = N5862 & N5867;
  assign N3011 = N5862 & N5868;
  assign N3010 = N5863 & N5885;
  assign N3009 = N5863 & N5886;
  assign N3008 = N5863 & N5887;
  assign N3007 = N5863 & N5864;
  assign N3006 = N5863 & N5865;
  assign N3005 = N5863 & N5866;
  assign N3004 = N5863 & N5867;
  assign N3003 = N5863 & N5868;
  assign N5869 = addr_i[3] & addr_i[4];
  assign N5870 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N5871 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N5872 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N5873 = addr_i[5] & N5869;
  assign N5874 = addr_i[5] & N5870;
  assign N5875 = addr_i[5] & N5871;
  assign N5876 = addr_i[5] & N5872;
  assign N5877 = N5825 & N5869;
  assign N5878 = N5825 & N5870;
  assign N5879 = N5825 & N5871;
  assign N5880 = N5825 & N5872;
  assign N5881 = addr_i[0] & addr_i[1];
  assign N5882 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N5883 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N5884 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N5885 = addr_i[2] & N5881;
  assign N5886 = addr_i[2] & N5882;
  assign N5887 = addr_i[2] & N5883;
  assign N5888 = addr_i[2] & N5884;
  assign N5889 = N5830 & N5881;
  assign N5890 = N5830 & N5882;
  assign N5891 = N5830 & N5883;
  assign N5892 = N5830 & N5884;
  assign N3186 = N5873 & N5885;
  assign N3185 = N5873 & N5886;
  assign N3184 = N5873 & N5887;
  assign N3183 = N5873 & N5888;
  assign N3182 = N5873 & N5889;
  assign N3181 = N5873 & N5890;
  assign N3180 = N5873 & N5891;
  assign N3179 = N5873 & N5892;
  assign N3178 = N5874 & N5885;
  assign N3177 = N5874 & N5886;
  assign N3176 = N5874 & N5887;
  assign N3175 = N5874 & N5888;
  assign N3174 = N5874 & N5889;
  assign N3173 = N5874 & N5890;
  assign N3172 = N5874 & N5891;
  assign N3171 = N5874 & N5892;
  assign N3170 = N5875 & N5885;
  assign N3169 = N5875 & N5886;
  assign N3168 = N5875 & N5887;
  assign N3167 = N5875 & N5888;
  assign N3166 = N5875 & N5889;
  assign N3165 = N5875 & N5890;
  assign N3164 = N5875 & N5891;
  assign N3163 = N5875 & N5892;
  assign N3162 = N5876 & N5885;
  assign N3161 = N5876 & N5886;
  assign N3160 = N5876 & N5887;
  assign N3159 = N5876 & N5888;
  assign N3158 = N5876 & N5889;
  assign N3157 = N5876 & N5890;
  assign N3156 = N5876 & N5891;
  assign N3155 = N5876 & N5892;
  assign N3154 = N5877 & N5885;
  assign N3153 = N5877 & N5886;
  assign N3152 = N5877 & N5887;
  assign N3151 = N5877 & N5888;
  assign N3150 = N5877 & N5889;
  assign N3149 = N5877 & N5890;
  assign N3148 = N5877 & N5891;
  assign N3147 = N5877 & N5892;
  assign N3146 = N5878 & N5885;
  assign N3145 = N5878 & N5886;
  assign N3144 = N5878 & N5887;
  assign N3143 = N5878 & N5888;
  assign N3142 = N5878 & N5889;
  assign N3141 = N5878 & N5890;
  assign N3140 = N5878 & N5891;
  assign N3139 = N5878 & N5892;
  assign N3138 = N5879 & N5885;
  assign N3137 = N5879 & N5886;
  assign N3136 = N5879 & N5887;
  assign N3135 = N5879 & N5888;
  assign N3134 = N5879 & N5889;
  assign N3133 = N5879 & N5890;
  assign N3132 = N5879 & N5891;
  assign N3131 = N5879 & N5892;
  assign N3130 = N5880 & N5885;
  assign N3129 = N5880 & N5886;
  assign N3128 = N5880 & N5887;
  assign N3127 = N5880 & N5888;
  assign N3126 = N5880 & N5889;
  assign N3125 = N5880 & N5890;
  assign N3124 = N5880 & N5891;
  assign N3123 = N5880 & N5892;
  assign { N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182 } = (N8)? { N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N3159, N878, N877, N876, N875, N388, N387, N386, N874, N1220, N1219, N1218, N1217, N385, N384, N383, N873, N1212, N1211, N1210, N1209, N382, N381, N380, N872, N1204, N1203, N1202, N1201, N379, N378, N377, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N181)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247 } = (N9)? { N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N3159, N878, N877, N876, N875, N388, N387, N386, N874, N1220, N1219, N1218, N1217, N385, N384, N383, N873, N1212, N1211, N1210, N1209, N382, N381, N380, N872, N1204, N1203, N1202, N1201, N379, N378, N377, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N246)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312 } = (N10)? { N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N3159, N878, N877, N876, N875, N388, N387, N386, N874, N1220, N1219, N1218, N1217, N385, N384, N383, N873, N1212, N1211, N1210, N1209, N382, N381, N380, N872, N1204, N1203, N1202, N1201, N379, N378, N377, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N311)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416 } = (N11)? { N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N3159, N878, N877, N876, N875, N388, N387, N386, N874, N1220, N1219, N1218, N1217, N385, N384, N383, N873, N1212, N1211, N1210, N1209, N382, N381, N380, N872, N1204, N1203, N1202, N1201, N379, N378, N377, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N376)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = w_mask_i[3];
  assign { N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481 } = (N12)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N480)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[4];
  assign { N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546 } = (N13)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N545)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[5];
  assign { N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611 } = (N14)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N610)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[6];
  assign { N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676 } = (N15)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N675)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = w_mask_i[7];
  assign { N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741 } = (N16)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N740)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = w_mask_i[8];
  assign { N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806 } = (N17)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N805)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = w_mask_i[9];
  assign { N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885 } = (N18)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N870)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = w_mask_i[10];
  assign { N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950 } = (N19)? { N1344, N1343, N1342, N1341, N1127, N1126, N1125, N1124, N1336, N1335, N1334, N1333, N1123, N1122, N1121, N1120, N1328, N1327, N1326, N1325, N1119, N1118, N1117, N1116, N1320, N1319, N1318, N3039, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                            (N949)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = w_mask_i[11];
  assign { N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015 } = (N20)? { N1344, N1343, N1342, N1341, N1127, N1126, N1125, N1124, N1336, N1335, N1334, N1333, N1123, N1122, N1121, N1120, N1328, N1327, N1326, N1325, N1119, N1118, N1117, N1116, N1320, N1319, N1318, N3039, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1014)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = w_mask_i[12];
  assign { N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128 } = (N21)? { N1344, N1343, N1342, N1341, N1127, N1126, N1125, N1124, N1336, N1335, N1334, N1333, N1123, N1122, N1121, N1120, N1328, N1327, N1326, N1325, N1119, N1118, N1117, N1116, N1320, N1319, N1318, N3039, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1079)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = w_mask_i[13];
  assign { N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241 } = (N22)? { N1344, N1343, N1342, N1341, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N1333, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N1325, N1232, N1231, N1230, N1229, N1320, N1319, N1318, N3039, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1192)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = w_mask_i[14];
  assign { N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345 } = (N23)? { N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N3039, N1742, N1741, N1740, N1739, N1317, N1316, N1315, N1738, N3150, N3149, N3148, N3147, N1314, N1313, N1312, N1737, N3142, N3141, N3140, N3139, N1311, N1310, N1309, N1736, N3134, N3133, N3132, N3131, N1308, N1307, N1306, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1305)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N23 = w_mask_i[15];
  assign { N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410 } = (N24)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1409)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N24 = w_mask_i[16];
  assign { N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475 } = (N25)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1474)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = w_mask_i[17];
  assign { N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540 } = (N26)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1539)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = w_mask_i[18];
  assign { N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605 } = (N27)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1604)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N27 = w_mask_i[19];
  assign { N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670 } = (N28)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1669)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N28 = w_mask_i[20];
  assign { N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749 } = (N29)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1734)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = w_mask_i[21];
  assign { N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814 } = (N30)? { N2209, N2208, N2207, N2206, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N2198, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N2190, N2032, N2031, N2030, N2029, N2185, N2184, N2183, N2919, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N2017, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N2013, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N2009, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1813)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N30 = w_mask_i[22];
  assign { N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879 } = (N31)? { N2209, N2208, N2207, N2206, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N2198, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N2190, N2032, N2031, N2030, N2029, N2185, N2184, N2183, N2919, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N2017, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N2013, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N2009, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1878)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N31 = w_mask_i[23];
  assign { N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944 } = (N32)? { N2209, N2208, N2207, N2206, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N2198, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N2190, N2032, N2031, N2030, N2029, N2185, N2184, N2183, N2919, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N2017, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N2013, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N2009, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1943)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = w_mask_i[24];
  assign { N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041 } = (N33)? { N2209, N2208, N2207, N2206, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N2198, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N2190, N2032, N2031, N2030, N2029, N2185, N2184, N2183, N2919, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N2017, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N2013, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N2009, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2008)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = w_mask_i[25];
  assign { N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106 } = (N34)? { N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2919, N2542, N2541, N2540, N2539, N2182, N2181, N2180, N2538, N3030, N3029, N3028, N3027, N2179, N2178, N2177, N2537, N3022, N3021, N3020, N3019, N2176, N2175, N2174, N2536, N3014, N3013, N3012, N3011, N2173, N2172, N2171, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2105)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34 = w_mask_i[26];
  assign { N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210 } = (N35)? { N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2919, N2542, N2541, N2540, N2539, N2182, N2181, N2180, N2538, N3030, N3029, N3028, N3027, N2179, N2178, N2177, N2537, N3022, N3021, N3020, N3019, N2176, N2175, N2174, N2536, N3014, N3013, N3012, N3011, N2173, N2172, N2171, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2170)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N35 = w_mask_i[27];
  assign { N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275 } = (N36)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2274)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N36 = w_mask_i[28];
  assign { N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340 } = (N37)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2339)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N37 = w_mask_i[29];
  assign { N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405 } = (N38)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2404)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N38 = w_mask_i[30];
  assign { N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470 } = (N39)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2469)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N39 = w_mask_i[31];
  assign { N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543 } = (N40)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = w_mask_i[32];
  assign { N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608 } = (N41)? { N3186, N3185, N3184, N2817, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2816, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2815, N3046, N3045, N3044, N3043, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N3034, N3033, N3032, N2806, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2805, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2804, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2803, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2607)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N41 = w_mask_i[33];
  assign { N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673 } = (N42)? { N3186, N3185, N3184, N2817, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2816, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2815, N3046, N3045, N3044, N3043, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N3034, N3033, N3032, N2806, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2805, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2804, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2803, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2672)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N42 = w_mask_i[34];
  assign { N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738 } = (N43)? { N3186, N3185, N3184, N2817, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2816, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2815, N3046, N3045, N3044, N3043, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N3034, N3033, N3032, N2806, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2805, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2804, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2803, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2737)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N43 = w_mask_i[35];
  assign { N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818 } = (N44)? { N3186, N3185, N3184, N2817, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2816, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2815, N3046, N3045, N3044, N3043, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N3034, N3033, N3032, N2806, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2805, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2804, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2803, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2802)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N44 = w_mask_i[36];
  assign { N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938 } = (N45)? { N3186, N3185, N3184, N2937, N2936, N2935, N2934, N2933, N3178, N3177, N3176, N2932, N2931, N2930, N2929, N2928, N3170, N3169, N3168, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2882)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N45 = w_mask_i[37];
  assign { N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058 } = (N46)? { N3186, N3185, N3184, N3057, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N3052, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3002)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N46 = w_mask_i[38];
  assign { N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N3226, N3225, N3224, N3223, N3222, N3221, N3220, N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187 } = (N47)? { N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3122)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N47 = w_mask_i[39];
  assign { N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721, N5720, N5719, N5718, N5717, N5716, N5715, N5714, N5713, N5712, N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, N5691, N5690, N5689, N5688, N5687, N5686, N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, N5676, N5675, N5674, N5673, N5672, N5671, N5670, N5669, N5668, N5667, N5666, N5665, N5664, N5663, N5662, N5661, N5660, N5659, N5658, N5657, N5656, N5655, N5654, N5653, N5652, N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642, N5641, N5640, N5639, N5638, N5637, N5636, N5635, N5634, N5633, N5632, N5631, N5630, N5629, N5628, N5627, N5626, N5625, N5624, N5623, N5622, N5621, N5620, N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589, N5588, N5587, N5586, N5585, N5584, N5583, N5582, N5581, N5580, N5579, N5578, N5577, N5576, N5575, N5574, N5573, N5572, N5571, N5570, N5569, N5568, N5567, N5566, N5565, N5564, N5563, N5562, N5561, N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524, N5523, N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459, N5458, N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432, N5431, N5430, N5429, N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419, N5418, N5417, N5416, N5415, N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, N4849, N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360, N4359, N4358, N4357, N4356, N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4127, N4126, N4125, N4124, N4123, N4122, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086, N4085, N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074, N4073, N4072, N4071, N4070, N4069, N4068, N4067, N4066, N4065, N4064, N4063, N4062, N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251 } = (N48)? { N3250, N3121, N3001, N2881, N2801, N2736, N2671, N2606, N2533, N2468, N2403, N2338, N2273, N2169, N2104, N2007, N1942, N1877, N1812, N1733, N1668, N1603, N1538, N1473, N1408, N1304, N1191, N1078, N1013, N948, N869, N804, N739, N674, N609, N544, N479, N375, N310, N245, N3249, N3120, N3000, N2880, N2800, N2735, N2670, N2605, N2532, N2467, N2402, N2337, N2272, N2168, N2103, N2006, N1941, N1876, N1811, N1732, N1667, N1602, N1537, N1472, N1407, N1303, N1190, N1077, N1012, N947, N868, N803, N738, N673, N608, N543, N478, N374, N309, N244, N3248, N3119, N2999, N2879, N2799, N2734, N2669, N2604, N2531, N2466, N2401, N2336, N2271, N2167, N2102, N2005, N1940, N1875, N1810, N1731, N1666, N1601, N1536, N1471, N1406, N1302, N1189, N1076, N1011, N946, N867, N802, N737, N672, N607, N542, N477, N373, N308, N243, N3247, N3118, N2998, N2878, N2798, N2733, N2668, N2603, N2530, N2465, N2400, N2335, N2270, N2166, N2101, N2004, N1939, N1874, N1809, N1730, N1665, N1600, N1535, N1470, N1405, N1301, N1188, N1075, N1010, N945, N866, N801, N736, N671, N606, N541, N476, N372, N307, N242, N3246, N3117, N2997, N2877, N2797, N2732, N2667, N2602, N2529, N2464, N2399, N2334, N2269, N2165, N2100, N2003, N1938, N1873, N1808, N1729, N1664, N1599, N1534, N1469, N1404, N1300, N1187, N1074, N1009, N944, N865, N800, N735, N670, N605, N540, N475, N371, N306, N241, N3245, N3116, N2996, N2876, N2796, N2731, N2666, N2601, N2528, N2463, N2398, N2333, N2268, N2164, N2099, N2002, N1937, N1872, N1807, N1728, N1663, N1598, N1533, N1468, N1403, N1299, N1186, N1073, N1008, N943, N864, N799, N734, N669, N604, N539, N474, N370, N305, N240, N3244, N3115, N2995, N2875, N2795, N2730, N2665, N2600, N2527, N2462, N2397, N2332, N2267, N2163, N2098, N2001, N1936, N1871, N1806, N1727, N1662, N1597, N1532, N1467, N1402, N1298, N1185, N1072, N1007, N942, N863, N798, N733, N668, N603, N538, N473, N369, N304, N239, N3243, N3114, N2994, N2874, N2794, N2729, N2664, N2599, N2526, N2461, N2396, N2331, N2266, N2162, N2097, N2000, N1935, N1870, N1805, N1726, N1661, N1596, N1531, N1466, N1401, N1297, N1184, N1071, N1006, N941, N862, N797, N732, N667, N602, N537, N472, N368, N303, N238, N3242, N3113, N2993, N2873, N2793, N2728, N2663, N2598, N2525, N2460, N2395, N2330, N2265, N2161, N2096, N1999, N1934, N1869, N1804, N1725, N1660, N1595, N1530, N1465, N1400, N1296, N1183, N1070, N1005, N940, N861, N796, N731, N666, N601, N536, N471, N367, N302, N237, N3241, N3112, N2992, N2872, N2792, N2727, N2662, N2597, N2524, N2459, N2394, N2329, N2264, N2160, N2095, N1998, N1933, N1868, N1803, N1724, N1659, N1594, N1529, N1464, N1399, N1295, N1182, N1069, N1004, N939, N860, N795, N730, N665, N600, N535, N470, N366, N301, N236, N3240, N3111, N2991, N2871, N2791, N2726, N2661, N2596, N2523, N2458, N2393, N2328, N2263, N2159, N2094, N1997, N1932, N1867, N1802, N1723, N1658, N1593, N1528, N1463, N1398, N1294, N1181, N1068, N1003, N938, N859, N794, N729, N664, N599, N534, N469, N365, N300, N235, N3239, N3110, N2990, N2870, N2790, N2725, N2660, N2595, N2522, N2457, N2392, N2327, N2262, N2158, N2093, N1996, N1931, N1866, N1801, N1722, N1657, N1592, N1527, N1462, N1397, N1293, N1180, N1067, N1002, N937, N858, N793, N728, N663, N598, N533, N468, N364, N299, N234, N3238, N3109, N2989, N2869, N2789, N2724, N2659, N2594, N2521, N2456, N2391, N2326, N2261, N2157, N2092, N1995, N1930, N1865, N1800, N1721, N1656, N1591, N1526, N1461, N1396, N1292, N1179, N1066, N1001, N936, N857, N792, N727, N662, N597, N532, N467, N363, N298, N233, N3237, N3108, N2988, N2868, N2788, N2723, N2658, N2593, N2520, N2455, N2390, N2325, N2260, N2156, N2091, N1994, N1929, N1864, N1799, N1720, N1655, N1590, N1525, N1460, N1395, N1291, N1178, N1065, N1000, N935, N856, N791, N726, N661, N596, N531, N466, N362, N297, N232, N3236, N3107, N2987, N2867, N2787, N2722, N2657, N2592, N2519, N2454, N2389, N2324, N2259, N2155, N2090, N1993, N1928, N1863, N1798, N1719, N1654, N1589, N1524, N1459, N1394, N1290, N1177, N1064, N999, N934, N855, N790, N725, N660, N595, N530, N465, N361, N296, N231, N3235, N3106, N2986, N2866, N2786, N2721, N2656, N2591, N2518, N2453, N2388, N2323, N2258, N2154, N2089, N1992, N1927, N1862, N1797, N1718, N1653, N1588, N1523, N1458, N1393, N1289, N1176, N1063, N998, N933, N854, N789, N724, N659, N594, N529, N464, N360, N295, N230, N3234, N3105, N2985, N2865, N2785, N2720, N2655, N2590, N2517, N2452, N2387, N2322, N2257, N2153, N2088, N1991, N1926, N1861, N1796, N1717, N1652, N1587, N1522, N1457, N1392, N1288, N1175, N1062, N997, N932, N853, N788, N723, N658, N593, N528, N463, N359, N294, N229, N3233, N3104, N2984, N2864, N2784, N2719, N2654, N2589, N2516, N2451, N2386, N2321, N2256, N2152, N2087, N1990, N1925, N1860, N1795, N1716, N1651, N1586, N1521, N1456, N1391, N1287, N1174, N1061, N996, N931, N852, N787, N722, N657, N592, N527, N462, N358, N293, N228, N3232, N3103, N2983, N2863, N2783, N2718, N2653, N2588, N2515, N2450, N2385, N2320, N2255, N2151, N2086, N1989, N1924, N1859, N1794, N1715, N1650, N1585, N1520, N1455, N1390, N1286, N1173, N1060, N995, N930, N851, N786, N721, N656, N591, N526, N461, N357, N292, N227, N3231, N3102, N2982, N2862, N2782, N2717, N2652, N2587, N2514, N2449, N2384, N2319, N2254, N2150, N2085, N1988, N1923, N1858, N1793, N1714, N1649, N1584, N1519, N1454, N1389, N1285, N1172, N1059, N994, N929, N850, N785, N720, N655, N590, N525, N460, N356, N291, N226, N3230, N3101, N2981, N2861, N2781, N2716, N2651, N2586, N2513, N2448, N2383, N2318, N2253, N2149, N2084, N1987, N1922, N1857, N1792, N1713, N1648, N1583, N1518, N1453, N1388, N1284, N1171, N1058, N993, N928, N849, N784, N719, N654, N589, N524, N459, N355, N290, N225, N3229, N3100, N2980, N2860, N2780, N2715, N2650, N2585, N2512, N2447, N2382, N2317, N2252, N2148, N2083, N1986, N1921, N1856, N1791, N1712, N1647, N1582, N1517, N1452, N1387, N1283, N1170, N1057, N992, N927, N848, N783, N718, N653, N588, N523, N458, N354, N289, N224, N3228, N3099, N2979, N2859, N2779, N2714, N2649, N2584, N2511, N2446, N2381, N2316, N2251, N2147, N2082, N1985, N1920, N1855, N1790, N1711, N1646, N1581, N1516, N1451, N1386, N1282, N1169, N1056, N991, N926, N847, N782, N717, N652, N587, N522, N457, N353, N288, N223, N3227, N3098, N2978, N2858, N2778, N2713, N2648, N2583, N2510, N2445, N2380, N2315, N2250, N2146, N2081, N1984, N1919, N1854, N1789, N1710, N1645, N1580, N1515, N1450, N1385, N1281, N1168, N1055, N990, N925, N846, N781, N716, N651, N586, N521, N456, N352, N287, N222, N3226, N3097, N2977, N2857, N2777, N2712, N2647, N2582, N2509, N2444, N2379, N2314, N2249, N2145, N2080, N1983, N1918, N1853, N1788, N1709, N1644, N1579, N1514, N1449, N1384, N1280, N1167, N1054, N989, N924, N845, N780, N715, N650, N585, N520, N455, N351, N286, N221, N3225, N3096, N2976, N2856, N2776, N2711, N2646, N2581, N2508, N2443, N2378, N2313, N2248, N2144, N2079, N1982, N1917, N1852, N1787, N1708, N1643, N1578, N1513, N1448, N1383, N1279, N1166, N1053, N988, N923, N844, N779, N714, N649, N584, N519, N454, N350, N285, N220, N3224, N3095, N2975, N2855, N2775, N2710, N2645, N2580, N2507, N2442, N2377, N2312, N2247, N2143, N2078, N1981, N1916, N1851, N1786, N1707, N1642, N1577, N1512, N1447, N1382, N1278, N1165, N1052, N987, N922, N843, N778, N713, N648, N583, N518, N453, N349, N284, N219, N3223, N3094, N2974, N2854, N2774, N2709, N2644, N2579, N2506, N2441, N2376, N2311, N2246, N2142, N2077, N1980, N1915, N1850, N1785, N1706, N1641, N1576, N1511, N1446, N1381, N1277, N1164, N1051, N986, N921, N842, N777, N712, N647, N582, N517, N452, N348, N283, N218, N3222, N3093, N2973, N2853, N2773, N2708, N2643, N2578, N2505, N2440, N2375, N2310, N2245, N2141, N2076, N1979, N1914, N1849, N1784, N1705, N1640, N1575, N1510, N1445, N1380, N1276, N1163, N1050, N985, N920, N841, N776, N711, N646, N581, N516, N451, N347, N282, N217, N3221, N3092, N2972, N2852, N2772, N2707, N2642, N2577, N2504, N2439, N2374, N2309, N2244, N2140, N2075, N1978, N1913, N1848, N1783, N1704, N1639, N1574, N1509, N1444, N1379, N1275, N1162, N1049, N984, N919, N840, N775, N710, N645, N580, N515, N450, N346, N281, N216, N3220, N3091, N2971, N2851, N2771, N2706, N2641, N2576, N2503, N2438, N2373, N2308, N2243, N2139, N2074, N1977, N1912, N1847, N1782, N1703, N1638, N1573, N1508, N1443, N1378, N1274, N1161, N1048, N983, N918, N839, N774, N709, N644, N579, N514, N449, N345, N280, N215, N3219, N3090, N2970, N2850, N2770, N2705, N2640, N2575, N2502, N2437, N2372, N2307, N2242, N2138, N2073, N1976, N1911, N1846, N1781, N1702, N1637, N1572, N1507, N1442, N1377, N1273, N1160, N1047, N982, N917, N838, N773, N708, N643, N578, N513, N448, N344, N279, N214, N3218, N3089, N2969, N2849, N2769, N2704, N2639, N2574, N2501, N2436, N2371, N2306, N2241, N2137, N2072, N1975, N1910, N1845, N1780, N1701, N1636, N1571, N1506, N1441, N1376, N1272, N1159, N1046, N981, N916, N837, N772, N707, N642, N577, N512, N447, N343, N278, N213, N3217, N3088, N2968, N2848, N2768, N2703, N2638, N2573, N2500, N2435, N2370, N2305, N2240, N2136, N2071, N1974, N1909, N1844, N1779, N1700, N1635, N1570, N1505, N1440, N1375, N1271, N1158, N1045, N980, N915, N836, N771, N706, N641, N576, N511, N446, N342, N277, N212, N3216, N3087, N2967, N2847, N2767, N2702, N2637, N2572, N2499, N2434, N2369, N2304, N2239, N2135, N2070, N1973, N1908, N1843, N1778, N1699, N1634, N1569, N1504, N1439, N1374, N1270, N1157, N1044, N979, N914, N835, N770, N705, N640, N575, N510, N445, N341, N276, N211, N3215, N3086, N2966, N2846, N2766, N2701, N2636, N2571, N2498, N2433, N2368, N2303, N2238, N2134, N2069, N1972, N1907, N1842, N1777, N1698, N1633, N1568, N1503, N1438, N1373, N1269, N1156, N1043, N978, N913, N834, N769, N704, N639, N574, N509, N444, N340, N275, N210, N3214, N3085, N2965, N2845, N2765, N2700, N2635, N2570, N2497, N2432, N2367, N2302, N2237, N2133, N2068, N1971, N1906, N1841, N1776, N1697, N1632, N1567, N1502, N1437, N1372, N1268, N1155, N1042, N977, N912, N833, N768, N703, N638, N573, N508, N443, N339, N274, N209, N3213, N3084, N2964, N2844, N2764, N2699, N2634, N2569, N2496, N2431, N2366, N2301, N2236, N2132, N2067, N1970, N1905, N1840, N1775, N1696, N1631, N1566, N1501, N1436, N1371, N1267, N1154, N1041, N976, N911, N832, N767, N702, N637, N572, N507, N442, N338, N273, N208, N3212, N3083, N2963, N2843, N2763, N2698, N2633, N2568, N2495, N2430, N2365, N2300, N2235, N2131, N2066, N1969, N1904, N1839, N1774, N1695, N1630, N1565, N1500, N1435, N1370, N1266, N1153, N1040, N975, N910, N831, N766, N701, N636, N571, N506, N441, N337, N272, N207, N3211, N3082, N2962, N2842, N2762, N2697, N2632, N2567, N2494, N2429, N2364, N2299, N2234, N2130, N2065, N1968, N1903, N1838, N1773, N1694, N1629, N1564, N1499, N1434, N1369, N1265, N1152, N1039, N974, N909, N830, N765, N700, N635, N570, N505, N440, N336, N271, N206, N3210, N3081, N2961, N2841, N2761, N2696, N2631, N2566, N2493, N2428, N2363, N2298, N2233, N2129, N2064, N1967, N1902, N1837, N1772, N1693, N1628, N1563, N1498, N1433, N1368, N1264, N1151, N1038, N973, N908, N829, N764, N699, N634, N569, N504, N439, N335, N270, N205, N3209, N3080, N2960, N2840, N2760, N2695, N2630, N2565, N2492, N2427, N2362, N2297, N2232, N2128, N2063, N1966, N1901, N1836, N1771, N1692, N1627, N1562, N1497, N1432, N1367, N1263, N1150, N1037, N972, N907, N828, N763, N698, N633, N568, N503, N438, N334, N269, N204, N3208, N3079, N2959, N2839, N2759, N2694, N2629, N2564, N2491, N2426, N2361, N2296, N2231, N2127, N2062, N1965, N1900, N1835, N1770, N1691, N1626, N1561, N1496, N1431, N1366, N1262, N1149, N1036, N971, N906, N827, N762, N697, N632, N567, N502, N437, N333, N268, N203, N3207, N3078, N2958, N2838, N2758, N2693, N2628, N2563, N2490, N2425, N2360, N2295, N2230, N2126, N2061, N1964, N1899, N1834, N1769, N1690, N1625, N1560, N1495, N1430, N1365, N1261, N1148, N1035, N970, N905, N826, N761, N696, N631, N566, N501, N436, N332, N267, N202, N3206, N3077, N2957, N2837, N2757, N2692, N2627, N2562, N2489, N2424, N2359, N2294, N2229, N2125, N2060, N1963, N1898, N1833, N1768, N1689, N1624, N1559, N1494, N1429, N1364, N1260, N1147, N1034, N969, N904, N825, N760, N695, N630, N565, N500, N435, N331, N266, N201, N3205, N3076, N2956, N2836, N2756, N2691, N2626, N2561, N2488, N2423, N2358, N2293, N2228, N2124, N2059, N1962, N1897, N1832, N1767, N1688, N1623, N1558, N1493, N1428, N1363, N1259, N1146, N1033, N968, N903, N824, N759, N694, N629, N564, N499, N434, N330, N265, N200, N3204, N3075, N2955, N2835, N2755, N2690, N2625, N2560, N2487, N2422, N2357, N2292, N2227, N2123, N2058, N1961, N1896, N1831, N1766, N1687, N1622, N1557, N1492, N1427, N1362, N1258, N1145, N1032, N967, N902, N823, N758, N693, N628, N563, N498, N433, N329, N264, N199, N3203, N3074, N2954, N2834, N2754, N2689, N2624, N2559, N2486, N2421, N2356, N2291, N2226, N2122, N2057, N1960, N1895, N1830, N1765, N1686, N1621, N1556, N1491, N1426, N1361, N1257, N1144, N1031, N966, N901, N822, N757, N692, N627, N562, N497, N432, N328, N263, N198, N3202, N3073, N2953, N2833, N2753, N2688, N2623, N2558, N2485, N2420, N2355, N2290, N2225, N2121, N2056, N1959, N1894, N1829, N1764, N1685, N1620, N1555, N1490, N1425, N1360, N1256, N1143, N1030, N965, N900, N821, N756, N691, N626, N561, N496, N431, N327, N262, N197, N3201, N3072, N2952, N2832, N2752, N2687, N2622, N2557, N2484, N2419, N2354, N2289, N2224, N2120, N2055, N1958, N1893, N1828, N1763, N1684, N1619, N1554, N1489, N1424, N1359, N1255, N1142, N1029, N964, N899, N820, N755, N690, N625, N560, N495, N430, N326, N261, N196, N3200, N3071, N2951, N2831, N2751, N2686, N2621, N2556, N2483, N2418, N2353, N2288, N2223, N2119, N2054, N1957, N1892, N1827, N1762, N1683, N1618, N1553, N1488, N1423, N1358, N1254, N1141, N1028, N963, N898, N819, N754, N689, N624, N559, N494, N429, N325, N260, N195, N3199, N3070, N2950, N2830, N2750, N2685, N2620, N2555, N2482, N2417, N2352, N2287, N2222, N2118, N2053, N1956, N1891, N1826, N1761, N1682, N1617, N1552, N1487, N1422, N1357, N1253, N1140, N1027, N962, N897, N818, N753, N688, N623, N558, N493, N428, N324, N259, N194, N3198, N3069, N2949, N2829, N2749, N2684, N2619, N2554, N2481, N2416, N2351, N2286, N2221, N2117, N2052, N1955, N1890, N1825, N1760, N1681, N1616, N1551, N1486, N1421, N1356, N1252, N1139, N1026, N961, N896, N817, N752, N687, N622, N557, N492, N427, N323, N258, N193, N3197, N3068, N2948, N2828, N2748, N2683, N2618, N2553, N2480, N2415, N2350, N2285, N2220, N2116, N2051, N1954, N1889, N1824, N1759, N1680, N1615, N1550, N1485, N1420, N1355, N1251, N1138, N1025, N960, N895, N816, N751, N686, N621, N556, N491, N426, N322, N257, N192, N3196, N3067, N2947, N2827, N2747, N2682, N2617, N2552, N2479, N2414, N2349, N2284, N2219, N2115, N2050, N1953, N1888, N1823, N1758, N1679, N1614, N1549, N1484, N1419, N1354, N1250, N1137, N1024, N959, N894, N815, N750, N685, N620, N555, N490, N425, N321, N256, N191, N3195, N3066, N2946, N2826, N2746, N2681, N2616, N2551, N2478, N2413, N2348, N2283, N2218, N2114, N2049, N1952, N1887, N1822, N1757, N1678, N1613, N1548, N1483, N1418, N1353, N1249, N1136, N1023, N958, N893, N814, N749, N684, N619, N554, N489, N424, N320, N255, N190, N3194, N3065, N2945, N2825, N2745, N2680, N2615, N2550, N2477, N2412, N2347, N2282, N2217, N2113, N2048, N1951, N1886, N1821, N1756, N1677, N1612, N1547, N1482, N1417, N1352, N1248, N1135, N1022, N957, N892, N813, N748, N683, N618, N553, N488, N423, N319, N254, N189, N3193, N3064, N2944, N2824, N2744, N2679, N2614, N2549, N2476, N2411, N2346, N2281, N2216, N2112, N2047, N1950, N1885, N1820, N1755, N1676, N1611, N1546, N1481, N1416, N1351, N1247, N1134, N1021, N956, N891, N812, N747, N682, N617, N552, N487, N422, N318, N253, N188, N3192, N3063, N2943, N2823, N2743, N2678, N2613, N2548, N2475, N2410, N2345, N2280, N2215, N2111, N2046, N1949, N1884, N1819, N1754, N1675, N1610, N1545, N1480, N1415, N1350, N1246, N1133, N1020, N955, N890, N811, N746, N681, N616, N551, N486, N421, N317, N252, N187, N3191, N3062, N2942, N2822, N2742, N2677, N2612, N2547, N2474, N2409, N2344, N2279, N2214, N2110, N2045, N1948, N1883, N1818, N1753, N1674, N1609, N1544, N1479, N1414, N1349, N1245, N1132, N1019, N954, N889, N810, N745, N680, N615, N550, N485, N420, N316, N251, N186, N3190, N3061, N2941, N2821, N2741, N2676, N2611, N2546, N2473, N2408, N2343, N2278, N2213, N2109, N2044, N1947, N1882, N1817, N1752, N1673, N1608, N1543, N1478, N1413, N1348, N1244, N1131, N1018, N953, N888, N809, N744, N679, N614, N549, N484, N419, N315, N250, N185, N3189, N3060, N2940, N2820, N2740, N2675, N2610, N2545, N2472, N2407, N2342, N2277, N2212, N2108, N2043, N1946, N1881, N1816, N1751, N1672, N1607, N1542, N1477, N1412, N1347, N1243, N1130, N1017, N952, N887, N808, N743, N678, N613, N548, N483, N418, N314, N249, N184, N3188, N3059, N2939, N2819, N2739, N2674, N2609, N2544, N2471, N2406, N2341, N2276, N2211, N2107, N2042, N1945, N1880, N1815, N1750, N1671, N1606, N1541, N1476, N1411, N1346, N1242, N1129, N1016, N951, N886, N807, N742, N677, N612, N547, N482, N417, N313, N248, N183, N3187, N3058, N2938, N2818, N2738, N2673, N2608, N2543, N2470, N2405, N2340, N2275, N2210, N2106, N2041, N1944, N1879, N1814, N1749, N1670, N1605, N1540, N1475, N1410, N1345, N1241, N1128, N1015, N950, N885, N806, N741, N676, N611, N546, N481, N416, N312, N247, N182 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N180)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = N179;
  assign read_en = v_i & N5893;
  assign N5893 = ~w_i;
  assign N49 = ~addr_r[0];
  assign N50 = ~addr_r[1];
  assign N51 = N49 & N50;
  assign N52 = N49 & addr_r[1];
  assign N53 = addr_r[0] & N50;
  assign N54 = addr_r[0] & addr_r[1];
  assign N55 = ~addr_r[2];
  assign N56 = N51 & N55;
  assign N57 = N51 & addr_r[2];
  assign N58 = N53 & N55;
  assign N59 = N53 & addr_r[2];
  assign N60 = N52 & N55;
  assign N61 = N52 & addr_r[2];
  assign N62 = N54 & N55;
  assign N63 = N54 & addr_r[2];
  assign N64 = ~addr_r[3];
  assign N65 = N56 & N64;
  assign N66 = N56 & addr_r[3];
  assign N67 = N58 & N64;
  assign N68 = N58 & addr_r[3];
  assign N69 = N60 & N64;
  assign N70 = N60 & addr_r[3];
  assign N71 = N62 & N64;
  assign N72 = N62 & addr_r[3];
  assign N73 = N57 & N64;
  assign N74 = N57 & addr_r[3];
  assign N75 = N59 & N64;
  assign N76 = N59 & addr_r[3];
  assign N77 = N61 & N64;
  assign N78 = N61 & addr_r[3];
  assign N79 = N63 & N64;
  assign N80 = N63 & addr_r[3];
  assign N81 = ~addr_r[4];
  assign N82 = N65 & N81;
  assign N83 = N65 & addr_r[4];
  assign N84 = N67 & N81;
  assign N85 = N67 & addr_r[4];
  assign N86 = N69 & N81;
  assign N87 = N69 & addr_r[4];
  assign N88 = N71 & N81;
  assign N89 = N71 & addr_r[4];
  assign N90 = N73 & N81;
  assign N91 = N73 & addr_r[4];
  assign N92 = N75 & N81;
  assign N93 = N75 & addr_r[4];
  assign N94 = N77 & N81;
  assign N95 = N77 & addr_r[4];
  assign N96 = N79 & N81;
  assign N97 = N79 & addr_r[4];
  assign N98 = N66 & N81;
  assign N99 = N66 & addr_r[4];
  assign N100 = N68 & N81;
  assign N101 = N68 & addr_r[4];
  assign N102 = N70 & N81;
  assign N103 = N70 & addr_r[4];
  assign N104 = N72 & N81;
  assign N105 = N72 & addr_r[4];
  assign N106 = N74 & N81;
  assign N107 = N74 & addr_r[4];
  assign N108 = N76 & N81;
  assign N109 = N76 & addr_r[4];
  assign N110 = N78 & N81;
  assign N111 = N78 & addr_r[4];
  assign N112 = N80 & N81;
  assign N113 = N80 & addr_r[4];
  assign N114 = ~addr_r[5];
  assign N115 = N82 & N114;
  assign N116 = N82 & addr_r[5];
  assign N117 = N84 & N114;
  assign N118 = N84 & addr_r[5];
  assign N119 = N86 & N114;
  assign N120 = N86 & addr_r[5];
  assign N121 = N88 & N114;
  assign N122 = N88 & addr_r[5];
  assign N123 = N90 & N114;
  assign N124 = N90 & addr_r[5];
  assign N125 = N92 & N114;
  assign N126 = N92 & addr_r[5];
  assign N127 = N94 & N114;
  assign N128 = N94 & addr_r[5];
  assign N129 = N96 & N114;
  assign N130 = N96 & addr_r[5];
  assign N131 = N98 & N114;
  assign N132 = N98 & addr_r[5];
  assign N133 = N100 & N114;
  assign N134 = N100 & addr_r[5];
  assign N135 = N102 & N114;
  assign N136 = N102 & addr_r[5];
  assign N137 = N104 & N114;
  assign N138 = N104 & addr_r[5];
  assign N139 = N106 & N114;
  assign N140 = N106 & addr_r[5];
  assign N141 = N108 & N114;
  assign N142 = N108 & addr_r[5];
  assign N143 = N110 & N114;
  assign N144 = N110 & addr_r[5];
  assign N145 = N112 & N114;
  assign N146 = N112 & addr_r[5];
  assign N147 = N83 & N114;
  assign N148 = N83 & addr_r[5];
  assign N149 = N85 & N114;
  assign N150 = N85 & addr_r[5];
  assign N151 = N87 & N114;
  assign N152 = N87 & addr_r[5];
  assign N153 = N89 & N114;
  assign N154 = N89 & addr_r[5];
  assign N155 = N91 & N114;
  assign N156 = N91 & addr_r[5];
  assign N157 = N93 & N114;
  assign N158 = N93 & addr_r[5];
  assign N159 = N95 & N114;
  assign N160 = N95 & addr_r[5];
  assign N161 = N97 & N114;
  assign N162 = N97 & addr_r[5];
  assign N163 = N99 & N114;
  assign N164 = N99 & addr_r[5];
  assign N165 = N101 & N114;
  assign N166 = N101 & addr_r[5];
  assign N167 = N103 & N114;
  assign N168 = N103 & addr_r[5];
  assign N169 = N105 & N114;
  assign N170 = N105 & addr_r[5];
  assign N171 = N107 & N114;
  assign N172 = N107 & addr_r[5];
  assign N173 = N109 & N114;
  assign N174 = N109 & addr_r[5];
  assign N175 = N111 & N114;
  assign N176 = N111 & addr_r[5];
  assign N177 = N113 & N114;
  assign N178 = N113 & addr_r[5];
  assign N179 = v_i & w_i;
  assign N180 = ~N179;
  assign N181 = ~w_mask_i[0];
  assign N246 = ~w_mask_i[1];
  assign N311 = ~w_mask_i[2];
  assign N376 = ~w_mask_i[3];
  assign N480 = ~w_mask_i[4];
  assign N545 = ~w_mask_i[5];
  assign N610 = ~w_mask_i[6];
  assign N675 = ~w_mask_i[7];
  assign N740 = ~w_mask_i[8];
  assign N805 = ~w_mask_i[9];
  assign N870 = ~w_mask_i[10];
  assign N949 = ~w_mask_i[11];
  assign N1014 = ~w_mask_i[12];
  assign N1079 = ~w_mask_i[13];
  assign N1192 = ~w_mask_i[14];
  assign N1305 = ~w_mask_i[15];
  assign N1409 = ~w_mask_i[16];
  assign N1474 = ~w_mask_i[17];
  assign N1539 = ~w_mask_i[18];
  assign N1604 = ~w_mask_i[19];
  assign N1669 = ~w_mask_i[20];
  assign N1734 = ~w_mask_i[21];
  assign N1813 = ~w_mask_i[22];
  assign N1878 = ~w_mask_i[23];
  assign N1943 = ~w_mask_i[24];
  assign N2008 = ~w_mask_i[25];
  assign N2105 = ~w_mask_i[26];
  assign N2170 = ~w_mask_i[27];
  assign N2274 = ~w_mask_i[28];
  assign N2339 = ~w_mask_i[29];
  assign N2404 = ~w_mask_i[30];
  assign N2469 = ~w_mask_i[31];
  assign N2534 = ~w_mask_i[32];
  assign N2607 = ~w_mask_i[33];
  assign N2672 = ~w_mask_i[34];
  assign N2737 = ~w_mask_i[35];
  assign N2802 = ~w_mask_i[36];
  assign N2882 = ~w_mask_i[37];
  assign N3002 = ~w_mask_i[38];
  assign N3122 = ~w_mask_i[39];

  always @(posedge clk_i) begin
    if(1'b1) begin
      { addr_r[5:0] } <= { addr_i[5:0] };
    end 
    if(N5810) begin
      { mem[2559:2559] } <= { data_i[39:39] };
    end 
    if(N5809) begin
      { mem[2558:2558] } <= { data_i[38:38] };
    end 
    if(N5808) begin
      { mem[2557:2557] } <= { data_i[37:37] };
    end 
    if(N5807) begin
      { mem[2556:2556] } <= { data_i[36:36] };
    end 
    if(N5806) begin
      { mem[2555:2555] } <= { data_i[35:35] };
    end 
    if(N5805) begin
      { mem[2554:2554] } <= { data_i[34:34] };
    end 
    if(N5804) begin
      { mem[2553:2553] } <= { data_i[33:33] };
    end 
    if(N5803) begin
      { mem[2552:2552] } <= { data_i[32:32] };
    end 
    if(N5802) begin
      { mem[2551:2551] } <= { data_i[31:31] };
    end 
    if(N5801) begin
      { mem[2550:2550] } <= { data_i[30:30] };
    end 
    if(N5800) begin
      { mem[2549:2549] } <= { data_i[29:29] };
    end 
    if(N5799) begin
      { mem[2548:2548] } <= { data_i[28:28] };
    end 
    if(N5798) begin
      { mem[2547:2547] } <= { data_i[27:27] };
    end 
    if(N5797) begin
      { mem[2546:2546] } <= { data_i[26:26] };
    end 
    if(N5796) begin
      { mem[2545:2545] } <= { data_i[25:25] };
    end 
    if(N5795) begin
      { mem[2544:2544] } <= { data_i[24:24] };
    end 
    if(N5794) begin
      { mem[2543:2543] } <= { data_i[23:23] };
    end 
    if(N5793) begin
      { mem[2542:2542] } <= { data_i[22:22] };
    end 
    if(N5792) begin
      { mem[2541:2541] } <= { data_i[21:21] };
    end 
    if(N5791) begin
      { mem[2540:2540] } <= { data_i[20:20] };
    end 
    if(N5790) begin
      { mem[2539:2539] } <= { data_i[19:19] };
    end 
    if(N5789) begin
      { mem[2538:2538] } <= { data_i[18:18] };
    end 
    if(N5788) begin
      { mem[2537:2537] } <= { data_i[17:17] };
    end 
    if(N5787) begin
      { mem[2536:2536] } <= { data_i[16:16] };
    end 
    if(N5786) begin
      { mem[2535:2535] } <= { data_i[15:15] };
    end 
    if(N5785) begin
      { mem[2534:2534] } <= { data_i[14:14] };
    end 
    if(N5784) begin
      { mem[2533:2533] } <= { data_i[13:13] };
    end 
    if(N5783) begin
      { mem[2532:2532] } <= { data_i[12:12] };
    end 
    if(N5782) begin
      { mem[2531:2531] } <= { data_i[11:11] };
    end 
    if(N5781) begin
      { mem[2530:2530] } <= { data_i[10:10] };
    end 
    if(N5780) begin
      { mem[2529:2529] } <= { data_i[9:9] };
    end 
    if(N5779) begin
      { mem[2528:2528] } <= { data_i[8:8] };
    end 
    if(N5778) begin
      { mem[2527:2527] } <= { data_i[7:7] };
    end 
    if(N5777) begin
      { mem[2526:2526] } <= { data_i[6:6] };
    end 
    if(N5776) begin
      { mem[2525:2525] } <= { data_i[5:5] };
    end 
    if(N5775) begin
      { mem[2524:2524] } <= { data_i[4:4] };
    end 
    if(N5774) begin
      { mem[2523:2523] } <= { data_i[3:3] };
    end 
    if(N5773) begin
      { mem[2522:2522] } <= { data_i[2:2] };
    end 
    if(N5772) begin
      { mem[2521:2521] } <= { data_i[1:1] };
    end 
    if(N5771) begin
      { mem[2520:2520] } <= { data_i[0:0] };
    end 
    if(N5770) begin
      { mem[2519:2519] } <= { data_i[39:39] };
    end 
    if(N5769) begin
      { mem[2518:2518] } <= { data_i[38:38] };
    end 
    if(N5768) begin
      { mem[2517:2517] } <= { data_i[37:37] };
    end 
    if(N5767) begin
      { mem[2516:2516] } <= { data_i[36:36] };
    end 
    if(N5766) begin
      { mem[2515:2515] } <= { data_i[35:35] };
    end 
    if(N5765) begin
      { mem[2514:2514] } <= { data_i[34:34] };
    end 
    if(N5764) begin
      { mem[2513:2513] } <= { data_i[33:33] };
    end 
    if(N5763) begin
      { mem[2512:2512] } <= { data_i[32:32] };
    end 
    if(N5762) begin
      { mem[2511:2511] } <= { data_i[31:31] };
    end 
    if(N5761) begin
      { mem[2510:2510] } <= { data_i[30:30] };
    end 
    if(N5760) begin
      { mem[2509:2509] } <= { data_i[29:29] };
    end 
    if(N5759) begin
      { mem[2508:2508] } <= { data_i[28:28] };
    end 
    if(N5758) begin
      { mem[2507:2507] } <= { data_i[27:27] };
    end 
    if(N5757) begin
      { mem[2506:2506] } <= { data_i[26:26] };
    end 
    if(N5756) begin
      { mem[2505:2505] } <= { data_i[25:25] };
    end 
    if(N5755) begin
      { mem[2504:2504] } <= { data_i[24:24] };
    end 
    if(N5754) begin
      { mem[2503:2503] } <= { data_i[23:23] };
    end 
    if(N5753) begin
      { mem[2502:2502] } <= { data_i[22:22] };
    end 
    if(N5752) begin
      { mem[2501:2501] } <= { data_i[21:21] };
    end 
    if(N5751) begin
      { mem[2500:2500] } <= { data_i[20:20] };
    end 
    if(N5750) begin
      { mem[2499:2499] } <= { data_i[19:19] };
    end 
    if(N5749) begin
      { mem[2498:2498] } <= { data_i[18:18] };
    end 
    if(N5748) begin
      { mem[2497:2497] } <= { data_i[17:17] };
    end 
    if(N5747) begin
      { mem[2496:2496] } <= { data_i[16:16] };
    end 
    if(N5746) begin
      { mem[2495:2495] } <= { data_i[15:15] };
    end 
    if(N5745) begin
      { mem[2494:2494] } <= { data_i[14:14] };
    end 
    if(N5744) begin
      { mem[2493:2493] } <= { data_i[13:13] };
    end 
    if(N5743) begin
      { mem[2492:2492] } <= { data_i[12:12] };
    end 
    if(N5742) begin
      { mem[2491:2491] } <= { data_i[11:11] };
    end 
    if(N5741) begin
      { mem[2490:2490] } <= { data_i[10:10] };
    end 
    if(N5740) begin
      { mem[2489:2489] } <= { data_i[9:9] };
    end 
    if(N5739) begin
      { mem[2488:2488] } <= { data_i[8:8] };
    end 
    if(N5738) begin
      { mem[2487:2487] } <= { data_i[7:7] };
    end 
    if(N5737) begin
      { mem[2486:2486] } <= { data_i[6:6] };
    end 
    if(N5736) begin
      { mem[2485:2485] } <= { data_i[5:5] };
    end 
    if(N5735) begin
      { mem[2484:2484] } <= { data_i[4:4] };
    end 
    if(N5734) begin
      { mem[2483:2483] } <= { data_i[3:3] };
    end 
    if(N5733) begin
      { mem[2482:2482] } <= { data_i[2:2] };
    end 
    if(N5732) begin
      { mem[2481:2481] } <= { data_i[1:1] };
    end 
    if(N5731) begin
      { mem[2480:2480] } <= { data_i[0:0] };
    end 
    if(N5730) begin
      { mem[2479:2479] } <= { data_i[39:39] };
    end 
    if(N5729) begin
      { mem[2478:2478] } <= { data_i[38:38] };
    end 
    if(N5728) begin
      { mem[2477:2477] } <= { data_i[37:37] };
    end 
    if(N5727) begin
      { mem[2476:2476] } <= { data_i[36:36] };
    end 
    if(N5726) begin
      { mem[2475:2475] } <= { data_i[35:35] };
    end 
    if(N5725) begin
      { mem[2474:2474] } <= { data_i[34:34] };
    end 
    if(N5724) begin
      { mem[2473:2473] } <= { data_i[33:33] };
    end 
    if(N5723) begin
      { mem[2472:2472] } <= { data_i[32:32] };
    end 
    if(N5722) begin
      { mem[2471:2471] } <= { data_i[31:31] };
    end 
    if(N5721) begin
      { mem[2470:2470] } <= { data_i[30:30] };
    end 
    if(N5720) begin
      { mem[2469:2469] } <= { data_i[29:29] };
    end 
    if(N5719) begin
      { mem[2468:2468] } <= { data_i[28:28] };
    end 
    if(N5718) begin
      { mem[2467:2467] } <= { data_i[27:27] };
    end 
    if(N5717) begin
      { mem[2466:2466] } <= { data_i[26:26] };
    end 
    if(N5716) begin
      { mem[2465:2465] } <= { data_i[25:25] };
    end 
    if(N5715) begin
      { mem[2464:2464] } <= { data_i[24:24] };
    end 
    if(N5714) begin
      { mem[2463:2463] } <= { data_i[23:23] };
    end 
    if(N5713) begin
      { mem[2462:2462] } <= { data_i[22:22] };
    end 
    if(N5712) begin
      { mem[2461:2461] } <= { data_i[21:21] };
    end 
    if(N5711) begin
      { mem[2460:2460] } <= { data_i[20:20] };
    end 
    if(N5710) begin
      { mem[2459:2459] } <= { data_i[19:19] };
    end 
    if(N5709) begin
      { mem[2458:2458] } <= { data_i[18:18] };
    end 
    if(N5708) begin
      { mem[2457:2457] } <= { data_i[17:17] };
    end 
    if(N5707) begin
      { mem[2456:2456] } <= { data_i[16:16] };
    end 
    if(N5706) begin
      { mem[2455:2455] } <= { data_i[15:15] };
    end 
    if(N5705) begin
      { mem[2454:2454] } <= { data_i[14:14] };
    end 
    if(N5704) begin
      { mem[2453:2453] } <= { data_i[13:13] };
    end 
    if(N5703) begin
      { mem[2452:2452] } <= { data_i[12:12] };
    end 
    if(N5702) begin
      { mem[2451:2451] } <= { data_i[11:11] };
    end 
    if(N5701) begin
      { mem[2450:2450] } <= { data_i[10:10] };
    end 
    if(N5700) begin
      { mem[2449:2449] } <= { data_i[9:9] };
    end 
    if(N5699) begin
      { mem[2448:2448] } <= { data_i[8:8] };
    end 
    if(N5698) begin
      { mem[2447:2447] } <= { data_i[7:7] };
    end 
    if(N5697) begin
      { mem[2446:2446] } <= { data_i[6:6] };
    end 
    if(N5696) begin
      { mem[2445:2445] } <= { data_i[5:5] };
    end 
    if(N5695) begin
      { mem[2444:2444] } <= { data_i[4:4] };
    end 
    if(N5694) begin
      { mem[2443:2443] } <= { data_i[3:3] };
    end 
    if(N5693) begin
      { mem[2442:2442] } <= { data_i[2:2] };
    end 
    if(N5692) begin
      { mem[2441:2441] } <= { data_i[1:1] };
    end 
    if(N5691) begin
      { mem[2440:2440] } <= { data_i[0:0] };
    end 
    if(N5690) begin
      { mem[2439:2439] } <= { data_i[39:39] };
    end 
    if(N5689) begin
      { mem[2438:2438] } <= { data_i[38:38] };
    end 
    if(N5688) begin
      { mem[2437:2437] } <= { data_i[37:37] };
    end 
    if(N5687) begin
      { mem[2436:2436] } <= { data_i[36:36] };
    end 
    if(N5686) begin
      { mem[2435:2435] } <= { data_i[35:35] };
    end 
    if(N5685) begin
      { mem[2434:2434] } <= { data_i[34:34] };
    end 
    if(N5684) begin
      { mem[2433:2433] } <= { data_i[33:33] };
    end 
    if(N5683) begin
      { mem[2432:2432] } <= { data_i[32:32] };
    end 
    if(N5682) begin
      { mem[2431:2431] } <= { data_i[31:31] };
    end 
    if(N5681) begin
      { mem[2430:2430] } <= { data_i[30:30] };
    end 
    if(N5680) begin
      { mem[2429:2429] } <= { data_i[29:29] };
    end 
    if(N5679) begin
      { mem[2428:2428] } <= { data_i[28:28] };
    end 
    if(N5678) begin
      { mem[2427:2427] } <= { data_i[27:27] };
    end 
    if(N5677) begin
      { mem[2426:2426] } <= { data_i[26:26] };
    end 
    if(N5676) begin
      { mem[2425:2425] } <= { data_i[25:25] };
    end 
    if(N5675) begin
      { mem[2424:2424] } <= { data_i[24:24] };
    end 
    if(N5674) begin
      { mem[2423:2423] } <= { data_i[23:23] };
    end 
    if(N5673) begin
      { mem[2422:2422] } <= { data_i[22:22] };
    end 
    if(N5672) begin
      { mem[2421:2421] } <= { data_i[21:21] };
    end 
    if(N5671) begin
      { mem[2420:2420] } <= { data_i[20:20] };
    end 
    if(N5670) begin
      { mem[2419:2419] } <= { data_i[19:19] };
    end 
    if(N5669) begin
      { mem[2418:2418] } <= { data_i[18:18] };
    end 
    if(N5668) begin
      { mem[2417:2417] } <= { data_i[17:17] };
    end 
    if(N5667) begin
      { mem[2416:2416] } <= { data_i[16:16] };
    end 
    if(N5666) begin
      { mem[2415:2415] } <= { data_i[15:15] };
    end 
    if(N5665) begin
      { mem[2414:2414] } <= { data_i[14:14] };
    end 
    if(N5664) begin
      { mem[2413:2413] } <= { data_i[13:13] };
    end 
    if(N5663) begin
      { mem[2412:2412] } <= { data_i[12:12] };
    end 
    if(N5662) begin
      { mem[2411:2411] } <= { data_i[11:11] };
    end 
    if(N5661) begin
      { mem[2410:2410] } <= { data_i[10:10] };
    end 
    if(N5660) begin
      { mem[2409:2409] } <= { data_i[9:9] };
    end 
    if(N5659) begin
      { mem[2408:2408] } <= { data_i[8:8] };
    end 
    if(N5658) begin
      { mem[2407:2407] } <= { data_i[7:7] };
    end 
    if(N5657) begin
      { mem[2406:2406] } <= { data_i[6:6] };
    end 
    if(N5656) begin
      { mem[2405:2405] } <= { data_i[5:5] };
    end 
    if(N5655) begin
      { mem[2404:2404] } <= { data_i[4:4] };
    end 
    if(N5654) begin
      { mem[2403:2403] } <= { data_i[3:3] };
    end 
    if(N5653) begin
      { mem[2402:2402] } <= { data_i[2:2] };
    end 
    if(N5652) begin
      { mem[2401:2401] } <= { data_i[1:1] };
    end 
    if(N5651) begin
      { mem[2400:2400] } <= { data_i[0:0] };
    end 
    if(N5650) begin
      { mem[2399:2399] } <= { data_i[39:39] };
    end 
    if(N5649) begin
      { mem[2398:2398] } <= { data_i[38:38] };
    end 
    if(N5648) begin
      { mem[2397:2397] } <= { data_i[37:37] };
    end 
    if(N5647) begin
      { mem[2396:2396] } <= { data_i[36:36] };
    end 
    if(N5646) begin
      { mem[2395:2395] } <= { data_i[35:35] };
    end 
    if(N5645) begin
      { mem[2394:2394] } <= { data_i[34:34] };
    end 
    if(N5644) begin
      { mem[2393:2393] } <= { data_i[33:33] };
    end 
    if(N5643) begin
      { mem[2392:2392] } <= { data_i[32:32] };
    end 
    if(N5642) begin
      { mem[2391:2391] } <= { data_i[31:31] };
    end 
    if(N5641) begin
      { mem[2390:2390] } <= { data_i[30:30] };
    end 
    if(N5640) begin
      { mem[2389:2389] } <= { data_i[29:29] };
    end 
    if(N5639) begin
      { mem[2388:2388] } <= { data_i[28:28] };
    end 
    if(N5638) begin
      { mem[2387:2387] } <= { data_i[27:27] };
    end 
    if(N5637) begin
      { mem[2386:2386] } <= { data_i[26:26] };
    end 
    if(N5636) begin
      { mem[2385:2385] } <= { data_i[25:25] };
    end 
    if(N5635) begin
      { mem[2384:2384] } <= { data_i[24:24] };
    end 
    if(N5634) begin
      { mem[2383:2383] } <= { data_i[23:23] };
    end 
    if(N5633) begin
      { mem[2382:2382] } <= { data_i[22:22] };
    end 
    if(N5632) begin
      { mem[2381:2381] } <= { data_i[21:21] };
    end 
    if(N5631) begin
      { mem[2380:2380] } <= { data_i[20:20] };
    end 
    if(N5630) begin
      { mem[2379:2379] } <= { data_i[19:19] };
    end 
    if(N5629) begin
      { mem[2378:2378] } <= { data_i[18:18] };
    end 
    if(N5628) begin
      { mem[2377:2377] } <= { data_i[17:17] };
    end 
    if(N5627) begin
      { mem[2376:2376] } <= { data_i[16:16] };
    end 
    if(N5626) begin
      { mem[2375:2375] } <= { data_i[15:15] };
    end 
    if(N5625) begin
      { mem[2374:2374] } <= { data_i[14:14] };
    end 
    if(N5624) begin
      { mem[2373:2373] } <= { data_i[13:13] };
    end 
    if(N5623) begin
      { mem[2372:2372] } <= { data_i[12:12] };
    end 
    if(N5622) begin
      { mem[2371:2371] } <= { data_i[11:11] };
    end 
    if(N5621) begin
      { mem[2370:2370] } <= { data_i[10:10] };
    end 
    if(N5620) begin
      { mem[2369:2369] } <= { data_i[9:9] };
    end 
    if(N5619) begin
      { mem[2368:2368] } <= { data_i[8:8] };
    end 
    if(N5618) begin
      { mem[2367:2367] } <= { data_i[7:7] };
    end 
    if(N5617) begin
      { mem[2366:2366] } <= { data_i[6:6] };
    end 
    if(N5616) begin
      { mem[2365:2365] } <= { data_i[5:5] };
    end 
    if(N5615) begin
      { mem[2364:2364] } <= { data_i[4:4] };
    end 
    if(N5614) begin
      { mem[2363:2363] } <= { data_i[3:3] };
    end 
    if(N5613) begin
      { mem[2362:2362] } <= { data_i[2:2] };
    end 
    if(N5612) begin
      { mem[2361:2361] } <= { data_i[1:1] };
    end 
    if(N5611) begin
      { mem[2360:2360] } <= { data_i[0:0] };
    end 
    if(N5610) begin
      { mem[2359:2359] } <= { data_i[39:39] };
    end 
    if(N5609) begin
      { mem[2358:2358] } <= { data_i[38:38] };
    end 
    if(N5608) begin
      { mem[2357:2357] } <= { data_i[37:37] };
    end 
    if(N5607) begin
      { mem[2356:2356] } <= { data_i[36:36] };
    end 
    if(N5606) begin
      { mem[2355:2355] } <= { data_i[35:35] };
    end 
    if(N5605) begin
      { mem[2354:2354] } <= { data_i[34:34] };
    end 
    if(N5604) begin
      { mem[2353:2353] } <= { data_i[33:33] };
    end 
    if(N5603) begin
      { mem[2352:2352] } <= { data_i[32:32] };
    end 
    if(N5602) begin
      { mem[2351:2351] } <= { data_i[31:31] };
    end 
    if(N5601) begin
      { mem[2350:2350] } <= { data_i[30:30] };
    end 
    if(N5600) begin
      { mem[2349:2349] } <= { data_i[29:29] };
    end 
    if(N5599) begin
      { mem[2348:2348] } <= { data_i[28:28] };
    end 
    if(N5598) begin
      { mem[2347:2347] } <= { data_i[27:27] };
    end 
    if(N5597) begin
      { mem[2346:2346] } <= { data_i[26:26] };
    end 
    if(N5596) begin
      { mem[2345:2345] } <= { data_i[25:25] };
    end 
    if(N5595) begin
      { mem[2344:2344] } <= { data_i[24:24] };
    end 
    if(N5594) begin
      { mem[2343:2343] } <= { data_i[23:23] };
    end 
    if(N5593) begin
      { mem[2342:2342] } <= { data_i[22:22] };
    end 
    if(N5592) begin
      { mem[2341:2341] } <= { data_i[21:21] };
    end 
    if(N5591) begin
      { mem[2340:2340] } <= { data_i[20:20] };
    end 
    if(N5590) begin
      { mem[2339:2339] } <= { data_i[19:19] };
    end 
    if(N5589) begin
      { mem[2338:2338] } <= { data_i[18:18] };
    end 
    if(N5588) begin
      { mem[2337:2337] } <= { data_i[17:17] };
    end 
    if(N5587) begin
      { mem[2336:2336] } <= { data_i[16:16] };
    end 
    if(N5586) begin
      { mem[2335:2335] } <= { data_i[15:15] };
    end 
    if(N5585) begin
      { mem[2334:2334] } <= { data_i[14:14] };
    end 
    if(N5584) begin
      { mem[2333:2333] } <= { data_i[13:13] };
    end 
    if(N5583) begin
      { mem[2332:2332] } <= { data_i[12:12] };
    end 
    if(N5582) begin
      { mem[2331:2331] } <= { data_i[11:11] };
    end 
    if(N5581) begin
      { mem[2330:2330] } <= { data_i[10:10] };
    end 
    if(N5580) begin
      { mem[2329:2329] } <= { data_i[9:9] };
    end 
    if(N5579) begin
      { mem[2328:2328] } <= { data_i[8:8] };
    end 
    if(N5578) begin
      { mem[2327:2327] } <= { data_i[7:7] };
    end 
    if(N5577) begin
      { mem[2326:2326] } <= { data_i[6:6] };
    end 
    if(N5576) begin
      { mem[2325:2325] } <= { data_i[5:5] };
    end 
    if(N5575) begin
      { mem[2324:2324] } <= { data_i[4:4] };
    end 
    if(N5574) begin
      { mem[2323:2323] } <= { data_i[3:3] };
    end 
    if(N5573) begin
      { mem[2322:2322] } <= { data_i[2:2] };
    end 
    if(N5572) begin
      { mem[2321:2321] } <= { data_i[1:1] };
    end 
    if(N5571) begin
      { mem[2320:2320] } <= { data_i[0:0] };
    end 
    if(N5570) begin
      { mem[2319:2319] } <= { data_i[39:39] };
    end 
    if(N5569) begin
      { mem[2318:2318] } <= { data_i[38:38] };
    end 
    if(N5568) begin
      { mem[2317:2317] } <= { data_i[37:37] };
    end 
    if(N5567) begin
      { mem[2316:2316] } <= { data_i[36:36] };
    end 
    if(N5566) begin
      { mem[2315:2315] } <= { data_i[35:35] };
    end 
    if(N5565) begin
      { mem[2314:2314] } <= { data_i[34:34] };
    end 
    if(N5564) begin
      { mem[2313:2313] } <= { data_i[33:33] };
    end 
    if(N5563) begin
      { mem[2312:2312] } <= { data_i[32:32] };
    end 
    if(N5562) begin
      { mem[2311:2311] } <= { data_i[31:31] };
    end 
    if(N5561) begin
      { mem[2310:2310] } <= { data_i[30:30] };
    end 
    if(N5560) begin
      { mem[2309:2309] } <= { data_i[29:29] };
    end 
    if(N5559) begin
      { mem[2308:2308] } <= { data_i[28:28] };
    end 
    if(N5558) begin
      { mem[2307:2307] } <= { data_i[27:27] };
    end 
    if(N5557) begin
      { mem[2306:2306] } <= { data_i[26:26] };
    end 
    if(N5556) begin
      { mem[2305:2305] } <= { data_i[25:25] };
    end 
    if(N5555) begin
      { mem[2304:2304] } <= { data_i[24:24] };
    end 
    if(N5554) begin
      { mem[2303:2303] } <= { data_i[23:23] };
    end 
    if(N5553) begin
      { mem[2302:2302] } <= { data_i[22:22] };
    end 
    if(N5552) begin
      { mem[2301:2301] } <= { data_i[21:21] };
    end 
    if(N5551) begin
      { mem[2300:2300] } <= { data_i[20:20] };
    end 
    if(N5550) begin
      { mem[2299:2299] } <= { data_i[19:19] };
    end 
    if(N5549) begin
      { mem[2298:2298] } <= { data_i[18:18] };
    end 
    if(N5548) begin
      { mem[2297:2297] } <= { data_i[17:17] };
    end 
    if(N5547) begin
      { mem[2296:2296] } <= { data_i[16:16] };
    end 
    if(N5546) begin
      { mem[2295:2295] } <= { data_i[15:15] };
    end 
    if(N5545) begin
      { mem[2294:2294] } <= { data_i[14:14] };
    end 
    if(N5544) begin
      { mem[2293:2293] } <= { data_i[13:13] };
    end 
    if(N5543) begin
      { mem[2292:2292] } <= { data_i[12:12] };
    end 
    if(N5542) begin
      { mem[2291:2291] } <= { data_i[11:11] };
    end 
    if(N5541) begin
      { mem[2290:2290] } <= { data_i[10:10] };
    end 
    if(N5540) begin
      { mem[2289:2289] } <= { data_i[9:9] };
    end 
    if(N5539) begin
      { mem[2288:2288] } <= { data_i[8:8] };
    end 
    if(N5538) begin
      { mem[2287:2287] } <= { data_i[7:7] };
    end 
    if(N5537) begin
      { mem[2286:2286] } <= { data_i[6:6] };
    end 
    if(N5536) begin
      { mem[2285:2285] } <= { data_i[5:5] };
    end 
    if(N5535) begin
      { mem[2284:2284] } <= { data_i[4:4] };
    end 
    if(N5534) begin
      { mem[2283:2283] } <= { data_i[3:3] };
    end 
    if(N5533) begin
      { mem[2282:2282] } <= { data_i[2:2] };
    end 
    if(N5532) begin
      { mem[2281:2281] } <= { data_i[1:1] };
    end 
    if(N5531) begin
      { mem[2280:2280] } <= { data_i[0:0] };
    end 
    if(N5530) begin
      { mem[2279:2279] } <= { data_i[39:39] };
    end 
    if(N5529) begin
      { mem[2278:2278] } <= { data_i[38:38] };
    end 
    if(N5528) begin
      { mem[2277:2277] } <= { data_i[37:37] };
    end 
    if(N5527) begin
      { mem[2276:2276] } <= { data_i[36:36] };
    end 
    if(N5526) begin
      { mem[2275:2275] } <= { data_i[35:35] };
    end 
    if(N5525) begin
      { mem[2274:2274] } <= { data_i[34:34] };
    end 
    if(N5524) begin
      { mem[2273:2273] } <= { data_i[33:33] };
    end 
    if(N5523) begin
      { mem[2272:2272] } <= { data_i[32:32] };
    end 
    if(N5522) begin
      { mem[2271:2271] } <= { data_i[31:31] };
    end 
    if(N5521) begin
      { mem[2270:2270] } <= { data_i[30:30] };
    end 
    if(N5520) begin
      { mem[2269:2269] } <= { data_i[29:29] };
    end 
    if(N5519) begin
      { mem[2268:2268] } <= { data_i[28:28] };
    end 
    if(N5518) begin
      { mem[2267:2267] } <= { data_i[27:27] };
    end 
    if(N5517) begin
      { mem[2266:2266] } <= { data_i[26:26] };
    end 
    if(N5516) begin
      { mem[2265:2265] } <= { data_i[25:25] };
    end 
    if(N5515) begin
      { mem[2264:2264] } <= { data_i[24:24] };
    end 
    if(N5514) begin
      { mem[2263:2263] } <= { data_i[23:23] };
    end 
    if(N5513) begin
      { mem[2262:2262] } <= { data_i[22:22] };
    end 
    if(N5512) begin
      { mem[2261:2261] } <= { data_i[21:21] };
    end 
    if(N5511) begin
      { mem[2260:2260] } <= { data_i[20:20] };
    end 
    if(N5510) begin
      { mem[2259:2259] } <= { data_i[19:19] };
    end 
    if(N5509) begin
      { mem[2258:2258] } <= { data_i[18:18] };
    end 
    if(N5508) begin
      { mem[2257:2257] } <= { data_i[17:17] };
    end 
    if(N5507) begin
      { mem[2256:2256] } <= { data_i[16:16] };
    end 
    if(N5506) begin
      { mem[2255:2255] } <= { data_i[15:15] };
    end 
    if(N5505) begin
      { mem[2254:2254] } <= { data_i[14:14] };
    end 
    if(N5504) begin
      { mem[2253:2253] } <= { data_i[13:13] };
    end 
    if(N5503) begin
      { mem[2252:2252] } <= { data_i[12:12] };
    end 
    if(N5502) begin
      { mem[2251:2251] } <= { data_i[11:11] };
    end 
    if(N5501) begin
      { mem[2250:2250] } <= { data_i[10:10] };
    end 
    if(N5500) begin
      { mem[2249:2249] } <= { data_i[9:9] };
    end 
    if(N5499) begin
      { mem[2248:2248] } <= { data_i[8:8] };
    end 
    if(N5498) begin
      { mem[2247:2247] } <= { data_i[7:7] };
    end 
    if(N5497) begin
      { mem[2246:2246] } <= { data_i[6:6] };
    end 
    if(N5496) begin
      { mem[2245:2245] } <= { data_i[5:5] };
    end 
    if(N5495) begin
      { mem[2244:2244] } <= { data_i[4:4] };
    end 
    if(N5494) begin
      { mem[2243:2243] } <= { data_i[3:3] };
    end 
    if(N5493) begin
      { mem[2242:2242] } <= { data_i[2:2] };
    end 
    if(N5492) begin
      { mem[2241:2241] } <= { data_i[1:1] };
    end 
    if(N5491) begin
      { mem[2240:2240] } <= { data_i[0:0] };
    end 
    if(N5490) begin
      { mem[2239:2239] } <= { data_i[39:39] };
    end 
    if(N5489) begin
      { mem[2238:2238] } <= { data_i[38:38] };
    end 
    if(N5488) begin
      { mem[2237:2237] } <= { data_i[37:37] };
    end 
    if(N5487) begin
      { mem[2236:2236] } <= { data_i[36:36] };
    end 
    if(N5486) begin
      { mem[2235:2235] } <= { data_i[35:35] };
    end 
    if(N5485) begin
      { mem[2234:2234] } <= { data_i[34:34] };
    end 
    if(N5484) begin
      { mem[2233:2233] } <= { data_i[33:33] };
    end 
    if(N5483) begin
      { mem[2232:2232] } <= { data_i[32:32] };
    end 
    if(N5482) begin
      { mem[2231:2231] } <= { data_i[31:31] };
    end 
    if(N5481) begin
      { mem[2230:2230] } <= { data_i[30:30] };
    end 
    if(N5480) begin
      { mem[2229:2229] } <= { data_i[29:29] };
    end 
    if(N5479) begin
      { mem[2228:2228] } <= { data_i[28:28] };
    end 
    if(N5478) begin
      { mem[2227:2227] } <= { data_i[27:27] };
    end 
    if(N5477) begin
      { mem[2226:2226] } <= { data_i[26:26] };
    end 
    if(N5476) begin
      { mem[2225:2225] } <= { data_i[25:25] };
    end 
    if(N5475) begin
      { mem[2224:2224] } <= { data_i[24:24] };
    end 
    if(N5474) begin
      { mem[2223:2223] } <= { data_i[23:23] };
    end 
    if(N5473) begin
      { mem[2222:2222] } <= { data_i[22:22] };
    end 
    if(N5472) begin
      { mem[2221:2221] } <= { data_i[21:21] };
    end 
    if(N5471) begin
      { mem[2220:2220] } <= { data_i[20:20] };
    end 
    if(N5470) begin
      { mem[2219:2219] } <= { data_i[19:19] };
    end 
    if(N5469) begin
      { mem[2218:2218] } <= { data_i[18:18] };
    end 
    if(N5468) begin
      { mem[2217:2217] } <= { data_i[17:17] };
    end 
    if(N5467) begin
      { mem[2216:2216] } <= { data_i[16:16] };
    end 
    if(N5466) begin
      { mem[2215:2215] } <= { data_i[15:15] };
    end 
    if(N5465) begin
      { mem[2214:2214] } <= { data_i[14:14] };
    end 
    if(N5464) begin
      { mem[2213:2213] } <= { data_i[13:13] };
    end 
    if(N5463) begin
      { mem[2212:2212] } <= { data_i[12:12] };
    end 
    if(N5462) begin
      { mem[2211:2211] } <= { data_i[11:11] };
    end 
    if(N5461) begin
      { mem[2210:2210] } <= { data_i[10:10] };
    end 
    if(N5460) begin
      { mem[2209:2209] } <= { data_i[9:9] };
    end 
    if(N5459) begin
      { mem[2208:2208] } <= { data_i[8:8] };
    end 
    if(N5458) begin
      { mem[2207:2207] } <= { data_i[7:7] };
    end 
    if(N5457) begin
      { mem[2206:2206] } <= { data_i[6:6] };
    end 
    if(N5456) begin
      { mem[2205:2205] } <= { data_i[5:5] };
    end 
    if(N5455) begin
      { mem[2204:2204] } <= { data_i[4:4] };
    end 
    if(N5454) begin
      { mem[2203:2203] } <= { data_i[3:3] };
    end 
    if(N5453) begin
      { mem[2202:2202] } <= { data_i[2:2] };
    end 
    if(N5452) begin
      { mem[2201:2201] } <= { data_i[1:1] };
    end 
    if(N5451) begin
      { mem[2200:2200] } <= { data_i[0:0] };
    end 
    if(N5450) begin
      { mem[2199:2199] } <= { data_i[39:39] };
    end 
    if(N5449) begin
      { mem[2198:2198] } <= { data_i[38:38] };
    end 
    if(N5448) begin
      { mem[2197:2197] } <= { data_i[37:37] };
    end 
    if(N5447) begin
      { mem[2196:2196] } <= { data_i[36:36] };
    end 
    if(N5446) begin
      { mem[2195:2195] } <= { data_i[35:35] };
    end 
    if(N5445) begin
      { mem[2194:2194] } <= { data_i[34:34] };
    end 
    if(N5444) begin
      { mem[2193:2193] } <= { data_i[33:33] };
    end 
    if(N5443) begin
      { mem[2192:2192] } <= { data_i[32:32] };
    end 
    if(N5442) begin
      { mem[2191:2191] } <= { data_i[31:31] };
    end 
    if(N5441) begin
      { mem[2190:2190] } <= { data_i[30:30] };
    end 
    if(N5440) begin
      { mem[2189:2189] } <= { data_i[29:29] };
    end 
    if(N5439) begin
      { mem[2188:2188] } <= { data_i[28:28] };
    end 
    if(N5438) begin
      { mem[2187:2187] } <= { data_i[27:27] };
    end 
    if(N5437) begin
      { mem[2186:2186] } <= { data_i[26:26] };
    end 
    if(N5436) begin
      { mem[2185:2185] } <= { data_i[25:25] };
    end 
    if(N5435) begin
      { mem[2184:2184] } <= { data_i[24:24] };
    end 
    if(N5434) begin
      { mem[2183:2183] } <= { data_i[23:23] };
    end 
    if(N5433) begin
      { mem[2182:2182] } <= { data_i[22:22] };
    end 
    if(N5432) begin
      { mem[2181:2181] } <= { data_i[21:21] };
    end 
    if(N5431) begin
      { mem[2180:2180] } <= { data_i[20:20] };
    end 
    if(N5430) begin
      { mem[2179:2179] } <= { data_i[19:19] };
    end 
    if(N5429) begin
      { mem[2178:2178] } <= { data_i[18:18] };
    end 
    if(N5428) begin
      { mem[2177:2177] } <= { data_i[17:17] };
    end 
    if(N5427) begin
      { mem[2176:2176] } <= { data_i[16:16] };
    end 
    if(N5426) begin
      { mem[2175:2175] } <= { data_i[15:15] };
    end 
    if(N5425) begin
      { mem[2174:2174] } <= { data_i[14:14] };
    end 
    if(N5424) begin
      { mem[2173:2173] } <= { data_i[13:13] };
    end 
    if(N5423) begin
      { mem[2172:2172] } <= { data_i[12:12] };
    end 
    if(N5422) begin
      { mem[2171:2171] } <= { data_i[11:11] };
    end 
    if(N5421) begin
      { mem[2170:2170] } <= { data_i[10:10] };
    end 
    if(N5420) begin
      { mem[2169:2169] } <= { data_i[9:9] };
    end 
    if(N5419) begin
      { mem[2168:2168] } <= { data_i[8:8] };
    end 
    if(N5418) begin
      { mem[2167:2167] } <= { data_i[7:7] };
    end 
    if(N5417) begin
      { mem[2166:2166] } <= { data_i[6:6] };
    end 
    if(N5416) begin
      { mem[2165:2165] } <= { data_i[5:5] };
    end 
    if(N5415) begin
      { mem[2164:2164] } <= { data_i[4:4] };
    end 
    if(N5414) begin
      { mem[2163:2163] } <= { data_i[3:3] };
    end 
    if(N5413) begin
      { mem[2162:2162] } <= { data_i[2:2] };
    end 
    if(N5412) begin
      { mem[2161:2161] } <= { data_i[1:1] };
    end 
    if(N5411) begin
      { mem[2160:2160] } <= { data_i[0:0] };
    end 
    if(N5410) begin
      { mem[2159:2159] } <= { data_i[39:39] };
    end 
    if(N5409) begin
      { mem[2158:2158] } <= { data_i[38:38] };
    end 
    if(N5408) begin
      { mem[2157:2157] } <= { data_i[37:37] };
    end 
    if(N5407) begin
      { mem[2156:2156] } <= { data_i[36:36] };
    end 
    if(N5406) begin
      { mem[2155:2155] } <= { data_i[35:35] };
    end 
    if(N5405) begin
      { mem[2154:2154] } <= { data_i[34:34] };
    end 
    if(N5404) begin
      { mem[2153:2153] } <= { data_i[33:33] };
    end 
    if(N5403) begin
      { mem[2152:2152] } <= { data_i[32:32] };
    end 
    if(N5402) begin
      { mem[2151:2151] } <= { data_i[31:31] };
    end 
    if(N5401) begin
      { mem[2150:2150] } <= { data_i[30:30] };
    end 
    if(N5400) begin
      { mem[2149:2149] } <= { data_i[29:29] };
    end 
    if(N5399) begin
      { mem[2148:2148] } <= { data_i[28:28] };
    end 
    if(N5398) begin
      { mem[2147:2147] } <= { data_i[27:27] };
    end 
    if(N5397) begin
      { mem[2146:2146] } <= { data_i[26:26] };
    end 
    if(N5396) begin
      { mem[2145:2145] } <= { data_i[25:25] };
    end 
    if(N5395) begin
      { mem[2144:2144] } <= { data_i[24:24] };
    end 
    if(N5394) begin
      { mem[2143:2143] } <= { data_i[23:23] };
    end 
    if(N5393) begin
      { mem[2142:2142] } <= { data_i[22:22] };
    end 
    if(N5392) begin
      { mem[2141:2141] } <= { data_i[21:21] };
    end 
    if(N5391) begin
      { mem[2140:2140] } <= { data_i[20:20] };
    end 
    if(N5390) begin
      { mem[2139:2139] } <= { data_i[19:19] };
    end 
    if(N5389) begin
      { mem[2138:2138] } <= { data_i[18:18] };
    end 
    if(N5388) begin
      { mem[2137:2137] } <= { data_i[17:17] };
    end 
    if(N5387) begin
      { mem[2136:2136] } <= { data_i[16:16] };
    end 
    if(N5386) begin
      { mem[2135:2135] } <= { data_i[15:15] };
    end 
    if(N5385) begin
      { mem[2134:2134] } <= { data_i[14:14] };
    end 
    if(N5384) begin
      { mem[2133:2133] } <= { data_i[13:13] };
    end 
    if(N5383) begin
      { mem[2132:2132] } <= { data_i[12:12] };
    end 
    if(N5382) begin
      { mem[2131:2131] } <= { data_i[11:11] };
    end 
    if(N5381) begin
      { mem[2130:2130] } <= { data_i[10:10] };
    end 
    if(N5380) begin
      { mem[2129:2129] } <= { data_i[9:9] };
    end 
    if(N5379) begin
      { mem[2128:2128] } <= { data_i[8:8] };
    end 
    if(N5378) begin
      { mem[2127:2127] } <= { data_i[7:7] };
    end 
    if(N5377) begin
      { mem[2126:2126] } <= { data_i[6:6] };
    end 
    if(N5376) begin
      { mem[2125:2125] } <= { data_i[5:5] };
    end 
    if(N5375) begin
      { mem[2124:2124] } <= { data_i[4:4] };
    end 
    if(N5374) begin
      { mem[2123:2123] } <= { data_i[3:3] };
    end 
    if(N5373) begin
      { mem[2122:2122] } <= { data_i[2:2] };
    end 
    if(N5372) begin
      { mem[2121:2121] } <= { data_i[1:1] };
    end 
    if(N5371) begin
      { mem[2120:2120] } <= { data_i[0:0] };
    end 
    if(N5370) begin
      { mem[2119:2119] } <= { data_i[39:39] };
    end 
    if(N5369) begin
      { mem[2118:2118] } <= { data_i[38:38] };
    end 
    if(N5368) begin
      { mem[2117:2117] } <= { data_i[37:37] };
    end 
    if(N5367) begin
      { mem[2116:2116] } <= { data_i[36:36] };
    end 
    if(N5366) begin
      { mem[2115:2115] } <= { data_i[35:35] };
    end 
    if(N5365) begin
      { mem[2114:2114] } <= { data_i[34:34] };
    end 
    if(N5364) begin
      { mem[2113:2113] } <= { data_i[33:33] };
    end 
    if(N5363) begin
      { mem[2112:2112] } <= { data_i[32:32] };
    end 
    if(N5362) begin
      { mem[2111:2111] } <= { data_i[31:31] };
    end 
    if(N5361) begin
      { mem[2110:2110] } <= { data_i[30:30] };
    end 
    if(N5360) begin
      { mem[2109:2109] } <= { data_i[29:29] };
    end 
    if(N5359) begin
      { mem[2108:2108] } <= { data_i[28:28] };
    end 
    if(N5358) begin
      { mem[2107:2107] } <= { data_i[27:27] };
    end 
    if(N5357) begin
      { mem[2106:2106] } <= { data_i[26:26] };
    end 
    if(N5356) begin
      { mem[2105:2105] } <= { data_i[25:25] };
    end 
    if(N5355) begin
      { mem[2104:2104] } <= { data_i[24:24] };
    end 
    if(N5354) begin
      { mem[2103:2103] } <= { data_i[23:23] };
    end 
    if(N5353) begin
      { mem[2102:2102] } <= { data_i[22:22] };
    end 
    if(N5352) begin
      { mem[2101:2101] } <= { data_i[21:21] };
    end 
    if(N5351) begin
      { mem[2100:2100] } <= { data_i[20:20] };
    end 
    if(N5350) begin
      { mem[2099:2099] } <= { data_i[19:19] };
    end 
    if(N5349) begin
      { mem[2098:2098] } <= { data_i[18:18] };
    end 
    if(N5348) begin
      { mem[2097:2097] } <= { data_i[17:17] };
    end 
    if(N5347) begin
      { mem[2096:2096] } <= { data_i[16:16] };
    end 
    if(N5346) begin
      { mem[2095:2095] } <= { data_i[15:15] };
    end 
    if(N5345) begin
      { mem[2094:2094] } <= { data_i[14:14] };
    end 
    if(N5344) begin
      { mem[2093:2093] } <= { data_i[13:13] };
    end 
    if(N5343) begin
      { mem[2092:2092] } <= { data_i[12:12] };
    end 
    if(N5342) begin
      { mem[2091:2091] } <= { data_i[11:11] };
    end 
    if(N5341) begin
      { mem[2090:2090] } <= { data_i[10:10] };
    end 
    if(N5340) begin
      { mem[2089:2089] } <= { data_i[9:9] };
    end 
    if(N5339) begin
      { mem[2088:2088] } <= { data_i[8:8] };
    end 
    if(N5338) begin
      { mem[2087:2087] } <= { data_i[7:7] };
    end 
    if(N5337) begin
      { mem[2086:2086] } <= { data_i[6:6] };
    end 
    if(N5336) begin
      { mem[2085:2085] } <= { data_i[5:5] };
    end 
    if(N5335) begin
      { mem[2084:2084] } <= { data_i[4:4] };
    end 
    if(N5334) begin
      { mem[2083:2083] } <= { data_i[3:3] };
    end 
    if(N5333) begin
      { mem[2082:2082] } <= { data_i[2:2] };
    end 
    if(N5332) begin
      { mem[2081:2081] } <= { data_i[1:1] };
    end 
    if(N5331) begin
      { mem[2080:2080] } <= { data_i[0:0] };
    end 
    if(N5330) begin
      { mem[2079:2079] } <= { data_i[39:39] };
    end 
    if(N5329) begin
      { mem[2078:2078] } <= { data_i[38:38] };
    end 
    if(N5328) begin
      { mem[2077:2077] } <= { data_i[37:37] };
    end 
    if(N5327) begin
      { mem[2076:2076] } <= { data_i[36:36] };
    end 
    if(N5326) begin
      { mem[2075:2075] } <= { data_i[35:35] };
    end 
    if(N5325) begin
      { mem[2074:2074] } <= { data_i[34:34] };
    end 
    if(N5324) begin
      { mem[2073:2073] } <= { data_i[33:33] };
    end 
    if(N5323) begin
      { mem[2072:2072] } <= { data_i[32:32] };
    end 
    if(N5322) begin
      { mem[2071:2071] } <= { data_i[31:31] };
    end 
    if(N5321) begin
      { mem[2070:2070] } <= { data_i[30:30] };
    end 
    if(N5320) begin
      { mem[2069:2069] } <= { data_i[29:29] };
    end 
    if(N5319) begin
      { mem[2068:2068] } <= { data_i[28:28] };
    end 
    if(N5318) begin
      { mem[2067:2067] } <= { data_i[27:27] };
    end 
    if(N5317) begin
      { mem[2066:2066] } <= { data_i[26:26] };
    end 
    if(N5316) begin
      { mem[2065:2065] } <= { data_i[25:25] };
    end 
    if(N5315) begin
      { mem[2064:2064] } <= { data_i[24:24] };
    end 
    if(N5314) begin
      { mem[2063:2063] } <= { data_i[23:23] };
    end 
    if(N5313) begin
      { mem[2062:2062] } <= { data_i[22:22] };
    end 
    if(N5312) begin
      { mem[2061:2061] } <= { data_i[21:21] };
    end 
    if(N5311) begin
      { mem[2060:2060] } <= { data_i[20:20] };
    end 
    if(N5310) begin
      { mem[2059:2059] } <= { data_i[19:19] };
    end 
    if(N5309) begin
      { mem[2058:2058] } <= { data_i[18:18] };
    end 
    if(N5308) begin
      { mem[2057:2057] } <= { data_i[17:17] };
    end 
    if(N5307) begin
      { mem[2056:2056] } <= { data_i[16:16] };
    end 
    if(N5306) begin
      { mem[2055:2055] } <= { data_i[15:15] };
    end 
    if(N5305) begin
      { mem[2054:2054] } <= { data_i[14:14] };
    end 
    if(N5304) begin
      { mem[2053:2053] } <= { data_i[13:13] };
    end 
    if(N5303) begin
      { mem[2052:2052] } <= { data_i[12:12] };
    end 
    if(N5302) begin
      { mem[2051:2051] } <= { data_i[11:11] };
    end 
    if(N5301) begin
      { mem[2050:2050] } <= { data_i[10:10] };
    end 
    if(N5300) begin
      { mem[2049:2049] } <= { data_i[9:9] };
    end 
    if(N5299) begin
      { mem[2048:2048] } <= { data_i[8:8] };
    end 
    if(N5298) begin
      { mem[2047:2047] } <= { data_i[7:7] };
    end 
    if(N5297) begin
      { mem[2046:2046] } <= { data_i[6:6] };
    end 
    if(N5296) begin
      { mem[2045:2045] } <= { data_i[5:5] };
    end 
    if(N5295) begin
      { mem[2044:2044] } <= { data_i[4:4] };
    end 
    if(N5294) begin
      { mem[2043:2043] } <= { data_i[3:3] };
    end 
    if(N5293) begin
      { mem[2042:2042] } <= { data_i[2:2] };
    end 
    if(N5292) begin
      { mem[2041:2041] } <= { data_i[1:1] };
    end 
    if(N5291) begin
      { mem[2040:2040] } <= { data_i[0:0] };
    end 
    if(N5290) begin
      { mem[2039:2039] } <= { data_i[39:39] };
    end 
    if(N5289) begin
      { mem[2038:2038] } <= { data_i[38:38] };
    end 
    if(N5288) begin
      { mem[2037:2037] } <= { data_i[37:37] };
    end 
    if(N5287) begin
      { mem[2036:2036] } <= { data_i[36:36] };
    end 
    if(N5286) begin
      { mem[2035:2035] } <= { data_i[35:35] };
    end 
    if(N5285) begin
      { mem[2034:2034] } <= { data_i[34:34] };
    end 
    if(N5284) begin
      { mem[2033:2033] } <= { data_i[33:33] };
    end 
    if(N5283) begin
      { mem[2032:2032] } <= { data_i[32:32] };
    end 
    if(N5282) begin
      { mem[2031:2031] } <= { data_i[31:31] };
    end 
    if(N5281) begin
      { mem[2030:2030] } <= { data_i[30:30] };
    end 
    if(N5280) begin
      { mem[2029:2029] } <= { data_i[29:29] };
    end 
    if(N5279) begin
      { mem[2028:2028] } <= { data_i[28:28] };
    end 
    if(N5278) begin
      { mem[2027:2027] } <= { data_i[27:27] };
    end 
    if(N5277) begin
      { mem[2026:2026] } <= { data_i[26:26] };
    end 
    if(N5276) begin
      { mem[2025:2025] } <= { data_i[25:25] };
    end 
    if(N5275) begin
      { mem[2024:2024] } <= { data_i[24:24] };
    end 
    if(N5274) begin
      { mem[2023:2023] } <= { data_i[23:23] };
    end 
    if(N5273) begin
      { mem[2022:2022] } <= { data_i[22:22] };
    end 
    if(N5272) begin
      { mem[2021:2021] } <= { data_i[21:21] };
    end 
    if(N5271) begin
      { mem[2020:2020] } <= { data_i[20:20] };
    end 
    if(N5270) begin
      { mem[2019:2019] } <= { data_i[19:19] };
    end 
    if(N5269) begin
      { mem[2018:2018] } <= { data_i[18:18] };
    end 
    if(N5268) begin
      { mem[2017:2017] } <= { data_i[17:17] };
    end 
    if(N5267) begin
      { mem[2016:2016] } <= { data_i[16:16] };
    end 
    if(N5266) begin
      { mem[2015:2015] } <= { data_i[15:15] };
    end 
    if(N5265) begin
      { mem[2014:2014] } <= { data_i[14:14] };
    end 
    if(N5264) begin
      { mem[2013:2013] } <= { data_i[13:13] };
    end 
    if(N5263) begin
      { mem[2012:2012] } <= { data_i[12:12] };
    end 
    if(N5262) begin
      { mem[2011:2011] } <= { data_i[11:11] };
    end 
    if(N5261) begin
      { mem[2010:2010] } <= { data_i[10:10] };
    end 
    if(N5260) begin
      { mem[2009:2009] } <= { data_i[9:9] };
    end 
    if(N5259) begin
      { mem[2008:2008] } <= { data_i[8:8] };
    end 
    if(N5258) begin
      { mem[2007:2007] } <= { data_i[7:7] };
    end 
    if(N5257) begin
      { mem[2006:2006] } <= { data_i[6:6] };
    end 
    if(N5256) begin
      { mem[2005:2005] } <= { data_i[5:5] };
    end 
    if(N5255) begin
      { mem[2004:2004] } <= { data_i[4:4] };
    end 
    if(N5254) begin
      { mem[2003:2003] } <= { data_i[3:3] };
    end 
    if(N5253) begin
      { mem[2002:2002] } <= { data_i[2:2] };
    end 
    if(N5252) begin
      { mem[2001:2001] } <= { data_i[1:1] };
    end 
    if(N5251) begin
      { mem[2000:2000] } <= { data_i[0:0] };
    end 
    if(N5250) begin
      { mem[1999:1999] } <= { data_i[39:39] };
    end 
    if(N5249) begin
      { mem[1998:1998] } <= { data_i[38:38] };
    end 
    if(N5248) begin
      { mem[1997:1997] } <= { data_i[37:37] };
    end 
    if(N5247) begin
      { mem[1996:1996] } <= { data_i[36:36] };
    end 
    if(N5246) begin
      { mem[1995:1995] } <= { data_i[35:35] };
    end 
    if(N5245) begin
      { mem[1994:1994] } <= { data_i[34:34] };
    end 
    if(N5244) begin
      { mem[1993:1993] } <= { data_i[33:33] };
    end 
    if(N5243) begin
      { mem[1992:1992] } <= { data_i[32:32] };
    end 
    if(N5242) begin
      { mem[1991:1991] } <= { data_i[31:31] };
    end 
    if(N5241) begin
      { mem[1990:1990] } <= { data_i[30:30] };
    end 
    if(N5240) begin
      { mem[1989:1989] } <= { data_i[29:29] };
    end 
    if(N5239) begin
      { mem[1988:1988] } <= { data_i[28:28] };
    end 
    if(N5238) begin
      { mem[1987:1987] } <= { data_i[27:27] };
    end 
    if(N5237) begin
      { mem[1986:1986] } <= { data_i[26:26] };
    end 
    if(N5236) begin
      { mem[1985:1985] } <= { data_i[25:25] };
    end 
    if(N5235) begin
      { mem[1984:1984] } <= { data_i[24:24] };
    end 
    if(N5234) begin
      { mem[1983:1983] } <= { data_i[23:23] };
    end 
    if(N5233) begin
      { mem[1982:1982] } <= { data_i[22:22] };
    end 
    if(N5232) begin
      { mem[1981:1981] } <= { data_i[21:21] };
    end 
    if(N5231) begin
      { mem[1980:1980] } <= { data_i[20:20] };
    end 
    if(N5230) begin
      { mem[1979:1979] } <= { data_i[19:19] };
    end 
    if(N5229) begin
      { mem[1978:1978] } <= { data_i[18:18] };
    end 
    if(N5228) begin
      { mem[1977:1977] } <= { data_i[17:17] };
    end 
    if(N5227) begin
      { mem[1976:1976] } <= { data_i[16:16] };
    end 
    if(N5226) begin
      { mem[1975:1975] } <= { data_i[15:15] };
    end 
    if(N5225) begin
      { mem[1974:1974] } <= { data_i[14:14] };
    end 
    if(N5224) begin
      { mem[1973:1973] } <= { data_i[13:13] };
    end 
    if(N5223) begin
      { mem[1972:1972] } <= { data_i[12:12] };
    end 
    if(N5222) begin
      { mem[1971:1971] } <= { data_i[11:11] };
    end 
    if(N5221) begin
      { mem[1970:1970] } <= { data_i[10:10] };
    end 
    if(N5220) begin
      { mem[1969:1969] } <= { data_i[9:9] };
    end 
    if(N5219) begin
      { mem[1968:1968] } <= { data_i[8:8] };
    end 
    if(N5218) begin
      { mem[1967:1967] } <= { data_i[7:7] };
    end 
    if(N5217) begin
      { mem[1966:1966] } <= { data_i[6:6] };
    end 
    if(N5216) begin
      { mem[1965:1965] } <= { data_i[5:5] };
    end 
    if(N5215) begin
      { mem[1964:1964] } <= { data_i[4:4] };
    end 
    if(N5214) begin
      { mem[1963:1963] } <= { data_i[3:3] };
    end 
    if(N5213) begin
      { mem[1962:1962] } <= { data_i[2:2] };
    end 
    if(N5212) begin
      { mem[1961:1961] } <= { data_i[1:1] };
    end 
    if(N5211) begin
      { mem[1960:1960] } <= { data_i[0:0] };
    end 
    if(N5210) begin
      { mem[1959:1959] } <= { data_i[39:39] };
    end 
    if(N5209) begin
      { mem[1958:1958] } <= { data_i[38:38] };
    end 
    if(N5208) begin
      { mem[1957:1957] } <= { data_i[37:37] };
    end 
    if(N5207) begin
      { mem[1956:1956] } <= { data_i[36:36] };
    end 
    if(N5206) begin
      { mem[1955:1955] } <= { data_i[35:35] };
    end 
    if(N5205) begin
      { mem[1954:1954] } <= { data_i[34:34] };
    end 
    if(N5204) begin
      { mem[1953:1953] } <= { data_i[33:33] };
    end 
    if(N5203) begin
      { mem[1952:1952] } <= { data_i[32:32] };
    end 
    if(N5202) begin
      { mem[1951:1951] } <= { data_i[31:31] };
    end 
    if(N5201) begin
      { mem[1950:1950] } <= { data_i[30:30] };
    end 
    if(N5200) begin
      { mem[1949:1949] } <= { data_i[29:29] };
    end 
    if(N5199) begin
      { mem[1948:1948] } <= { data_i[28:28] };
    end 
    if(N5198) begin
      { mem[1947:1947] } <= { data_i[27:27] };
    end 
    if(N5197) begin
      { mem[1946:1946] } <= { data_i[26:26] };
    end 
    if(N5196) begin
      { mem[1945:1945] } <= { data_i[25:25] };
    end 
    if(N5195) begin
      { mem[1944:1944] } <= { data_i[24:24] };
    end 
    if(N5194) begin
      { mem[1943:1943] } <= { data_i[23:23] };
    end 
    if(N5193) begin
      { mem[1942:1942] } <= { data_i[22:22] };
    end 
    if(N5192) begin
      { mem[1941:1941] } <= { data_i[21:21] };
    end 
    if(N5191) begin
      { mem[1940:1940] } <= { data_i[20:20] };
    end 
    if(N5190) begin
      { mem[1939:1939] } <= { data_i[19:19] };
    end 
    if(N5189) begin
      { mem[1938:1938] } <= { data_i[18:18] };
    end 
    if(N5188) begin
      { mem[1937:1937] } <= { data_i[17:17] };
    end 
    if(N5187) begin
      { mem[1936:1936] } <= { data_i[16:16] };
    end 
    if(N5186) begin
      { mem[1935:1935] } <= { data_i[15:15] };
    end 
    if(N5185) begin
      { mem[1934:1934] } <= { data_i[14:14] };
    end 
    if(N5184) begin
      { mem[1933:1933] } <= { data_i[13:13] };
    end 
    if(N5183) begin
      { mem[1932:1932] } <= { data_i[12:12] };
    end 
    if(N5182) begin
      { mem[1931:1931] } <= { data_i[11:11] };
    end 
    if(N5181) begin
      { mem[1930:1930] } <= { data_i[10:10] };
    end 
    if(N5180) begin
      { mem[1929:1929] } <= { data_i[9:9] };
    end 
    if(N5179) begin
      { mem[1928:1928] } <= { data_i[8:8] };
    end 
    if(N5178) begin
      { mem[1927:1927] } <= { data_i[7:7] };
    end 
    if(N5177) begin
      { mem[1926:1926] } <= { data_i[6:6] };
    end 
    if(N5176) begin
      { mem[1925:1925] } <= { data_i[5:5] };
    end 
    if(N5175) begin
      { mem[1924:1924] } <= { data_i[4:4] };
    end 
    if(N5174) begin
      { mem[1923:1923] } <= { data_i[3:3] };
    end 
    if(N5173) begin
      { mem[1922:1922] } <= { data_i[2:2] };
    end 
    if(N5172) begin
      { mem[1921:1921] } <= { data_i[1:1] };
    end 
    if(N5171) begin
      { mem[1920:1920] } <= { data_i[0:0] };
    end 
    if(N5170) begin
      { mem[1919:1919] } <= { data_i[39:39] };
    end 
    if(N5169) begin
      { mem[1918:1918] } <= { data_i[38:38] };
    end 
    if(N5168) begin
      { mem[1917:1917] } <= { data_i[37:37] };
    end 
    if(N5167) begin
      { mem[1916:1916] } <= { data_i[36:36] };
    end 
    if(N5166) begin
      { mem[1915:1915] } <= { data_i[35:35] };
    end 
    if(N5165) begin
      { mem[1914:1914] } <= { data_i[34:34] };
    end 
    if(N5164) begin
      { mem[1913:1913] } <= { data_i[33:33] };
    end 
    if(N5163) begin
      { mem[1912:1912] } <= { data_i[32:32] };
    end 
    if(N5162) begin
      { mem[1911:1911] } <= { data_i[31:31] };
    end 
    if(N5161) begin
      { mem[1910:1910] } <= { data_i[30:30] };
    end 
    if(N5160) begin
      { mem[1909:1909] } <= { data_i[29:29] };
    end 
    if(N5159) begin
      { mem[1908:1908] } <= { data_i[28:28] };
    end 
    if(N5158) begin
      { mem[1907:1907] } <= { data_i[27:27] };
    end 
    if(N5157) begin
      { mem[1906:1906] } <= { data_i[26:26] };
    end 
    if(N5156) begin
      { mem[1905:1905] } <= { data_i[25:25] };
    end 
    if(N5155) begin
      { mem[1904:1904] } <= { data_i[24:24] };
    end 
    if(N5154) begin
      { mem[1903:1903] } <= { data_i[23:23] };
    end 
    if(N5153) begin
      { mem[1902:1902] } <= { data_i[22:22] };
    end 
    if(N5152) begin
      { mem[1901:1901] } <= { data_i[21:21] };
    end 
    if(N5151) begin
      { mem[1900:1900] } <= { data_i[20:20] };
    end 
    if(N5150) begin
      { mem[1899:1899] } <= { data_i[19:19] };
    end 
    if(N5149) begin
      { mem[1898:1898] } <= { data_i[18:18] };
    end 
    if(N5148) begin
      { mem[1897:1897] } <= { data_i[17:17] };
    end 
    if(N5147) begin
      { mem[1896:1896] } <= { data_i[16:16] };
    end 
    if(N5146) begin
      { mem[1895:1895] } <= { data_i[15:15] };
    end 
    if(N5145) begin
      { mem[1894:1894] } <= { data_i[14:14] };
    end 
    if(N5144) begin
      { mem[1893:1893] } <= { data_i[13:13] };
    end 
    if(N5143) begin
      { mem[1892:1892] } <= { data_i[12:12] };
    end 
    if(N5142) begin
      { mem[1891:1891] } <= { data_i[11:11] };
    end 
    if(N5141) begin
      { mem[1890:1890] } <= { data_i[10:10] };
    end 
    if(N5140) begin
      { mem[1889:1889] } <= { data_i[9:9] };
    end 
    if(N5139) begin
      { mem[1888:1888] } <= { data_i[8:8] };
    end 
    if(N5138) begin
      { mem[1887:1887] } <= { data_i[7:7] };
    end 
    if(N5137) begin
      { mem[1886:1886] } <= { data_i[6:6] };
    end 
    if(N5136) begin
      { mem[1885:1885] } <= { data_i[5:5] };
    end 
    if(N5135) begin
      { mem[1884:1884] } <= { data_i[4:4] };
    end 
    if(N5134) begin
      { mem[1883:1883] } <= { data_i[3:3] };
    end 
    if(N5133) begin
      { mem[1882:1882] } <= { data_i[2:2] };
    end 
    if(N5132) begin
      { mem[1881:1881] } <= { data_i[1:1] };
    end 
    if(N5131) begin
      { mem[1880:1880] } <= { data_i[0:0] };
    end 
    if(N5130) begin
      { mem[1879:1879] } <= { data_i[39:39] };
    end 
    if(N5129) begin
      { mem[1878:1878] } <= { data_i[38:38] };
    end 
    if(N5128) begin
      { mem[1877:1877] } <= { data_i[37:37] };
    end 
    if(N5127) begin
      { mem[1876:1876] } <= { data_i[36:36] };
    end 
    if(N5126) begin
      { mem[1875:1875] } <= { data_i[35:35] };
    end 
    if(N5125) begin
      { mem[1874:1874] } <= { data_i[34:34] };
    end 
    if(N5124) begin
      { mem[1873:1873] } <= { data_i[33:33] };
    end 
    if(N5123) begin
      { mem[1872:1872] } <= { data_i[32:32] };
    end 
    if(N5122) begin
      { mem[1871:1871] } <= { data_i[31:31] };
    end 
    if(N5121) begin
      { mem[1870:1870] } <= { data_i[30:30] };
    end 
    if(N5120) begin
      { mem[1869:1869] } <= { data_i[29:29] };
    end 
    if(N5119) begin
      { mem[1868:1868] } <= { data_i[28:28] };
    end 
    if(N5118) begin
      { mem[1867:1867] } <= { data_i[27:27] };
    end 
    if(N5117) begin
      { mem[1866:1866] } <= { data_i[26:26] };
    end 
    if(N5116) begin
      { mem[1865:1865] } <= { data_i[25:25] };
    end 
    if(N5115) begin
      { mem[1864:1864] } <= { data_i[24:24] };
    end 
    if(N5114) begin
      { mem[1863:1863] } <= { data_i[23:23] };
    end 
    if(N5113) begin
      { mem[1862:1862] } <= { data_i[22:22] };
    end 
    if(N5112) begin
      { mem[1861:1861] } <= { data_i[21:21] };
    end 
    if(N5111) begin
      { mem[1860:1860] } <= { data_i[20:20] };
    end 
    if(N5110) begin
      { mem[1859:1859] } <= { data_i[19:19] };
    end 
    if(N5109) begin
      { mem[1858:1858] } <= { data_i[18:18] };
    end 
    if(N5108) begin
      { mem[1857:1857] } <= { data_i[17:17] };
    end 
    if(N5107) begin
      { mem[1856:1856] } <= { data_i[16:16] };
    end 
    if(N5106) begin
      { mem[1855:1855] } <= { data_i[15:15] };
    end 
    if(N5105) begin
      { mem[1854:1854] } <= { data_i[14:14] };
    end 
    if(N5104) begin
      { mem[1853:1853] } <= { data_i[13:13] };
    end 
    if(N5103) begin
      { mem[1852:1852] } <= { data_i[12:12] };
    end 
    if(N5102) begin
      { mem[1851:1851] } <= { data_i[11:11] };
    end 
    if(N5101) begin
      { mem[1850:1850] } <= { data_i[10:10] };
    end 
    if(N5100) begin
      { mem[1849:1849] } <= { data_i[9:9] };
    end 
    if(N5099) begin
      { mem[1848:1848] } <= { data_i[8:8] };
    end 
    if(N5098) begin
      { mem[1847:1847] } <= { data_i[7:7] };
    end 
    if(N5097) begin
      { mem[1846:1846] } <= { data_i[6:6] };
    end 
    if(N5096) begin
      { mem[1845:1845] } <= { data_i[5:5] };
    end 
    if(N5095) begin
      { mem[1844:1844] } <= { data_i[4:4] };
    end 
    if(N5094) begin
      { mem[1843:1843] } <= { data_i[3:3] };
    end 
    if(N5093) begin
      { mem[1842:1842] } <= { data_i[2:2] };
    end 
    if(N5092) begin
      { mem[1841:1841] } <= { data_i[1:1] };
    end 
    if(N5091) begin
      { mem[1840:1840] } <= { data_i[0:0] };
    end 
    if(N5090) begin
      { mem[1839:1839] } <= { data_i[39:39] };
    end 
    if(N5089) begin
      { mem[1838:1838] } <= { data_i[38:38] };
    end 
    if(N5088) begin
      { mem[1837:1837] } <= { data_i[37:37] };
    end 
    if(N5087) begin
      { mem[1836:1836] } <= { data_i[36:36] };
    end 
    if(N5086) begin
      { mem[1835:1835] } <= { data_i[35:35] };
    end 
    if(N5085) begin
      { mem[1834:1834] } <= { data_i[34:34] };
    end 
    if(N5084) begin
      { mem[1833:1833] } <= { data_i[33:33] };
    end 
    if(N5083) begin
      { mem[1832:1832] } <= { data_i[32:32] };
    end 
    if(N5082) begin
      { mem[1831:1831] } <= { data_i[31:31] };
    end 
    if(N5081) begin
      { mem[1830:1830] } <= { data_i[30:30] };
    end 
    if(N5080) begin
      { mem[1829:1829] } <= { data_i[29:29] };
    end 
    if(N5079) begin
      { mem[1828:1828] } <= { data_i[28:28] };
    end 
    if(N5078) begin
      { mem[1827:1827] } <= { data_i[27:27] };
    end 
    if(N5077) begin
      { mem[1826:1826] } <= { data_i[26:26] };
    end 
    if(N5076) begin
      { mem[1825:1825] } <= { data_i[25:25] };
    end 
    if(N5075) begin
      { mem[1824:1824] } <= { data_i[24:24] };
    end 
    if(N5074) begin
      { mem[1823:1823] } <= { data_i[23:23] };
    end 
    if(N5073) begin
      { mem[1822:1822] } <= { data_i[22:22] };
    end 
    if(N5072) begin
      { mem[1821:1821] } <= { data_i[21:21] };
    end 
    if(N5071) begin
      { mem[1820:1820] } <= { data_i[20:20] };
    end 
    if(N5070) begin
      { mem[1819:1819] } <= { data_i[19:19] };
    end 
    if(N5069) begin
      { mem[1818:1818] } <= { data_i[18:18] };
    end 
    if(N5068) begin
      { mem[1817:1817] } <= { data_i[17:17] };
    end 
    if(N5067) begin
      { mem[1816:1816] } <= { data_i[16:16] };
    end 
    if(N5066) begin
      { mem[1815:1815] } <= { data_i[15:15] };
    end 
    if(N5065) begin
      { mem[1814:1814] } <= { data_i[14:14] };
    end 
    if(N5064) begin
      { mem[1813:1813] } <= { data_i[13:13] };
    end 
    if(N5063) begin
      { mem[1812:1812] } <= { data_i[12:12] };
    end 
    if(N5062) begin
      { mem[1811:1811] } <= { data_i[11:11] };
    end 
    if(N5061) begin
      { mem[1810:1810] } <= { data_i[10:10] };
    end 
    if(N5060) begin
      { mem[1809:1809] } <= { data_i[9:9] };
    end 
    if(N5059) begin
      { mem[1808:1808] } <= { data_i[8:8] };
    end 
    if(N5058) begin
      { mem[1807:1807] } <= { data_i[7:7] };
    end 
    if(N5057) begin
      { mem[1806:1806] } <= { data_i[6:6] };
    end 
    if(N5056) begin
      { mem[1805:1805] } <= { data_i[5:5] };
    end 
    if(N5055) begin
      { mem[1804:1804] } <= { data_i[4:4] };
    end 
    if(N5054) begin
      { mem[1803:1803] } <= { data_i[3:3] };
    end 
    if(N5053) begin
      { mem[1802:1802] } <= { data_i[2:2] };
    end 
    if(N5052) begin
      { mem[1801:1801] } <= { data_i[1:1] };
    end 
    if(N5051) begin
      { mem[1800:1800] } <= { data_i[0:0] };
    end 
    if(N5050) begin
      { mem[1799:1799] } <= { data_i[39:39] };
    end 
    if(N5049) begin
      { mem[1798:1798] } <= { data_i[38:38] };
    end 
    if(N5048) begin
      { mem[1797:1797] } <= { data_i[37:37] };
    end 
    if(N5047) begin
      { mem[1796:1796] } <= { data_i[36:36] };
    end 
    if(N5046) begin
      { mem[1795:1795] } <= { data_i[35:35] };
    end 
    if(N5045) begin
      { mem[1794:1794] } <= { data_i[34:34] };
    end 
    if(N5044) begin
      { mem[1793:1793] } <= { data_i[33:33] };
    end 
    if(N5043) begin
      { mem[1792:1792] } <= { data_i[32:32] };
    end 
    if(N5042) begin
      { mem[1791:1791] } <= { data_i[31:31] };
    end 
    if(N5041) begin
      { mem[1790:1790] } <= { data_i[30:30] };
    end 
    if(N5040) begin
      { mem[1789:1789] } <= { data_i[29:29] };
    end 
    if(N5039) begin
      { mem[1788:1788] } <= { data_i[28:28] };
    end 
    if(N5038) begin
      { mem[1787:1787] } <= { data_i[27:27] };
    end 
    if(N5037) begin
      { mem[1786:1786] } <= { data_i[26:26] };
    end 
    if(N5036) begin
      { mem[1785:1785] } <= { data_i[25:25] };
    end 
    if(N5035) begin
      { mem[1784:1784] } <= { data_i[24:24] };
    end 
    if(N5034) begin
      { mem[1783:1783] } <= { data_i[23:23] };
    end 
    if(N5033) begin
      { mem[1782:1782] } <= { data_i[22:22] };
    end 
    if(N5032) begin
      { mem[1781:1781] } <= { data_i[21:21] };
    end 
    if(N5031) begin
      { mem[1780:1780] } <= { data_i[20:20] };
    end 
    if(N5030) begin
      { mem[1779:1779] } <= { data_i[19:19] };
    end 
    if(N5029) begin
      { mem[1778:1778] } <= { data_i[18:18] };
    end 
    if(N5028) begin
      { mem[1777:1777] } <= { data_i[17:17] };
    end 
    if(N5027) begin
      { mem[1776:1776] } <= { data_i[16:16] };
    end 
    if(N5026) begin
      { mem[1775:1775] } <= { data_i[15:15] };
    end 
    if(N5025) begin
      { mem[1774:1774] } <= { data_i[14:14] };
    end 
    if(N5024) begin
      { mem[1773:1773] } <= { data_i[13:13] };
    end 
    if(N5023) begin
      { mem[1772:1772] } <= { data_i[12:12] };
    end 
    if(N5022) begin
      { mem[1771:1771] } <= { data_i[11:11] };
    end 
    if(N5021) begin
      { mem[1770:1770] } <= { data_i[10:10] };
    end 
    if(N5020) begin
      { mem[1769:1769] } <= { data_i[9:9] };
    end 
    if(N5019) begin
      { mem[1768:1768] } <= { data_i[8:8] };
    end 
    if(N5018) begin
      { mem[1767:1767] } <= { data_i[7:7] };
    end 
    if(N5017) begin
      { mem[1766:1766] } <= { data_i[6:6] };
    end 
    if(N5016) begin
      { mem[1765:1765] } <= { data_i[5:5] };
    end 
    if(N5015) begin
      { mem[1764:1764] } <= { data_i[4:4] };
    end 
    if(N5014) begin
      { mem[1763:1763] } <= { data_i[3:3] };
    end 
    if(N5013) begin
      { mem[1762:1762] } <= { data_i[2:2] };
    end 
    if(N5012) begin
      { mem[1761:1761] } <= { data_i[1:1] };
    end 
    if(N5011) begin
      { mem[1760:1760] } <= { data_i[0:0] };
    end 
    if(N5010) begin
      { mem[1759:1759] } <= { data_i[39:39] };
    end 
    if(N5009) begin
      { mem[1758:1758] } <= { data_i[38:38] };
    end 
    if(N5008) begin
      { mem[1757:1757] } <= { data_i[37:37] };
    end 
    if(N5007) begin
      { mem[1756:1756] } <= { data_i[36:36] };
    end 
    if(N5006) begin
      { mem[1755:1755] } <= { data_i[35:35] };
    end 
    if(N5005) begin
      { mem[1754:1754] } <= { data_i[34:34] };
    end 
    if(N5004) begin
      { mem[1753:1753] } <= { data_i[33:33] };
    end 
    if(N5003) begin
      { mem[1752:1752] } <= { data_i[32:32] };
    end 
    if(N5002) begin
      { mem[1751:1751] } <= { data_i[31:31] };
    end 
    if(N5001) begin
      { mem[1750:1750] } <= { data_i[30:30] };
    end 
    if(N5000) begin
      { mem[1749:1749] } <= { data_i[29:29] };
    end 
    if(N4999) begin
      { mem[1748:1748] } <= { data_i[28:28] };
    end 
    if(N4998) begin
      { mem[1747:1747] } <= { data_i[27:27] };
    end 
    if(N4997) begin
      { mem[1746:1746] } <= { data_i[26:26] };
    end 
    if(N4996) begin
      { mem[1745:1745] } <= { data_i[25:25] };
    end 
    if(N4995) begin
      { mem[1744:1744] } <= { data_i[24:24] };
    end 
    if(N4994) begin
      { mem[1743:1743] } <= { data_i[23:23] };
    end 
    if(N4993) begin
      { mem[1742:1742] } <= { data_i[22:22] };
    end 
    if(N4992) begin
      { mem[1741:1741] } <= { data_i[21:21] };
    end 
    if(N4991) begin
      { mem[1740:1740] } <= { data_i[20:20] };
    end 
    if(N4990) begin
      { mem[1739:1739] } <= { data_i[19:19] };
    end 
    if(N4989) begin
      { mem[1738:1738] } <= { data_i[18:18] };
    end 
    if(N4988) begin
      { mem[1737:1737] } <= { data_i[17:17] };
    end 
    if(N4987) begin
      { mem[1736:1736] } <= { data_i[16:16] };
    end 
    if(N4986) begin
      { mem[1735:1735] } <= { data_i[15:15] };
    end 
    if(N4985) begin
      { mem[1734:1734] } <= { data_i[14:14] };
    end 
    if(N4984) begin
      { mem[1733:1733] } <= { data_i[13:13] };
    end 
    if(N4983) begin
      { mem[1732:1732] } <= { data_i[12:12] };
    end 
    if(N4982) begin
      { mem[1731:1731] } <= { data_i[11:11] };
    end 
    if(N4981) begin
      { mem[1730:1730] } <= { data_i[10:10] };
    end 
    if(N4980) begin
      { mem[1729:1729] } <= { data_i[9:9] };
    end 
    if(N4979) begin
      { mem[1728:1728] } <= { data_i[8:8] };
    end 
    if(N4978) begin
      { mem[1727:1727] } <= { data_i[7:7] };
    end 
    if(N4977) begin
      { mem[1726:1726] } <= { data_i[6:6] };
    end 
    if(N4976) begin
      { mem[1725:1725] } <= { data_i[5:5] };
    end 
    if(N4975) begin
      { mem[1724:1724] } <= { data_i[4:4] };
    end 
    if(N4974) begin
      { mem[1723:1723] } <= { data_i[3:3] };
    end 
    if(N4973) begin
      { mem[1722:1722] } <= { data_i[2:2] };
    end 
    if(N4972) begin
      { mem[1721:1721] } <= { data_i[1:1] };
    end 
    if(N4971) begin
      { mem[1720:1720] } <= { data_i[0:0] };
    end 
    if(N4970) begin
      { mem[1719:1719] } <= { data_i[39:39] };
    end 
    if(N4969) begin
      { mem[1718:1718] } <= { data_i[38:38] };
    end 
    if(N4968) begin
      { mem[1717:1717] } <= { data_i[37:37] };
    end 
    if(N4967) begin
      { mem[1716:1716] } <= { data_i[36:36] };
    end 
    if(N4966) begin
      { mem[1715:1715] } <= { data_i[35:35] };
    end 
    if(N4965) begin
      { mem[1714:1714] } <= { data_i[34:34] };
    end 
    if(N4964) begin
      { mem[1713:1713] } <= { data_i[33:33] };
    end 
    if(N4963) begin
      { mem[1712:1712] } <= { data_i[32:32] };
    end 
    if(N4962) begin
      { mem[1711:1711] } <= { data_i[31:31] };
    end 
    if(N4961) begin
      { mem[1710:1710] } <= { data_i[30:30] };
    end 
    if(N4960) begin
      { mem[1709:1709] } <= { data_i[29:29] };
    end 
    if(N4959) begin
      { mem[1708:1708] } <= { data_i[28:28] };
    end 
    if(N4958) begin
      { mem[1707:1707] } <= { data_i[27:27] };
    end 
    if(N4957) begin
      { mem[1706:1706] } <= { data_i[26:26] };
    end 
    if(N4956) begin
      { mem[1705:1705] } <= { data_i[25:25] };
    end 
    if(N4955) begin
      { mem[1704:1704] } <= { data_i[24:24] };
    end 
    if(N4954) begin
      { mem[1703:1703] } <= { data_i[23:23] };
    end 
    if(N4953) begin
      { mem[1702:1702] } <= { data_i[22:22] };
    end 
    if(N4952) begin
      { mem[1701:1701] } <= { data_i[21:21] };
    end 
    if(N4951) begin
      { mem[1700:1700] } <= { data_i[20:20] };
    end 
    if(N4950) begin
      { mem[1699:1699] } <= { data_i[19:19] };
    end 
    if(N4949) begin
      { mem[1698:1698] } <= { data_i[18:18] };
    end 
    if(N4948) begin
      { mem[1697:1697] } <= { data_i[17:17] };
    end 
    if(N4947) begin
      { mem[1696:1696] } <= { data_i[16:16] };
    end 
    if(N4946) begin
      { mem[1695:1695] } <= { data_i[15:15] };
    end 
    if(N4945) begin
      { mem[1694:1694] } <= { data_i[14:14] };
    end 
    if(N4944) begin
      { mem[1693:1693] } <= { data_i[13:13] };
    end 
    if(N4943) begin
      { mem[1692:1692] } <= { data_i[12:12] };
    end 
    if(N4942) begin
      { mem[1691:1691] } <= { data_i[11:11] };
    end 
    if(N4941) begin
      { mem[1690:1690] } <= { data_i[10:10] };
    end 
    if(N4940) begin
      { mem[1689:1689] } <= { data_i[9:9] };
    end 
    if(N4939) begin
      { mem[1688:1688] } <= { data_i[8:8] };
    end 
    if(N4938) begin
      { mem[1687:1687] } <= { data_i[7:7] };
    end 
    if(N4937) begin
      { mem[1686:1686] } <= { data_i[6:6] };
    end 
    if(N4936) begin
      { mem[1685:1685] } <= { data_i[5:5] };
    end 
    if(N4935) begin
      { mem[1684:1684] } <= { data_i[4:4] };
    end 
    if(N4934) begin
      { mem[1683:1683] } <= { data_i[3:3] };
    end 
    if(N4933) begin
      { mem[1682:1682] } <= { data_i[2:2] };
    end 
    if(N4932) begin
      { mem[1681:1681] } <= { data_i[1:1] };
    end 
    if(N4931) begin
      { mem[1680:1680] } <= { data_i[0:0] };
    end 
    if(N4930) begin
      { mem[1679:1679] } <= { data_i[39:39] };
    end 
    if(N4929) begin
      { mem[1678:1678] } <= { data_i[38:38] };
    end 
    if(N4928) begin
      { mem[1677:1677] } <= { data_i[37:37] };
    end 
    if(N4927) begin
      { mem[1676:1676] } <= { data_i[36:36] };
    end 
    if(N4926) begin
      { mem[1675:1675] } <= { data_i[35:35] };
    end 
    if(N4925) begin
      { mem[1674:1674] } <= { data_i[34:34] };
    end 
    if(N4924) begin
      { mem[1673:1673] } <= { data_i[33:33] };
    end 
    if(N4923) begin
      { mem[1672:1672] } <= { data_i[32:32] };
    end 
    if(N4922) begin
      { mem[1671:1671] } <= { data_i[31:31] };
    end 
    if(N4921) begin
      { mem[1670:1670] } <= { data_i[30:30] };
    end 
    if(N4920) begin
      { mem[1669:1669] } <= { data_i[29:29] };
    end 
    if(N4919) begin
      { mem[1668:1668] } <= { data_i[28:28] };
    end 
    if(N4918) begin
      { mem[1667:1667] } <= { data_i[27:27] };
    end 
    if(N4917) begin
      { mem[1666:1666] } <= { data_i[26:26] };
    end 
    if(N4916) begin
      { mem[1665:1665] } <= { data_i[25:25] };
    end 
    if(N4915) begin
      { mem[1664:1664] } <= { data_i[24:24] };
    end 
    if(N4914) begin
      { mem[1663:1663] } <= { data_i[23:23] };
    end 
    if(N4913) begin
      { mem[1662:1662] } <= { data_i[22:22] };
    end 
    if(N4912) begin
      { mem[1661:1661] } <= { data_i[21:21] };
    end 
    if(N4911) begin
      { mem[1660:1660] } <= { data_i[20:20] };
    end 
    if(N4910) begin
      { mem[1659:1659] } <= { data_i[19:19] };
    end 
    if(N4909) begin
      { mem[1658:1658] } <= { data_i[18:18] };
    end 
    if(N4908) begin
      { mem[1657:1657] } <= { data_i[17:17] };
    end 
    if(N4907) begin
      { mem[1656:1656] } <= { data_i[16:16] };
    end 
    if(N4906) begin
      { mem[1655:1655] } <= { data_i[15:15] };
    end 
    if(N4905) begin
      { mem[1654:1654] } <= { data_i[14:14] };
    end 
    if(N4904) begin
      { mem[1653:1653] } <= { data_i[13:13] };
    end 
    if(N4903) begin
      { mem[1652:1652] } <= { data_i[12:12] };
    end 
    if(N4902) begin
      { mem[1651:1651] } <= { data_i[11:11] };
    end 
    if(N4901) begin
      { mem[1650:1650] } <= { data_i[10:10] };
    end 
    if(N4900) begin
      { mem[1649:1649] } <= { data_i[9:9] };
    end 
    if(N4899) begin
      { mem[1648:1648] } <= { data_i[8:8] };
    end 
    if(N4898) begin
      { mem[1647:1647] } <= { data_i[7:7] };
    end 
    if(N4897) begin
      { mem[1646:1646] } <= { data_i[6:6] };
    end 
    if(N4896) begin
      { mem[1645:1645] } <= { data_i[5:5] };
    end 
    if(N4895) begin
      { mem[1644:1644] } <= { data_i[4:4] };
    end 
    if(N4894) begin
      { mem[1643:1643] } <= { data_i[3:3] };
    end 
    if(N4893) begin
      { mem[1642:1642] } <= { data_i[2:2] };
    end 
    if(N4892) begin
      { mem[1641:1641] } <= { data_i[1:1] };
    end 
    if(N4891) begin
      { mem[1640:1640] } <= { data_i[0:0] };
    end 
    if(N4890) begin
      { mem[1639:1639] } <= { data_i[39:39] };
    end 
    if(N4889) begin
      { mem[1638:1638] } <= { data_i[38:38] };
    end 
    if(N4888) begin
      { mem[1637:1637] } <= { data_i[37:37] };
    end 
    if(N4887) begin
      { mem[1636:1636] } <= { data_i[36:36] };
    end 
    if(N4886) begin
      { mem[1635:1635] } <= { data_i[35:35] };
    end 
    if(N4885) begin
      { mem[1634:1634] } <= { data_i[34:34] };
    end 
    if(N4884) begin
      { mem[1633:1633] } <= { data_i[33:33] };
    end 
    if(N4883) begin
      { mem[1632:1632] } <= { data_i[32:32] };
    end 
    if(N4882) begin
      { mem[1631:1631] } <= { data_i[31:31] };
    end 
    if(N4881) begin
      { mem[1630:1630] } <= { data_i[30:30] };
    end 
    if(N4880) begin
      { mem[1629:1629] } <= { data_i[29:29] };
    end 
    if(N4879) begin
      { mem[1628:1628] } <= { data_i[28:28] };
    end 
    if(N4878) begin
      { mem[1627:1627] } <= { data_i[27:27] };
    end 
    if(N4877) begin
      { mem[1626:1626] } <= { data_i[26:26] };
    end 
    if(N4876) begin
      { mem[1625:1625] } <= { data_i[25:25] };
    end 
    if(N4875) begin
      { mem[1624:1624] } <= { data_i[24:24] };
    end 
    if(N4874) begin
      { mem[1623:1623] } <= { data_i[23:23] };
    end 
    if(N4873) begin
      { mem[1622:1622] } <= { data_i[22:22] };
    end 
    if(N4872) begin
      { mem[1621:1621] } <= { data_i[21:21] };
    end 
    if(N4871) begin
      { mem[1620:1620] } <= { data_i[20:20] };
    end 
    if(N4870) begin
      { mem[1619:1619] } <= { data_i[19:19] };
    end 
    if(N4869) begin
      { mem[1618:1618] } <= { data_i[18:18] };
    end 
    if(N4868) begin
      { mem[1617:1617] } <= { data_i[17:17] };
    end 
    if(N4867) begin
      { mem[1616:1616] } <= { data_i[16:16] };
    end 
    if(N4866) begin
      { mem[1615:1615] } <= { data_i[15:15] };
    end 
    if(N4865) begin
      { mem[1614:1614] } <= { data_i[14:14] };
    end 
    if(N4864) begin
      { mem[1613:1613] } <= { data_i[13:13] };
    end 
    if(N4863) begin
      { mem[1612:1612] } <= { data_i[12:12] };
    end 
    if(N4862) begin
      { mem[1611:1611] } <= { data_i[11:11] };
    end 
    if(N4861) begin
      { mem[1610:1610] } <= { data_i[10:10] };
    end 
    if(N4860) begin
      { mem[1609:1609] } <= { data_i[9:9] };
    end 
    if(N4859) begin
      { mem[1608:1608] } <= { data_i[8:8] };
    end 
    if(N4858) begin
      { mem[1607:1607] } <= { data_i[7:7] };
    end 
    if(N4857) begin
      { mem[1606:1606] } <= { data_i[6:6] };
    end 
    if(N4856) begin
      { mem[1605:1605] } <= { data_i[5:5] };
    end 
    if(N4855) begin
      { mem[1604:1604] } <= { data_i[4:4] };
    end 
    if(N4854) begin
      { mem[1603:1603] } <= { data_i[3:3] };
    end 
    if(N4853) begin
      { mem[1602:1602] } <= { data_i[2:2] };
    end 
    if(N4852) begin
      { mem[1601:1601] } <= { data_i[1:1] };
    end 
    if(N4851) begin
      { mem[1600:1600] } <= { data_i[0:0] };
    end 
    if(N4850) begin
      { mem[1599:1599] } <= { data_i[39:39] };
    end 
    if(N4849) begin
      { mem[1598:1598] } <= { data_i[38:38] };
    end 
    if(N4848) begin
      { mem[1597:1597] } <= { data_i[37:37] };
    end 
    if(N4847) begin
      { mem[1596:1596] } <= { data_i[36:36] };
    end 
    if(N4846) begin
      { mem[1595:1595] } <= { data_i[35:35] };
    end 
    if(N4845) begin
      { mem[1594:1594] } <= { data_i[34:34] };
    end 
    if(N4844) begin
      { mem[1593:1593] } <= { data_i[33:33] };
    end 
    if(N4843) begin
      { mem[1592:1592] } <= { data_i[32:32] };
    end 
    if(N4842) begin
      { mem[1591:1591] } <= { data_i[31:31] };
    end 
    if(N4841) begin
      { mem[1590:1590] } <= { data_i[30:30] };
    end 
    if(N4840) begin
      { mem[1589:1589] } <= { data_i[29:29] };
    end 
    if(N4839) begin
      { mem[1588:1588] } <= { data_i[28:28] };
    end 
    if(N4838) begin
      { mem[1587:1587] } <= { data_i[27:27] };
    end 
    if(N4837) begin
      { mem[1586:1586] } <= { data_i[26:26] };
    end 
    if(N4836) begin
      { mem[1585:1585] } <= { data_i[25:25] };
    end 
    if(N4835) begin
      { mem[1584:1584] } <= { data_i[24:24] };
    end 
    if(N4834) begin
      { mem[1583:1583] } <= { data_i[23:23] };
    end 
    if(N4833) begin
      { mem[1582:1582] } <= { data_i[22:22] };
    end 
    if(N4832) begin
      { mem[1581:1581] } <= { data_i[21:21] };
    end 
    if(N4831) begin
      { mem[1580:1580] } <= { data_i[20:20] };
    end 
    if(N4830) begin
      { mem[1579:1579] } <= { data_i[19:19] };
    end 
    if(N4829) begin
      { mem[1578:1578] } <= { data_i[18:18] };
    end 
    if(N4828) begin
      { mem[1577:1577] } <= { data_i[17:17] };
    end 
    if(N4827) begin
      { mem[1576:1576] } <= { data_i[16:16] };
    end 
    if(N4826) begin
      { mem[1575:1575] } <= { data_i[15:15] };
    end 
    if(N4825) begin
      { mem[1574:1574] } <= { data_i[14:14] };
    end 
    if(N4824) begin
      { mem[1573:1573] } <= { data_i[13:13] };
    end 
    if(N4823) begin
      { mem[1572:1572] } <= { data_i[12:12] };
    end 
    if(N4822) begin
      { mem[1571:1571] } <= { data_i[11:11] };
    end 
    if(N4821) begin
      { mem[1570:1570] } <= { data_i[10:10] };
    end 
    if(N4820) begin
      { mem[1569:1569] } <= { data_i[9:9] };
    end 
    if(N4819) begin
      { mem[1568:1568] } <= { data_i[8:8] };
    end 
    if(N4818) begin
      { mem[1567:1567] } <= { data_i[7:7] };
    end 
    if(N4817) begin
      { mem[1566:1566] } <= { data_i[6:6] };
    end 
    if(N4816) begin
      { mem[1565:1565] } <= { data_i[5:5] };
    end 
    if(N4815) begin
      { mem[1564:1564] } <= { data_i[4:4] };
    end 
    if(N4814) begin
      { mem[1563:1563] } <= { data_i[3:3] };
    end 
    if(N4813) begin
      { mem[1562:1562] } <= { data_i[2:2] };
    end 
    if(N4812) begin
      { mem[1561:1561] } <= { data_i[1:1] };
    end 
    if(N4811) begin
      { mem[1560:1560] } <= { data_i[0:0] };
    end 
    if(N4810) begin
      { mem[1559:1559] } <= { data_i[39:39] };
    end 
    if(N4809) begin
      { mem[1558:1558] } <= { data_i[38:38] };
    end 
    if(N4808) begin
      { mem[1557:1557] } <= { data_i[37:37] };
    end 
    if(N4807) begin
      { mem[1556:1556] } <= { data_i[36:36] };
    end 
    if(N4806) begin
      { mem[1555:1555] } <= { data_i[35:35] };
    end 
    if(N4805) begin
      { mem[1554:1554] } <= { data_i[34:34] };
    end 
    if(N4804) begin
      { mem[1553:1553] } <= { data_i[33:33] };
    end 
    if(N4803) begin
      { mem[1552:1552] } <= { data_i[32:32] };
    end 
    if(N4802) begin
      { mem[1551:1551] } <= { data_i[31:31] };
    end 
    if(N4801) begin
      { mem[1550:1550] } <= { data_i[30:30] };
    end 
    if(N4800) begin
      { mem[1549:1549] } <= { data_i[29:29] };
    end 
    if(N4799) begin
      { mem[1548:1548] } <= { data_i[28:28] };
    end 
    if(N4798) begin
      { mem[1547:1547] } <= { data_i[27:27] };
    end 
    if(N4797) begin
      { mem[1546:1546] } <= { data_i[26:26] };
    end 
    if(N4796) begin
      { mem[1545:1545] } <= { data_i[25:25] };
    end 
    if(N4795) begin
      { mem[1544:1544] } <= { data_i[24:24] };
    end 
    if(N4794) begin
      { mem[1543:1543] } <= { data_i[23:23] };
    end 
    if(N4793) begin
      { mem[1542:1542] } <= { data_i[22:22] };
    end 
    if(N4792) begin
      { mem[1541:1541] } <= { data_i[21:21] };
    end 
    if(N4791) begin
      { mem[1540:1540] } <= { data_i[20:20] };
    end 
    if(N4790) begin
      { mem[1539:1539] } <= { data_i[19:19] };
    end 
    if(N4789) begin
      { mem[1538:1538] } <= { data_i[18:18] };
    end 
    if(N4788) begin
      { mem[1537:1537] } <= { data_i[17:17] };
    end 
    if(N4787) begin
      { mem[1536:1536] } <= { data_i[16:16] };
    end 
    if(N4786) begin
      { mem[1535:1535] } <= { data_i[15:15] };
    end 
    if(N4785) begin
      { mem[1534:1534] } <= { data_i[14:14] };
    end 
    if(N4784) begin
      { mem[1533:1533] } <= { data_i[13:13] };
    end 
    if(N4783) begin
      { mem[1532:1532] } <= { data_i[12:12] };
    end 
    if(N4782) begin
      { mem[1531:1531] } <= { data_i[11:11] };
    end 
    if(N4781) begin
      { mem[1530:1530] } <= { data_i[10:10] };
    end 
    if(N4780) begin
      { mem[1529:1529] } <= { data_i[9:9] };
    end 
    if(N4779) begin
      { mem[1528:1528] } <= { data_i[8:8] };
    end 
    if(N4778) begin
      { mem[1527:1527] } <= { data_i[7:7] };
    end 
    if(N4777) begin
      { mem[1526:1526] } <= { data_i[6:6] };
    end 
    if(N4776) begin
      { mem[1525:1525] } <= { data_i[5:5] };
    end 
    if(N4775) begin
      { mem[1524:1524] } <= { data_i[4:4] };
    end 
    if(N4774) begin
      { mem[1523:1523] } <= { data_i[3:3] };
    end 
    if(N4773) begin
      { mem[1522:1522] } <= { data_i[2:2] };
    end 
    if(N4772) begin
      { mem[1521:1521] } <= { data_i[1:1] };
    end 
    if(N4771) begin
      { mem[1520:1520] } <= { data_i[0:0] };
    end 
    if(N4770) begin
      { mem[1519:1519] } <= { data_i[39:39] };
    end 
    if(N4769) begin
      { mem[1518:1518] } <= { data_i[38:38] };
    end 
    if(N4768) begin
      { mem[1517:1517] } <= { data_i[37:37] };
    end 
    if(N4767) begin
      { mem[1516:1516] } <= { data_i[36:36] };
    end 
    if(N4766) begin
      { mem[1515:1515] } <= { data_i[35:35] };
    end 
    if(N4765) begin
      { mem[1514:1514] } <= { data_i[34:34] };
    end 
    if(N4764) begin
      { mem[1513:1513] } <= { data_i[33:33] };
    end 
    if(N4763) begin
      { mem[1512:1512] } <= { data_i[32:32] };
    end 
    if(N4762) begin
      { mem[1511:1511] } <= { data_i[31:31] };
    end 
    if(N4761) begin
      { mem[1510:1510] } <= { data_i[30:30] };
    end 
    if(N4760) begin
      { mem[1509:1509] } <= { data_i[29:29] };
    end 
    if(N4759) begin
      { mem[1508:1508] } <= { data_i[28:28] };
    end 
    if(N4758) begin
      { mem[1507:1507] } <= { data_i[27:27] };
    end 
    if(N4757) begin
      { mem[1506:1506] } <= { data_i[26:26] };
    end 
    if(N4756) begin
      { mem[1505:1505] } <= { data_i[25:25] };
    end 
    if(N4755) begin
      { mem[1504:1504] } <= { data_i[24:24] };
    end 
    if(N4754) begin
      { mem[1503:1503] } <= { data_i[23:23] };
    end 
    if(N4753) begin
      { mem[1502:1502] } <= { data_i[22:22] };
    end 
    if(N4752) begin
      { mem[1501:1501] } <= { data_i[21:21] };
    end 
    if(N4751) begin
      { mem[1500:1500] } <= { data_i[20:20] };
    end 
    if(N4750) begin
      { mem[1499:1499] } <= { data_i[19:19] };
    end 
    if(N4749) begin
      { mem[1498:1498] } <= { data_i[18:18] };
    end 
    if(N4748) begin
      { mem[1497:1497] } <= { data_i[17:17] };
    end 
    if(N4747) begin
      { mem[1496:1496] } <= { data_i[16:16] };
    end 
    if(N4746) begin
      { mem[1495:1495] } <= { data_i[15:15] };
    end 
    if(N4745) begin
      { mem[1494:1494] } <= { data_i[14:14] };
    end 
    if(N4744) begin
      { mem[1493:1493] } <= { data_i[13:13] };
    end 
    if(N4743) begin
      { mem[1492:1492] } <= { data_i[12:12] };
    end 
    if(N4742) begin
      { mem[1491:1491] } <= { data_i[11:11] };
    end 
    if(N4741) begin
      { mem[1490:1490] } <= { data_i[10:10] };
    end 
    if(N4740) begin
      { mem[1489:1489] } <= { data_i[9:9] };
    end 
    if(N4739) begin
      { mem[1488:1488] } <= { data_i[8:8] };
    end 
    if(N4738) begin
      { mem[1487:1487] } <= { data_i[7:7] };
    end 
    if(N4737) begin
      { mem[1486:1486] } <= { data_i[6:6] };
    end 
    if(N4736) begin
      { mem[1485:1485] } <= { data_i[5:5] };
    end 
    if(N4735) begin
      { mem[1484:1484] } <= { data_i[4:4] };
    end 
    if(N4734) begin
      { mem[1483:1483] } <= { data_i[3:3] };
    end 
    if(N4733) begin
      { mem[1482:1482] } <= { data_i[2:2] };
    end 
    if(N4732) begin
      { mem[1481:1481] } <= { data_i[1:1] };
    end 
    if(N4731) begin
      { mem[1480:1480] } <= { data_i[0:0] };
    end 
    if(N4730) begin
      { mem[1479:1479] } <= { data_i[39:39] };
    end 
    if(N4729) begin
      { mem[1478:1478] } <= { data_i[38:38] };
    end 
    if(N4728) begin
      { mem[1477:1477] } <= { data_i[37:37] };
    end 
    if(N4727) begin
      { mem[1476:1476] } <= { data_i[36:36] };
    end 
    if(N4726) begin
      { mem[1475:1475] } <= { data_i[35:35] };
    end 
    if(N4725) begin
      { mem[1474:1474] } <= { data_i[34:34] };
    end 
    if(N4724) begin
      { mem[1473:1473] } <= { data_i[33:33] };
    end 
    if(N4723) begin
      { mem[1472:1472] } <= { data_i[32:32] };
    end 
    if(N4722) begin
      { mem[1471:1471] } <= { data_i[31:31] };
    end 
    if(N4721) begin
      { mem[1470:1470] } <= { data_i[30:30] };
    end 
    if(N4720) begin
      { mem[1469:1469] } <= { data_i[29:29] };
    end 
    if(N4719) begin
      { mem[1468:1468] } <= { data_i[28:28] };
    end 
    if(N4718) begin
      { mem[1467:1467] } <= { data_i[27:27] };
    end 
    if(N4717) begin
      { mem[1466:1466] } <= { data_i[26:26] };
    end 
    if(N4716) begin
      { mem[1465:1465] } <= { data_i[25:25] };
    end 
    if(N4715) begin
      { mem[1464:1464] } <= { data_i[24:24] };
    end 
    if(N4714) begin
      { mem[1463:1463] } <= { data_i[23:23] };
    end 
    if(N4713) begin
      { mem[1462:1462] } <= { data_i[22:22] };
    end 
    if(N4712) begin
      { mem[1461:1461] } <= { data_i[21:21] };
    end 
    if(N4711) begin
      { mem[1460:1460] } <= { data_i[20:20] };
    end 
    if(N4710) begin
      { mem[1459:1459] } <= { data_i[19:19] };
    end 
    if(N4709) begin
      { mem[1458:1458] } <= { data_i[18:18] };
    end 
    if(N4708) begin
      { mem[1457:1457] } <= { data_i[17:17] };
    end 
    if(N4707) begin
      { mem[1456:1456] } <= { data_i[16:16] };
    end 
    if(N4706) begin
      { mem[1455:1455] } <= { data_i[15:15] };
    end 
    if(N4705) begin
      { mem[1454:1454] } <= { data_i[14:14] };
    end 
    if(N4704) begin
      { mem[1453:1453] } <= { data_i[13:13] };
    end 
    if(N4703) begin
      { mem[1452:1452] } <= { data_i[12:12] };
    end 
    if(N4702) begin
      { mem[1451:1451] } <= { data_i[11:11] };
    end 
    if(N4701) begin
      { mem[1450:1450] } <= { data_i[10:10] };
    end 
    if(N4700) begin
      { mem[1449:1449] } <= { data_i[9:9] };
    end 
    if(N4699) begin
      { mem[1448:1448] } <= { data_i[8:8] };
    end 
    if(N4698) begin
      { mem[1447:1447] } <= { data_i[7:7] };
    end 
    if(N4697) begin
      { mem[1446:1446] } <= { data_i[6:6] };
    end 
    if(N4696) begin
      { mem[1445:1445] } <= { data_i[5:5] };
    end 
    if(N4695) begin
      { mem[1444:1444] } <= { data_i[4:4] };
    end 
    if(N4694) begin
      { mem[1443:1443] } <= { data_i[3:3] };
    end 
    if(N4693) begin
      { mem[1442:1442] } <= { data_i[2:2] };
    end 
    if(N4692) begin
      { mem[1441:1441] } <= { data_i[1:1] };
    end 
    if(N4691) begin
      { mem[1440:1440] } <= { data_i[0:0] };
    end 
    if(N4690) begin
      { mem[1439:1439] } <= { data_i[39:39] };
    end 
    if(N4689) begin
      { mem[1438:1438] } <= { data_i[38:38] };
    end 
    if(N4688) begin
      { mem[1437:1437] } <= { data_i[37:37] };
    end 
    if(N4687) begin
      { mem[1436:1436] } <= { data_i[36:36] };
    end 
    if(N4686) begin
      { mem[1435:1435] } <= { data_i[35:35] };
    end 
    if(N4685) begin
      { mem[1434:1434] } <= { data_i[34:34] };
    end 
    if(N4684) begin
      { mem[1433:1433] } <= { data_i[33:33] };
    end 
    if(N4683) begin
      { mem[1432:1432] } <= { data_i[32:32] };
    end 
    if(N4682) begin
      { mem[1431:1431] } <= { data_i[31:31] };
    end 
    if(N4681) begin
      { mem[1430:1430] } <= { data_i[30:30] };
    end 
    if(N4680) begin
      { mem[1429:1429] } <= { data_i[29:29] };
    end 
    if(N4679) begin
      { mem[1428:1428] } <= { data_i[28:28] };
    end 
    if(N4678) begin
      { mem[1427:1427] } <= { data_i[27:27] };
    end 
    if(N4677) begin
      { mem[1426:1426] } <= { data_i[26:26] };
    end 
    if(N4676) begin
      { mem[1425:1425] } <= { data_i[25:25] };
    end 
    if(N4675) begin
      { mem[1424:1424] } <= { data_i[24:24] };
    end 
    if(N4674) begin
      { mem[1423:1423] } <= { data_i[23:23] };
    end 
    if(N4673) begin
      { mem[1422:1422] } <= { data_i[22:22] };
    end 
    if(N4672) begin
      { mem[1421:1421] } <= { data_i[21:21] };
    end 
    if(N4671) begin
      { mem[1420:1420] } <= { data_i[20:20] };
    end 
    if(N4670) begin
      { mem[1419:1419] } <= { data_i[19:19] };
    end 
    if(N4669) begin
      { mem[1418:1418] } <= { data_i[18:18] };
    end 
    if(N4668) begin
      { mem[1417:1417] } <= { data_i[17:17] };
    end 
    if(N4667) begin
      { mem[1416:1416] } <= { data_i[16:16] };
    end 
    if(N4666) begin
      { mem[1415:1415] } <= { data_i[15:15] };
    end 
    if(N4665) begin
      { mem[1414:1414] } <= { data_i[14:14] };
    end 
    if(N4664) begin
      { mem[1413:1413] } <= { data_i[13:13] };
    end 
    if(N4663) begin
      { mem[1412:1412] } <= { data_i[12:12] };
    end 
    if(N4662) begin
      { mem[1411:1411] } <= { data_i[11:11] };
    end 
    if(N4661) begin
      { mem[1410:1410] } <= { data_i[10:10] };
    end 
    if(N4660) begin
      { mem[1409:1409] } <= { data_i[9:9] };
    end 
    if(N4659) begin
      { mem[1408:1408] } <= { data_i[8:8] };
    end 
    if(N4658) begin
      { mem[1407:1407] } <= { data_i[7:7] };
    end 
    if(N4657) begin
      { mem[1406:1406] } <= { data_i[6:6] };
    end 
    if(N4656) begin
      { mem[1405:1405] } <= { data_i[5:5] };
    end 
    if(N4655) begin
      { mem[1404:1404] } <= { data_i[4:4] };
    end 
    if(N4654) begin
      { mem[1403:1403] } <= { data_i[3:3] };
    end 
    if(N4653) begin
      { mem[1402:1402] } <= { data_i[2:2] };
    end 
    if(N4652) begin
      { mem[1401:1401] } <= { data_i[1:1] };
    end 
    if(N4651) begin
      { mem[1400:1400] } <= { data_i[0:0] };
    end 
    if(N4650) begin
      { mem[1399:1399] } <= { data_i[39:39] };
    end 
    if(N4649) begin
      { mem[1398:1398] } <= { data_i[38:38] };
    end 
    if(N4648) begin
      { mem[1397:1397] } <= { data_i[37:37] };
    end 
    if(N4647) begin
      { mem[1396:1396] } <= { data_i[36:36] };
    end 
    if(N4646) begin
      { mem[1395:1395] } <= { data_i[35:35] };
    end 
    if(N4645) begin
      { mem[1394:1394] } <= { data_i[34:34] };
    end 
    if(N4644) begin
      { mem[1393:1393] } <= { data_i[33:33] };
    end 
    if(N4643) begin
      { mem[1392:1392] } <= { data_i[32:32] };
    end 
    if(N4642) begin
      { mem[1391:1391] } <= { data_i[31:31] };
    end 
    if(N4641) begin
      { mem[1390:1390] } <= { data_i[30:30] };
    end 
    if(N4640) begin
      { mem[1389:1389] } <= { data_i[29:29] };
    end 
    if(N4639) begin
      { mem[1388:1388] } <= { data_i[28:28] };
    end 
    if(N4638) begin
      { mem[1387:1387] } <= { data_i[27:27] };
    end 
    if(N4637) begin
      { mem[1386:1386] } <= { data_i[26:26] };
    end 
    if(N4636) begin
      { mem[1385:1385] } <= { data_i[25:25] };
    end 
    if(N4635) begin
      { mem[1384:1384] } <= { data_i[24:24] };
    end 
    if(N4634) begin
      { mem[1383:1383] } <= { data_i[23:23] };
    end 
    if(N4633) begin
      { mem[1382:1382] } <= { data_i[22:22] };
    end 
    if(N4632) begin
      { mem[1381:1381] } <= { data_i[21:21] };
    end 
    if(N4631) begin
      { mem[1380:1380] } <= { data_i[20:20] };
    end 
    if(N4630) begin
      { mem[1379:1379] } <= { data_i[19:19] };
    end 
    if(N4629) begin
      { mem[1378:1378] } <= { data_i[18:18] };
    end 
    if(N4628) begin
      { mem[1377:1377] } <= { data_i[17:17] };
    end 
    if(N4627) begin
      { mem[1376:1376] } <= { data_i[16:16] };
    end 
    if(N4626) begin
      { mem[1375:1375] } <= { data_i[15:15] };
    end 
    if(N4625) begin
      { mem[1374:1374] } <= { data_i[14:14] };
    end 
    if(N4624) begin
      { mem[1373:1373] } <= { data_i[13:13] };
    end 
    if(N4623) begin
      { mem[1372:1372] } <= { data_i[12:12] };
    end 
    if(N4622) begin
      { mem[1371:1371] } <= { data_i[11:11] };
    end 
    if(N4621) begin
      { mem[1370:1370] } <= { data_i[10:10] };
    end 
    if(N4620) begin
      { mem[1369:1369] } <= { data_i[9:9] };
    end 
    if(N4619) begin
      { mem[1368:1368] } <= { data_i[8:8] };
    end 
    if(N4618) begin
      { mem[1367:1367] } <= { data_i[7:7] };
    end 
    if(N4617) begin
      { mem[1366:1366] } <= { data_i[6:6] };
    end 
    if(N4616) begin
      { mem[1365:1365] } <= { data_i[5:5] };
    end 
    if(N4615) begin
      { mem[1364:1364] } <= { data_i[4:4] };
    end 
    if(N4614) begin
      { mem[1363:1363] } <= { data_i[3:3] };
    end 
    if(N4613) begin
      { mem[1362:1362] } <= { data_i[2:2] };
    end 
    if(N4612) begin
      { mem[1361:1361] } <= { data_i[1:1] };
    end 
    if(N4611) begin
      { mem[1360:1360] } <= { data_i[0:0] };
    end 
    if(N4610) begin
      { mem[1359:1359] } <= { data_i[39:39] };
    end 
    if(N4609) begin
      { mem[1358:1358] } <= { data_i[38:38] };
    end 
    if(N4608) begin
      { mem[1357:1357] } <= { data_i[37:37] };
    end 
    if(N4607) begin
      { mem[1356:1356] } <= { data_i[36:36] };
    end 
    if(N4606) begin
      { mem[1355:1355] } <= { data_i[35:35] };
    end 
    if(N4605) begin
      { mem[1354:1354] } <= { data_i[34:34] };
    end 
    if(N4604) begin
      { mem[1353:1353] } <= { data_i[33:33] };
    end 
    if(N4603) begin
      { mem[1352:1352] } <= { data_i[32:32] };
    end 
    if(N4602) begin
      { mem[1351:1351] } <= { data_i[31:31] };
    end 
    if(N4601) begin
      { mem[1350:1350] } <= { data_i[30:30] };
    end 
    if(N4600) begin
      { mem[1349:1349] } <= { data_i[29:29] };
    end 
    if(N4599) begin
      { mem[1348:1348] } <= { data_i[28:28] };
    end 
    if(N4598) begin
      { mem[1347:1347] } <= { data_i[27:27] };
    end 
    if(N4597) begin
      { mem[1346:1346] } <= { data_i[26:26] };
    end 
    if(N4596) begin
      { mem[1345:1345] } <= { data_i[25:25] };
    end 
    if(N4595) begin
      { mem[1344:1344] } <= { data_i[24:24] };
    end 
    if(N4594) begin
      { mem[1343:1343] } <= { data_i[23:23] };
    end 
    if(N4593) begin
      { mem[1342:1342] } <= { data_i[22:22] };
    end 
    if(N4592) begin
      { mem[1341:1341] } <= { data_i[21:21] };
    end 
    if(N4591) begin
      { mem[1340:1340] } <= { data_i[20:20] };
    end 
    if(N4590) begin
      { mem[1339:1339] } <= { data_i[19:19] };
    end 
    if(N4589) begin
      { mem[1338:1338] } <= { data_i[18:18] };
    end 
    if(N4588) begin
      { mem[1337:1337] } <= { data_i[17:17] };
    end 
    if(N4587) begin
      { mem[1336:1336] } <= { data_i[16:16] };
    end 
    if(N4586) begin
      { mem[1335:1335] } <= { data_i[15:15] };
    end 
    if(N4585) begin
      { mem[1334:1334] } <= { data_i[14:14] };
    end 
    if(N4584) begin
      { mem[1333:1333] } <= { data_i[13:13] };
    end 
    if(N4583) begin
      { mem[1332:1332] } <= { data_i[12:12] };
    end 
    if(N4582) begin
      { mem[1331:1331] } <= { data_i[11:11] };
    end 
    if(N4581) begin
      { mem[1330:1330] } <= { data_i[10:10] };
    end 
    if(N4580) begin
      { mem[1329:1329] } <= { data_i[9:9] };
    end 
    if(N4579) begin
      { mem[1328:1328] } <= { data_i[8:8] };
    end 
    if(N4578) begin
      { mem[1327:1327] } <= { data_i[7:7] };
    end 
    if(N4577) begin
      { mem[1326:1326] } <= { data_i[6:6] };
    end 
    if(N4576) begin
      { mem[1325:1325] } <= { data_i[5:5] };
    end 
    if(N4575) begin
      { mem[1324:1324] } <= { data_i[4:4] };
    end 
    if(N4574) begin
      { mem[1323:1323] } <= { data_i[3:3] };
    end 
    if(N4573) begin
      { mem[1322:1322] } <= { data_i[2:2] };
    end 
    if(N4572) begin
      { mem[1321:1321] } <= { data_i[1:1] };
    end 
    if(N4571) begin
      { mem[1320:1320] } <= { data_i[0:0] };
    end 
    if(N4570) begin
      { mem[1319:1319] } <= { data_i[39:39] };
    end 
    if(N4569) begin
      { mem[1318:1318] } <= { data_i[38:38] };
    end 
    if(N4568) begin
      { mem[1317:1317] } <= { data_i[37:37] };
    end 
    if(N4567) begin
      { mem[1316:1316] } <= { data_i[36:36] };
    end 
    if(N4566) begin
      { mem[1315:1315] } <= { data_i[35:35] };
    end 
    if(N4565) begin
      { mem[1314:1314] } <= { data_i[34:34] };
    end 
    if(N4564) begin
      { mem[1313:1313] } <= { data_i[33:33] };
    end 
    if(N4563) begin
      { mem[1312:1312] } <= { data_i[32:32] };
    end 
    if(N4562) begin
      { mem[1311:1311] } <= { data_i[31:31] };
    end 
    if(N4561) begin
      { mem[1310:1310] } <= { data_i[30:30] };
    end 
    if(N4560) begin
      { mem[1309:1309] } <= { data_i[29:29] };
    end 
    if(N4559) begin
      { mem[1308:1308] } <= { data_i[28:28] };
    end 
    if(N4558) begin
      { mem[1307:1307] } <= { data_i[27:27] };
    end 
    if(N4557) begin
      { mem[1306:1306] } <= { data_i[26:26] };
    end 
    if(N4556) begin
      { mem[1305:1305] } <= { data_i[25:25] };
    end 
    if(N4555) begin
      { mem[1304:1304] } <= { data_i[24:24] };
    end 
    if(N4554) begin
      { mem[1303:1303] } <= { data_i[23:23] };
    end 
    if(N4553) begin
      { mem[1302:1302] } <= { data_i[22:22] };
    end 
    if(N4552) begin
      { mem[1301:1301] } <= { data_i[21:21] };
    end 
    if(N4551) begin
      { mem[1300:1300] } <= { data_i[20:20] };
    end 
    if(N4550) begin
      { mem[1299:1299] } <= { data_i[19:19] };
    end 
    if(N4549) begin
      { mem[1298:1298] } <= { data_i[18:18] };
    end 
    if(N4548) begin
      { mem[1297:1297] } <= { data_i[17:17] };
    end 
    if(N4547) begin
      { mem[1296:1296] } <= { data_i[16:16] };
    end 
    if(N4546) begin
      { mem[1295:1295] } <= { data_i[15:15] };
    end 
    if(N4545) begin
      { mem[1294:1294] } <= { data_i[14:14] };
    end 
    if(N4544) begin
      { mem[1293:1293] } <= { data_i[13:13] };
    end 
    if(N4543) begin
      { mem[1292:1292] } <= { data_i[12:12] };
    end 
    if(N4542) begin
      { mem[1291:1291] } <= { data_i[11:11] };
    end 
    if(N4541) begin
      { mem[1290:1290] } <= { data_i[10:10] };
    end 
    if(N4540) begin
      { mem[1289:1289] } <= { data_i[9:9] };
    end 
    if(N4539) begin
      { mem[1288:1288] } <= { data_i[8:8] };
    end 
    if(N4538) begin
      { mem[1287:1287] } <= { data_i[7:7] };
    end 
    if(N4537) begin
      { mem[1286:1286] } <= { data_i[6:6] };
    end 
    if(N4536) begin
      { mem[1285:1285] } <= { data_i[5:5] };
    end 
    if(N4535) begin
      { mem[1284:1284] } <= { data_i[4:4] };
    end 
    if(N4534) begin
      { mem[1283:1283] } <= { data_i[3:3] };
    end 
    if(N4533) begin
      { mem[1282:1282] } <= { data_i[2:2] };
    end 
    if(N4532) begin
      { mem[1281:1281] } <= { data_i[1:1] };
    end 
    if(N4531) begin
      { mem[1280:1280] } <= { data_i[0:0] };
    end 
    if(N4530) begin
      { mem[1279:1279] } <= { data_i[39:39] };
    end 
    if(N4529) begin
      { mem[1278:1278] } <= { data_i[38:38] };
    end 
    if(N4528) begin
      { mem[1277:1277] } <= { data_i[37:37] };
    end 
    if(N4527) begin
      { mem[1276:1276] } <= { data_i[36:36] };
    end 
    if(N4526) begin
      { mem[1275:1275] } <= { data_i[35:35] };
    end 
    if(N4525) begin
      { mem[1274:1274] } <= { data_i[34:34] };
    end 
    if(N4524) begin
      { mem[1273:1273] } <= { data_i[33:33] };
    end 
    if(N4523) begin
      { mem[1272:1272] } <= { data_i[32:32] };
    end 
    if(N4522) begin
      { mem[1271:1271] } <= { data_i[31:31] };
    end 
    if(N4521) begin
      { mem[1270:1270] } <= { data_i[30:30] };
    end 
    if(N4520) begin
      { mem[1269:1269] } <= { data_i[29:29] };
    end 
    if(N4519) begin
      { mem[1268:1268] } <= { data_i[28:28] };
    end 
    if(N4518) begin
      { mem[1267:1267] } <= { data_i[27:27] };
    end 
    if(N4517) begin
      { mem[1266:1266] } <= { data_i[26:26] };
    end 
    if(N4516) begin
      { mem[1265:1265] } <= { data_i[25:25] };
    end 
    if(N4515) begin
      { mem[1264:1264] } <= { data_i[24:24] };
    end 
    if(N4514) begin
      { mem[1263:1263] } <= { data_i[23:23] };
    end 
    if(N4513) begin
      { mem[1262:1262] } <= { data_i[22:22] };
    end 
    if(N4512) begin
      { mem[1261:1261] } <= { data_i[21:21] };
    end 
    if(N4511) begin
      { mem[1260:1260] } <= { data_i[20:20] };
    end 
    if(N4510) begin
      { mem[1259:1259] } <= { data_i[19:19] };
    end 
    if(N4509) begin
      { mem[1258:1258] } <= { data_i[18:18] };
    end 
    if(N4508) begin
      { mem[1257:1257] } <= { data_i[17:17] };
    end 
    if(N4507) begin
      { mem[1256:1256] } <= { data_i[16:16] };
    end 
    if(N4506) begin
      { mem[1255:1255] } <= { data_i[15:15] };
    end 
    if(N4505) begin
      { mem[1254:1254] } <= { data_i[14:14] };
    end 
    if(N4504) begin
      { mem[1253:1253] } <= { data_i[13:13] };
    end 
    if(N4503) begin
      { mem[1252:1252] } <= { data_i[12:12] };
    end 
    if(N4502) begin
      { mem[1251:1251] } <= { data_i[11:11] };
    end 
    if(N4501) begin
      { mem[1250:1250] } <= { data_i[10:10] };
    end 
    if(N4500) begin
      { mem[1249:1249] } <= { data_i[9:9] };
    end 
    if(N4499) begin
      { mem[1248:1248] } <= { data_i[8:8] };
    end 
    if(N4498) begin
      { mem[1247:1247] } <= { data_i[7:7] };
    end 
    if(N4497) begin
      { mem[1246:1246] } <= { data_i[6:6] };
    end 
    if(N4496) begin
      { mem[1245:1245] } <= { data_i[5:5] };
    end 
    if(N4495) begin
      { mem[1244:1244] } <= { data_i[4:4] };
    end 
    if(N4494) begin
      { mem[1243:1243] } <= { data_i[3:3] };
    end 
    if(N4493) begin
      { mem[1242:1242] } <= { data_i[2:2] };
    end 
    if(N4492) begin
      { mem[1241:1241] } <= { data_i[1:1] };
    end 
    if(N4491) begin
      { mem[1240:1240] } <= { data_i[0:0] };
    end 
    if(N4490) begin
      { mem[1239:1239] } <= { data_i[39:39] };
    end 
    if(N4489) begin
      { mem[1238:1238] } <= { data_i[38:38] };
    end 
    if(N4488) begin
      { mem[1237:1237] } <= { data_i[37:37] };
    end 
    if(N4487) begin
      { mem[1236:1236] } <= { data_i[36:36] };
    end 
    if(N4486) begin
      { mem[1235:1235] } <= { data_i[35:35] };
    end 
    if(N4485) begin
      { mem[1234:1234] } <= { data_i[34:34] };
    end 
    if(N4484) begin
      { mem[1233:1233] } <= { data_i[33:33] };
    end 
    if(N4483) begin
      { mem[1232:1232] } <= { data_i[32:32] };
    end 
    if(N4482) begin
      { mem[1231:1231] } <= { data_i[31:31] };
    end 
    if(N4481) begin
      { mem[1230:1230] } <= { data_i[30:30] };
    end 
    if(N4480) begin
      { mem[1229:1229] } <= { data_i[29:29] };
    end 
    if(N4479) begin
      { mem[1228:1228] } <= { data_i[28:28] };
    end 
    if(N4478) begin
      { mem[1227:1227] } <= { data_i[27:27] };
    end 
    if(N4477) begin
      { mem[1226:1226] } <= { data_i[26:26] };
    end 
    if(N4476) begin
      { mem[1225:1225] } <= { data_i[25:25] };
    end 
    if(N4475) begin
      { mem[1224:1224] } <= { data_i[24:24] };
    end 
    if(N4474) begin
      { mem[1223:1223] } <= { data_i[23:23] };
    end 
    if(N4473) begin
      { mem[1222:1222] } <= { data_i[22:22] };
    end 
    if(N4472) begin
      { mem[1221:1221] } <= { data_i[21:21] };
    end 
    if(N4471) begin
      { mem[1220:1220] } <= { data_i[20:20] };
    end 
    if(N4470) begin
      { mem[1219:1219] } <= { data_i[19:19] };
    end 
    if(N4469) begin
      { mem[1218:1218] } <= { data_i[18:18] };
    end 
    if(N4468) begin
      { mem[1217:1217] } <= { data_i[17:17] };
    end 
    if(N4467) begin
      { mem[1216:1216] } <= { data_i[16:16] };
    end 
    if(N4466) begin
      { mem[1215:1215] } <= { data_i[15:15] };
    end 
    if(N4465) begin
      { mem[1214:1214] } <= { data_i[14:14] };
    end 
    if(N4464) begin
      { mem[1213:1213] } <= { data_i[13:13] };
    end 
    if(N4463) begin
      { mem[1212:1212] } <= { data_i[12:12] };
    end 
    if(N4462) begin
      { mem[1211:1211] } <= { data_i[11:11] };
    end 
    if(N4461) begin
      { mem[1210:1210] } <= { data_i[10:10] };
    end 
    if(N4460) begin
      { mem[1209:1209] } <= { data_i[9:9] };
    end 
    if(N4459) begin
      { mem[1208:1208] } <= { data_i[8:8] };
    end 
    if(N4458) begin
      { mem[1207:1207] } <= { data_i[7:7] };
    end 
    if(N4457) begin
      { mem[1206:1206] } <= { data_i[6:6] };
    end 
    if(N4456) begin
      { mem[1205:1205] } <= { data_i[5:5] };
    end 
    if(N4455) begin
      { mem[1204:1204] } <= { data_i[4:4] };
    end 
    if(N4454) begin
      { mem[1203:1203] } <= { data_i[3:3] };
    end 
    if(N4453) begin
      { mem[1202:1202] } <= { data_i[2:2] };
    end 
    if(N4452) begin
      { mem[1201:1201] } <= { data_i[1:1] };
    end 
    if(N4451) begin
      { mem[1200:1200] } <= { data_i[0:0] };
    end 
    if(N4450) begin
      { mem[1199:1199] } <= { data_i[39:39] };
    end 
    if(N4449) begin
      { mem[1198:1198] } <= { data_i[38:38] };
    end 
    if(N4448) begin
      { mem[1197:1197] } <= { data_i[37:37] };
    end 
    if(N4447) begin
      { mem[1196:1196] } <= { data_i[36:36] };
    end 
    if(N4446) begin
      { mem[1195:1195] } <= { data_i[35:35] };
    end 
    if(N4445) begin
      { mem[1194:1194] } <= { data_i[34:34] };
    end 
    if(N4444) begin
      { mem[1193:1193] } <= { data_i[33:33] };
    end 
    if(N4443) begin
      { mem[1192:1192] } <= { data_i[32:32] };
    end 
    if(N4442) begin
      { mem[1191:1191] } <= { data_i[31:31] };
    end 
    if(N4441) begin
      { mem[1190:1190] } <= { data_i[30:30] };
    end 
    if(N4440) begin
      { mem[1189:1189] } <= { data_i[29:29] };
    end 
    if(N4439) begin
      { mem[1188:1188] } <= { data_i[28:28] };
    end 
    if(N4438) begin
      { mem[1187:1187] } <= { data_i[27:27] };
    end 
    if(N4437) begin
      { mem[1186:1186] } <= { data_i[26:26] };
    end 
    if(N4436) begin
      { mem[1185:1185] } <= { data_i[25:25] };
    end 
    if(N4435) begin
      { mem[1184:1184] } <= { data_i[24:24] };
    end 
    if(N4434) begin
      { mem[1183:1183] } <= { data_i[23:23] };
    end 
    if(N4433) begin
      { mem[1182:1182] } <= { data_i[22:22] };
    end 
    if(N4432) begin
      { mem[1181:1181] } <= { data_i[21:21] };
    end 
    if(N4431) begin
      { mem[1180:1180] } <= { data_i[20:20] };
    end 
    if(N4430) begin
      { mem[1179:1179] } <= { data_i[19:19] };
    end 
    if(N4429) begin
      { mem[1178:1178] } <= { data_i[18:18] };
    end 
    if(N4428) begin
      { mem[1177:1177] } <= { data_i[17:17] };
    end 
    if(N4427) begin
      { mem[1176:1176] } <= { data_i[16:16] };
    end 
    if(N4426) begin
      { mem[1175:1175] } <= { data_i[15:15] };
    end 
    if(N4425) begin
      { mem[1174:1174] } <= { data_i[14:14] };
    end 
    if(N4424) begin
      { mem[1173:1173] } <= { data_i[13:13] };
    end 
    if(N4423) begin
      { mem[1172:1172] } <= { data_i[12:12] };
    end 
    if(N4422) begin
      { mem[1171:1171] } <= { data_i[11:11] };
    end 
    if(N4421) begin
      { mem[1170:1170] } <= { data_i[10:10] };
    end 
    if(N4420) begin
      { mem[1169:1169] } <= { data_i[9:9] };
    end 
    if(N4419) begin
      { mem[1168:1168] } <= { data_i[8:8] };
    end 
    if(N4418) begin
      { mem[1167:1167] } <= { data_i[7:7] };
    end 
    if(N4417) begin
      { mem[1166:1166] } <= { data_i[6:6] };
    end 
    if(N4416) begin
      { mem[1165:1165] } <= { data_i[5:5] };
    end 
    if(N4415) begin
      { mem[1164:1164] } <= { data_i[4:4] };
    end 
    if(N4414) begin
      { mem[1163:1163] } <= { data_i[3:3] };
    end 
    if(N4413) begin
      { mem[1162:1162] } <= { data_i[2:2] };
    end 
    if(N4412) begin
      { mem[1161:1161] } <= { data_i[1:1] };
    end 
    if(N4411) begin
      { mem[1160:1160] } <= { data_i[0:0] };
    end 
    if(N4410) begin
      { mem[1159:1159] } <= { data_i[39:39] };
    end 
    if(N4409) begin
      { mem[1158:1158] } <= { data_i[38:38] };
    end 
    if(N4408) begin
      { mem[1157:1157] } <= { data_i[37:37] };
    end 
    if(N4407) begin
      { mem[1156:1156] } <= { data_i[36:36] };
    end 
    if(N4406) begin
      { mem[1155:1155] } <= { data_i[35:35] };
    end 
    if(N4405) begin
      { mem[1154:1154] } <= { data_i[34:34] };
    end 
    if(N4404) begin
      { mem[1153:1153] } <= { data_i[33:33] };
    end 
    if(N4403) begin
      { mem[1152:1152] } <= { data_i[32:32] };
    end 
    if(N4402) begin
      { mem[1151:1151] } <= { data_i[31:31] };
    end 
    if(N4401) begin
      { mem[1150:1150] } <= { data_i[30:30] };
    end 
    if(N4400) begin
      { mem[1149:1149] } <= { data_i[29:29] };
    end 
    if(N4399) begin
      { mem[1148:1148] } <= { data_i[28:28] };
    end 
    if(N4398) begin
      { mem[1147:1147] } <= { data_i[27:27] };
    end 
    if(N4397) begin
      { mem[1146:1146] } <= { data_i[26:26] };
    end 
    if(N4396) begin
      { mem[1145:1145] } <= { data_i[25:25] };
    end 
    if(N4395) begin
      { mem[1144:1144] } <= { data_i[24:24] };
    end 
    if(N4394) begin
      { mem[1143:1143] } <= { data_i[23:23] };
    end 
    if(N4393) begin
      { mem[1142:1142] } <= { data_i[22:22] };
    end 
    if(N4392) begin
      { mem[1141:1141] } <= { data_i[21:21] };
    end 
    if(N4391) begin
      { mem[1140:1140] } <= { data_i[20:20] };
    end 
    if(N4390) begin
      { mem[1139:1139] } <= { data_i[19:19] };
    end 
    if(N4389) begin
      { mem[1138:1138] } <= { data_i[18:18] };
    end 
    if(N4388) begin
      { mem[1137:1137] } <= { data_i[17:17] };
    end 
    if(N4387) begin
      { mem[1136:1136] } <= { data_i[16:16] };
    end 
    if(N4386) begin
      { mem[1135:1135] } <= { data_i[15:15] };
    end 
    if(N4385) begin
      { mem[1134:1134] } <= { data_i[14:14] };
    end 
    if(N4384) begin
      { mem[1133:1133] } <= { data_i[13:13] };
    end 
    if(N4383) begin
      { mem[1132:1132] } <= { data_i[12:12] };
    end 
    if(N4382) begin
      { mem[1131:1131] } <= { data_i[11:11] };
    end 
    if(N4381) begin
      { mem[1130:1130] } <= { data_i[10:10] };
    end 
    if(N4380) begin
      { mem[1129:1129] } <= { data_i[9:9] };
    end 
    if(N4379) begin
      { mem[1128:1128] } <= { data_i[8:8] };
    end 
    if(N4378) begin
      { mem[1127:1127] } <= { data_i[7:7] };
    end 
    if(N4377) begin
      { mem[1126:1126] } <= { data_i[6:6] };
    end 
    if(N4376) begin
      { mem[1125:1125] } <= { data_i[5:5] };
    end 
    if(N4375) begin
      { mem[1124:1124] } <= { data_i[4:4] };
    end 
    if(N4374) begin
      { mem[1123:1123] } <= { data_i[3:3] };
    end 
    if(N4373) begin
      { mem[1122:1122] } <= { data_i[2:2] };
    end 
    if(N4372) begin
      { mem[1121:1121] } <= { data_i[1:1] };
    end 
    if(N4371) begin
      { mem[1120:1120] } <= { data_i[0:0] };
    end 
    if(N4370) begin
      { mem[1119:1119] } <= { data_i[39:39] };
    end 
    if(N4369) begin
      { mem[1118:1118] } <= { data_i[38:38] };
    end 
    if(N4368) begin
      { mem[1117:1117] } <= { data_i[37:37] };
    end 
    if(N4367) begin
      { mem[1116:1116] } <= { data_i[36:36] };
    end 
    if(N4366) begin
      { mem[1115:1115] } <= { data_i[35:35] };
    end 
    if(N4365) begin
      { mem[1114:1114] } <= { data_i[34:34] };
    end 
    if(N4364) begin
      { mem[1113:1113] } <= { data_i[33:33] };
    end 
    if(N4363) begin
      { mem[1112:1112] } <= { data_i[32:32] };
    end 
    if(N4362) begin
      { mem[1111:1111] } <= { data_i[31:31] };
    end 
    if(N4361) begin
      { mem[1110:1110] } <= { data_i[30:30] };
    end 
    if(N4360) begin
      { mem[1109:1109] } <= { data_i[29:29] };
    end 
    if(N4359) begin
      { mem[1108:1108] } <= { data_i[28:28] };
    end 
    if(N4358) begin
      { mem[1107:1107] } <= { data_i[27:27] };
    end 
    if(N4357) begin
      { mem[1106:1106] } <= { data_i[26:26] };
    end 
    if(N4356) begin
      { mem[1105:1105] } <= { data_i[25:25] };
    end 
    if(N4355) begin
      { mem[1104:1104] } <= { data_i[24:24] };
    end 
    if(N4354) begin
      { mem[1103:1103] } <= { data_i[23:23] };
    end 
    if(N4353) begin
      { mem[1102:1102] } <= { data_i[22:22] };
    end 
    if(N4352) begin
      { mem[1101:1101] } <= { data_i[21:21] };
    end 
    if(N4351) begin
      { mem[1100:1100] } <= { data_i[20:20] };
    end 
    if(N4350) begin
      { mem[1099:1099] } <= { data_i[19:19] };
    end 
    if(N4349) begin
      { mem[1098:1098] } <= { data_i[18:18] };
    end 
    if(N4348) begin
      { mem[1097:1097] } <= { data_i[17:17] };
    end 
    if(N4347) begin
      { mem[1096:1096] } <= { data_i[16:16] };
    end 
    if(N4346) begin
      { mem[1095:1095] } <= { data_i[15:15] };
    end 
    if(N4345) begin
      { mem[1094:1094] } <= { data_i[14:14] };
    end 
    if(N4344) begin
      { mem[1093:1093] } <= { data_i[13:13] };
    end 
    if(N4343) begin
      { mem[1092:1092] } <= { data_i[12:12] };
    end 
    if(N4342) begin
      { mem[1091:1091] } <= { data_i[11:11] };
    end 
    if(N4341) begin
      { mem[1090:1090] } <= { data_i[10:10] };
    end 
    if(N4340) begin
      { mem[1089:1089] } <= { data_i[9:9] };
    end 
    if(N4339) begin
      { mem[1088:1088] } <= { data_i[8:8] };
    end 
    if(N4338) begin
      { mem[1087:1087] } <= { data_i[7:7] };
    end 
    if(N4337) begin
      { mem[1086:1086] } <= { data_i[6:6] };
    end 
    if(N4336) begin
      { mem[1085:1085] } <= { data_i[5:5] };
    end 
    if(N4335) begin
      { mem[1084:1084] } <= { data_i[4:4] };
    end 
    if(N4334) begin
      { mem[1083:1083] } <= { data_i[3:3] };
    end 
    if(N4333) begin
      { mem[1082:1082] } <= { data_i[2:2] };
    end 
    if(N4332) begin
      { mem[1081:1081] } <= { data_i[1:1] };
    end 
    if(N4331) begin
      { mem[1080:1080] } <= { data_i[0:0] };
    end 
    if(N4330) begin
      { mem[1079:1079] } <= { data_i[39:39] };
    end 
    if(N4329) begin
      { mem[1078:1078] } <= { data_i[38:38] };
    end 
    if(N4328) begin
      { mem[1077:1077] } <= { data_i[37:37] };
    end 
    if(N4327) begin
      { mem[1076:1076] } <= { data_i[36:36] };
    end 
    if(N4326) begin
      { mem[1075:1075] } <= { data_i[35:35] };
    end 
    if(N4325) begin
      { mem[1074:1074] } <= { data_i[34:34] };
    end 
    if(N4324) begin
      { mem[1073:1073] } <= { data_i[33:33] };
    end 
    if(N4323) begin
      { mem[1072:1072] } <= { data_i[32:32] };
    end 
    if(N4322) begin
      { mem[1071:1071] } <= { data_i[31:31] };
    end 
    if(N4321) begin
      { mem[1070:1070] } <= { data_i[30:30] };
    end 
    if(N4320) begin
      { mem[1069:1069] } <= { data_i[29:29] };
    end 
    if(N4319) begin
      { mem[1068:1068] } <= { data_i[28:28] };
    end 
    if(N4318) begin
      { mem[1067:1067] } <= { data_i[27:27] };
    end 
    if(N4317) begin
      { mem[1066:1066] } <= { data_i[26:26] };
    end 
    if(N4316) begin
      { mem[1065:1065] } <= { data_i[25:25] };
    end 
    if(N4315) begin
      { mem[1064:1064] } <= { data_i[24:24] };
    end 
    if(N4314) begin
      { mem[1063:1063] } <= { data_i[23:23] };
    end 
    if(N4313) begin
      { mem[1062:1062] } <= { data_i[22:22] };
    end 
    if(N4312) begin
      { mem[1061:1061] } <= { data_i[21:21] };
    end 
    if(N4311) begin
      { mem[1060:1060] } <= { data_i[20:20] };
    end 
    if(N4310) begin
      { mem[1059:1059] } <= { data_i[19:19] };
    end 
    if(N4309) begin
      { mem[1058:1058] } <= { data_i[18:18] };
    end 
    if(N4308) begin
      { mem[1057:1057] } <= { data_i[17:17] };
    end 
    if(N4307) begin
      { mem[1056:1056] } <= { data_i[16:16] };
    end 
    if(N4306) begin
      { mem[1055:1055] } <= { data_i[15:15] };
    end 
    if(N4305) begin
      { mem[1054:1054] } <= { data_i[14:14] };
    end 
    if(N4304) begin
      { mem[1053:1053] } <= { data_i[13:13] };
    end 
    if(N4303) begin
      { mem[1052:1052] } <= { data_i[12:12] };
    end 
    if(N4302) begin
      { mem[1051:1051] } <= { data_i[11:11] };
    end 
    if(N4301) begin
      { mem[1050:1050] } <= { data_i[10:10] };
    end 
    if(N4300) begin
      { mem[1049:1049] } <= { data_i[9:9] };
    end 
    if(N4299) begin
      { mem[1048:1048] } <= { data_i[8:8] };
    end 
    if(N4298) begin
      { mem[1047:1047] } <= { data_i[7:7] };
    end 
    if(N4297) begin
      { mem[1046:1046] } <= { data_i[6:6] };
    end 
    if(N4296) begin
      { mem[1045:1045] } <= { data_i[5:5] };
    end 
    if(N4295) begin
      { mem[1044:1044] } <= { data_i[4:4] };
    end 
    if(N4294) begin
      { mem[1043:1043] } <= { data_i[3:3] };
    end 
    if(N4293) begin
      { mem[1042:1042] } <= { data_i[2:2] };
    end 
    if(N4292) begin
      { mem[1041:1041] } <= { data_i[1:1] };
    end 
    if(N4291) begin
      { mem[1040:1040] } <= { data_i[0:0] };
    end 
    if(N4290) begin
      { mem[1039:1039] } <= { data_i[39:39] };
    end 
    if(N4289) begin
      { mem[1038:1038] } <= { data_i[38:38] };
    end 
    if(N4288) begin
      { mem[1037:1037] } <= { data_i[37:37] };
    end 
    if(N4287) begin
      { mem[1036:1036] } <= { data_i[36:36] };
    end 
    if(N4286) begin
      { mem[1035:1035] } <= { data_i[35:35] };
    end 
    if(N4285) begin
      { mem[1034:1034] } <= { data_i[34:34] };
    end 
    if(N4284) begin
      { mem[1033:1033] } <= { data_i[33:33] };
    end 
    if(N4283) begin
      { mem[1032:1032] } <= { data_i[32:32] };
    end 
    if(N4282) begin
      { mem[1031:1031] } <= { data_i[31:31] };
    end 
    if(N4281) begin
      { mem[1030:1030] } <= { data_i[30:30] };
    end 
    if(N4280) begin
      { mem[1029:1029] } <= { data_i[29:29] };
    end 
    if(N4279) begin
      { mem[1028:1028] } <= { data_i[28:28] };
    end 
    if(N4278) begin
      { mem[1027:1027] } <= { data_i[27:27] };
    end 
    if(N4277) begin
      { mem[1026:1026] } <= { data_i[26:26] };
    end 
    if(N4276) begin
      { mem[1025:1025] } <= { data_i[25:25] };
    end 
    if(N4275) begin
      { mem[1024:1024] } <= { data_i[24:24] };
    end 
    if(N4274) begin
      { mem[1023:1023] } <= { data_i[23:23] };
    end 
    if(N4273) begin
      { mem[1022:1022] } <= { data_i[22:22] };
    end 
    if(N4272) begin
      { mem[1021:1021] } <= { data_i[21:21] };
    end 
    if(N4271) begin
      { mem[1020:1020] } <= { data_i[20:20] };
    end 
    if(N4270) begin
      { mem[1019:1019] } <= { data_i[19:19] };
    end 
    if(N4269) begin
      { mem[1018:1018] } <= { data_i[18:18] };
    end 
    if(N4268) begin
      { mem[1017:1017] } <= { data_i[17:17] };
    end 
    if(N4267) begin
      { mem[1016:1016] } <= { data_i[16:16] };
    end 
    if(N4266) begin
      { mem[1015:1015] } <= { data_i[15:15] };
    end 
    if(N4265) begin
      { mem[1014:1014] } <= { data_i[14:14] };
    end 
    if(N4264) begin
      { mem[1013:1013] } <= { data_i[13:13] };
    end 
    if(N4263) begin
      { mem[1012:1012] } <= { data_i[12:12] };
    end 
    if(N4262) begin
      { mem[1011:1011] } <= { data_i[11:11] };
    end 
    if(N4261) begin
      { mem[1010:1010] } <= { data_i[10:10] };
    end 
    if(N4260) begin
      { mem[1009:1009] } <= { data_i[9:9] };
    end 
    if(N4259) begin
      { mem[1008:1008] } <= { data_i[8:8] };
    end 
    if(N4258) begin
      { mem[1007:1007] } <= { data_i[7:7] };
    end 
    if(N4257) begin
      { mem[1006:1006] } <= { data_i[6:6] };
    end 
    if(N4256) begin
      { mem[1005:1005] } <= { data_i[5:5] };
    end 
    if(N4255) begin
      { mem[1004:1004] } <= { data_i[4:4] };
    end 
    if(N4254) begin
      { mem[1003:1003] } <= { data_i[3:3] };
    end 
    if(N4253) begin
      { mem[1002:1002] } <= { data_i[2:2] };
    end 
    if(N4252) begin
      { mem[1001:1001] } <= { data_i[1:1] };
    end 
    if(N4251) begin
      { mem[1000:1000] } <= { data_i[0:0] };
    end 
    if(N4250) begin
      { mem[999:999] } <= { data_i[39:39] };
    end 
    if(N4249) begin
      { mem[998:998] } <= { data_i[38:38] };
    end 
    if(N4248) begin
      { mem[997:997] } <= { data_i[37:37] };
    end 
    if(N4247) begin
      { mem[996:996] } <= { data_i[36:36] };
    end 
    if(N4246) begin
      { mem[995:995] } <= { data_i[35:35] };
    end 
    if(N4245) begin
      { mem[994:994] } <= { data_i[34:34] };
    end 
    if(N4244) begin
      { mem[993:993] } <= { data_i[33:33] };
    end 
    if(N4243) begin
      { mem[992:992] } <= { data_i[32:32] };
    end 
    if(N4242) begin
      { mem[991:991] } <= { data_i[31:31] };
    end 
    if(N4241) begin
      { mem[990:990] } <= { data_i[30:30] };
    end 
    if(N4240) begin
      { mem[989:989] } <= { data_i[29:29] };
    end 
    if(N4239) begin
      { mem[988:988] } <= { data_i[28:28] };
    end 
    if(N4238) begin
      { mem[987:987] } <= { data_i[27:27] };
    end 
    if(N4237) begin
      { mem[986:986] } <= { data_i[26:26] };
    end 
    if(N4236) begin
      { mem[985:985] } <= { data_i[25:25] };
    end 
    if(N4235) begin
      { mem[984:984] } <= { data_i[24:24] };
    end 
    if(N4234) begin
      { mem[983:983] } <= { data_i[23:23] };
    end 
    if(N4233) begin
      { mem[982:982] } <= { data_i[22:22] };
    end 
    if(N4232) begin
      { mem[981:981] } <= { data_i[21:21] };
    end 
    if(N4231) begin
      { mem[980:980] } <= { data_i[20:20] };
    end 
    if(N4230) begin
      { mem[979:979] } <= { data_i[19:19] };
    end 
    if(N4229) begin
      { mem[978:978] } <= { data_i[18:18] };
    end 
    if(N4228) begin
      { mem[977:977] } <= { data_i[17:17] };
    end 
    if(N4227) begin
      { mem[976:976] } <= { data_i[16:16] };
    end 
    if(N4226) begin
      { mem[975:975] } <= { data_i[15:15] };
    end 
    if(N4225) begin
      { mem[974:974] } <= { data_i[14:14] };
    end 
    if(N4224) begin
      { mem[973:973] } <= { data_i[13:13] };
    end 
    if(N4223) begin
      { mem[972:972] } <= { data_i[12:12] };
    end 
    if(N4222) begin
      { mem[971:971] } <= { data_i[11:11] };
    end 
    if(N4221) begin
      { mem[970:970] } <= { data_i[10:10] };
    end 
    if(N4220) begin
      { mem[969:969] } <= { data_i[9:9] };
    end 
    if(N4219) begin
      { mem[968:968] } <= { data_i[8:8] };
    end 
    if(N4218) begin
      { mem[967:967] } <= { data_i[7:7] };
    end 
    if(N4217) begin
      { mem[966:966] } <= { data_i[6:6] };
    end 
    if(N4216) begin
      { mem[965:965] } <= { data_i[5:5] };
    end 
    if(N4215) begin
      { mem[964:964] } <= { data_i[4:4] };
    end 
    if(N4214) begin
      { mem[963:963] } <= { data_i[3:3] };
    end 
    if(N4213) begin
      { mem[962:962] } <= { data_i[2:2] };
    end 
    if(N4212) begin
      { mem[961:961] } <= { data_i[1:1] };
    end 
    if(N4211) begin
      { mem[960:960] } <= { data_i[0:0] };
    end 
    if(N4210) begin
      { mem[959:959] } <= { data_i[39:39] };
    end 
    if(N4209) begin
      { mem[958:958] } <= { data_i[38:38] };
    end 
    if(N4208) begin
      { mem[957:957] } <= { data_i[37:37] };
    end 
    if(N4207) begin
      { mem[956:956] } <= { data_i[36:36] };
    end 
    if(N4206) begin
      { mem[955:955] } <= { data_i[35:35] };
    end 
    if(N4205) begin
      { mem[954:954] } <= { data_i[34:34] };
    end 
    if(N4204) begin
      { mem[953:953] } <= { data_i[33:33] };
    end 
    if(N4203) begin
      { mem[952:952] } <= { data_i[32:32] };
    end 
    if(N4202) begin
      { mem[951:951] } <= { data_i[31:31] };
    end 
    if(N4201) begin
      { mem[950:950] } <= { data_i[30:30] };
    end 
    if(N4200) begin
      { mem[949:949] } <= { data_i[29:29] };
    end 
    if(N4199) begin
      { mem[948:948] } <= { data_i[28:28] };
    end 
    if(N4198) begin
      { mem[947:947] } <= { data_i[27:27] };
    end 
    if(N4197) begin
      { mem[946:946] } <= { data_i[26:26] };
    end 
    if(N4196) begin
      { mem[945:945] } <= { data_i[25:25] };
    end 
    if(N4195) begin
      { mem[944:944] } <= { data_i[24:24] };
    end 
    if(N4194) begin
      { mem[943:943] } <= { data_i[23:23] };
    end 
    if(N4193) begin
      { mem[942:942] } <= { data_i[22:22] };
    end 
    if(N4192) begin
      { mem[941:941] } <= { data_i[21:21] };
    end 
    if(N4191) begin
      { mem[940:940] } <= { data_i[20:20] };
    end 
    if(N4190) begin
      { mem[939:939] } <= { data_i[19:19] };
    end 
    if(N4189) begin
      { mem[938:938] } <= { data_i[18:18] };
    end 
    if(N4188) begin
      { mem[937:937] } <= { data_i[17:17] };
    end 
    if(N4187) begin
      { mem[936:936] } <= { data_i[16:16] };
    end 
    if(N4186) begin
      { mem[935:935] } <= { data_i[15:15] };
    end 
    if(N4185) begin
      { mem[934:934] } <= { data_i[14:14] };
    end 
    if(N4184) begin
      { mem[933:933] } <= { data_i[13:13] };
    end 
    if(N4183) begin
      { mem[932:932] } <= { data_i[12:12] };
    end 
    if(N4182) begin
      { mem[931:931] } <= { data_i[11:11] };
    end 
    if(N4181) begin
      { mem[930:930] } <= { data_i[10:10] };
    end 
    if(N4180) begin
      { mem[929:929] } <= { data_i[9:9] };
    end 
    if(N4179) begin
      { mem[928:928] } <= { data_i[8:8] };
    end 
    if(N4178) begin
      { mem[927:927] } <= { data_i[7:7] };
    end 
    if(N4177) begin
      { mem[926:926] } <= { data_i[6:6] };
    end 
    if(N4176) begin
      { mem[925:925] } <= { data_i[5:5] };
    end 
    if(N4175) begin
      { mem[924:924] } <= { data_i[4:4] };
    end 
    if(N4174) begin
      { mem[923:923] } <= { data_i[3:3] };
    end 
    if(N4173) begin
      { mem[922:922] } <= { data_i[2:2] };
    end 
    if(N4172) begin
      { mem[921:921] } <= { data_i[1:1] };
    end 
    if(N4171) begin
      { mem[920:920] } <= { data_i[0:0] };
    end 
    if(N4170) begin
      { mem[919:919] } <= { data_i[39:39] };
    end 
    if(N4169) begin
      { mem[918:918] } <= { data_i[38:38] };
    end 
    if(N4168) begin
      { mem[917:917] } <= { data_i[37:37] };
    end 
    if(N4167) begin
      { mem[916:916] } <= { data_i[36:36] };
    end 
    if(N4166) begin
      { mem[915:915] } <= { data_i[35:35] };
    end 
    if(N4165) begin
      { mem[914:914] } <= { data_i[34:34] };
    end 
    if(N4164) begin
      { mem[913:913] } <= { data_i[33:33] };
    end 
    if(N4163) begin
      { mem[912:912] } <= { data_i[32:32] };
    end 
    if(N4162) begin
      { mem[911:911] } <= { data_i[31:31] };
    end 
    if(N4161) begin
      { mem[910:910] } <= { data_i[30:30] };
    end 
    if(N4160) begin
      { mem[909:909] } <= { data_i[29:29] };
    end 
    if(N4159) begin
      { mem[908:908] } <= { data_i[28:28] };
    end 
    if(N4158) begin
      { mem[907:907] } <= { data_i[27:27] };
    end 
    if(N4157) begin
      { mem[906:906] } <= { data_i[26:26] };
    end 
    if(N4156) begin
      { mem[905:905] } <= { data_i[25:25] };
    end 
    if(N4155) begin
      { mem[904:904] } <= { data_i[24:24] };
    end 
    if(N4154) begin
      { mem[903:903] } <= { data_i[23:23] };
    end 
    if(N4153) begin
      { mem[902:902] } <= { data_i[22:22] };
    end 
    if(N4152) begin
      { mem[901:901] } <= { data_i[21:21] };
    end 
    if(N4151) begin
      { mem[900:900] } <= { data_i[20:20] };
    end 
    if(N4150) begin
      { mem[899:899] } <= { data_i[19:19] };
    end 
    if(N4149) begin
      { mem[898:898] } <= { data_i[18:18] };
    end 
    if(N4148) begin
      { mem[897:897] } <= { data_i[17:17] };
    end 
    if(N4147) begin
      { mem[896:896] } <= { data_i[16:16] };
    end 
    if(N4146) begin
      { mem[895:895] } <= { data_i[15:15] };
    end 
    if(N4145) begin
      { mem[894:894] } <= { data_i[14:14] };
    end 
    if(N4144) begin
      { mem[893:893] } <= { data_i[13:13] };
    end 
    if(N4143) begin
      { mem[892:892] } <= { data_i[12:12] };
    end 
    if(N4142) begin
      { mem[891:891] } <= { data_i[11:11] };
    end 
    if(N4141) begin
      { mem[890:890] } <= { data_i[10:10] };
    end 
    if(N4140) begin
      { mem[889:889] } <= { data_i[9:9] };
    end 
    if(N4139) begin
      { mem[888:888] } <= { data_i[8:8] };
    end 
    if(N4138) begin
      { mem[887:887] } <= { data_i[7:7] };
    end 
    if(N4137) begin
      { mem[886:886] } <= { data_i[6:6] };
    end 
    if(N4136) begin
      { mem[885:885] } <= { data_i[5:5] };
    end 
    if(N4135) begin
      { mem[884:884] } <= { data_i[4:4] };
    end 
    if(N4134) begin
      { mem[883:883] } <= { data_i[3:3] };
    end 
    if(N4133) begin
      { mem[882:882] } <= { data_i[2:2] };
    end 
    if(N4132) begin
      { mem[881:881] } <= { data_i[1:1] };
    end 
    if(N4131) begin
      { mem[880:880] } <= { data_i[0:0] };
    end 
    if(N4130) begin
      { mem[879:879] } <= { data_i[39:39] };
    end 
    if(N4129) begin
      { mem[878:878] } <= { data_i[38:38] };
    end 
    if(N4128) begin
      { mem[877:877] } <= { data_i[37:37] };
    end 
    if(N4127) begin
      { mem[876:876] } <= { data_i[36:36] };
    end 
    if(N4126) begin
      { mem[875:875] } <= { data_i[35:35] };
    end 
    if(N4125) begin
      { mem[874:874] } <= { data_i[34:34] };
    end 
    if(N4124) begin
      { mem[873:873] } <= { data_i[33:33] };
    end 
    if(N4123) begin
      { mem[872:872] } <= { data_i[32:32] };
    end 
    if(N4122) begin
      { mem[871:871] } <= { data_i[31:31] };
    end 
    if(N4121) begin
      { mem[870:870] } <= { data_i[30:30] };
    end 
    if(N4120) begin
      { mem[869:869] } <= { data_i[29:29] };
    end 
    if(N4119) begin
      { mem[868:868] } <= { data_i[28:28] };
    end 
    if(N4118) begin
      { mem[867:867] } <= { data_i[27:27] };
    end 
    if(N4117) begin
      { mem[866:866] } <= { data_i[26:26] };
    end 
    if(N4116) begin
      { mem[865:865] } <= { data_i[25:25] };
    end 
    if(N4115) begin
      { mem[864:864] } <= { data_i[24:24] };
    end 
    if(N4114) begin
      { mem[863:863] } <= { data_i[23:23] };
    end 
    if(N4113) begin
      { mem[862:862] } <= { data_i[22:22] };
    end 
    if(N4112) begin
      { mem[861:861] } <= { data_i[21:21] };
    end 
    if(N4111) begin
      { mem[860:860] } <= { data_i[20:20] };
    end 
    if(N4110) begin
      { mem[859:859] } <= { data_i[19:19] };
    end 
    if(N4109) begin
      { mem[858:858] } <= { data_i[18:18] };
    end 
    if(N4108) begin
      { mem[857:857] } <= { data_i[17:17] };
    end 
    if(N4107) begin
      { mem[856:856] } <= { data_i[16:16] };
    end 
    if(N4106) begin
      { mem[855:855] } <= { data_i[15:15] };
    end 
    if(N4105) begin
      { mem[854:854] } <= { data_i[14:14] };
    end 
    if(N4104) begin
      { mem[853:853] } <= { data_i[13:13] };
    end 
    if(N4103) begin
      { mem[852:852] } <= { data_i[12:12] };
    end 
    if(N4102) begin
      { mem[851:851] } <= { data_i[11:11] };
    end 
    if(N4101) begin
      { mem[850:850] } <= { data_i[10:10] };
    end 
    if(N4100) begin
      { mem[849:849] } <= { data_i[9:9] };
    end 
    if(N4099) begin
      { mem[848:848] } <= { data_i[8:8] };
    end 
    if(N4098) begin
      { mem[847:847] } <= { data_i[7:7] };
    end 
    if(N4097) begin
      { mem[846:846] } <= { data_i[6:6] };
    end 
    if(N4096) begin
      { mem[845:845] } <= { data_i[5:5] };
    end 
    if(N4095) begin
      { mem[844:844] } <= { data_i[4:4] };
    end 
    if(N4094) begin
      { mem[843:843] } <= { data_i[3:3] };
    end 
    if(N4093) begin
      { mem[842:842] } <= { data_i[2:2] };
    end 
    if(N4092) begin
      { mem[841:841] } <= { data_i[1:1] };
    end 
    if(N4091) begin
      { mem[840:840] } <= { data_i[0:0] };
    end 
    if(N4090) begin
      { mem[839:839] } <= { data_i[39:39] };
    end 
    if(N4089) begin
      { mem[838:838] } <= { data_i[38:38] };
    end 
    if(N4088) begin
      { mem[837:837] } <= { data_i[37:37] };
    end 
    if(N4087) begin
      { mem[836:836] } <= { data_i[36:36] };
    end 
    if(N4086) begin
      { mem[835:835] } <= { data_i[35:35] };
    end 
    if(N4085) begin
      { mem[834:834] } <= { data_i[34:34] };
    end 
    if(N4084) begin
      { mem[833:833] } <= { data_i[33:33] };
    end 
    if(N4083) begin
      { mem[832:832] } <= { data_i[32:32] };
    end 
    if(N4082) begin
      { mem[831:831] } <= { data_i[31:31] };
    end 
    if(N4081) begin
      { mem[830:830] } <= { data_i[30:30] };
    end 
    if(N4080) begin
      { mem[829:829] } <= { data_i[29:29] };
    end 
    if(N4079) begin
      { mem[828:828] } <= { data_i[28:28] };
    end 
    if(N4078) begin
      { mem[827:827] } <= { data_i[27:27] };
    end 
    if(N4077) begin
      { mem[826:826] } <= { data_i[26:26] };
    end 
    if(N4076) begin
      { mem[825:825] } <= { data_i[25:25] };
    end 
    if(N4075) begin
      { mem[824:824] } <= { data_i[24:24] };
    end 
    if(N4074) begin
      { mem[823:823] } <= { data_i[23:23] };
    end 
    if(N4073) begin
      { mem[822:822] } <= { data_i[22:22] };
    end 
    if(N4072) begin
      { mem[821:821] } <= { data_i[21:21] };
    end 
    if(N4071) begin
      { mem[820:820] } <= { data_i[20:20] };
    end 
    if(N4070) begin
      { mem[819:819] } <= { data_i[19:19] };
    end 
    if(N4069) begin
      { mem[818:818] } <= { data_i[18:18] };
    end 
    if(N4068) begin
      { mem[817:817] } <= { data_i[17:17] };
    end 
    if(N4067) begin
      { mem[816:816] } <= { data_i[16:16] };
    end 
    if(N4066) begin
      { mem[815:815] } <= { data_i[15:15] };
    end 
    if(N4065) begin
      { mem[814:814] } <= { data_i[14:14] };
    end 
    if(N4064) begin
      { mem[813:813] } <= { data_i[13:13] };
    end 
    if(N4063) begin
      { mem[812:812] } <= { data_i[12:12] };
    end 
    if(N4062) begin
      { mem[811:811] } <= { data_i[11:11] };
    end 
    if(N4061) begin
      { mem[810:810] } <= { data_i[10:10] };
    end 
    if(N4060) begin
      { mem[809:809] } <= { data_i[9:9] };
    end 
    if(N4059) begin
      { mem[808:808] } <= { data_i[8:8] };
    end 
    if(N4058) begin
      { mem[807:807] } <= { data_i[7:7] };
    end 
    if(N4057) begin
      { mem[806:806] } <= { data_i[6:6] };
    end 
    if(N4056) begin
      { mem[805:805] } <= { data_i[5:5] };
    end 
    if(N4055) begin
      { mem[804:804] } <= { data_i[4:4] };
    end 
    if(N4054) begin
      { mem[803:803] } <= { data_i[3:3] };
    end 
    if(N4053) begin
      { mem[802:802] } <= { data_i[2:2] };
    end 
    if(N4052) begin
      { mem[801:801] } <= { data_i[1:1] };
    end 
    if(N4051) begin
      { mem[800:800] } <= { data_i[0:0] };
    end 
    if(N4050) begin
      { mem[799:799] } <= { data_i[39:39] };
    end 
    if(N4049) begin
      { mem[798:798] } <= { data_i[38:38] };
    end 
    if(N4048) begin
      { mem[797:797] } <= { data_i[37:37] };
    end 
    if(N4047) begin
      { mem[796:796] } <= { data_i[36:36] };
    end 
    if(N4046) begin
      { mem[795:795] } <= { data_i[35:35] };
    end 
    if(N4045) begin
      { mem[794:794] } <= { data_i[34:34] };
    end 
    if(N4044) begin
      { mem[793:793] } <= { data_i[33:33] };
    end 
    if(N4043) begin
      { mem[792:792] } <= { data_i[32:32] };
    end 
    if(N4042) begin
      { mem[791:791] } <= { data_i[31:31] };
    end 
    if(N4041) begin
      { mem[790:790] } <= { data_i[30:30] };
    end 
    if(N4040) begin
      { mem[789:789] } <= { data_i[29:29] };
    end 
    if(N4039) begin
      { mem[788:788] } <= { data_i[28:28] };
    end 
    if(N4038) begin
      { mem[787:787] } <= { data_i[27:27] };
    end 
    if(N4037) begin
      { mem[786:786] } <= { data_i[26:26] };
    end 
    if(N4036) begin
      { mem[785:785] } <= { data_i[25:25] };
    end 
    if(N4035) begin
      { mem[784:784] } <= { data_i[24:24] };
    end 
    if(N4034) begin
      { mem[783:783] } <= { data_i[23:23] };
    end 
    if(N4033) begin
      { mem[782:782] } <= { data_i[22:22] };
    end 
    if(N4032) begin
      { mem[781:781] } <= { data_i[21:21] };
    end 
    if(N4031) begin
      { mem[780:780] } <= { data_i[20:20] };
    end 
    if(N4030) begin
      { mem[779:779] } <= { data_i[19:19] };
    end 
    if(N4029) begin
      { mem[778:778] } <= { data_i[18:18] };
    end 
    if(N4028) begin
      { mem[777:777] } <= { data_i[17:17] };
    end 
    if(N4027) begin
      { mem[776:776] } <= { data_i[16:16] };
    end 
    if(N4026) begin
      { mem[775:775] } <= { data_i[15:15] };
    end 
    if(N4025) begin
      { mem[774:774] } <= { data_i[14:14] };
    end 
    if(N4024) begin
      { mem[773:773] } <= { data_i[13:13] };
    end 
    if(N4023) begin
      { mem[772:772] } <= { data_i[12:12] };
    end 
    if(N4022) begin
      { mem[771:771] } <= { data_i[11:11] };
    end 
    if(N4021) begin
      { mem[770:770] } <= { data_i[10:10] };
    end 
    if(N4020) begin
      { mem[769:769] } <= { data_i[9:9] };
    end 
    if(N4019) begin
      { mem[768:768] } <= { data_i[8:8] };
    end 
    if(N4018) begin
      { mem[767:767] } <= { data_i[7:7] };
    end 
    if(N4017) begin
      { mem[766:766] } <= { data_i[6:6] };
    end 
    if(N4016) begin
      { mem[765:765] } <= { data_i[5:5] };
    end 
    if(N4015) begin
      { mem[764:764] } <= { data_i[4:4] };
    end 
    if(N4014) begin
      { mem[763:763] } <= { data_i[3:3] };
    end 
    if(N4013) begin
      { mem[762:762] } <= { data_i[2:2] };
    end 
    if(N4012) begin
      { mem[761:761] } <= { data_i[1:1] };
    end 
    if(N4011) begin
      { mem[760:760] } <= { data_i[0:0] };
    end 
    if(N4010) begin
      { mem[759:759] } <= { data_i[39:39] };
    end 
    if(N4009) begin
      { mem[758:758] } <= { data_i[38:38] };
    end 
    if(N4008) begin
      { mem[757:757] } <= { data_i[37:37] };
    end 
    if(N4007) begin
      { mem[756:756] } <= { data_i[36:36] };
    end 
    if(N4006) begin
      { mem[755:755] } <= { data_i[35:35] };
    end 
    if(N4005) begin
      { mem[754:754] } <= { data_i[34:34] };
    end 
    if(N4004) begin
      { mem[753:753] } <= { data_i[33:33] };
    end 
    if(N4003) begin
      { mem[752:752] } <= { data_i[32:32] };
    end 
    if(N4002) begin
      { mem[751:751] } <= { data_i[31:31] };
    end 
    if(N4001) begin
      { mem[750:750] } <= { data_i[30:30] };
    end 
    if(N4000) begin
      { mem[749:749] } <= { data_i[29:29] };
    end 
    if(N3999) begin
      { mem[748:748] } <= { data_i[28:28] };
    end 
    if(N3998) begin
      { mem[747:747] } <= { data_i[27:27] };
    end 
    if(N3997) begin
      { mem[746:746] } <= { data_i[26:26] };
    end 
    if(N3996) begin
      { mem[745:745] } <= { data_i[25:25] };
    end 
    if(N3995) begin
      { mem[744:744] } <= { data_i[24:24] };
    end 
    if(N3994) begin
      { mem[743:743] } <= { data_i[23:23] };
    end 
    if(N3993) begin
      { mem[742:742] } <= { data_i[22:22] };
    end 
    if(N3992) begin
      { mem[741:741] } <= { data_i[21:21] };
    end 
    if(N3991) begin
      { mem[740:740] } <= { data_i[20:20] };
    end 
    if(N3990) begin
      { mem[739:739] } <= { data_i[19:19] };
    end 
    if(N3989) begin
      { mem[738:738] } <= { data_i[18:18] };
    end 
    if(N3988) begin
      { mem[737:737] } <= { data_i[17:17] };
    end 
    if(N3987) begin
      { mem[736:736] } <= { data_i[16:16] };
    end 
    if(N3986) begin
      { mem[735:735] } <= { data_i[15:15] };
    end 
    if(N3985) begin
      { mem[734:734] } <= { data_i[14:14] };
    end 
    if(N3984) begin
      { mem[733:733] } <= { data_i[13:13] };
    end 
    if(N3983) begin
      { mem[732:732] } <= { data_i[12:12] };
    end 
    if(N3982) begin
      { mem[731:731] } <= { data_i[11:11] };
    end 
    if(N3981) begin
      { mem[730:730] } <= { data_i[10:10] };
    end 
    if(N3980) begin
      { mem[729:729] } <= { data_i[9:9] };
    end 
    if(N3979) begin
      { mem[728:728] } <= { data_i[8:8] };
    end 
    if(N3978) begin
      { mem[727:727] } <= { data_i[7:7] };
    end 
    if(N3977) begin
      { mem[726:726] } <= { data_i[6:6] };
    end 
    if(N3976) begin
      { mem[725:725] } <= { data_i[5:5] };
    end 
    if(N3975) begin
      { mem[724:724] } <= { data_i[4:4] };
    end 
    if(N3974) begin
      { mem[723:723] } <= { data_i[3:3] };
    end 
    if(N3973) begin
      { mem[722:722] } <= { data_i[2:2] };
    end 
    if(N3972) begin
      { mem[721:721] } <= { data_i[1:1] };
    end 
    if(N3971) begin
      { mem[720:720] } <= { data_i[0:0] };
    end 
    if(N3970) begin
      { mem[719:719] } <= { data_i[39:39] };
    end 
    if(N3969) begin
      { mem[718:718] } <= { data_i[38:38] };
    end 
    if(N3968) begin
      { mem[717:717] } <= { data_i[37:37] };
    end 
    if(N3967) begin
      { mem[716:716] } <= { data_i[36:36] };
    end 
    if(N3966) begin
      { mem[715:715] } <= { data_i[35:35] };
    end 
    if(N3965) begin
      { mem[714:714] } <= { data_i[34:34] };
    end 
    if(N3964) begin
      { mem[713:713] } <= { data_i[33:33] };
    end 
    if(N3963) begin
      { mem[712:712] } <= { data_i[32:32] };
    end 
    if(N3962) begin
      { mem[711:711] } <= { data_i[31:31] };
    end 
    if(N3961) begin
      { mem[710:710] } <= { data_i[30:30] };
    end 
    if(N3960) begin
      { mem[709:709] } <= { data_i[29:29] };
    end 
    if(N3959) begin
      { mem[708:708] } <= { data_i[28:28] };
    end 
    if(N3958) begin
      { mem[707:707] } <= { data_i[27:27] };
    end 
    if(N3957) begin
      { mem[706:706] } <= { data_i[26:26] };
    end 
    if(N3956) begin
      { mem[705:705] } <= { data_i[25:25] };
    end 
    if(N3955) begin
      { mem[704:704] } <= { data_i[24:24] };
    end 
    if(N3954) begin
      { mem[703:703] } <= { data_i[23:23] };
    end 
    if(N3953) begin
      { mem[702:702] } <= { data_i[22:22] };
    end 
    if(N3952) begin
      { mem[701:701] } <= { data_i[21:21] };
    end 
    if(N3951) begin
      { mem[700:700] } <= { data_i[20:20] };
    end 
    if(N3950) begin
      { mem[699:699] } <= { data_i[19:19] };
    end 
    if(N3949) begin
      { mem[698:698] } <= { data_i[18:18] };
    end 
    if(N3948) begin
      { mem[697:697] } <= { data_i[17:17] };
    end 
    if(N3947) begin
      { mem[696:696] } <= { data_i[16:16] };
    end 
    if(N3946) begin
      { mem[695:695] } <= { data_i[15:15] };
    end 
    if(N3945) begin
      { mem[694:694] } <= { data_i[14:14] };
    end 
    if(N3944) begin
      { mem[693:693] } <= { data_i[13:13] };
    end 
    if(N3943) begin
      { mem[692:692] } <= { data_i[12:12] };
    end 
    if(N3942) begin
      { mem[691:691] } <= { data_i[11:11] };
    end 
    if(N3941) begin
      { mem[690:690] } <= { data_i[10:10] };
    end 
    if(N3940) begin
      { mem[689:689] } <= { data_i[9:9] };
    end 
    if(N3939) begin
      { mem[688:688] } <= { data_i[8:8] };
    end 
    if(N3938) begin
      { mem[687:687] } <= { data_i[7:7] };
    end 
    if(N3937) begin
      { mem[686:686] } <= { data_i[6:6] };
    end 
    if(N3936) begin
      { mem[685:685] } <= { data_i[5:5] };
    end 
    if(N3935) begin
      { mem[684:684] } <= { data_i[4:4] };
    end 
    if(N3934) begin
      { mem[683:683] } <= { data_i[3:3] };
    end 
    if(N3933) begin
      { mem[682:682] } <= { data_i[2:2] };
    end 
    if(N3932) begin
      { mem[681:681] } <= { data_i[1:1] };
    end 
    if(N3931) begin
      { mem[680:680] } <= { data_i[0:0] };
    end 
    if(N3930) begin
      { mem[679:679] } <= { data_i[39:39] };
    end 
    if(N3929) begin
      { mem[678:678] } <= { data_i[38:38] };
    end 
    if(N3928) begin
      { mem[677:677] } <= { data_i[37:37] };
    end 
    if(N3927) begin
      { mem[676:676] } <= { data_i[36:36] };
    end 
    if(N3926) begin
      { mem[675:675] } <= { data_i[35:35] };
    end 
    if(N3925) begin
      { mem[674:674] } <= { data_i[34:34] };
    end 
    if(N3924) begin
      { mem[673:673] } <= { data_i[33:33] };
    end 
    if(N3923) begin
      { mem[672:672] } <= { data_i[32:32] };
    end 
    if(N3922) begin
      { mem[671:671] } <= { data_i[31:31] };
    end 
    if(N3921) begin
      { mem[670:670] } <= { data_i[30:30] };
    end 
    if(N3920) begin
      { mem[669:669] } <= { data_i[29:29] };
    end 
    if(N3919) begin
      { mem[668:668] } <= { data_i[28:28] };
    end 
    if(N3918) begin
      { mem[667:667] } <= { data_i[27:27] };
    end 
    if(N3917) begin
      { mem[666:666] } <= { data_i[26:26] };
    end 
    if(N3916) begin
      { mem[665:665] } <= { data_i[25:25] };
    end 
    if(N3915) begin
      { mem[664:664] } <= { data_i[24:24] };
    end 
    if(N3914) begin
      { mem[663:663] } <= { data_i[23:23] };
    end 
    if(N3913) begin
      { mem[662:662] } <= { data_i[22:22] };
    end 
    if(N3912) begin
      { mem[661:661] } <= { data_i[21:21] };
    end 
    if(N3911) begin
      { mem[660:660] } <= { data_i[20:20] };
    end 
    if(N3910) begin
      { mem[659:659] } <= { data_i[19:19] };
    end 
    if(N3909) begin
      { mem[658:658] } <= { data_i[18:18] };
    end 
    if(N3908) begin
      { mem[657:657] } <= { data_i[17:17] };
    end 
    if(N3907) begin
      { mem[656:656] } <= { data_i[16:16] };
    end 
    if(N3906) begin
      { mem[655:655] } <= { data_i[15:15] };
    end 
    if(N3905) begin
      { mem[654:654] } <= { data_i[14:14] };
    end 
    if(N3904) begin
      { mem[653:653] } <= { data_i[13:13] };
    end 
    if(N3903) begin
      { mem[652:652] } <= { data_i[12:12] };
    end 
    if(N3902) begin
      { mem[651:651] } <= { data_i[11:11] };
    end 
    if(N3901) begin
      { mem[650:650] } <= { data_i[10:10] };
    end 
    if(N3900) begin
      { mem[649:649] } <= { data_i[9:9] };
    end 
    if(N3899) begin
      { mem[648:648] } <= { data_i[8:8] };
    end 
    if(N3898) begin
      { mem[647:647] } <= { data_i[7:7] };
    end 
    if(N3897) begin
      { mem[646:646] } <= { data_i[6:6] };
    end 
    if(N3896) begin
      { mem[645:645] } <= { data_i[5:5] };
    end 
    if(N3895) begin
      { mem[644:644] } <= { data_i[4:4] };
    end 
    if(N3894) begin
      { mem[643:643] } <= { data_i[3:3] };
    end 
    if(N3893) begin
      { mem[642:642] } <= { data_i[2:2] };
    end 
    if(N3892) begin
      { mem[641:641] } <= { data_i[1:1] };
    end 
    if(N3891) begin
      { mem[640:640] } <= { data_i[0:0] };
    end 
    if(N3890) begin
      { mem[639:639] } <= { data_i[39:39] };
    end 
    if(N3889) begin
      { mem[638:638] } <= { data_i[38:38] };
    end 
    if(N3888) begin
      { mem[637:637] } <= { data_i[37:37] };
    end 
    if(N3887) begin
      { mem[636:636] } <= { data_i[36:36] };
    end 
    if(N3886) begin
      { mem[635:635] } <= { data_i[35:35] };
    end 
    if(N3885) begin
      { mem[634:634] } <= { data_i[34:34] };
    end 
    if(N3884) begin
      { mem[633:633] } <= { data_i[33:33] };
    end 
    if(N3883) begin
      { mem[632:632] } <= { data_i[32:32] };
    end 
    if(N3882) begin
      { mem[631:631] } <= { data_i[31:31] };
    end 
    if(N3881) begin
      { mem[630:630] } <= { data_i[30:30] };
    end 
    if(N3880) begin
      { mem[629:629] } <= { data_i[29:29] };
    end 
    if(N3879) begin
      { mem[628:628] } <= { data_i[28:28] };
    end 
    if(N3878) begin
      { mem[627:627] } <= { data_i[27:27] };
    end 
    if(N3877) begin
      { mem[626:626] } <= { data_i[26:26] };
    end 
    if(N3876) begin
      { mem[625:625] } <= { data_i[25:25] };
    end 
    if(N3875) begin
      { mem[624:624] } <= { data_i[24:24] };
    end 
    if(N3874) begin
      { mem[623:623] } <= { data_i[23:23] };
    end 
    if(N3873) begin
      { mem[622:622] } <= { data_i[22:22] };
    end 
    if(N3872) begin
      { mem[621:621] } <= { data_i[21:21] };
    end 
    if(N3871) begin
      { mem[620:620] } <= { data_i[20:20] };
    end 
    if(N3870) begin
      { mem[619:619] } <= { data_i[19:19] };
    end 
    if(N3869) begin
      { mem[618:618] } <= { data_i[18:18] };
    end 
    if(N3868) begin
      { mem[617:617] } <= { data_i[17:17] };
    end 
    if(N3867) begin
      { mem[616:616] } <= { data_i[16:16] };
    end 
    if(N3866) begin
      { mem[615:615] } <= { data_i[15:15] };
    end 
    if(N3865) begin
      { mem[614:614] } <= { data_i[14:14] };
    end 
    if(N3864) begin
      { mem[613:613] } <= { data_i[13:13] };
    end 
    if(N3863) begin
      { mem[612:612] } <= { data_i[12:12] };
    end 
    if(N3862) begin
      { mem[611:611] } <= { data_i[11:11] };
    end 
    if(N3861) begin
      { mem[610:610] } <= { data_i[10:10] };
    end 
    if(N3860) begin
      { mem[609:609] } <= { data_i[9:9] };
    end 
    if(N3859) begin
      { mem[608:608] } <= { data_i[8:8] };
    end 
    if(N3858) begin
      { mem[607:607] } <= { data_i[7:7] };
    end 
    if(N3857) begin
      { mem[606:606] } <= { data_i[6:6] };
    end 
    if(N3856) begin
      { mem[605:605] } <= { data_i[5:5] };
    end 
    if(N3855) begin
      { mem[604:604] } <= { data_i[4:4] };
    end 
    if(N3854) begin
      { mem[603:603] } <= { data_i[3:3] };
    end 
    if(N3853) begin
      { mem[602:602] } <= { data_i[2:2] };
    end 
    if(N3852) begin
      { mem[601:601] } <= { data_i[1:1] };
    end 
    if(N3851) begin
      { mem[600:600] } <= { data_i[0:0] };
    end 
    if(N3850) begin
      { mem[599:599] } <= { data_i[39:39] };
    end 
    if(N3849) begin
      { mem[598:598] } <= { data_i[38:38] };
    end 
    if(N3848) begin
      { mem[597:597] } <= { data_i[37:37] };
    end 
    if(N3847) begin
      { mem[596:596] } <= { data_i[36:36] };
    end 
    if(N3846) begin
      { mem[595:595] } <= { data_i[35:35] };
    end 
    if(N3845) begin
      { mem[594:594] } <= { data_i[34:34] };
    end 
    if(N3844) begin
      { mem[593:593] } <= { data_i[33:33] };
    end 
    if(N3843) begin
      { mem[592:592] } <= { data_i[32:32] };
    end 
    if(N3842) begin
      { mem[591:591] } <= { data_i[31:31] };
    end 
    if(N3841) begin
      { mem[590:590] } <= { data_i[30:30] };
    end 
    if(N3840) begin
      { mem[589:589] } <= { data_i[29:29] };
    end 
    if(N3839) begin
      { mem[588:588] } <= { data_i[28:28] };
    end 
    if(N3838) begin
      { mem[587:587] } <= { data_i[27:27] };
    end 
    if(N3837) begin
      { mem[586:586] } <= { data_i[26:26] };
    end 
    if(N3836) begin
      { mem[585:585] } <= { data_i[25:25] };
    end 
    if(N3835) begin
      { mem[584:584] } <= { data_i[24:24] };
    end 
    if(N3834) begin
      { mem[583:583] } <= { data_i[23:23] };
    end 
    if(N3833) begin
      { mem[582:582] } <= { data_i[22:22] };
    end 
    if(N3832) begin
      { mem[581:581] } <= { data_i[21:21] };
    end 
    if(N3831) begin
      { mem[580:580] } <= { data_i[20:20] };
    end 
    if(N3830) begin
      { mem[579:579] } <= { data_i[19:19] };
    end 
    if(N3829) begin
      { mem[578:578] } <= { data_i[18:18] };
    end 
    if(N3828) begin
      { mem[577:577] } <= { data_i[17:17] };
    end 
    if(N3827) begin
      { mem[576:576] } <= { data_i[16:16] };
    end 
    if(N3826) begin
      { mem[575:575] } <= { data_i[15:15] };
    end 
    if(N3825) begin
      { mem[574:574] } <= { data_i[14:14] };
    end 
    if(N3824) begin
      { mem[573:573] } <= { data_i[13:13] };
    end 
    if(N3823) begin
      { mem[572:572] } <= { data_i[12:12] };
    end 
    if(N3822) begin
      { mem[571:571] } <= { data_i[11:11] };
    end 
    if(N3821) begin
      { mem[570:570] } <= { data_i[10:10] };
    end 
    if(N3820) begin
      { mem[569:569] } <= { data_i[9:9] };
    end 
    if(N3819) begin
      { mem[568:568] } <= { data_i[8:8] };
    end 
    if(N3818) begin
      { mem[567:567] } <= { data_i[7:7] };
    end 
    if(N3817) begin
      { mem[566:566] } <= { data_i[6:6] };
    end 
    if(N3816) begin
      { mem[565:565] } <= { data_i[5:5] };
    end 
    if(N3815) begin
      { mem[564:564] } <= { data_i[4:4] };
    end 
    if(N3814) begin
      { mem[563:563] } <= { data_i[3:3] };
    end 
    if(N3813) begin
      { mem[562:562] } <= { data_i[2:2] };
    end 
    if(N3812) begin
      { mem[561:561] } <= { data_i[1:1] };
    end 
    if(N3811) begin
      { mem[560:560] } <= { data_i[0:0] };
    end 
    if(N3810) begin
      { mem[559:559] } <= { data_i[39:39] };
    end 
    if(N3809) begin
      { mem[558:558] } <= { data_i[38:38] };
    end 
    if(N3808) begin
      { mem[557:557] } <= { data_i[37:37] };
    end 
    if(N3807) begin
      { mem[556:556] } <= { data_i[36:36] };
    end 
    if(N3806) begin
      { mem[555:555] } <= { data_i[35:35] };
    end 
    if(N3805) begin
      { mem[554:554] } <= { data_i[34:34] };
    end 
    if(N3804) begin
      { mem[553:553] } <= { data_i[33:33] };
    end 
    if(N3803) begin
      { mem[552:552] } <= { data_i[32:32] };
    end 
    if(N3802) begin
      { mem[551:551] } <= { data_i[31:31] };
    end 
    if(N3801) begin
      { mem[550:550] } <= { data_i[30:30] };
    end 
    if(N3800) begin
      { mem[549:549] } <= { data_i[29:29] };
    end 
    if(N3799) begin
      { mem[548:548] } <= { data_i[28:28] };
    end 
    if(N3798) begin
      { mem[547:547] } <= { data_i[27:27] };
    end 
    if(N3797) begin
      { mem[546:546] } <= { data_i[26:26] };
    end 
    if(N3796) begin
      { mem[545:545] } <= { data_i[25:25] };
    end 
    if(N3795) begin
      { mem[544:544] } <= { data_i[24:24] };
    end 
    if(N3794) begin
      { mem[543:543] } <= { data_i[23:23] };
    end 
    if(N3793) begin
      { mem[542:542] } <= { data_i[22:22] };
    end 
    if(N3792) begin
      { mem[541:541] } <= { data_i[21:21] };
    end 
    if(N3791) begin
      { mem[540:540] } <= { data_i[20:20] };
    end 
    if(N3790) begin
      { mem[539:539] } <= { data_i[19:19] };
    end 
    if(N3789) begin
      { mem[538:538] } <= { data_i[18:18] };
    end 
    if(N3788) begin
      { mem[537:537] } <= { data_i[17:17] };
    end 
    if(N3787) begin
      { mem[536:536] } <= { data_i[16:16] };
    end 
    if(N3786) begin
      { mem[535:535] } <= { data_i[15:15] };
    end 
    if(N3785) begin
      { mem[534:534] } <= { data_i[14:14] };
    end 
    if(N3784) begin
      { mem[533:533] } <= { data_i[13:13] };
    end 
    if(N3783) begin
      { mem[532:532] } <= { data_i[12:12] };
    end 
    if(N3782) begin
      { mem[531:531] } <= { data_i[11:11] };
    end 
    if(N3781) begin
      { mem[530:530] } <= { data_i[10:10] };
    end 
    if(N3780) begin
      { mem[529:529] } <= { data_i[9:9] };
    end 
    if(N3779) begin
      { mem[528:528] } <= { data_i[8:8] };
    end 
    if(N3778) begin
      { mem[527:527] } <= { data_i[7:7] };
    end 
    if(N3777) begin
      { mem[526:526] } <= { data_i[6:6] };
    end 
    if(N3776) begin
      { mem[525:525] } <= { data_i[5:5] };
    end 
    if(N3775) begin
      { mem[524:524] } <= { data_i[4:4] };
    end 
    if(N3774) begin
      { mem[523:523] } <= { data_i[3:3] };
    end 
    if(N3773) begin
      { mem[522:522] } <= { data_i[2:2] };
    end 
    if(N3772) begin
      { mem[521:521] } <= { data_i[1:1] };
    end 
    if(N3771) begin
      { mem[520:520] } <= { data_i[0:0] };
    end 
    if(N3770) begin
      { mem[519:519] } <= { data_i[39:39] };
    end 
    if(N3769) begin
      { mem[518:518] } <= { data_i[38:38] };
    end 
    if(N3768) begin
      { mem[517:517] } <= { data_i[37:37] };
    end 
    if(N3767) begin
      { mem[516:516] } <= { data_i[36:36] };
    end 
    if(N3766) begin
      { mem[515:515] } <= { data_i[35:35] };
    end 
    if(N3765) begin
      { mem[514:514] } <= { data_i[34:34] };
    end 
    if(N3764) begin
      { mem[513:513] } <= { data_i[33:33] };
    end 
    if(N3763) begin
      { mem[512:512] } <= { data_i[32:32] };
    end 
    if(N3762) begin
      { mem[511:511] } <= { data_i[31:31] };
    end 
    if(N3761) begin
      { mem[510:510] } <= { data_i[30:30] };
    end 
    if(N3760) begin
      { mem[509:509] } <= { data_i[29:29] };
    end 
    if(N3759) begin
      { mem[508:508] } <= { data_i[28:28] };
    end 
    if(N3758) begin
      { mem[507:507] } <= { data_i[27:27] };
    end 
    if(N3757) begin
      { mem[506:506] } <= { data_i[26:26] };
    end 
    if(N3756) begin
      { mem[505:505] } <= { data_i[25:25] };
    end 
    if(N3755) begin
      { mem[504:504] } <= { data_i[24:24] };
    end 
    if(N3754) begin
      { mem[503:503] } <= { data_i[23:23] };
    end 
    if(N3753) begin
      { mem[502:502] } <= { data_i[22:22] };
    end 
    if(N3752) begin
      { mem[501:501] } <= { data_i[21:21] };
    end 
    if(N3751) begin
      { mem[500:500] } <= { data_i[20:20] };
    end 
    if(N3750) begin
      { mem[499:499] } <= { data_i[19:19] };
    end 
    if(N3749) begin
      { mem[498:498] } <= { data_i[18:18] };
    end 
    if(N3748) begin
      { mem[497:497] } <= { data_i[17:17] };
    end 
    if(N3747) begin
      { mem[496:496] } <= { data_i[16:16] };
    end 
    if(N3746) begin
      { mem[495:495] } <= { data_i[15:15] };
    end 
    if(N3745) begin
      { mem[494:494] } <= { data_i[14:14] };
    end 
    if(N3744) begin
      { mem[493:493] } <= { data_i[13:13] };
    end 
    if(N3743) begin
      { mem[492:492] } <= { data_i[12:12] };
    end 
    if(N3742) begin
      { mem[491:491] } <= { data_i[11:11] };
    end 
    if(N3741) begin
      { mem[490:490] } <= { data_i[10:10] };
    end 
    if(N3740) begin
      { mem[489:489] } <= { data_i[9:9] };
    end 
    if(N3739) begin
      { mem[488:488] } <= { data_i[8:8] };
    end 
    if(N3738) begin
      { mem[487:487] } <= { data_i[7:7] };
    end 
    if(N3737) begin
      { mem[486:486] } <= { data_i[6:6] };
    end 
    if(N3736) begin
      { mem[485:485] } <= { data_i[5:5] };
    end 
    if(N3735) begin
      { mem[484:484] } <= { data_i[4:4] };
    end 
    if(N3734) begin
      { mem[483:483] } <= { data_i[3:3] };
    end 
    if(N3733) begin
      { mem[482:482] } <= { data_i[2:2] };
    end 
    if(N3732) begin
      { mem[481:481] } <= { data_i[1:1] };
    end 
    if(N3731) begin
      { mem[480:480] } <= { data_i[0:0] };
    end 
    if(N3730) begin
      { mem[479:479] } <= { data_i[39:39] };
    end 
    if(N3729) begin
      { mem[478:478] } <= { data_i[38:38] };
    end 
    if(N3728) begin
      { mem[477:477] } <= { data_i[37:37] };
    end 
    if(N3727) begin
      { mem[476:476] } <= { data_i[36:36] };
    end 
    if(N3726) begin
      { mem[475:475] } <= { data_i[35:35] };
    end 
    if(N3725) begin
      { mem[474:474] } <= { data_i[34:34] };
    end 
    if(N3724) begin
      { mem[473:473] } <= { data_i[33:33] };
    end 
    if(N3723) begin
      { mem[472:472] } <= { data_i[32:32] };
    end 
    if(N3722) begin
      { mem[471:471] } <= { data_i[31:31] };
    end 
    if(N3721) begin
      { mem[470:470] } <= { data_i[30:30] };
    end 
    if(N3720) begin
      { mem[469:469] } <= { data_i[29:29] };
    end 
    if(N3719) begin
      { mem[468:468] } <= { data_i[28:28] };
    end 
    if(N3718) begin
      { mem[467:467] } <= { data_i[27:27] };
    end 
    if(N3717) begin
      { mem[466:466] } <= { data_i[26:26] };
    end 
    if(N3716) begin
      { mem[465:465] } <= { data_i[25:25] };
    end 
    if(N3715) begin
      { mem[464:464] } <= { data_i[24:24] };
    end 
    if(N3714) begin
      { mem[463:463] } <= { data_i[23:23] };
    end 
    if(N3713) begin
      { mem[462:462] } <= { data_i[22:22] };
    end 
    if(N3712) begin
      { mem[461:461] } <= { data_i[21:21] };
    end 
    if(N3711) begin
      { mem[460:460] } <= { data_i[20:20] };
    end 
    if(N3710) begin
      { mem[459:459] } <= { data_i[19:19] };
    end 
    if(N3709) begin
      { mem[458:458] } <= { data_i[18:18] };
    end 
    if(N3708) begin
      { mem[457:457] } <= { data_i[17:17] };
    end 
    if(N3707) begin
      { mem[456:456] } <= { data_i[16:16] };
    end 
    if(N3706) begin
      { mem[455:455] } <= { data_i[15:15] };
    end 
    if(N3705) begin
      { mem[454:454] } <= { data_i[14:14] };
    end 
    if(N3704) begin
      { mem[453:453] } <= { data_i[13:13] };
    end 
    if(N3703) begin
      { mem[452:452] } <= { data_i[12:12] };
    end 
    if(N3702) begin
      { mem[451:451] } <= { data_i[11:11] };
    end 
    if(N3701) begin
      { mem[450:450] } <= { data_i[10:10] };
    end 
    if(N3700) begin
      { mem[449:449] } <= { data_i[9:9] };
    end 
    if(N3699) begin
      { mem[448:448] } <= { data_i[8:8] };
    end 
    if(N3698) begin
      { mem[447:447] } <= { data_i[7:7] };
    end 
    if(N3697) begin
      { mem[446:446] } <= { data_i[6:6] };
    end 
    if(N3696) begin
      { mem[445:445] } <= { data_i[5:5] };
    end 
    if(N3695) begin
      { mem[444:444] } <= { data_i[4:4] };
    end 
    if(N3694) begin
      { mem[443:443] } <= { data_i[3:3] };
    end 
    if(N3693) begin
      { mem[442:442] } <= { data_i[2:2] };
    end 
    if(N3692) begin
      { mem[441:441] } <= { data_i[1:1] };
    end 
    if(N3691) begin
      { mem[440:440] } <= { data_i[0:0] };
    end 
    if(N3690) begin
      { mem[439:439] } <= { data_i[39:39] };
    end 
    if(N3689) begin
      { mem[438:438] } <= { data_i[38:38] };
    end 
    if(N3688) begin
      { mem[437:437] } <= { data_i[37:37] };
    end 
    if(N3687) begin
      { mem[436:436] } <= { data_i[36:36] };
    end 
    if(N3686) begin
      { mem[435:435] } <= { data_i[35:35] };
    end 
    if(N3685) begin
      { mem[434:434] } <= { data_i[34:34] };
    end 
    if(N3684) begin
      { mem[433:433] } <= { data_i[33:33] };
    end 
    if(N3683) begin
      { mem[432:432] } <= { data_i[32:32] };
    end 
    if(N3682) begin
      { mem[431:431] } <= { data_i[31:31] };
    end 
    if(N3681) begin
      { mem[430:430] } <= { data_i[30:30] };
    end 
    if(N3680) begin
      { mem[429:429] } <= { data_i[29:29] };
    end 
    if(N3679) begin
      { mem[428:428] } <= { data_i[28:28] };
    end 
    if(N3678) begin
      { mem[427:427] } <= { data_i[27:27] };
    end 
    if(N3677) begin
      { mem[426:426] } <= { data_i[26:26] };
    end 
    if(N3676) begin
      { mem[425:425] } <= { data_i[25:25] };
    end 
    if(N3675) begin
      { mem[424:424] } <= { data_i[24:24] };
    end 
    if(N3674) begin
      { mem[423:423] } <= { data_i[23:23] };
    end 
    if(N3673) begin
      { mem[422:422] } <= { data_i[22:22] };
    end 
    if(N3672) begin
      { mem[421:421] } <= { data_i[21:21] };
    end 
    if(N3671) begin
      { mem[420:420] } <= { data_i[20:20] };
    end 
    if(N3670) begin
      { mem[419:419] } <= { data_i[19:19] };
    end 
    if(N3669) begin
      { mem[418:418] } <= { data_i[18:18] };
    end 
    if(N3668) begin
      { mem[417:417] } <= { data_i[17:17] };
    end 
    if(N3667) begin
      { mem[416:416] } <= { data_i[16:16] };
    end 
    if(N3666) begin
      { mem[415:415] } <= { data_i[15:15] };
    end 
    if(N3665) begin
      { mem[414:414] } <= { data_i[14:14] };
    end 
    if(N3664) begin
      { mem[413:413] } <= { data_i[13:13] };
    end 
    if(N3663) begin
      { mem[412:412] } <= { data_i[12:12] };
    end 
    if(N3662) begin
      { mem[411:411] } <= { data_i[11:11] };
    end 
    if(N3661) begin
      { mem[410:410] } <= { data_i[10:10] };
    end 
    if(N3660) begin
      { mem[409:409] } <= { data_i[9:9] };
    end 
    if(N3659) begin
      { mem[408:408] } <= { data_i[8:8] };
    end 
    if(N3658) begin
      { mem[407:407] } <= { data_i[7:7] };
    end 
    if(N3657) begin
      { mem[406:406] } <= { data_i[6:6] };
    end 
    if(N3656) begin
      { mem[405:405] } <= { data_i[5:5] };
    end 
    if(N3655) begin
      { mem[404:404] } <= { data_i[4:4] };
    end 
    if(N3654) begin
      { mem[403:403] } <= { data_i[3:3] };
    end 
    if(N3653) begin
      { mem[402:402] } <= { data_i[2:2] };
    end 
    if(N3652) begin
      { mem[401:401] } <= { data_i[1:1] };
    end 
    if(N3651) begin
      { mem[400:400] } <= { data_i[0:0] };
    end 
    if(N3650) begin
      { mem[399:399] } <= { data_i[39:39] };
    end 
    if(N3649) begin
      { mem[398:398] } <= { data_i[38:38] };
    end 
    if(N3648) begin
      { mem[397:397] } <= { data_i[37:37] };
    end 
    if(N3647) begin
      { mem[396:396] } <= { data_i[36:36] };
    end 
    if(N3646) begin
      { mem[395:395] } <= { data_i[35:35] };
    end 
    if(N3645) begin
      { mem[394:394] } <= { data_i[34:34] };
    end 
    if(N3644) begin
      { mem[393:393] } <= { data_i[33:33] };
    end 
    if(N3643) begin
      { mem[392:392] } <= { data_i[32:32] };
    end 
    if(N3642) begin
      { mem[391:391] } <= { data_i[31:31] };
    end 
    if(N3641) begin
      { mem[390:390] } <= { data_i[30:30] };
    end 
    if(N3640) begin
      { mem[389:389] } <= { data_i[29:29] };
    end 
    if(N3639) begin
      { mem[388:388] } <= { data_i[28:28] };
    end 
    if(N3638) begin
      { mem[387:387] } <= { data_i[27:27] };
    end 
    if(N3637) begin
      { mem[386:386] } <= { data_i[26:26] };
    end 
    if(N3636) begin
      { mem[385:385] } <= { data_i[25:25] };
    end 
    if(N3635) begin
      { mem[384:384] } <= { data_i[24:24] };
    end 
    if(N3634) begin
      { mem[383:383] } <= { data_i[23:23] };
    end 
    if(N3633) begin
      { mem[382:382] } <= { data_i[22:22] };
    end 
    if(N3632) begin
      { mem[381:381] } <= { data_i[21:21] };
    end 
    if(N3631) begin
      { mem[380:380] } <= { data_i[20:20] };
    end 
    if(N3630) begin
      { mem[379:379] } <= { data_i[19:19] };
    end 
    if(N3629) begin
      { mem[378:378] } <= { data_i[18:18] };
    end 
    if(N3628) begin
      { mem[377:377] } <= { data_i[17:17] };
    end 
    if(N3627) begin
      { mem[376:376] } <= { data_i[16:16] };
    end 
    if(N3626) begin
      { mem[375:375] } <= { data_i[15:15] };
    end 
    if(N3625) begin
      { mem[374:374] } <= { data_i[14:14] };
    end 
    if(N3624) begin
      { mem[373:373] } <= { data_i[13:13] };
    end 
    if(N3623) begin
      { mem[372:372] } <= { data_i[12:12] };
    end 
    if(N3622) begin
      { mem[371:371] } <= { data_i[11:11] };
    end 
    if(N3621) begin
      { mem[370:370] } <= { data_i[10:10] };
    end 
    if(N3620) begin
      { mem[369:369] } <= { data_i[9:9] };
    end 
    if(N3619) begin
      { mem[368:368] } <= { data_i[8:8] };
    end 
    if(N3618) begin
      { mem[367:367] } <= { data_i[7:7] };
    end 
    if(N3617) begin
      { mem[366:366] } <= { data_i[6:6] };
    end 
    if(N3616) begin
      { mem[365:365] } <= { data_i[5:5] };
    end 
    if(N3615) begin
      { mem[364:364] } <= { data_i[4:4] };
    end 
    if(N3614) begin
      { mem[363:363] } <= { data_i[3:3] };
    end 
    if(N3613) begin
      { mem[362:362] } <= { data_i[2:2] };
    end 
    if(N3612) begin
      { mem[361:361] } <= { data_i[1:1] };
    end 
    if(N3611) begin
      { mem[360:360] } <= { data_i[0:0] };
    end 
    if(N3610) begin
      { mem[359:359] } <= { data_i[39:39] };
    end 
    if(N3609) begin
      { mem[358:358] } <= { data_i[38:38] };
    end 
    if(N3608) begin
      { mem[357:357] } <= { data_i[37:37] };
    end 
    if(N3607) begin
      { mem[356:356] } <= { data_i[36:36] };
    end 
    if(N3606) begin
      { mem[355:355] } <= { data_i[35:35] };
    end 
    if(N3605) begin
      { mem[354:354] } <= { data_i[34:34] };
    end 
    if(N3604) begin
      { mem[353:353] } <= { data_i[33:33] };
    end 
    if(N3603) begin
      { mem[352:352] } <= { data_i[32:32] };
    end 
    if(N3602) begin
      { mem[351:351] } <= { data_i[31:31] };
    end 
    if(N3601) begin
      { mem[350:350] } <= { data_i[30:30] };
    end 
    if(N3600) begin
      { mem[349:349] } <= { data_i[29:29] };
    end 
    if(N3599) begin
      { mem[348:348] } <= { data_i[28:28] };
    end 
    if(N3598) begin
      { mem[347:347] } <= { data_i[27:27] };
    end 
    if(N3597) begin
      { mem[346:346] } <= { data_i[26:26] };
    end 
    if(N3596) begin
      { mem[345:345] } <= { data_i[25:25] };
    end 
    if(N3595) begin
      { mem[344:344] } <= { data_i[24:24] };
    end 
    if(N3594) begin
      { mem[343:343] } <= { data_i[23:23] };
    end 
    if(N3593) begin
      { mem[342:342] } <= { data_i[22:22] };
    end 
    if(N3592) begin
      { mem[341:341] } <= { data_i[21:21] };
    end 
    if(N3591) begin
      { mem[340:340] } <= { data_i[20:20] };
    end 
    if(N3590) begin
      { mem[339:339] } <= { data_i[19:19] };
    end 
    if(N3589) begin
      { mem[338:338] } <= { data_i[18:18] };
    end 
    if(N3588) begin
      { mem[337:337] } <= { data_i[17:17] };
    end 
    if(N3587) begin
      { mem[336:336] } <= { data_i[16:16] };
    end 
    if(N3586) begin
      { mem[335:335] } <= { data_i[15:15] };
    end 
    if(N3585) begin
      { mem[334:334] } <= { data_i[14:14] };
    end 
    if(N3584) begin
      { mem[333:333] } <= { data_i[13:13] };
    end 
    if(N3583) begin
      { mem[332:332] } <= { data_i[12:12] };
    end 
    if(N3582) begin
      { mem[331:331] } <= { data_i[11:11] };
    end 
    if(N3581) begin
      { mem[330:330] } <= { data_i[10:10] };
    end 
    if(N3580) begin
      { mem[329:329] } <= { data_i[9:9] };
    end 
    if(N3579) begin
      { mem[328:328] } <= { data_i[8:8] };
    end 
    if(N3578) begin
      { mem[327:327] } <= { data_i[7:7] };
    end 
    if(N3577) begin
      { mem[326:326] } <= { data_i[6:6] };
    end 
    if(N3576) begin
      { mem[325:325] } <= { data_i[5:5] };
    end 
    if(N3575) begin
      { mem[324:324] } <= { data_i[4:4] };
    end 
    if(N3574) begin
      { mem[323:323] } <= { data_i[3:3] };
    end 
    if(N3573) begin
      { mem[322:322] } <= { data_i[2:2] };
    end 
    if(N3572) begin
      { mem[321:321] } <= { data_i[1:1] };
    end 
    if(N3571) begin
      { mem[320:320] } <= { data_i[0:0] };
    end 
    if(N3570) begin
      { mem[319:319] } <= { data_i[39:39] };
    end 
    if(N3569) begin
      { mem[318:318] } <= { data_i[38:38] };
    end 
    if(N3568) begin
      { mem[317:317] } <= { data_i[37:37] };
    end 
    if(N3567) begin
      { mem[316:316] } <= { data_i[36:36] };
    end 
    if(N3566) begin
      { mem[315:315] } <= { data_i[35:35] };
    end 
    if(N3565) begin
      { mem[314:314] } <= { data_i[34:34] };
    end 
    if(N3564) begin
      { mem[313:313] } <= { data_i[33:33] };
    end 
    if(N3563) begin
      { mem[312:312] } <= { data_i[32:32] };
    end 
    if(N3562) begin
      { mem[311:311] } <= { data_i[31:31] };
    end 
    if(N3561) begin
      { mem[310:310] } <= { data_i[30:30] };
    end 
    if(N3560) begin
      { mem[309:309] } <= { data_i[29:29] };
    end 
    if(N3559) begin
      { mem[308:308] } <= { data_i[28:28] };
    end 
    if(N3558) begin
      { mem[307:307] } <= { data_i[27:27] };
    end 
    if(N3557) begin
      { mem[306:306] } <= { data_i[26:26] };
    end 
    if(N3556) begin
      { mem[305:305] } <= { data_i[25:25] };
    end 
    if(N3555) begin
      { mem[304:304] } <= { data_i[24:24] };
    end 
    if(N3554) begin
      { mem[303:303] } <= { data_i[23:23] };
    end 
    if(N3553) begin
      { mem[302:302] } <= { data_i[22:22] };
    end 
    if(N3552) begin
      { mem[301:301] } <= { data_i[21:21] };
    end 
    if(N3551) begin
      { mem[300:300] } <= { data_i[20:20] };
    end 
    if(N3550) begin
      { mem[299:299] } <= { data_i[19:19] };
    end 
    if(N3549) begin
      { mem[298:298] } <= { data_i[18:18] };
    end 
    if(N3548) begin
      { mem[297:297] } <= { data_i[17:17] };
    end 
    if(N3547) begin
      { mem[296:296] } <= { data_i[16:16] };
    end 
    if(N3546) begin
      { mem[295:295] } <= { data_i[15:15] };
    end 
    if(N3545) begin
      { mem[294:294] } <= { data_i[14:14] };
    end 
    if(N3544) begin
      { mem[293:293] } <= { data_i[13:13] };
    end 
    if(N3543) begin
      { mem[292:292] } <= { data_i[12:12] };
    end 
    if(N3542) begin
      { mem[291:291] } <= { data_i[11:11] };
    end 
    if(N3541) begin
      { mem[290:290] } <= { data_i[10:10] };
    end 
    if(N3540) begin
      { mem[289:289] } <= { data_i[9:9] };
    end 
    if(N3539) begin
      { mem[288:288] } <= { data_i[8:8] };
    end 
    if(N3538) begin
      { mem[287:287] } <= { data_i[7:7] };
    end 
    if(N3537) begin
      { mem[286:286] } <= { data_i[6:6] };
    end 
    if(N3536) begin
      { mem[285:285] } <= { data_i[5:5] };
    end 
    if(N3535) begin
      { mem[284:284] } <= { data_i[4:4] };
    end 
    if(N3534) begin
      { mem[283:283] } <= { data_i[3:3] };
    end 
    if(N3533) begin
      { mem[282:282] } <= { data_i[2:2] };
    end 
    if(N3532) begin
      { mem[281:281] } <= { data_i[1:1] };
    end 
    if(N3531) begin
      { mem[280:280] } <= { data_i[0:0] };
    end 
    if(N3530) begin
      { mem[279:279] } <= { data_i[39:39] };
    end 
    if(N3529) begin
      { mem[278:278] } <= { data_i[38:38] };
    end 
    if(N3528) begin
      { mem[277:277] } <= { data_i[37:37] };
    end 
    if(N3527) begin
      { mem[276:276] } <= { data_i[36:36] };
    end 
    if(N3526) begin
      { mem[275:275] } <= { data_i[35:35] };
    end 
    if(N3525) begin
      { mem[274:274] } <= { data_i[34:34] };
    end 
    if(N3524) begin
      { mem[273:273] } <= { data_i[33:33] };
    end 
    if(N3523) begin
      { mem[272:272] } <= { data_i[32:32] };
    end 
    if(N3522) begin
      { mem[271:271] } <= { data_i[31:31] };
    end 
    if(N3521) begin
      { mem[270:270] } <= { data_i[30:30] };
    end 
    if(N3520) begin
      { mem[269:269] } <= { data_i[29:29] };
    end 
    if(N3519) begin
      { mem[268:268] } <= { data_i[28:28] };
    end 
    if(N3518) begin
      { mem[267:267] } <= { data_i[27:27] };
    end 
    if(N3517) begin
      { mem[266:266] } <= { data_i[26:26] };
    end 
    if(N3516) begin
      { mem[265:265] } <= { data_i[25:25] };
    end 
    if(N3515) begin
      { mem[264:264] } <= { data_i[24:24] };
    end 
    if(N3514) begin
      { mem[263:263] } <= { data_i[23:23] };
    end 
    if(N3513) begin
      { mem[262:262] } <= { data_i[22:22] };
    end 
    if(N3512) begin
      { mem[261:261] } <= { data_i[21:21] };
    end 
    if(N3511) begin
      { mem[260:260] } <= { data_i[20:20] };
    end 
    if(N3510) begin
      { mem[259:259] } <= { data_i[19:19] };
    end 
    if(N3509) begin
      { mem[258:258] } <= { data_i[18:18] };
    end 
    if(N3508) begin
      { mem[257:257] } <= { data_i[17:17] };
    end 
    if(N3507) begin
      { mem[256:256] } <= { data_i[16:16] };
    end 
    if(N3506) begin
      { mem[255:255] } <= { data_i[15:15] };
    end 
    if(N3505) begin
      { mem[254:254] } <= { data_i[14:14] };
    end 
    if(N3504) begin
      { mem[253:253] } <= { data_i[13:13] };
    end 
    if(N3503) begin
      { mem[252:252] } <= { data_i[12:12] };
    end 
    if(N3502) begin
      { mem[251:251] } <= { data_i[11:11] };
    end 
    if(N3501) begin
      { mem[250:250] } <= { data_i[10:10] };
    end 
    if(N3500) begin
      { mem[249:249] } <= { data_i[9:9] };
    end 
    if(N3499) begin
      { mem[248:248] } <= { data_i[8:8] };
    end 
    if(N3498) begin
      { mem[247:247] } <= { data_i[7:7] };
    end 
    if(N3497) begin
      { mem[246:246] } <= { data_i[6:6] };
    end 
    if(N3496) begin
      { mem[245:245] } <= { data_i[5:5] };
    end 
    if(N3495) begin
      { mem[244:244] } <= { data_i[4:4] };
    end 
    if(N3494) begin
      { mem[243:243] } <= { data_i[3:3] };
    end 
    if(N3493) begin
      { mem[242:242] } <= { data_i[2:2] };
    end 
    if(N3492) begin
      { mem[241:241] } <= { data_i[1:1] };
    end 
    if(N3491) begin
      { mem[240:240] } <= { data_i[0:0] };
    end 
    if(N3490) begin
      { mem[239:239] } <= { data_i[39:39] };
    end 
    if(N3489) begin
      { mem[238:238] } <= { data_i[38:38] };
    end 
    if(N3488) begin
      { mem[237:237] } <= { data_i[37:37] };
    end 
    if(N3487) begin
      { mem[236:236] } <= { data_i[36:36] };
    end 
    if(N3486) begin
      { mem[235:235] } <= { data_i[35:35] };
    end 
    if(N3485) begin
      { mem[234:234] } <= { data_i[34:34] };
    end 
    if(N3484) begin
      { mem[233:233] } <= { data_i[33:33] };
    end 
    if(N3483) begin
      { mem[232:232] } <= { data_i[32:32] };
    end 
    if(N3482) begin
      { mem[231:231] } <= { data_i[31:31] };
    end 
    if(N3481) begin
      { mem[230:230] } <= { data_i[30:30] };
    end 
    if(N3480) begin
      { mem[229:229] } <= { data_i[29:29] };
    end 
    if(N3479) begin
      { mem[228:228] } <= { data_i[28:28] };
    end 
    if(N3478) begin
      { mem[227:227] } <= { data_i[27:27] };
    end 
    if(N3477) begin
      { mem[226:226] } <= { data_i[26:26] };
    end 
    if(N3476) begin
      { mem[225:225] } <= { data_i[25:25] };
    end 
    if(N3475) begin
      { mem[224:224] } <= { data_i[24:24] };
    end 
    if(N3474) begin
      { mem[223:223] } <= { data_i[23:23] };
    end 
    if(N3473) begin
      { mem[222:222] } <= { data_i[22:22] };
    end 
    if(N3472) begin
      { mem[221:221] } <= { data_i[21:21] };
    end 
    if(N3471) begin
      { mem[220:220] } <= { data_i[20:20] };
    end 
    if(N3470) begin
      { mem[219:219] } <= { data_i[19:19] };
    end 
    if(N3469) begin
      { mem[218:218] } <= { data_i[18:18] };
    end 
    if(N3468) begin
      { mem[217:217] } <= { data_i[17:17] };
    end 
    if(N3467) begin
      { mem[216:216] } <= { data_i[16:16] };
    end 
    if(N3466) begin
      { mem[215:215] } <= { data_i[15:15] };
    end 
    if(N3465) begin
      { mem[214:214] } <= { data_i[14:14] };
    end 
    if(N3464) begin
      { mem[213:213] } <= { data_i[13:13] };
    end 
    if(N3463) begin
      { mem[212:212] } <= { data_i[12:12] };
    end 
    if(N3462) begin
      { mem[211:211] } <= { data_i[11:11] };
    end 
    if(N3461) begin
      { mem[210:210] } <= { data_i[10:10] };
    end 
    if(N3460) begin
      { mem[209:209] } <= { data_i[9:9] };
    end 
    if(N3459) begin
      { mem[208:208] } <= { data_i[8:8] };
    end 
    if(N3458) begin
      { mem[207:207] } <= { data_i[7:7] };
    end 
    if(N3457) begin
      { mem[206:206] } <= { data_i[6:6] };
    end 
    if(N3456) begin
      { mem[205:205] } <= { data_i[5:5] };
    end 
    if(N3455) begin
      { mem[204:204] } <= { data_i[4:4] };
    end 
    if(N3454) begin
      { mem[203:203] } <= { data_i[3:3] };
    end 
    if(N3453) begin
      { mem[202:202] } <= { data_i[2:2] };
    end 
    if(N3452) begin
      { mem[201:201] } <= { data_i[1:1] };
    end 
    if(N3451) begin
      { mem[200:200] } <= { data_i[0:0] };
    end 
    if(N3450) begin
      { mem[199:199] } <= { data_i[39:39] };
    end 
    if(N3449) begin
      { mem[198:198] } <= { data_i[38:38] };
    end 
    if(N3448) begin
      { mem[197:197] } <= { data_i[37:37] };
    end 
    if(N3447) begin
      { mem[196:196] } <= { data_i[36:36] };
    end 
    if(N3446) begin
      { mem[195:195] } <= { data_i[35:35] };
    end 
    if(N3445) begin
      { mem[194:194] } <= { data_i[34:34] };
    end 
    if(N3444) begin
      { mem[193:193] } <= { data_i[33:33] };
    end 
    if(N3443) begin
      { mem[192:192] } <= { data_i[32:32] };
    end 
    if(N3442) begin
      { mem[191:191] } <= { data_i[31:31] };
    end 
    if(N3441) begin
      { mem[190:190] } <= { data_i[30:30] };
    end 
    if(N3440) begin
      { mem[189:189] } <= { data_i[29:29] };
    end 
    if(N3439) begin
      { mem[188:188] } <= { data_i[28:28] };
    end 
    if(N3438) begin
      { mem[187:187] } <= { data_i[27:27] };
    end 
    if(N3437) begin
      { mem[186:186] } <= { data_i[26:26] };
    end 
    if(N3436) begin
      { mem[185:185] } <= { data_i[25:25] };
    end 
    if(N3435) begin
      { mem[184:184] } <= { data_i[24:24] };
    end 
    if(N3434) begin
      { mem[183:183] } <= { data_i[23:23] };
    end 
    if(N3433) begin
      { mem[182:182] } <= { data_i[22:22] };
    end 
    if(N3432) begin
      { mem[181:181] } <= { data_i[21:21] };
    end 
    if(N3431) begin
      { mem[180:180] } <= { data_i[20:20] };
    end 
    if(N3430) begin
      { mem[179:179] } <= { data_i[19:19] };
    end 
    if(N3429) begin
      { mem[178:178] } <= { data_i[18:18] };
    end 
    if(N3428) begin
      { mem[177:177] } <= { data_i[17:17] };
    end 
    if(N3427) begin
      { mem[176:176] } <= { data_i[16:16] };
    end 
    if(N3426) begin
      { mem[175:175] } <= { data_i[15:15] };
    end 
    if(N3425) begin
      { mem[174:174] } <= { data_i[14:14] };
    end 
    if(N3424) begin
      { mem[173:173] } <= { data_i[13:13] };
    end 
    if(N3423) begin
      { mem[172:172] } <= { data_i[12:12] };
    end 
    if(N3422) begin
      { mem[171:171] } <= { data_i[11:11] };
    end 
    if(N3421) begin
      { mem[170:170] } <= { data_i[10:10] };
    end 
    if(N3420) begin
      { mem[169:169] } <= { data_i[9:9] };
    end 
    if(N3419) begin
      { mem[168:168] } <= { data_i[8:8] };
    end 
    if(N3418) begin
      { mem[167:167] } <= { data_i[7:7] };
    end 
    if(N3417) begin
      { mem[166:166] } <= { data_i[6:6] };
    end 
    if(N3416) begin
      { mem[165:165] } <= { data_i[5:5] };
    end 
    if(N3415) begin
      { mem[164:164] } <= { data_i[4:4] };
    end 
    if(N3414) begin
      { mem[163:163] } <= { data_i[3:3] };
    end 
    if(N3413) begin
      { mem[162:162] } <= { data_i[2:2] };
    end 
    if(N3412) begin
      { mem[161:161] } <= { data_i[1:1] };
    end 
    if(N3411) begin
      { mem[160:160] } <= { data_i[0:0] };
    end 
    if(N3410) begin
      { mem[159:159] } <= { data_i[39:39] };
    end 
    if(N3409) begin
      { mem[158:158] } <= { data_i[38:38] };
    end 
    if(N3408) begin
      { mem[157:157] } <= { data_i[37:37] };
    end 
    if(N3407) begin
      { mem[156:156] } <= { data_i[36:36] };
    end 
    if(N3406) begin
      { mem[155:155] } <= { data_i[35:35] };
    end 
    if(N3405) begin
      { mem[154:154] } <= { data_i[34:34] };
    end 
    if(N3404) begin
      { mem[153:153] } <= { data_i[33:33] };
    end 
    if(N3403) begin
      { mem[152:152] } <= { data_i[32:32] };
    end 
    if(N3402) begin
      { mem[151:151] } <= { data_i[31:31] };
    end 
    if(N3401) begin
      { mem[150:150] } <= { data_i[30:30] };
    end 
    if(N3400) begin
      { mem[149:149] } <= { data_i[29:29] };
    end 
    if(N3399) begin
      { mem[148:148] } <= { data_i[28:28] };
    end 
    if(N3398) begin
      { mem[147:147] } <= { data_i[27:27] };
    end 
    if(N3397) begin
      { mem[146:146] } <= { data_i[26:26] };
    end 
    if(N3396) begin
      { mem[145:145] } <= { data_i[25:25] };
    end 
    if(N3395) begin
      { mem[144:144] } <= { data_i[24:24] };
    end 
    if(N3394) begin
      { mem[143:143] } <= { data_i[23:23] };
    end 
    if(N3393) begin
      { mem[142:142] } <= { data_i[22:22] };
    end 
    if(N3392) begin
      { mem[141:141] } <= { data_i[21:21] };
    end 
    if(N3391) begin
      { mem[140:140] } <= { data_i[20:20] };
    end 
    if(N3390) begin
      { mem[139:139] } <= { data_i[19:19] };
    end 
    if(N3389) begin
      { mem[138:138] } <= { data_i[18:18] };
    end 
    if(N3388) begin
      { mem[137:137] } <= { data_i[17:17] };
    end 
    if(N3387) begin
      { mem[136:136] } <= { data_i[16:16] };
    end 
    if(N3386) begin
      { mem[135:135] } <= { data_i[15:15] };
    end 
    if(N3385) begin
      { mem[134:134] } <= { data_i[14:14] };
    end 
    if(N3384) begin
      { mem[133:133] } <= { data_i[13:13] };
    end 
    if(N3383) begin
      { mem[132:132] } <= { data_i[12:12] };
    end 
    if(N3382) begin
      { mem[131:131] } <= { data_i[11:11] };
    end 
    if(N3381) begin
      { mem[130:130] } <= { data_i[10:10] };
    end 
    if(N3380) begin
      { mem[129:129] } <= { data_i[9:9] };
    end 
    if(N3379) begin
      { mem[128:128] } <= { data_i[8:8] };
    end 
    if(N3378) begin
      { mem[127:127] } <= { data_i[7:7] };
    end 
    if(N3377) begin
      { mem[126:126] } <= { data_i[6:6] };
    end 
    if(N3376) begin
      { mem[125:125] } <= { data_i[5:5] };
    end 
    if(N3375) begin
      { mem[124:124] } <= { data_i[4:4] };
    end 
    if(N3374) begin
      { mem[123:123] } <= { data_i[3:3] };
    end 
    if(N3373) begin
      { mem[122:122] } <= { data_i[2:2] };
    end 
    if(N3372) begin
      { mem[121:121] } <= { data_i[1:1] };
    end 
    if(N3371) begin
      { mem[120:120] } <= { data_i[0:0] };
    end 
    if(N3370) begin
      { mem[119:119] } <= { data_i[39:39] };
    end 
    if(N3369) begin
      { mem[118:118] } <= { data_i[38:38] };
    end 
    if(N3368) begin
      { mem[117:117] } <= { data_i[37:37] };
    end 
    if(N3367) begin
      { mem[116:116] } <= { data_i[36:36] };
    end 
    if(N3366) begin
      { mem[115:115] } <= { data_i[35:35] };
    end 
    if(N3365) begin
      { mem[114:114] } <= { data_i[34:34] };
    end 
    if(N3364) begin
      { mem[113:113] } <= { data_i[33:33] };
    end 
    if(N3363) begin
      { mem[112:112] } <= { data_i[32:32] };
    end 
    if(N3362) begin
      { mem[111:111] } <= { data_i[31:31] };
    end 
    if(N3361) begin
      { mem[110:110] } <= { data_i[30:30] };
    end 
    if(N3360) begin
      { mem[109:109] } <= { data_i[29:29] };
    end 
    if(N3359) begin
      { mem[108:108] } <= { data_i[28:28] };
    end 
    if(N3358) begin
      { mem[107:107] } <= { data_i[27:27] };
    end 
    if(N3357) begin
      { mem[106:106] } <= { data_i[26:26] };
    end 
    if(N3356) begin
      { mem[105:105] } <= { data_i[25:25] };
    end 
    if(N3355) begin
      { mem[104:104] } <= { data_i[24:24] };
    end 
    if(N3354) begin
      { mem[103:103] } <= { data_i[23:23] };
    end 
    if(N3353) begin
      { mem[102:102] } <= { data_i[22:22] };
    end 
    if(N3352) begin
      { mem[101:101] } <= { data_i[21:21] };
    end 
    if(N3351) begin
      { mem[100:100] } <= { data_i[20:20] };
    end 
    if(N3350) begin
      { mem[99:99] } <= { data_i[19:19] };
    end 
    if(N3349) begin
      { mem[98:98] } <= { data_i[18:18] };
    end 
    if(N3348) begin
      { mem[97:97] } <= { data_i[17:17] };
    end 
    if(N3347) begin
      { mem[96:96] } <= { data_i[16:16] };
    end 
    if(N3346) begin
      { mem[95:95] } <= { data_i[15:15] };
    end 
    if(N3345) begin
      { mem[94:94] } <= { data_i[14:14] };
    end 
    if(N3344) begin
      { mem[93:93] } <= { data_i[13:13] };
    end 
    if(N3343) begin
      { mem[92:92] } <= { data_i[12:12] };
    end 
    if(N3342) begin
      { mem[91:91] } <= { data_i[11:11] };
    end 
    if(N3341) begin
      { mem[90:90] } <= { data_i[10:10] };
    end 
    if(N3340) begin
      { mem[89:89] } <= { data_i[9:9] };
    end 
    if(N3339) begin
      { mem[88:88] } <= { data_i[8:8] };
    end 
    if(N3338) begin
      { mem[87:87] } <= { data_i[7:7] };
    end 
    if(N3337) begin
      { mem[86:86] } <= { data_i[6:6] };
    end 
    if(N3336) begin
      { mem[85:85] } <= { data_i[5:5] };
    end 
    if(N3335) begin
      { mem[84:84] } <= { data_i[4:4] };
    end 
    if(N3334) begin
      { mem[83:83] } <= { data_i[3:3] };
    end 
    if(N3333) begin
      { mem[82:82] } <= { data_i[2:2] };
    end 
    if(N3332) begin
      { mem[81:81] } <= { data_i[1:1] };
    end 
    if(N3331) begin
      { mem[80:80] } <= { data_i[0:0] };
    end 
    if(N3330) begin
      { mem[79:79] } <= { data_i[39:39] };
    end 
    if(N3329) begin
      { mem[78:78] } <= { data_i[38:38] };
    end 
    if(N3328) begin
      { mem[77:77] } <= { data_i[37:37] };
    end 
    if(N3327) begin
      { mem[76:76] } <= { data_i[36:36] };
    end 
    if(N3326) begin
      { mem[75:75] } <= { data_i[35:35] };
    end 
    if(N3325) begin
      { mem[74:74] } <= { data_i[34:34] };
    end 
    if(N3324) begin
      { mem[73:73] } <= { data_i[33:33] };
    end 
    if(N3323) begin
      { mem[72:72] } <= { data_i[32:32] };
    end 
    if(N3322) begin
      { mem[71:71] } <= { data_i[31:31] };
    end 
    if(N3321) begin
      { mem[70:70] } <= { data_i[30:30] };
    end 
    if(N3320) begin
      { mem[69:69] } <= { data_i[29:29] };
    end 
    if(N3319) begin
      { mem[68:68] } <= { data_i[28:28] };
    end 
    if(N3318) begin
      { mem[67:67] } <= { data_i[27:27] };
    end 
    if(N3317) begin
      { mem[66:66] } <= { data_i[26:26] };
    end 
    if(N3316) begin
      { mem[65:65] } <= { data_i[25:25] };
    end 
    if(N3315) begin
      { mem[64:64] } <= { data_i[24:24] };
    end 
    if(N3314) begin
      { mem[63:63] } <= { data_i[23:23] };
    end 
    if(N3313) begin
      { mem[62:62] } <= { data_i[22:22] };
    end 
    if(N3312) begin
      { mem[61:61] } <= { data_i[21:21] };
    end 
    if(N3311) begin
      { mem[60:60] } <= { data_i[20:20] };
    end 
    if(N3310) begin
      { mem[59:59] } <= { data_i[19:19] };
    end 
    if(N3309) begin
      { mem[58:58] } <= { data_i[18:18] };
    end 
    if(N3308) begin
      { mem[57:57] } <= { data_i[17:17] };
    end 
    if(N3307) begin
      { mem[56:56] } <= { data_i[16:16] };
    end 
    if(N3306) begin
      { mem[55:55] } <= { data_i[15:15] };
    end 
    if(N3305) begin
      { mem[54:54] } <= { data_i[14:14] };
    end 
    if(N3304) begin
      { mem[53:53] } <= { data_i[13:13] };
    end 
    if(N3303) begin
      { mem[52:52] } <= { data_i[12:12] };
    end 
    if(N3302) begin
      { mem[51:51] } <= { data_i[11:11] };
    end 
    if(N3301) begin
      { mem[50:50] } <= { data_i[10:10] };
    end 
    if(N3300) begin
      { mem[49:49] } <= { data_i[9:9] };
    end 
    if(N3299) begin
      { mem[48:48] } <= { data_i[8:8] };
    end 
    if(N3298) begin
      { mem[47:47] } <= { data_i[7:7] };
    end 
    if(N3297) begin
      { mem[46:46] } <= { data_i[6:6] };
    end 
    if(N3296) begin
      { mem[45:45] } <= { data_i[5:5] };
    end 
    if(N3295) begin
      { mem[44:44] } <= { data_i[4:4] };
    end 
    if(N3294) begin
      { mem[43:43] } <= { data_i[3:3] };
    end 
    if(N3293) begin
      { mem[42:42] } <= { data_i[2:2] };
    end 
    if(N3292) begin
      { mem[41:41] } <= { data_i[1:1] };
    end 
    if(N3291) begin
      { mem[40:40] } <= { data_i[0:0] };
    end 
    if(N3290) begin
      { mem[39:39] } <= { data_i[39:39] };
    end 
    if(N3289) begin
      { mem[38:38] } <= { data_i[38:38] };
    end 
    if(N3288) begin
      { mem[37:37] } <= { data_i[37:37] };
    end 
    if(N3287) begin
      { mem[36:36] } <= { data_i[36:36] };
    end 
    if(N3286) begin
      { mem[35:35] } <= { data_i[35:35] };
    end 
    if(N3285) begin
      { mem[34:34] } <= { data_i[34:34] };
    end 
    if(N3284) begin
      { mem[33:33] } <= { data_i[33:33] };
    end 
    if(N3283) begin
      { mem[32:32] } <= { data_i[32:32] };
    end 
    if(N3282) begin
      { mem[31:31] } <= { data_i[31:31] };
    end 
    if(N3281) begin
      { mem[30:30] } <= { data_i[30:30] };
    end 
    if(N3280) begin
      { mem[29:29] } <= { data_i[29:29] };
    end 
    if(N3279) begin
      { mem[28:28] } <= { data_i[28:28] };
    end 
    if(N3278) begin
      { mem[27:27] } <= { data_i[27:27] };
    end 
    if(N3277) begin
      { mem[26:26] } <= { data_i[26:26] };
    end 
    if(N3276) begin
      { mem[25:25] } <= { data_i[25:25] };
    end 
    if(N3275) begin
      { mem[24:24] } <= { data_i[24:24] };
    end 
    if(N3274) begin
      { mem[23:23] } <= { data_i[23:23] };
    end 
    if(N3273) begin
      { mem[22:22] } <= { data_i[22:22] };
    end 
    if(N3272) begin
      { mem[21:21] } <= { data_i[21:21] };
    end 
    if(N3271) begin
      { mem[20:20] } <= { data_i[20:20] };
    end 
    if(N3270) begin
      { mem[19:19] } <= { data_i[19:19] };
    end 
    if(N3269) begin
      { mem[18:18] } <= { data_i[18:18] };
    end 
    if(N3268) begin
      { mem[17:17] } <= { data_i[17:17] };
    end 
    if(N3267) begin
      { mem[16:16] } <= { data_i[16:16] };
    end 
    if(N3266) begin
      { mem[15:15] } <= { data_i[15:15] };
    end 
    if(N3265) begin
      { mem[14:14] } <= { data_i[14:14] };
    end 
    if(N3264) begin
      { mem[13:13] } <= { data_i[13:13] };
    end 
    if(N3263) begin
      { mem[12:12] } <= { data_i[12:12] };
    end 
    if(N3262) begin
      { mem[11:11] } <= { data_i[11:11] };
    end 
    if(N3261) begin
      { mem[10:10] } <= { data_i[10:10] };
    end 
    if(N3260) begin
      { mem[9:9] } <= { data_i[9:9] };
    end 
    if(N3259) begin
      { mem[8:8] } <= { data_i[8:8] };
    end 
    if(N3258) begin
      { mem[7:7] } <= { data_i[7:7] };
    end 
    if(N3257) begin
      { mem[6:6] } <= { data_i[6:6] };
    end 
    if(N3256) begin
      { mem[5:5] } <= { data_i[5:5] };
    end 
    if(N3255) begin
      { mem[4:4] } <= { data_i[4:4] };
    end 
    if(N3254) begin
      { mem[3:3] } <= { data_i[3:3] };
    end 
    if(N3253) begin
      { mem[2:2] } <= { data_i[2:2] };
    end 
    if(N3252) begin
      { mem[1:1] } <= { data_i[1:1] };
    end 
    if(N3251) begin
      { mem[0:0] } <= { data_i[0:0] };
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p40_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [39:0] data_i;
  input [5:0] addr_i;
  input [39:0] w_mask_i;
  output [39:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [39:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p40_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_en_width_p8_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input en_i;
  reg [7:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[7:0] } <= { data_i[7:0] };
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p8
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input en_i;
  wire [7:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p8_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_synth_width_p8_els_p256_latch_last_read_p1
(
  clk_i,
  v_i,
  reset_i,
  data_i,
  addr_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [7:0] addr_i;
  output [7:0] data_o;
  input clk_i;
  input v_i;
  input reset_i;
  input w_i;
  wire [7:0] data_o,data_out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,read_en,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,llr_read_en_r,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,
  N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,
  N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,
  N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,
  N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,
  N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,
  N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,
  N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,
  N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095;
  reg [7:0] addr_r;
  reg [2047:0] mem;
  assign data_out[7] = (N277)? mem[7] : 
                       (N279)? mem[15] : 
                       (N281)? mem[23] : 
                       (N283)? mem[31] : 
                       (N285)? mem[39] : 
                       (N287)? mem[47] : 
                       (N289)? mem[55] : 
                       (N291)? mem[63] : 
                       (N293)? mem[71] : 
                       (N295)? mem[79] : 
                       (N297)? mem[87] : 
                       (N299)? mem[95] : 
                       (N301)? mem[103] : 
                       (N303)? mem[111] : 
                       (N305)? mem[119] : 
                       (N307)? mem[127] : 
                       (N309)? mem[135] : 
                       (N311)? mem[143] : 
                       (N313)? mem[151] : 
                       (N315)? mem[159] : 
                       (N317)? mem[167] : 
                       (N319)? mem[175] : 
                       (N321)? mem[183] : 
                       (N323)? mem[191] : 
                       (N325)? mem[199] : 
                       (N327)? mem[207] : 
                       (N329)? mem[215] : 
                       (N331)? mem[223] : 
                       (N333)? mem[231] : 
                       (N335)? mem[239] : 
                       (N337)? mem[247] : 
                       (N339)? mem[255] : 
                       (N341)? mem[263] : 
                       (N343)? mem[271] : 
                       (N345)? mem[279] : 
                       (N347)? mem[287] : 
                       (N349)? mem[295] : 
                       (N351)? mem[303] : 
                       (N353)? mem[311] : 
                       (N355)? mem[319] : 
                       (N357)? mem[327] : 
                       (N359)? mem[335] : 
                       (N361)? mem[343] : 
                       (N363)? mem[351] : 
                       (N365)? mem[359] : 
                       (N367)? mem[367] : 
                       (N369)? mem[375] : 
                       (N371)? mem[383] : 
                       (N373)? mem[391] : 
                       (N375)? mem[399] : 
                       (N377)? mem[407] : 
                       (N379)? mem[415] : 
                       (N381)? mem[423] : 
                       (N383)? mem[431] : 
                       (N385)? mem[439] : 
                       (N387)? mem[447] : 
                       (N389)? mem[455] : 
                       (N391)? mem[463] : 
                       (N393)? mem[471] : 
                       (N395)? mem[479] : 
                       (N397)? mem[487] : 
                       (N399)? mem[495] : 
                       (N401)? mem[503] : 
                       (N403)? mem[511] : 
                       (N405)? mem[519] : 
                       (N407)? mem[527] : 
                       (N409)? mem[535] : 
                       (N411)? mem[543] : 
                       (N413)? mem[551] : 
                       (N415)? mem[559] : 
                       (N417)? mem[567] : 
                       (N419)? mem[575] : 
                       (N421)? mem[583] : 
                       (N423)? mem[591] : 
                       (N425)? mem[599] : 
                       (N427)? mem[607] : 
                       (N429)? mem[615] : 
                       (N431)? mem[623] : 
                       (N433)? mem[631] : 
                       (N435)? mem[639] : 
                       (N437)? mem[647] : 
                       (N439)? mem[655] : 
                       (N441)? mem[663] : 
                       (N443)? mem[671] : 
                       (N445)? mem[679] : 
                       (N447)? mem[687] : 
                       (N449)? mem[695] : 
                       (N451)? mem[703] : 
                       (N453)? mem[711] : 
                       (N455)? mem[719] : 
                       (N457)? mem[727] : 
                       (N459)? mem[735] : 
                       (N461)? mem[743] : 
                       (N463)? mem[751] : 
                       (N465)? mem[759] : 
                       (N467)? mem[767] : 
                       (N469)? mem[775] : 
                       (N471)? mem[783] : 
                       (N473)? mem[791] : 
                       (N475)? mem[799] : 
                       (N477)? mem[807] : 
                       (N479)? mem[815] : 
                       (N481)? mem[823] : 
                       (N483)? mem[831] : 
                       (N485)? mem[839] : 
                       (N487)? mem[847] : 
                       (N489)? mem[855] : 
                       (N491)? mem[863] : 
                       (N493)? mem[871] : 
                       (N495)? mem[879] : 
                       (N497)? mem[887] : 
                       (N499)? mem[895] : 
                       (N501)? mem[903] : 
                       (N503)? mem[911] : 
                       (N505)? mem[919] : 
                       (N507)? mem[927] : 
                       (N509)? mem[935] : 
                       (N511)? mem[943] : 
                       (N513)? mem[951] : 
                       (N515)? mem[959] : 
                       (N517)? mem[967] : 
                       (N519)? mem[975] : 
                       (N521)? mem[983] : 
                       (N523)? mem[991] : 
                       (N525)? mem[999] : 
                       (N527)? mem[1007] : 
                       (N529)? mem[1015] : 
                       (N531)? mem[1023] : 
                       (N278)? mem[1031] : 
                       (N280)? mem[1039] : 
                       (N282)? mem[1047] : 
                       (N284)? mem[1055] : 
                       (N286)? mem[1063] : 
                       (N288)? mem[1071] : 
                       (N290)? mem[1079] : 
                       (N292)? mem[1087] : 
                       (N294)? mem[1095] : 
                       (N296)? mem[1103] : 
                       (N298)? mem[1111] : 
                       (N300)? mem[1119] : 
                       (N302)? mem[1127] : 
                       (N304)? mem[1135] : 
                       (N306)? mem[1143] : 
                       (N308)? mem[1151] : 
                       (N310)? mem[1159] : 
                       (N312)? mem[1167] : 
                       (N314)? mem[1175] : 
                       (N316)? mem[1183] : 
                       (N318)? mem[1191] : 
                       (N320)? mem[1199] : 
                       (N322)? mem[1207] : 
                       (N324)? mem[1215] : 
                       (N326)? mem[1223] : 
                       (N328)? mem[1231] : 
                       (N330)? mem[1239] : 
                       (N332)? mem[1247] : 
                       (N334)? mem[1255] : 
                       (N336)? mem[1263] : 
                       (N338)? mem[1271] : 
                       (N340)? mem[1279] : 
                       (N342)? mem[1287] : 
                       (N344)? mem[1295] : 
                       (N346)? mem[1303] : 
                       (N348)? mem[1311] : 
                       (N350)? mem[1319] : 
                       (N352)? mem[1327] : 
                       (N354)? mem[1335] : 
                       (N356)? mem[1343] : 
                       (N358)? mem[1351] : 
                       (N360)? mem[1359] : 
                       (N362)? mem[1367] : 
                       (N364)? mem[1375] : 
                       (N366)? mem[1383] : 
                       (N368)? mem[1391] : 
                       (N370)? mem[1399] : 
                       (N372)? mem[1407] : 
                       (N374)? mem[1415] : 
                       (N376)? mem[1423] : 
                       (N378)? mem[1431] : 
                       (N380)? mem[1439] : 
                       (N382)? mem[1447] : 
                       (N384)? mem[1455] : 
                       (N386)? mem[1463] : 
                       (N388)? mem[1471] : 
                       (N390)? mem[1479] : 
                       (N392)? mem[1487] : 
                       (N394)? mem[1495] : 
                       (N396)? mem[1503] : 
                       (N398)? mem[1511] : 
                       (N400)? mem[1519] : 
                       (N402)? mem[1527] : 
                       (N404)? mem[1535] : 
                       (N406)? mem[1543] : 
                       (N408)? mem[1551] : 
                       (N410)? mem[1559] : 
                       (N412)? mem[1567] : 
                       (N414)? mem[1575] : 
                       (N416)? mem[1583] : 
                       (N418)? mem[1591] : 
                       (N420)? mem[1599] : 
                       (N422)? mem[1607] : 
                       (N424)? mem[1615] : 
                       (N426)? mem[1623] : 
                       (N428)? mem[1631] : 
                       (N430)? mem[1639] : 
                       (N432)? mem[1647] : 
                       (N434)? mem[1655] : 
                       (N436)? mem[1663] : 
                       (N438)? mem[1671] : 
                       (N440)? mem[1679] : 
                       (N442)? mem[1687] : 
                       (N444)? mem[1695] : 
                       (N446)? mem[1703] : 
                       (N448)? mem[1711] : 
                       (N450)? mem[1719] : 
                       (N452)? mem[1727] : 
                       (N454)? mem[1735] : 
                       (N456)? mem[1743] : 
                       (N458)? mem[1751] : 
                       (N460)? mem[1759] : 
                       (N462)? mem[1767] : 
                       (N464)? mem[1775] : 
                       (N466)? mem[1783] : 
                       (N468)? mem[1791] : 
                       (N470)? mem[1799] : 
                       (N472)? mem[1807] : 
                       (N474)? mem[1815] : 
                       (N476)? mem[1823] : 
                       (N478)? mem[1831] : 
                       (N480)? mem[1839] : 
                       (N482)? mem[1847] : 
                       (N484)? mem[1855] : 
                       (N486)? mem[1863] : 
                       (N488)? mem[1871] : 
                       (N490)? mem[1879] : 
                       (N492)? mem[1887] : 
                       (N494)? mem[1895] : 
                       (N496)? mem[1903] : 
                       (N498)? mem[1911] : 
                       (N500)? mem[1919] : 
                       (N502)? mem[1927] : 
                       (N504)? mem[1935] : 
                       (N506)? mem[1943] : 
                       (N508)? mem[1951] : 
                       (N510)? mem[1959] : 
                       (N512)? mem[1967] : 
                       (N514)? mem[1975] : 
                       (N516)? mem[1983] : 
                       (N518)? mem[1991] : 
                       (N520)? mem[1999] : 
                       (N522)? mem[2007] : 
                       (N524)? mem[2015] : 
                       (N526)? mem[2023] : 
                       (N528)? mem[2031] : 
                       (N530)? mem[2039] : 
                       (N532)? mem[2047] : 1'b0;
  assign data_out[6] = (N277)? mem[6] : 
                       (N279)? mem[14] : 
                       (N281)? mem[22] : 
                       (N283)? mem[30] : 
                       (N285)? mem[38] : 
                       (N287)? mem[46] : 
                       (N289)? mem[54] : 
                       (N291)? mem[62] : 
                       (N293)? mem[70] : 
                       (N295)? mem[78] : 
                       (N297)? mem[86] : 
                       (N299)? mem[94] : 
                       (N301)? mem[102] : 
                       (N303)? mem[110] : 
                       (N305)? mem[118] : 
                       (N307)? mem[126] : 
                       (N309)? mem[134] : 
                       (N311)? mem[142] : 
                       (N313)? mem[150] : 
                       (N315)? mem[158] : 
                       (N317)? mem[166] : 
                       (N319)? mem[174] : 
                       (N321)? mem[182] : 
                       (N323)? mem[190] : 
                       (N325)? mem[198] : 
                       (N327)? mem[206] : 
                       (N329)? mem[214] : 
                       (N331)? mem[222] : 
                       (N333)? mem[230] : 
                       (N335)? mem[238] : 
                       (N337)? mem[246] : 
                       (N339)? mem[254] : 
                       (N341)? mem[262] : 
                       (N343)? mem[270] : 
                       (N345)? mem[278] : 
                       (N347)? mem[286] : 
                       (N349)? mem[294] : 
                       (N351)? mem[302] : 
                       (N353)? mem[310] : 
                       (N355)? mem[318] : 
                       (N357)? mem[326] : 
                       (N359)? mem[334] : 
                       (N361)? mem[342] : 
                       (N363)? mem[350] : 
                       (N365)? mem[358] : 
                       (N367)? mem[366] : 
                       (N369)? mem[374] : 
                       (N371)? mem[382] : 
                       (N373)? mem[390] : 
                       (N375)? mem[398] : 
                       (N377)? mem[406] : 
                       (N379)? mem[414] : 
                       (N381)? mem[422] : 
                       (N383)? mem[430] : 
                       (N385)? mem[438] : 
                       (N387)? mem[446] : 
                       (N389)? mem[454] : 
                       (N391)? mem[462] : 
                       (N393)? mem[470] : 
                       (N395)? mem[478] : 
                       (N397)? mem[486] : 
                       (N399)? mem[494] : 
                       (N401)? mem[502] : 
                       (N403)? mem[510] : 
                       (N405)? mem[518] : 
                       (N407)? mem[526] : 
                       (N409)? mem[534] : 
                       (N411)? mem[542] : 
                       (N413)? mem[550] : 
                       (N415)? mem[558] : 
                       (N417)? mem[566] : 
                       (N419)? mem[574] : 
                       (N421)? mem[582] : 
                       (N423)? mem[590] : 
                       (N425)? mem[598] : 
                       (N427)? mem[606] : 
                       (N429)? mem[614] : 
                       (N431)? mem[622] : 
                       (N433)? mem[630] : 
                       (N435)? mem[638] : 
                       (N437)? mem[646] : 
                       (N439)? mem[654] : 
                       (N441)? mem[662] : 
                       (N443)? mem[670] : 
                       (N445)? mem[678] : 
                       (N447)? mem[686] : 
                       (N449)? mem[694] : 
                       (N451)? mem[702] : 
                       (N453)? mem[710] : 
                       (N455)? mem[718] : 
                       (N457)? mem[726] : 
                       (N459)? mem[734] : 
                       (N461)? mem[742] : 
                       (N463)? mem[750] : 
                       (N465)? mem[758] : 
                       (N467)? mem[766] : 
                       (N469)? mem[774] : 
                       (N471)? mem[782] : 
                       (N473)? mem[790] : 
                       (N475)? mem[798] : 
                       (N477)? mem[806] : 
                       (N479)? mem[814] : 
                       (N481)? mem[822] : 
                       (N483)? mem[830] : 
                       (N485)? mem[838] : 
                       (N487)? mem[846] : 
                       (N489)? mem[854] : 
                       (N491)? mem[862] : 
                       (N493)? mem[870] : 
                       (N495)? mem[878] : 
                       (N497)? mem[886] : 
                       (N499)? mem[894] : 
                       (N501)? mem[902] : 
                       (N503)? mem[910] : 
                       (N505)? mem[918] : 
                       (N507)? mem[926] : 
                       (N509)? mem[934] : 
                       (N511)? mem[942] : 
                       (N513)? mem[950] : 
                       (N515)? mem[958] : 
                       (N517)? mem[966] : 
                       (N519)? mem[974] : 
                       (N521)? mem[982] : 
                       (N523)? mem[990] : 
                       (N525)? mem[998] : 
                       (N527)? mem[1006] : 
                       (N529)? mem[1014] : 
                       (N531)? mem[1022] : 
                       (N278)? mem[1030] : 
                       (N280)? mem[1038] : 
                       (N282)? mem[1046] : 
                       (N284)? mem[1054] : 
                       (N286)? mem[1062] : 
                       (N288)? mem[1070] : 
                       (N290)? mem[1078] : 
                       (N292)? mem[1086] : 
                       (N294)? mem[1094] : 
                       (N296)? mem[1102] : 
                       (N298)? mem[1110] : 
                       (N300)? mem[1118] : 
                       (N302)? mem[1126] : 
                       (N304)? mem[1134] : 
                       (N306)? mem[1142] : 
                       (N308)? mem[1150] : 
                       (N310)? mem[1158] : 
                       (N312)? mem[1166] : 
                       (N314)? mem[1174] : 
                       (N316)? mem[1182] : 
                       (N318)? mem[1190] : 
                       (N320)? mem[1198] : 
                       (N322)? mem[1206] : 
                       (N324)? mem[1214] : 
                       (N326)? mem[1222] : 
                       (N328)? mem[1230] : 
                       (N330)? mem[1238] : 
                       (N332)? mem[1246] : 
                       (N334)? mem[1254] : 
                       (N336)? mem[1262] : 
                       (N338)? mem[1270] : 
                       (N340)? mem[1278] : 
                       (N342)? mem[1286] : 
                       (N344)? mem[1294] : 
                       (N346)? mem[1302] : 
                       (N348)? mem[1310] : 
                       (N350)? mem[1318] : 
                       (N352)? mem[1326] : 
                       (N354)? mem[1334] : 
                       (N356)? mem[1342] : 
                       (N358)? mem[1350] : 
                       (N360)? mem[1358] : 
                       (N362)? mem[1366] : 
                       (N364)? mem[1374] : 
                       (N366)? mem[1382] : 
                       (N368)? mem[1390] : 
                       (N370)? mem[1398] : 
                       (N372)? mem[1406] : 
                       (N374)? mem[1414] : 
                       (N376)? mem[1422] : 
                       (N378)? mem[1430] : 
                       (N380)? mem[1438] : 
                       (N382)? mem[1446] : 
                       (N384)? mem[1454] : 
                       (N386)? mem[1462] : 
                       (N388)? mem[1470] : 
                       (N390)? mem[1478] : 
                       (N392)? mem[1486] : 
                       (N394)? mem[1494] : 
                       (N396)? mem[1502] : 
                       (N398)? mem[1510] : 
                       (N400)? mem[1518] : 
                       (N402)? mem[1526] : 
                       (N404)? mem[1534] : 
                       (N406)? mem[1542] : 
                       (N408)? mem[1550] : 
                       (N410)? mem[1558] : 
                       (N412)? mem[1566] : 
                       (N414)? mem[1574] : 
                       (N416)? mem[1582] : 
                       (N418)? mem[1590] : 
                       (N420)? mem[1598] : 
                       (N422)? mem[1606] : 
                       (N424)? mem[1614] : 
                       (N426)? mem[1622] : 
                       (N428)? mem[1630] : 
                       (N430)? mem[1638] : 
                       (N432)? mem[1646] : 
                       (N434)? mem[1654] : 
                       (N436)? mem[1662] : 
                       (N438)? mem[1670] : 
                       (N440)? mem[1678] : 
                       (N442)? mem[1686] : 
                       (N444)? mem[1694] : 
                       (N446)? mem[1702] : 
                       (N448)? mem[1710] : 
                       (N450)? mem[1718] : 
                       (N452)? mem[1726] : 
                       (N454)? mem[1734] : 
                       (N456)? mem[1742] : 
                       (N458)? mem[1750] : 
                       (N460)? mem[1758] : 
                       (N462)? mem[1766] : 
                       (N464)? mem[1774] : 
                       (N466)? mem[1782] : 
                       (N468)? mem[1790] : 
                       (N470)? mem[1798] : 
                       (N472)? mem[1806] : 
                       (N474)? mem[1814] : 
                       (N476)? mem[1822] : 
                       (N478)? mem[1830] : 
                       (N480)? mem[1838] : 
                       (N482)? mem[1846] : 
                       (N484)? mem[1854] : 
                       (N486)? mem[1862] : 
                       (N488)? mem[1870] : 
                       (N490)? mem[1878] : 
                       (N492)? mem[1886] : 
                       (N494)? mem[1894] : 
                       (N496)? mem[1902] : 
                       (N498)? mem[1910] : 
                       (N500)? mem[1918] : 
                       (N502)? mem[1926] : 
                       (N504)? mem[1934] : 
                       (N506)? mem[1942] : 
                       (N508)? mem[1950] : 
                       (N510)? mem[1958] : 
                       (N512)? mem[1966] : 
                       (N514)? mem[1974] : 
                       (N516)? mem[1982] : 
                       (N518)? mem[1990] : 
                       (N520)? mem[1998] : 
                       (N522)? mem[2006] : 
                       (N524)? mem[2014] : 
                       (N526)? mem[2022] : 
                       (N528)? mem[2030] : 
                       (N530)? mem[2038] : 
                       (N532)? mem[2046] : 1'b0;
  assign data_out[5] = (N277)? mem[5] : 
                       (N279)? mem[13] : 
                       (N281)? mem[21] : 
                       (N283)? mem[29] : 
                       (N285)? mem[37] : 
                       (N287)? mem[45] : 
                       (N289)? mem[53] : 
                       (N291)? mem[61] : 
                       (N293)? mem[69] : 
                       (N295)? mem[77] : 
                       (N297)? mem[85] : 
                       (N299)? mem[93] : 
                       (N301)? mem[101] : 
                       (N303)? mem[109] : 
                       (N305)? mem[117] : 
                       (N307)? mem[125] : 
                       (N309)? mem[133] : 
                       (N311)? mem[141] : 
                       (N313)? mem[149] : 
                       (N315)? mem[157] : 
                       (N317)? mem[165] : 
                       (N319)? mem[173] : 
                       (N321)? mem[181] : 
                       (N323)? mem[189] : 
                       (N325)? mem[197] : 
                       (N327)? mem[205] : 
                       (N329)? mem[213] : 
                       (N331)? mem[221] : 
                       (N333)? mem[229] : 
                       (N335)? mem[237] : 
                       (N337)? mem[245] : 
                       (N339)? mem[253] : 
                       (N341)? mem[261] : 
                       (N343)? mem[269] : 
                       (N345)? mem[277] : 
                       (N347)? mem[285] : 
                       (N349)? mem[293] : 
                       (N351)? mem[301] : 
                       (N353)? mem[309] : 
                       (N355)? mem[317] : 
                       (N357)? mem[325] : 
                       (N359)? mem[333] : 
                       (N361)? mem[341] : 
                       (N363)? mem[349] : 
                       (N365)? mem[357] : 
                       (N367)? mem[365] : 
                       (N369)? mem[373] : 
                       (N371)? mem[381] : 
                       (N373)? mem[389] : 
                       (N375)? mem[397] : 
                       (N377)? mem[405] : 
                       (N379)? mem[413] : 
                       (N381)? mem[421] : 
                       (N383)? mem[429] : 
                       (N385)? mem[437] : 
                       (N387)? mem[445] : 
                       (N389)? mem[453] : 
                       (N391)? mem[461] : 
                       (N393)? mem[469] : 
                       (N395)? mem[477] : 
                       (N397)? mem[485] : 
                       (N399)? mem[493] : 
                       (N401)? mem[501] : 
                       (N403)? mem[509] : 
                       (N405)? mem[517] : 
                       (N407)? mem[525] : 
                       (N409)? mem[533] : 
                       (N411)? mem[541] : 
                       (N413)? mem[549] : 
                       (N415)? mem[557] : 
                       (N417)? mem[565] : 
                       (N419)? mem[573] : 
                       (N421)? mem[581] : 
                       (N423)? mem[589] : 
                       (N425)? mem[597] : 
                       (N427)? mem[605] : 
                       (N429)? mem[613] : 
                       (N431)? mem[621] : 
                       (N433)? mem[629] : 
                       (N435)? mem[637] : 
                       (N437)? mem[645] : 
                       (N439)? mem[653] : 
                       (N441)? mem[661] : 
                       (N443)? mem[669] : 
                       (N445)? mem[677] : 
                       (N447)? mem[685] : 
                       (N449)? mem[693] : 
                       (N451)? mem[701] : 
                       (N453)? mem[709] : 
                       (N455)? mem[717] : 
                       (N457)? mem[725] : 
                       (N459)? mem[733] : 
                       (N461)? mem[741] : 
                       (N463)? mem[749] : 
                       (N465)? mem[757] : 
                       (N467)? mem[765] : 
                       (N469)? mem[773] : 
                       (N471)? mem[781] : 
                       (N473)? mem[789] : 
                       (N475)? mem[797] : 
                       (N477)? mem[805] : 
                       (N479)? mem[813] : 
                       (N481)? mem[821] : 
                       (N483)? mem[829] : 
                       (N485)? mem[837] : 
                       (N487)? mem[845] : 
                       (N489)? mem[853] : 
                       (N491)? mem[861] : 
                       (N493)? mem[869] : 
                       (N495)? mem[877] : 
                       (N497)? mem[885] : 
                       (N499)? mem[893] : 
                       (N501)? mem[901] : 
                       (N503)? mem[909] : 
                       (N505)? mem[917] : 
                       (N507)? mem[925] : 
                       (N509)? mem[933] : 
                       (N511)? mem[941] : 
                       (N513)? mem[949] : 
                       (N515)? mem[957] : 
                       (N517)? mem[965] : 
                       (N519)? mem[973] : 
                       (N521)? mem[981] : 
                       (N523)? mem[989] : 
                       (N525)? mem[997] : 
                       (N527)? mem[1005] : 
                       (N529)? mem[1013] : 
                       (N531)? mem[1021] : 
                       (N278)? mem[1029] : 
                       (N280)? mem[1037] : 
                       (N282)? mem[1045] : 
                       (N284)? mem[1053] : 
                       (N286)? mem[1061] : 
                       (N288)? mem[1069] : 
                       (N290)? mem[1077] : 
                       (N292)? mem[1085] : 
                       (N294)? mem[1093] : 
                       (N296)? mem[1101] : 
                       (N298)? mem[1109] : 
                       (N300)? mem[1117] : 
                       (N302)? mem[1125] : 
                       (N304)? mem[1133] : 
                       (N306)? mem[1141] : 
                       (N308)? mem[1149] : 
                       (N310)? mem[1157] : 
                       (N312)? mem[1165] : 
                       (N314)? mem[1173] : 
                       (N316)? mem[1181] : 
                       (N318)? mem[1189] : 
                       (N320)? mem[1197] : 
                       (N322)? mem[1205] : 
                       (N324)? mem[1213] : 
                       (N326)? mem[1221] : 
                       (N328)? mem[1229] : 
                       (N330)? mem[1237] : 
                       (N332)? mem[1245] : 
                       (N334)? mem[1253] : 
                       (N336)? mem[1261] : 
                       (N338)? mem[1269] : 
                       (N340)? mem[1277] : 
                       (N342)? mem[1285] : 
                       (N344)? mem[1293] : 
                       (N346)? mem[1301] : 
                       (N348)? mem[1309] : 
                       (N350)? mem[1317] : 
                       (N352)? mem[1325] : 
                       (N354)? mem[1333] : 
                       (N356)? mem[1341] : 
                       (N358)? mem[1349] : 
                       (N360)? mem[1357] : 
                       (N362)? mem[1365] : 
                       (N364)? mem[1373] : 
                       (N366)? mem[1381] : 
                       (N368)? mem[1389] : 
                       (N370)? mem[1397] : 
                       (N372)? mem[1405] : 
                       (N374)? mem[1413] : 
                       (N376)? mem[1421] : 
                       (N378)? mem[1429] : 
                       (N380)? mem[1437] : 
                       (N382)? mem[1445] : 
                       (N384)? mem[1453] : 
                       (N386)? mem[1461] : 
                       (N388)? mem[1469] : 
                       (N390)? mem[1477] : 
                       (N392)? mem[1485] : 
                       (N394)? mem[1493] : 
                       (N396)? mem[1501] : 
                       (N398)? mem[1509] : 
                       (N400)? mem[1517] : 
                       (N402)? mem[1525] : 
                       (N404)? mem[1533] : 
                       (N406)? mem[1541] : 
                       (N408)? mem[1549] : 
                       (N410)? mem[1557] : 
                       (N412)? mem[1565] : 
                       (N414)? mem[1573] : 
                       (N416)? mem[1581] : 
                       (N418)? mem[1589] : 
                       (N420)? mem[1597] : 
                       (N422)? mem[1605] : 
                       (N424)? mem[1613] : 
                       (N426)? mem[1621] : 
                       (N428)? mem[1629] : 
                       (N430)? mem[1637] : 
                       (N432)? mem[1645] : 
                       (N434)? mem[1653] : 
                       (N436)? mem[1661] : 
                       (N438)? mem[1669] : 
                       (N440)? mem[1677] : 
                       (N442)? mem[1685] : 
                       (N444)? mem[1693] : 
                       (N446)? mem[1701] : 
                       (N448)? mem[1709] : 
                       (N450)? mem[1717] : 
                       (N452)? mem[1725] : 
                       (N454)? mem[1733] : 
                       (N456)? mem[1741] : 
                       (N458)? mem[1749] : 
                       (N460)? mem[1757] : 
                       (N462)? mem[1765] : 
                       (N464)? mem[1773] : 
                       (N466)? mem[1781] : 
                       (N468)? mem[1789] : 
                       (N470)? mem[1797] : 
                       (N472)? mem[1805] : 
                       (N474)? mem[1813] : 
                       (N476)? mem[1821] : 
                       (N478)? mem[1829] : 
                       (N480)? mem[1837] : 
                       (N482)? mem[1845] : 
                       (N484)? mem[1853] : 
                       (N486)? mem[1861] : 
                       (N488)? mem[1869] : 
                       (N490)? mem[1877] : 
                       (N492)? mem[1885] : 
                       (N494)? mem[1893] : 
                       (N496)? mem[1901] : 
                       (N498)? mem[1909] : 
                       (N500)? mem[1917] : 
                       (N502)? mem[1925] : 
                       (N504)? mem[1933] : 
                       (N506)? mem[1941] : 
                       (N508)? mem[1949] : 
                       (N510)? mem[1957] : 
                       (N512)? mem[1965] : 
                       (N514)? mem[1973] : 
                       (N516)? mem[1981] : 
                       (N518)? mem[1989] : 
                       (N520)? mem[1997] : 
                       (N522)? mem[2005] : 
                       (N524)? mem[2013] : 
                       (N526)? mem[2021] : 
                       (N528)? mem[2029] : 
                       (N530)? mem[2037] : 
                       (N532)? mem[2045] : 1'b0;
  assign data_out[4] = (N277)? mem[4] : 
                       (N279)? mem[12] : 
                       (N281)? mem[20] : 
                       (N283)? mem[28] : 
                       (N285)? mem[36] : 
                       (N287)? mem[44] : 
                       (N289)? mem[52] : 
                       (N291)? mem[60] : 
                       (N293)? mem[68] : 
                       (N295)? mem[76] : 
                       (N297)? mem[84] : 
                       (N299)? mem[92] : 
                       (N301)? mem[100] : 
                       (N303)? mem[108] : 
                       (N305)? mem[116] : 
                       (N307)? mem[124] : 
                       (N309)? mem[132] : 
                       (N311)? mem[140] : 
                       (N313)? mem[148] : 
                       (N315)? mem[156] : 
                       (N317)? mem[164] : 
                       (N319)? mem[172] : 
                       (N321)? mem[180] : 
                       (N323)? mem[188] : 
                       (N325)? mem[196] : 
                       (N327)? mem[204] : 
                       (N329)? mem[212] : 
                       (N331)? mem[220] : 
                       (N333)? mem[228] : 
                       (N335)? mem[236] : 
                       (N337)? mem[244] : 
                       (N339)? mem[252] : 
                       (N341)? mem[260] : 
                       (N343)? mem[268] : 
                       (N345)? mem[276] : 
                       (N347)? mem[284] : 
                       (N349)? mem[292] : 
                       (N351)? mem[300] : 
                       (N353)? mem[308] : 
                       (N355)? mem[316] : 
                       (N357)? mem[324] : 
                       (N359)? mem[332] : 
                       (N361)? mem[340] : 
                       (N363)? mem[348] : 
                       (N365)? mem[356] : 
                       (N367)? mem[364] : 
                       (N369)? mem[372] : 
                       (N371)? mem[380] : 
                       (N373)? mem[388] : 
                       (N375)? mem[396] : 
                       (N377)? mem[404] : 
                       (N379)? mem[412] : 
                       (N381)? mem[420] : 
                       (N383)? mem[428] : 
                       (N385)? mem[436] : 
                       (N387)? mem[444] : 
                       (N389)? mem[452] : 
                       (N391)? mem[460] : 
                       (N393)? mem[468] : 
                       (N395)? mem[476] : 
                       (N397)? mem[484] : 
                       (N399)? mem[492] : 
                       (N401)? mem[500] : 
                       (N403)? mem[508] : 
                       (N405)? mem[516] : 
                       (N407)? mem[524] : 
                       (N409)? mem[532] : 
                       (N411)? mem[540] : 
                       (N413)? mem[548] : 
                       (N415)? mem[556] : 
                       (N417)? mem[564] : 
                       (N419)? mem[572] : 
                       (N421)? mem[580] : 
                       (N423)? mem[588] : 
                       (N425)? mem[596] : 
                       (N427)? mem[604] : 
                       (N429)? mem[612] : 
                       (N431)? mem[620] : 
                       (N433)? mem[628] : 
                       (N435)? mem[636] : 
                       (N437)? mem[644] : 
                       (N439)? mem[652] : 
                       (N441)? mem[660] : 
                       (N443)? mem[668] : 
                       (N445)? mem[676] : 
                       (N447)? mem[684] : 
                       (N449)? mem[692] : 
                       (N451)? mem[700] : 
                       (N453)? mem[708] : 
                       (N455)? mem[716] : 
                       (N457)? mem[724] : 
                       (N459)? mem[732] : 
                       (N461)? mem[740] : 
                       (N463)? mem[748] : 
                       (N465)? mem[756] : 
                       (N467)? mem[764] : 
                       (N469)? mem[772] : 
                       (N471)? mem[780] : 
                       (N473)? mem[788] : 
                       (N475)? mem[796] : 
                       (N477)? mem[804] : 
                       (N479)? mem[812] : 
                       (N481)? mem[820] : 
                       (N483)? mem[828] : 
                       (N485)? mem[836] : 
                       (N487)? mem[844] : 
                       (N489)? mem[852] : 
                       (N491)? mem[860] : 
                       (N493)? mem[868] : 
                       (N495)? mem[876] : 
                       (N497)? mem[884] : 
                       (N499)? mem[892] : 
                       (N501)? mem[900] : 
                       (N503)? mem[908] : 
                       (N505)? mem[916] : 
                       (N507)? mem[924] : 
                       (N509)? mem[932] : 
                       (N511)? mem[940] : 
                       (N513)? mem[948] : 
                       (N515)? mem[956] : 
                       (N517)? mem[964] : 
                       (N519)? mem[972] : 
                       (N521)? mem[980] : 
                       (N523)? mem[988] : 
                       (N525)? mem[996] : 
                       (N527)? mem[1004] : 
                       (N529)? mem[1012] : 
                       (N531)? mem[1020] : 
                       (N278)? mem[1028] : 
                       (N280)? mem[1036] : 
                       (N282)? mem[1044] : 
                       (N284)? mem[1052] : 
                       (N286)? mem[1060] : 
                       (N288)? mem[1068] : 
                       (N290)? mem[1076] : 
                       (N292)? mem[1084] : 
                       (N294)? mem[1092] : 
                       (N296)? mem[1100] : 
                       (N298)? mem[1108] : 
                       (N300)? mem[1116] : 
                       (N302)? mem[1124] : 
                       (N304)? mem[1132] : 
                       (N306)? mem[1140] : 
                       (N308)? mem[1148] : 
                       (N310)? mem[1156] : 
                       (N312)? mem[1164] : 
                       (N314)? mem[1172] : 
                       (N316)? mem[1180] : 
                       (N318)? mem[1188] : 
                       (N320)? mem[1196] : 
                       (N322)? mem[1204] : 
                       (N324)? mem[1212] : 
                       (N326)? mem[1220] : 
                       (N328)? mem[1228] : 
                       (N330)? mem[1236] : 
                       (N332)? mem[1244] : 
                       (N334)? mem[1252] : 
                       (N336)? mem[1260] : 
                       (N338)? mem[1268] : 
                       (N340)? mem[1276] : 
                       (N342)? mem[1284] : 
                       (N344)? mem[1292] : 
                       (N346)? mem[1300] : 
                       (N348)? mem[1308] : 
                       (N350)? mem[1316] : 
                       (N352)? mem[1324] : 
                       (N354)? mem[1332] : 
                       (N356)? mem[1340] : 
                       (N358)? mem[1348] : 
                       (N360)? mem[1356] : 
                       (N362)? mem[1364] : 
                       (N364)? mem[1372] : 
                       (N366)? mem[1380] : 
                       (N368)? mem[1388] : 
                       (N370)? mem[1396] : 
                       (N372)? mem[1404] : 
                       (N374)? mem[1412] : 
                       (N376)? mem[1420] : 
                       (N378)? mem[1428] : 
                       (N380)? mem[1436] : 
                       (N382)? mem[1444] : 
                       (N384)? mem[1452] : 
                       (N386)? mem[1460] : 
                       (N388)? mem[1468] : 
                       (N390)? mem[1476] : 
                       (N392)? mem[1484] : 
                       (N394)? mem[1492] : 
                       (N396)? mem[1500] : 
                       (N398)? mem[1508] : 
                       (N400)? mem[1516] : 
                       (N402)? mem[1524] : 
                       (N404)? mem[1532] : 
                       (N406)? mem[1540] : 
                       (N408)? mem[1548] : 
                       (N410)? mem[1556] : 
                       (N412)? mem[1564] : 
                       (N414)? mem[1572] : 
                       (N416)? mem[1580] : 
                       (N418)? mem[1588] : 
                       (N420)? mem[1596] : 
                       (N422)? mem[1604] : 
                       (N424)? mem[1612] : 
                       (N426)? mem[1620] : 
                       (N428)? mem[1628] : 
                       (N430)? mem[1636] : 
                       (N432)? mem[1644] : 
                       (N434)? mem[1652] : 
                       (N436)? mem[1660] : 
                       (N438)? mem[1668] : 
                       (N440)? mem[1676] : 
                       (N442)? mem[1684] : 
                       (N444)? mem[1692] : 
                       (N446)? mem[1700] : 
                       (N448)? mem[1708] : 
                       (N450)? mem[1716] : 
                       (N452)? mem[1724] : 
                       (N454)? mem[1732] : 
                       (N456)? mem[1740] : 
                       (N458)? mem[1748] : 
                       (N460)? mem[1756] : 
                       (N462)? mem[1764] : 
                       (N464)? mem[1772] : 
                       (N466)? mem[1780] : 
                       (N468)? mem[1788] : 
                       (N470)? mem[1796] : 
                       (N472)? mem[1804] : 
                       (N474)? mem[1812] : 
                       (N476)? mem[1820] : 
                       (N478)? mem[1828] : 
                       (N480)? mem[1836] : 
                       (N482)? mem[1844] : 
                       (N484)? mem[1852] : 
                       (N486)? mem[1860] : 
                       (N488)? mem[1868] : 
                       (N490)? mem[1876] : 
                       (N492)? mem[1884] : 
                       (N494)? mem[1892] : 
                       (N496)? mem[1900] : 
                       (N498)? mem[1908] : 
                       (N500)? mem[1916] : 
                       (N502)? mem[1924] : 
                       (N504)? mem[1932] : 
                       (N506)? mem[1940] : 
                       (N508)? mem[1948] : 
                       (N510)? mem[1956] : 
                       (N512)? mem[1964] : 
                       (N514)? mem[1972] : 
                       (N516)? mem[1980] : 
                       (N518)? mem[1988] : 
                       (N520)? mem[1996] : 
                       (N522)? mem[2004] : 
                       (N524)? mem[2012] : 
                       (N526)? mem[2020] : 
                       (N528)? mem[2028] : 
                       (N530)? mem[2036] : 
                       (N532)? mem[2044] : 1'b0;
  assign data_out[3] = (N277)? mem[3] : 
                       (N279)? mem[11] : 
                       (N281)? mem[19] : 
                       (N283)? mem[27] : 
                       (N285)? mem[35] : 
                       (N287)? mem[43] : 
                       (N289)? mem[51] : 
                       (N291)? mem[59] : 
                       (N293)? mem[67] : 
                       (N295)? mem[75] : 
                       (N297)? mem[83] : 
                       (N299)? mem[91] : 
                       (N301)? mem[99] : 
                       (N303)? mem[107] : 
                       (N305)? mem[115] : 
                       (N307)? mem[123] : 
                       (N309)? mem[131] : 
                       (N311)? mem[139] : 
                       (N313)? mem[147] : 
                       (N315)? mem[155] : 
                       (N317)? mem[163] : 
                       (N319)? mem[171] : 
                       (N321)? mem[179] : 
                       (N323)? mem[187] : 
                       (N325)? mem[195] : 
                       (N327)? mem[203] : 
                       (N329)? mem[211] : 
                       (N331)? mem[219] : 
                       (N333)? mem[227] : 
                       (N335)? mem[235] : 
                       (N337)? mem[243] : 
                       (N339)? mem[251] : 
                       (N341)? mem[259] : 
                       (N343)? mem[267] : 
                       (N345)? mem[275] : 
                       (N347)? mem[283] : 
                       (N349)? mem[291] : 
                       (N351)? mem[299] : 
                       (N353)? mem[307] : 
                       (N355)? mem[315] : 
                       (N357)? mem[323] : 
                       (N359)? mem[331] : 
                       (N361)? mem[339] : 
                       (N363)? mem[347] : 
                       (N365)? mem[355] : 
                       (N367)? mem[363] : 
                       (N369)? mem[371] : 
                       (N371)? mem[379] : 
                       (N373)? mem[387] : 
                       (N375)? mem[395] : 
                       (N377)? mem[403] : 
                       (N379)? mem[411] : 
                       (N381)? mem[419] : 
                       (N383)? mem[427] : 
                       (N385)? mem[435] : 
                       (N387)? mem[443] : 
                       (N389)? mem[451] : 
                       (N391)? mem[459] : 
                       (N393)? mem[467] : 
                       (N395)? mem[475] : 
                       (N397)? mem[483] : 
                       (N399)? mem[491] : 
                       (N401)? mem[499] : 
                       (N403)? mem[507] : 
                       (N405)? mem[515] : 
                       (N407)? mem[523] : 
                       (N409)? mem[531] : 
                       (N411)? mem[539] : 
                       (N413)? mem[547] : 
                       (N415)? mem[555] : 
                       (N417)? mem[563] : 
                       (N419)? mem[571] : 
                       (N421)? mem[579] : 
                       (N423)? mem[587] : 
                       (N425)? mem[595] : 
                       (N427)? mem[603] : 
                       (N429)? mem[611] : 
                       (N431)? mem[619] : 
                       (N433)? mem[627] : 
                       (N435)? mem[635] : 
                       (N437)? mem[643] : 
                       (N439)? mem[651] : 
                       (N441)? mem[659] : 
                       (N443)? mem[667] : 
                       (N445)? mem[675] : 
                       (N447)? mem[683] : 
                       (N449)? mem[691] : 
                       (N451)? mem[699] : 
                       (N453)? mem[707] : 
                       (N455)? mem[715] : 
                       (N457)? mem[723] : 
                       (N459)? mem[731] : 
                       (N461)? mem[739] : 
                       (N463)? mem[747] : 
                       (N465)? mem[755] : 
                       (N467)? mem[763] : 
                       (N469)? mem[771] : 
                       (N471)? mem[779] : 
                       (N473)? mem[787] : 
                       (N475)? mem[795] : 
                       (N477)? mem[803] : 
                       (N479)? mem[811] : 
                       (N481)? mem[819] : 
                       (N483)? mem[827] : 
                       (N485)? mem[835] : 
                       (N487)? mem[843] : 
                       (N489)? mem[851] : 
                       (N491)? mem[859] : 
                       (N493)? mem[867] : 
                       (N495)? mem[875] : 
                       (N497)? mem[883] : 
                       (N499)? mem[891] : 
                       (N501)? mem[899] : 
                       (N503)? mem[907] : 
                       (N505)? mem[915] : 
                       (N507)? mem[923] : 
                       (N509)? mem[931] : 
                       (N511)? mem[939] : 
                       (N513)? mem[947] : 
                       (N515)? mem[955] : 
                       (N517)? mem[963] : 
                       (N519)? mem[971] : 
                       (N521)? mem[979] : 
                       (N523)? mem[987] : 
                       (N525)? mem[995] : 
                       (N527)? mem[1003] : 
                       (N529)? mem[1011] : 
                       (N531)? mem[1019] : 
                       (N278)? mem[1027] : 
                       (N280)? mem[1035] : 
                       (N282)? mem[1043] : 
                       (N284)? mem[1051] : 
                       (N286)? mem[1059] : 
                       (N288)? mem[1067] : 
                       (N290)? mem[1075] : 
                       (N292)? mem[1083] : 
                       (N294)? mem[1091] : 
                       (N296)? mem[1099] : 
                       (N298)? mem[1107] : 
                       (N300)? mem[1115] : 
                       (N302)? mem[1123] : 
                       (N304)? mem[1131] : 
                       (N306)? mem[1139] : 
                       (N308)? mem[1147] : 
                       (N310)? mem[1155] : 
                       (N312)? mem[1163] : 
                       (N314)? mem[1171] : 
                       (N316)? mem[1179] : 
                       (N318)? mem[1187] : 
                       (N320)? mem[1195] : 
                       (N322)? mem[1203] : 
                       (N324)? mem[1211] : 
                       (N326)? mem[1219] : 
                       (N328)? mem[1227] : 
                       (N330)? mem[1235] : 
                       (N332)? mem[1243] : 
                       (N334)? mem[1251] : 
                       (N336)? mem[1259] : 
                       (N338)? mem[1267] : 
                       (N340)? mem[1275] : 
                       (N342)? mem[1283] : 
                       (N344)? mem[1291] : 
                       (N346)? mem[1299] : 
                       (N348)? mem[1307] : 
                       (N350)? mem[1315] : 
                       (N352)? mem[1323] : 
                       (N354)? mem[1331] : 
                       (N356)? mem[1339] : 
                       (N358)? mem[1347] : 
                       (N360)? mem[1355] : 
                       (N362)? mem[1363] : 
                       (N364)? mem[1371] : 
                       (N366)? mem[1379] : 
                       (N368)? mem[1387] : 
                       (N370)? mem[1395] : 
                       (N372)? mem[1403] : 
                       (N374)? mem[1411] : 
                       (N376)? mem[1419] : 
                       (N378)? mem[1427] : 
                       (N380)? mem[1435] : 
                       (N382)? mem[1443] : 
                       (N384)? mem[1451] : 
                       (N386)? mem[1459] : 
                       (N388)? mem[1467] : 
                       (N390)? mem[1475] : 
                       (N392)? mem[1483] : 
                       (N394)? mem[1491] : 
                       (N396)? mem[1499] : 
                       (N398)? mem[1507] : 
                       (N400)? mem[1515] : 
                       (N402)? mem[1523] : 
                       (N404)? mem[1531] : 
                       (N406)? mem[1539] : 
                       (N408)? mem[1547] : 
                       (N410)? mem[1555] : 
                       (N412)? mem[1563] : 
                       (N414)? mem[1571] : 
                       (N416)? mem[1579] : 
                       (N418)? mem[1587] : 
                       (N420)? mem[1595] : 
                       (N422)? mem[1603] : 
                       (N424)? mem[1611] : 
                       (N426)? mem[1619] : 
                       (N428)? mem[1627] : 
                       (N430)? mem[1635] : 
                       (N432)? mem[1643] : 
                       (N434)? mem[1651] : 
                       (N436)? mem[1659] : 
                       (N438)? mem[1667] : 
                       (N440)? mem[1675] : 
                       (N442)? mem[1683] : 
                       (N444)? mem[1691] : 
                       (N446)? mem[1699] : 
                       (N448)? mem[1707] : 
                       (N450)? mem[1715] : 
                       (N452)? mem[1723] : 
                       (N454)? mem[1731] : 
                       (N456)? mem[1739] : 
                       (N458)? mem[1747] : 
                       (N460)? mem[1755] : 
                       (N462)? mem[1763] : 
                       (N464)? mem[1771] : 
                       (N466)? mem[1779] : 
                       (N468)? mem[1787] : 
                       (N470)? mem[1795] : 
                       (N472)? mem[1803] : 
                       (N474)? mem[1811] : 
                       (N476)? mem[1819] : 
                       (N478)? mem[1827] : 
                       (N480)? mem[1835] : 
                       (N482)? mem[1843] : 
                       (N484)? mem[1851] : 
                       (N486)? mem[1859] : 
                       (N488)? mem[1867] : 
                       (N490)? mem[1875] : 
                       (N492)? mem[1883] : 
                       (N494)? mem[1891] : 
                       (N496)? mem[1899] : 
                       (N498)? mem[1907] : 
                       (N500)? mem[1915] : 
                       (N502)? mem[1923] : 
                       (N504)? mem[1931] : 
                       (N506)? mem[1939] : 
                       (N508)? mem[1947] : 
                       (N510)? mem[1955] : 
                       (N512)? mem[1963] : 
                       (N514)? mem[1971] : 
                       (N516)? mem[1979] : 
                       (N518)? mem[1987] : 
                       (N520)? mem[1995] : 
                       (N522)? mem[2003] : 
                       (N524)? mem[2011] : 
                       (N526)? mem[2019] : 
                       (N528)? mem[2027] : 
                       (N530)? mem[2035] : 
                       (N532)? mem[2043] : 1'b0;
  assign data_out[2] = (N277)? mem[2] : 
                       (N279)? mem[10] : 
                       (N281)? mem[18] : 
                       (N283)? mem[26] : 
                       (N285)? mem[34] : 
                       (N287)? mem[42] : 
                       (N289)? mem[50] : 
                       (N291)? mem[58] : 
                       (N293)? mem[66] : 
                       (N295)? mem[74] : 
                       (N297)? mem[82] : 
                       (N299)? mem[90] : 
                       (N301)? mem[98] : 
                       (N303)? mem[106] : 
                       (N305)? mem[114] : 
                       (N307)? mem[122] : 
                       (N309)? mem[130] : 
                       (N311)? mem[138] : 
                       (N313)? mem[146] : 
                       (N315)? mem[154] : 
                       (N317)? mem[162] : 
                       (N319)? mem[170] : 
                       (N321)? mem[178] : 
                       (N323)? mem[186] : 
                       (N325)? mem[194] : 
                       (N327)? mem[202] : 
                       (N329)? mem[210] : 
                       (N331)? mem[218] : 
                       (N333)? mem[226] : 
                       (N335)? mem[234] : 
                       (N337)? mem[242] : 
                       (N339)? mem[250] : 
                       (N341)? mem[258] : 
                       (N343)? mem[266] : 
                       (N345)? mem[274] : 
                       (N347)? mem[282] : 
                       (N349)? mem[290] : 
                       (N351)? mem[298] : 
                       (N353)? mem[306] : 
                       (N355)? mem[314] : 
                       (N357)? mem[322] : 
                       (N359)? mem[330] : 
                       (N361)? mem[338] : 
                       (N363)? mem[346] : 
                       (N365)? mem[354] : 
                       (N367)? mem[362] : 
                       (N369)? mem[370] : 
                       (N371)? mem[378] : 
                       (N373)? mem[386] : 
                       (N375)? mem[394] : 
                       (N377)? mem[402] : 
                       (N379)? mem[410] : 
                       (N381)? mem[418] : 
                       (N383)? mem[426] : 
                       (N385)? mem[434] : 
                       (N387)? mem[442] : 
                       (N389)? mem[450] : 
                       (N391)? mem[458] : 
                       (N393)? mem[466] : 
                       (N395)? mem[474] : 
                       (N397)? mem[482] : 
                       (N399)? mem[490] : 
                       (N401)? mem[498] : 
                       (N403)? mem[506] : 
                       (N405)? mem[514] : 
                       (N407)? mem[522] : 
                       (N409)? mem[530] : 
                       (N411)? mem[538] : 
                       (N413)? mem[546] : 
                       (N415)? mem[554] : 
                       (N417)? mem[562] : 
                       (N419)? mem[570] : 
                       (N421)? mem[578] : 
                       (N423)? mem[586] : 
                       (N425)? mem[594] : 
                       (N427)? mem[602] : 
                       (N429)? mem[610] : 
                       (N431)? mem[618] : 
                       (N433)? mem[626] : 
                       (N435)? mem[634] : 
                       (N437)? mem[642] : 
                       (N439)? mem[650] : 
                       (N441)? mem[658] : 
                       (N443)? mem[666] : 
                       (N445)? mem[674] : 
                       (N447)? mem[682] : 
                       (N449)? mem[690] : 
                       (N451)? mem[698] : 
                       (N453)? mem[706] : 
                       (N455)? mem[714] : 
                       (N457)? mem[722] : 
                       (N459)? mem[730] : 
                       (N461)? mem[738] : 
                       (N463)? mem[746] : 
                       (N465)? mem[754] : 
                       (N467)? mem[762] : 
                       (N469)? mem[770] : 
                       (N471)? mem[778] : 
                       (N473)? mem[786] : 
                       (N475)? mem[794] : 
                       (N477)? mem[802] : 
                       (N479)? mem[810] : 
                       (N481)? mem[818] : 
                       (N483)? mem[826] : 
                       (N485)? mem[834] : 
                       (N487)? mem[842] : 
                       (N489)? mem[850] : 
                       (N491)? mem[858] : 
                       (N493)? mem[866] : 
                       (N495)? mem[874] : 
                       (N497)? mem[882] : 
                       (N499)? mem[890] : 
                       (N501)? mem[898] : 
                       (N503)? mem[906] : 
                       (N505)? mem[914] : 
                       (N507)? mem[922] : 
                       (N509)? mem[930] : 
                       (N511)? mem[938] : 
                       (N513)? mem[946] : 
                       (N515)? mem[954] : 
                       (N517)? mem[962] : 
                       (N519)? mem[970] : 
                       (N521)? mem[978] : 
                       (N523)? mem[986] : 
                       (N525)? mem[994] : 
                       (N527)? mem[1002] : 
                       (N529)? mem[1010] : 
                       (N531)? mem[1018] : 
                       (N278)? mem[1026] : 
                       (N280)? mem[1034] : 
                       (N282)? mem[1042] : 
                       (N284)? mem[1050] : 
                       (N286)? mem[1058] : 
                       (N288)? mem[1066] : 
                       (N290)? mem[1074] : 
                       (N292)? mem[1082] : 
                       (N294)? mem[1090] : 
                       (N296)? mem[1098] : 
                       (N298)? mem[1106] : 
                       (N300)? mem[1114] : 
                       (N302)? mem[1122] : 
                       (N304)? mem[1130] : 
                       (N306)? mem[1138] : 
                       (N308)? mem[1146] : 
                       (N310)? mem[1154] : 
                       (N312)? mem[1162] : 
                       (N314)? mem[1170] : 
                       (N316)? mem[1178] : 
                       (N318)? mem[1186] : 
                       (N320)? mem[1194] : 
                       (N322)? mem[1202] : 
                       (N324)? mem[1210] : 
                       (N326)? mem[1218] : 
                       (N328)? mem[1226] : 
                       (N330)? mem[1234] : 
                       (N332)? mem[1242] : 
                       (N334)? mem[1250] : 
                       (N336)? mem[1258] : 
                       (N338)? mem[1266] : 
                       (N340)? mem[1274] : 
                       (N342)? mem[1282] : 
                       (N344)? mem[1290] : 
                       (N346)? mem[1298] : 
                       (N348)? mem[1306] : 
                       (N350)? mem[1314] : 
                       (N352)? mem[1322] : 
                       (N354)? mem[1330] : 
                       (N356)? mem[1338] : 
                       (N358)? mem[1346] : 
                       (N360)? mem[1354] : 
                       (N362)? mem[1362] : 
                       (N364)? mem[1370] : 
                       (N366)? mem[1378] : 
                       (N368)? mem[1386] : 
                       (N370)? mem[1394] : 
                       (N372)? mem[1402] : 
                       (N374)? mem[1410] : 
                       (N376)? mem[1418] : 
                       (N378)? mem[1426] : 
                       (N380)? mem[1434] : 
                       (N382)? mem[1442] : 
                       (N384)? mem[1450] : 
                       (N386)? mem[1458] : 
                       (N388)? mem[1466] : 
                       (N390)? mem[1474] : 
                       (N392)? mem[1482] : 
                       (N394)? mem[1490] : 
                       (N396)? mem[1498] : 
                       (N398)? mem[1506] : 
                       (N400)? mem[1514] : 
                       (N402)? mem[1522] : 
                       (N404)? mem[1530] : 
                       (N406)? mem[1538] : 
                       (N408)? mem[1546] : 
                       (N410)? mem[1554] : 
                       (N412)? mem[1562] : 
                       (N414)? mem[1570] : 
                       (N416)? mem[1578] : 
                       (N418)? mem[1586] : 
                       (N420)? mem[1594] : 
                       (N422)? mem[1602] : 
                       (N424)? mem[1610] : 
                       (N426)? mem[1618] : 
                       (N428)? mem[1626] : 
                       (N430)? mem[1634] : 
                       (N432)? mem[1642] : 
                       (N434)? mem[1650] : 
                       (N436)? mem[1658] : 
                       (N438)? mem[1666] : 
                       (N440)? mem[1674] : 
                       (N442)? mem[1682] : 
                       (N444)? mem[1690] : 
                       (N446)? mem[1698] : 
                       (N448)? mem[1706] : 
                       (N450)? mem[1714] : 
                       (N452)? mem[1722] : 
                       (N454)? mem[1730] : 
                       (N456)? mem[1738] : 
                       (N458)? mem[1746] : 
                       (N460)? mem[1754] : 
                       (N462)? mem[1762] : 
                       (N464)? mem[1770] : 
                       (N466)? mem[1778] : 
                       (N468)? mem[1786] : 
                       (N470)? mem[1794] : 
                       (N472)? mem[1802] : 
                       (N474)? mem[1810] : 
                       (N476)? mem[1818] : 
                       (N478)? mem[1826] : 
                       (N480)? mem[1834] : 
                       (N482)? mem[1842] : 
                       (N484)? mem[1850] : 
                       (N486)? mem[1858] : 
                       (N488)? mem[1866] : 
                       (N490)? mem[1874] : 
                       (N492)? mem[1882] : 
                       (N494)? mem[1890] : 
                       (N496)? mem[1898] : 
                       (N498)? mem[1906] : 
                       (N500)? mem[1914] : 
                       (N502)? mem[1922] : 
                       (N504)? mem[1930] : 
                       (N506)? mem[1938] : 
                       (N508)? mem[1946] : 
                       (N510)? mem[1954] : 
                       (N512)? mem[1962] : 
                       (N514)? mem[1970] : 
                       (N516)? mem[1978] : 
                       (N518)? mem[1986] : 
                       (N520)? mem[1994] : 
                       (N522)? mem[2002] : 
                       (N524)? mem[2010] : 
                       (N526)? mem[2018] : 
                       (N528)? mem[2026] : 
                       (N530)? mem[2034] : 
                       (N532)? mem[2042] : 1'b0;
  assign data_out[1] = (N277)? mem[1] : 
                       (N279)? mem[9] : 
                       (N281)? mem[17] : 
                       (N283)? mem[25] : 
                       (N285)? mem[33] : 
                       (N287)? mem[41] : 
                       (N289)? mem[49] : 
                       (N291)? mem[57] : 
                       (N293)? mem[65] : 
                       (N295)? mem[73] : 
                       (N297)? mem[81] : 
                       (N299)? mem[89] : 
                       (N301)? mem[97] : 
                       (N303)? mem[105] : 
                       (N305)? mem[113] : 
                       (N307)? mem[121] : 
                       (N309)? mem[129] : 
                       (N311)? mem[137] : 
                       (N313)? mem[145] : 
                       (N315)? mem[153] : 
                       (N317)? mem[161] : 
                       (N319)? mem[169] : 
                       (N321)? mem[177] : 
                       (N323)? mem[185] : 
                       (N325)? mem[193] : 
                       (N327)? mem[201] : 
                       (N329)? mem[209] : 
                       (N331)? mem[217] : 
                       (N333)? mem[225] : 
                       (N335)? mem[233] : 
                       (N337)? mem[241] : 
                       (N339)? mem[249] : 
                       (N341)? mem[257] : 
                       (N343)? mem[265] : 
                       (N345)? mem[273] : 
                       (N347)? mem[281] : 
                       (N349)? mem[289] : 
                       (N351)? mem[297] : 
                       (N353)? mem[305] : 
                       (N355)? mem[313] : 
                       (N357)? mem[321] : 
                       (N359)? mem[329] : 
                       (N361)? mem[337] : 
                       (N363)? mem[345] : 
                       (N365)? mem[353] : 
                       (N367)? mem[361] : 
                       (N369)? mem[369] : 
                       (N371)? mem[377] : 
                       (N373)? mem[385] : 
                       (N375)? mem[393] : 
                       (N377)? mem[401] : 
                       (N379)? mem[409] : 
                       (N381)? mem[417] : 
                       (N383)? mem[425] : 
                       (N385)? mem[433] : 
                       (N387)? mem[441] : 
                       (N389)? mem[449] : 
                       (N391)? mem[457] : 
                       (N393)? mem[465] : 
                       (N395)? mem[473] : 
                       (N397)? mem[481] : 
                       (N399)? mem[489] : 
                       (N401)? mem[497] : 
                       (N403)? mem[505] : 
                       (N405)? mem[513] : 
                       (N407)? mem[521] : 
                       (N409)? mem[529] : 
                       (N411)? mem[537] : 
                       (N413)? mem[545] : 
                       (N415)? mem[553] : 
                       (N417)? mem[561] : 
                       (N419)? mem[569] : 
                       (N421)? mem[577] : 
                       (N423)? mem[585] : 
                       (N425)? mem[593] : 
                       (N427)? mem[601] : 
                       (N429)? mem[609] : 
                       (N431)? mem[617] : 
                       (N433)? mem[625] : 
                       (N435)? mem[633] : 
                       (N437)? mem[641] : 
                       (N439)? mem[649] : 
                       (N441)? mem[657] : 
                       (N443)? mem[665] : 
                       (N445)? mem[673] : 
                       (N447)? mem[681] : 
                       (N449)? mem[689] : 
                       (N451)? mem[697] : 
                       (N453)? mem[705] : 
                       (N455)? mem[713] : 
                       (N457)? mem[721] : 
                       (N459)? mem[729] : 
                       (N461)? mem[737] : 
                       (N463)? mem[745] : 
                       (N465)? mem[753] : 
                       (N467)? mem[761] : 
                       (N469)? mem[769] : 
                       (N471)? mem[777] : 
                       (N473)? mem[785] : 
                       (N475)? mem[793] : 
                       (N477)? mem[801] : 
                       (N479)? mem[809] : 
                       (N481)? mem[817] : 
                       (N483)? mem[825] : 
                       (N485)? mem[833] : 
                       (N487)? mem[841] : 
                       (N489)? mem[849] : 
                       (N491)? mem[857] : 
                       (N493)? mem[865] : 
                       (N495)? mem[873] : 
                       (N497)? mem[881] : 
                       (N499)? mem[889] : 
                       (N501)? mem[897] : 
                       (N503)? mem[905] : 
                       (N505)? mem[913] : 
                       (N507)? mem[921] : 
                       (N509)? mem[929] : 
                       (N511)? mem[937] : 
                       (N513)? mem[945] : 
                       (N515)? mem[953] : 
                       (N517)? mem[961] : 
                       (N519)? mem[969] : 
                       (N521)? mem[977] : 
                       (N523)? mem[985] : 
                       (N525)? mem[993] : 
                       (N527)? mem[1001] : 
                       (N529)? mem[1009] : 
                       (N531)? mem[1017] : 
                       (N278)? mem[1025] : 
                       (N280)? mem[1033] : 
                       (N282)? mem[1041] : 
                       (N284)? mem[1049] : 
                       (N286)? mem[1057] : 
                       (N288)? mem[1065] : 
                       (N290)? mem[1073] : 
                       (N292)? mem[1081] : 
                       (N294)? mem[1089] : 
                       (N296)? mem[1097] : 
                       (N298)? mem[1105] : 
                       (N300)? mem[1113] : 
                       (N302)? mem[1121] : 
                       (N304)? mem[1129] : 
                       (N306)? mem[1137] : 
                       (N308)? mem[1145] : 
                       (N310)? mem[1153] : 
                       (N312)? mem[1161] : 
                       (N314)? mem[1169] : 
                       (N316)? mem[1177] : 
                       (N318)? mem[1185] : 
                       (N320)? mem[1193] : 
                       (N322)? mem[1201] : 
                       (N324)? mem[1209] : 
                       (N326)? mem[1217] : 
                       (N328)? mem[1225] : 
                       (N330)? mem[1233] : 
                       (N332)? mem[1241] : 
                       (N334)? mem[1249] : 
                       (N336)? mem[1257] : 
                       (N338)? mem[1265] : 
                       (N340)? mem[1273] : 
                       (N342)? mem[1281] : 
                       (N344)? mem[1289] : 
                       (N346)? mem[1297] : 
                       (N348)? mem[1305] : 
                       (N350)? mem[1313] : 
                       (N352)? mem[1321] : 
                       (N354)? mem[1329] : 
                       (N356)? mem[1337] : 
                       (N358)? mem[1345] : 
                       (N360)? mem[1353] : 
                       (N362)? mem[1361] : 
                       (N364)? mem[1369] : 
                       (N366)? mem[1377] : 
                       (N368)? mem[1385] : 
                       (N370)? mem[1393] : 
                       (N372)? mem[1401] : 
                       (N374)? mem[1409] : 
                       (N376)? mem[1417] : 
                       (N378)? mem[1425] : 
                       (N380)? mem[1433] : 
                       (N382)? mem[1441] : 
                       (N384)? mem[1449] : 
                       (N386)? mem[1457] : 
                       (N388)? mem[1465] : 
                       (N390)? mem[1473] : 
                       (N392)? mem[1481] : 
                       (N394)? mem[1489] : 
                       (N396)? mem[1497] : 
                       (N398)? mem[1505] : 
                       (N400)? mem[1513] : 
                       (N402)? mem[1521] : 
                       (N404)? mem[1529] : 
                       (N406)? mem[1537] : 
                       (N408)? mem[1545] : 
                       (N410)? mem[1553] : 
                       (N412)? mem[1561] : 
                       (N414)? mem[1569] : 
                       (N416)? mem[1577] : 
                       (N418)? mem[1585] : 
                       (N420)? mem[1593] : 
                       (N422)? mem[1601] : 
                       (N424)? mem[1609] : 
                       (N426)? mem[1617] : 
                       (N428)? mem[1625] : 
                       (N430)? mem[1633] : 
                       (N432)? mem[1641] : 
                       (N434)? mem[1649] : 
                       (N436)? mem[1657] : 
                       (N438)? mem[1665] : 
                       (N440)? mem[1673] : 
                       (N442)? mem[1681] : 
                       (N444)? mem[1689] : 
                       (N446)? mem[1697] : 
                       (N448)? mem[1705] : 
                       (N450)? mem[1713] : 
                       (N452)? mem[1721] : 
                       (N454)? mem[1729] : 
                       (N456)? mem[1737] : 
                       (N458)? mem[1745] : 
                       (N460)? mem[1753] : 
                       (N462)? mem[1761] : 
                       (N464)? mem[1769] : 
                       (N466)? mem[1777] : 
                       (N468)? mem[1785] : 
                       (N470)? mem[1793] : 
                       (N472)? mem[1801] : 
                       (N474)? mem[1809] : 
                       (N476)? mem[1817] : 
                       (N478)? mem[1825] : 
                       (N480)? mem[1833] : 
                       (N482)? mem[1841] : 
                       (N484)? mem[1849] : 
                       (N486)? mem[1857] : 
                       (N488)? mem[1865] : 
                       (N490)? mem[1873] : 
                       (N492)? mem[1881] : 
                       (N494)? mem[1889] : 
                       (N496)? mem[1897] : 
                       (N498)? mem[1905] : 
                       (N500)? mem[1913] : 
                       (N502)? mem[1921] : 
                       (N504)? mem[1929] : 
                       (N506)? mem[1937] : 
                       (N508)? mem[1945] : 
                       (N510)? mem[1953] : 
                       (N512)? mem[1961] : 
                       (N514)? mem[1969] : 
                       (N516)? mem[1977] : 
                       (N518)? mem[1985] : 
                       (N520)? mem[1993] : 
                       (N522)? mem[2001] : 
                       (N524)? mem[2009] : 
                       (N526)? mem[2017] : 
                       (N528)? mem[2025] : 
                       (N530)? mem[2033] : 
                       (N532)? mem[2041] : 1'b0;
  assign data_out[0] = (N277)? mem[0] : 
                       (N279)? mem[8] : 
                       (N281)? mem[16] : 
                       (N283)? mem[24] : 
                       (N285)? mem[32] : 
                       (N287)? mem[40] : 
                       (N289)? mem[48] : 
                       (N291)? mem[56] : 
                       (N293)? mem[64] : 
                       (N295)? mem[72] : 
                       (N297)? mem[80] : 
                       (N299)? mem[88] : 
                       (N301)? mem[96] : 
                       (N303)? mem[104] : 
                       (N305)? mem[112] : 
                       (N307)? mem[120] : 
                       (N309)? mem[128] : 
                       (N311)? mem[136] : 
                       (N313)? mem[144] : 
                       (N315)? mem[152] : 
                       (N317)? mem[160] : 
                       (N319)? mem[168] : 
                       (N321)? mem[176] : 
                       (N323)? mem[184] : 
                       (N325)? mem[192] : 
                       (N327)? mem[200] : 
                       (N329)? mem[208] : 
                       (N331)? mem[216] : 
                       (N333)? mem[224] : 
                       (N335)? mem[232] : 
                       (N337)? mem[240] : 
                       (N339)? mem[248] : 
                       (N341)? mem[256] : 
                       (N343)? mem[264] : 
                       (N345)? mem[272] : 
                       (N347)? mem[280] : 
                       (N349)? mem[288] : 
                       (N351)? mem[296] : 
                       (N353)? mem[304] : 
                       (N355)? mem[312] : 
                       (N357)? mem[320] : 
                       (N359)? mem[328] : 
                       (N361)? mem[336] : 
                       (N363)? mem[344] : 
                       (N365)? mem[352] : 
                       (N367)? mem[360] : 
                       (N369)? mem[368] : 
                       (N371)? mem[376] : 
                       (N373)? mem[384] : 
                       (N375)? mem[392] : 
                       (N377)? mem[400] : 
                       (N379)? mem[408] : 
                       (N381)? mem[416] : 
                       (N383)? mem[424] : 
                       (N385)? mem[432] : 
                       (N387)? mem[440] : 
                       (N389)? mem[448] : 
                       (N391)? mem[456] : 
                       (N393)? mem[464] : 
                       (N395)? mem[472] : 
                       (N397)? mem[480] : 
                       (N399)? mem[488] : 
                       (N401)? mem[496] : 
                       (N403)? mem[504] : 
                       (N405)? mem[512] : 
                       (N407)? mem[520] : 
                       (N409)? mem[528] : 
                       (N411)? mem[536] : 
                       (N413)? mem[544] : 
                       (N415)? mem[552] : 
                       (N417)? mem[560] : 
                       (N419)? mem[568] : 
                       (N421)? mem[576] : 
                       (N423)? mem[584] : 
                       (N425)? mem[592] : 
                       (N427)? mem[600] : 
                       (N429)? mem[608] : 
                       (N431)? mem[616] : 
                       (N433)? mem[624] : 
                       (N435)? mem[632] : 
                       (N437)? mem[640] : 
                       (N439)? mem[648] : 
                       (N441)? mem[656] : 
                       (N443)? mem[664] : 
                       (N445)? mem[672] : 
                       (N447)? mem[680] : 
                       (N449)? mem[688] : 
                       (N451)? mem[696] : 
                       (N453)? mem[704] : 
                       (N455)? mem[712] : 
                       (N457)? mem[720] : 
                       (N459)? mem[728] : 
                       (N461)? mem[736] : 
                       (N463)? mem[744] : 
                       (N465)? mem[752] : 
                       (N467)? mem[760] : 
                       (N469)? mem[768] : 
                       (N471)? mem[776] : 
                       (N473)? mem[784] : 
                       (N475)? mem[792] : 
                       (N477)? mem[800] : 
                       (N479)? mem[808] : 
                       (N481)? mem[816] : 
                       (N483)? mem[824] : 
                       (N485)? mem[832] : 
                       (N487)? mem[840] : 
                       (N489)? mem[848] : 
                       (N491)? mem[856] : 
                       (N493)? mem[864] : 
                       (N495)? mem[872] : 
                       (N497)? mem[880] : 
                       (N499)? mem[888] : 
                       (N501)? mem[896] : 
                       (N503)? mem[904] : 
                       (N505)? mem[912] : 
                       (N507)? mem[920] : 
                       (N509)? mem[928] : 
                       (N511)? mem[936] : 
                       (N513)? mem[944] : 
                       (N515)? mem[952] : 
                       (N517)? mem[960] : 
                       (N519)? mem[968] : 
                       (N521)? mem[976] : 
                       (N523)? mem[984] : 
                       (N525)? mem[992] : 
                       (N527)? mem[1000] : 
                       (N529)? mem[1008] : 
                       (N531)? mem[1016] : 
                       (N278)? mem[1024] : 
                       (N280)? mem[1032] : 
                       (N282)? mem[1040] : 
                       (N284)? mem[1048] : 
                       (N286)? mem[1056] : 
                       (N288)? mem[1064] : 
                       (N290)? mem[1072] : 
                       (N292)? mem[1080] : 
                       (N294)? mem[1088] : 
                       (N296)? mem[1096] : 
                       (N298)? mem[1104] : 
                       (N300)? mem[1112] : 
                       (N302)? mem[1120] : 
                       (N304)? mem[1128] : 
                       (N306)? mem[1136] : 
                       (N308)? mem[1144] : 
                       (N310)? mem[1152] : 
                       (N312)? mem[1160] : 
                       (N314)? mem[1168] : 
                       (N316)? mem[1176] : 
                       (N318)? mem[1184] : 
                       (N320)? mem[1192] : 
                       (N322)? mem[1200] : 
                       (N324)? mem[1208] : 
                       (N326)? mem[1216] : 
                       (N328)? mem[1224] : 
                       (N330)? mem[1232] : 
                       (N332)? mem[1240] : 
                       (N334)? mem[1248] : 
                       (N336)? mem[1256] : 
                       (N338)? mem[1264] : 
                       (N340)? mem[1272] : 
                       (N342)? mem[1280] : 
                       (N344)? mem[1288] : 
                       (N346)? mem[1296] : 
                       (N348)? mem[1304] : 
                       (N350)? mem[1312] : 
                       (N352)? mem[1320] : 
                       (N354)? mem[1328] : 
                       (N356)? mem[1336] : 
                       (N358)? mem[1344] : 
                       (N360)? mem[1352] : 
                       (N362)? mem[1360] : 
                       (N364)? mem[1368] : 
                       (N366)? mem[1376] : 
                       (N368)? mem[1384] : 
                       (N370)? mem[1392] : 
                       (N372)? mem[1400] : 
                       (N374)? mem[1408] : 
                       (N376)? mem[1416] : 
                       (N378)? mem[1424] : 
                       (N380)? mem[1432] : 
                       (N382)? mem[1440] : 
                       (N384)? mem[1448] : 
                       (N386)? mem[1456] : 
                       (N388)? mem[1464] : 
                       (N390)? mem[1472] : 
                       (N392)? mem[1480] : 
                       (N394)? mem[1488] : 
                       (N396)? mem[1496] : 
                       (N398)? mem[1504] : 
                       (N400)? mem[1512] : 
                       (N402)? mem[1520] : 
                       (N404)? mem[1528] : 
                       (N406)? mem[1536] : 
                       (N408)? mem[1544] : 
                       (N410)? mem[1552] : 
                       (N412)? mem[1560] : 
                       (N414)? mem[1568] : 
                       (N416)? mem[1576] : 
                       (N418)? mem[1584] : 
                       (N420)? mem[1592] : 
                       (N422)? mem[1600] : 
                       (N424)? mem[1608] : 
                       (N426)? mem[1616] : 
                       (N428)? mem[1624] : 
                       (N430)? mem[1632] : 
                       (N432)? mem[1640] : 
                       (N434)? mem[1648] : 
                       (N436)? mem[1656] : 
                       (N438)? mem[1664] : 
                       (N440)? mem[1672] : 
                       (N442)? mem[1680] : 
                       (N444)? mem[1688] : 
                       (N446)? mem[1696] : 
                       (N448)? mem[1704] : 
                       (N450)? mem[1712] : 
                       (N452)? mem[1720] : 
                       (N454)? mem[1728] : 
                       (N456)? mem[1736] : 
                       (N458)? mem[1744] : 
                       (N460)? mem[1752] : 
                       (N462)? mem[1760] : 
                       (N464)? mem[1768] : 
                       (N466)? mem[1776] : 
                       (N468)? mem[1784] : 
                       (N470)? mem[1792] : 
                       (N472)? mem[1800] : 
                       (N474)? mem[1808] : 
                       (N476)? mem[1816] : 
                       (N478)? mem[1824] : 
                       (N480)? mem[1832] : 
                       (N482)? mem[1840] : 
                       (N484)? mem[1848] : 
                       (N486)? mem[1856] : 
                       (N488)? mem[1864] : 
                       (N490)? mem[1872] : 
                       (N492)? mem[1880] : 
                       (N494)? mem[1888] : 
                       (N496)? mem[1896] : 
                       (N498)? mem[1904] : 
                       (N500)? mem[1912] : 
                       (N502)? mem[1920] : 
                       (N504)? mem[1928] : 
                       (N506)? mem[1936] : 
                       (N508)? mem[1944] : 
                       (N510)? mem[1952] : 
                       (N512)? mem[1960] : 
                       (N514)? mem[1968] : 
                       (N516)? mem[1976] : 
                       (N518)? mem[1984] : 
                       (N520)? mem[1992] : 
                       (N522)? mem[2000] : 
                       (N524)? mem[2008] : 
                       (N526)? mem[2016] : 
                       (N528)? mem[2024] : 
                       (N530)? mem[2032] : 
                       (N532)? mem[2040] : 1'b0;

  bsg_dff_width_p1
  llr_read_en_dff
  (
    .clk_i(clk_i),
    .data_i(read_en),
    .data_o(llr_read_en_r)
  );


  bsg_dff_en_bypass_width_p8
  llr_dff_bypass
  (
    .clk_i(clk_i),
    .en_i(llr_read_en_r),
    .data_i(data_out),
    .data_o(data_o)
  );

  assign N1047 = addr_i[6] & addr_i[7];
  assign N1048 = N0 & addr_i[7];
  assign N0 = ~addr_i[6];
  assign N1049 = addr_i[6] & N1;
  assign N1 = ~addr_i[7];
  assign N1050 = N2 & N3;
  assign N2 = ~addr_i[6];
  assign N3 = ~addr_i[7];
  assign N1051 = addr_i[4] & addr_i[5];
  assign N1052 = N4 & addr_i[5];
  assign N4 = ~addr_i[4];
  assign N1053 = addr_i[4] & N5;
  assign N5 = ~addr_i[5];
  assign N1054 = N6 & N7;
  assign N6 = ~addr_i[4];
  assign N7 = ~addr_i[5];
  assign N1055 = N1047 & N1051;
  assign N1056 = N1047 & N1052;
  assign N1057 = N1047 & N1053;
  assign N1058 = N1047 & N1054;
  assign N1059 = N1048 & N1051;
  assign N1060 = N1048 & N1052;
  assign N1061 = N1048 & N1053;
  assign N1062 = N1048 & N1054;
  assign N1063 = N1049 & N1051;
  assign N1064 = N1049 & N1052;
  assign N1065 = N1049 & N1053;
  assign N1066 = N1049 & N1054;
  assign N1067 = N1050 & N1051;
  assign N1068 = N1050 & N1052;
  assign N1069 = N1050 & N1053;
  assign N1070 = N1050 & N1054;
  assign N1071 = addr_i[2] & addr_i[3];
  assign N1072 = N8 & addr_i[3];
  assign N8 = ~addr_i[2];
  assign N1073 = addr_i[2] & N9;
  assign N9 = ~addr_i[3];
  assign N1074 = N10 & N11;
  assign N10 = ~addr_i[2];
  assign N11 = ~addr_i[3];
  assign N1075 = addr_i[0] & addr_i[1];
  assign N1076 = N12 & addr_i[1];
  assign N12 = ~addr_i[0];
  assign N1077 = addr_i[0] & N13;
  assign N13 = ~addr_i[1];
  assign N1078 = N14 & N15;
  assign N14 = ~addr_i[0];
  assign N15 = ~addr_i[1];
  assign N1079 = N1071 & N1075;
  assign N1080 = N1071 & N1076;
  assign N1081 = N1071 & N1077;
  assign N1082 = N1071 & N1078;
  assign N1083 = N1072 & N1075;
  assign N1084 = N1072 & N1076;
  assign N1085 = N1072 & N1077;
  assign N1086 = N1072 & N1078;
  assign N1087 = N1073 & N1075;
  assign N1088 = N1073 & N1076;
  assign N1089 = N1073 & N1077;
  assign N1090 = N1073 & N1078;
  assign N1091 = N1074 & N1075;
  assign N1092 = N1074 & N1076;
  assign N1093 = N1074 & N1077;
  assign N1094 = N1074 & N1078;
  assign N790 = N1055 & N1079;
  assign N789 = N1055 & N1080;
  assign N788 = N1055 & N1081;
  assign N787 = N1055 & N1082;
  assign N786 = N1055 & N1083;
  assign N785 = N1055 & N1084;
  assign N784 = N1055 & N1085;
  assign N783 = N1055 & N1086;
  assign N782 = N1055 & N1087;
  assign N781 = N1055 & N1088;
  assign N780 = N1055 & N1089;
  assign N779 = N1055 & N1090;
  assign N778 = N1055 & N1091;
  assign N777 = N1055 & N1092;
  assign N776 = N1055 & N1093;
  assign N775 = N1055 & N1094;
  assign N774 = N1056 & N1079;
  assign N773 = N1056 & N1080;
  assign N772 = N1056 & N1081;
  assign N771 = N1056 & N1082;
  assign N770 = N1056 & N1083;
  assign N769 = N1056 & N1084;
  assign N768 = N1056 & N1085;
  assign N767 = N1056 & N1086;
  assign N766 = N1056 & N1087;
  assign N765 = N1056 & N1088;
  assign N764 = N1056 & N1089;
  assign N763 = N1056 & N1090;
  assign N762 = N1056 & N1091;
  assign N761 = N1056 & N1092;
  assign N760 = N1056 & N1093;
  assign N759 = N1056 & N1094;
  assign N758 = N1057 & N1079;
  assign N757 = N1057 & N1080;
  assign N756 = N1057 & N1081;
  assign N755 = N1057 & N1082;
  assign N754 = N1057 & N1083;
  assign N753 = N1057 & N1084;
  assign N752 = N1057 & N1085;
  assign N751 = N1057 & N1086;
  assign N750 = N1057 & N1087;
  assign N749 = N1057 & N1088;
  assign N748 = N1057 & N1089;
  assign N747 = N1057 & N1090;
  assign N746 = N1057 & N1091;
  assign N745 = N1057 & N1092;
  assign N744 = N1057 & N1093;
  assign N743 = N1057 & N1094;
  assign N742 = N1058 & N1079;
  assign N741 = N1058 & N1080;
  assign N740 = N1058 & N1081;
  assign N739 = N1058 & N1082;
  assign N738 = N1058 & N1083;
  assign N737 = N1058 & N1084;
  assign N736 = N1058 & N1085;
  assign N735 = N1058 & N1086;
  assign N734 = N1058 & N1087;
  assign N733 = N1058 & N1088;
  assign N732 = N1058 & N1089;
  assign N731 = N1058 & N1090;
  assign N730 = N1058 & N1091;
  assign N729 = N1058 & N1092;
  assign N728 = N1058 & N1093;
  assign N727 = N1058 & N1094;
  assign N726 = N1059 & N1079;
  assign N725 = N1059 & N1080;
  assign N724 = N1059 & N1081;
  assign N723 = N1059 & N1082;
  assign N722 = N1059 & N1083;
  assign N721 = N1059 & N1084;
  assign N720 = N1059 & N1085;
  assign N719 = N1059 & N1086;
  assign N718 = N1059 & N1087;
  assign N717 = N1059 & N1088;
  assign N716 = N1059 & N1089;
  assign N715 = N1059 & N1090;
  assign N714 = N1059 & N1091;
  assign N713 = N1059 & N1092;
  assign N712 = N1059 & N1093;
  assign N711 = N1059 & N1094;
  assign N710 = N1060 & N1079;
  assign N709 = N1060 & N1080;
  assign N708 = N1060 & N1081;
  assign N707 = N1060 & N1082;
  assign N706 = N1060 & N1083;
  assign N705 = N1060 & N1084;
  assign N704 = N1060 & N1085;
  assign N703 = N1060 & N1086;
  assign N702 = N1060 & N1087;
  assign N701 = N1060 & N1088;
  assign N700 = N1060 & N1089;
  assign N699 = N1060 & N1090;
  assign N698 = N1060 & N1091;
  assign N697 = N1060 & N1092;
  assign N696 = N1060 & N1093;
  assign N695 = N1060 & N1094;
  assign N694 = N1061 & N1079;
  assign N693 = N1061 & N1080;
  assign N692 = N1061 & N1081;
  assign N691 = N1061 & N1082;
  assign N690 = N1061 & N1083;
  assign N689 = N1061 & N1084;
  assign N688 = N1061 & N1085;
  assign N687 = N1061 & N1086;
  assign N686 = N1061 & N1087;
  assign N685 = N1061 & N1088;
  assign N684 = N1061 & N1089;
  assign N683 = N1061 & N1090;
  assign N682 = N1061 & N1091;
  assign N681 = N1061 & N1092;
  assign N680 = N1061 & N1093;
  assign N679 = N1061 & N1094;
  assign N678 = N1062 & N1079;
  assign N677 = N1062 & N1080;
  assign N676 = N1062 & N1081;
  assign N675 = N1062 & N1082;
  assign N674 = N1062 & N1083;
  assign N673 = N1062 & N1084;
  assign N672 = N1062 & N1085;
  assign N671 = N1062 & N1086;
  assign N670 = N1062 & N1087;
  assign N669 = N1062 & N1088;
  assign N668 = N1062 & N1089;
  assign N667 = N1062 & N1090;
  assign N666 = N1062 & N1091;
  assign N665 = N1062 & N1092;
  assign N664 = N1062 & N1093;
  assign N663 = N1062 & N1094;
  assign N662 = N1063 & N1079;
  assign N661 = N1063 & N1080;
  assign N660 = N1063 & N1081;
  assign N659 = N1063 & N1082;
  assign N658 = N1063 & N1083;
  assign N657 = N1063 & N1084;
  assign N656 = N1063 & N1085;
  assign N655 = N1063 & N1086;
  assign N654 = N1063 & N1087;
  assign N653 = N1063 & N1088;
  assign N652 = N1063 & N1089;
  assign N651 = N1063 & N1090;
  assign N650 = N1063 & N1091;
  assign N649 = N1063 & N1092;
  assign N648 = N1063 & N1093;
  assign N647 = N1063 & N1094;
  assign N646 = N1064 & N1079;
  assign N645 = N1064 & N1080;
  assign N644 = N1064 & N1081;
  assign N643 = N1064 & N1082;
  assign N642 = N1064 & N1083;
  assign N641 = N1064 & N1084;
  assign N640 = N1064 & N1085;
  assign N639 = N1064 & N1086;
  assign N638 = N1064 & N1087;
  assign N637 = N1064 & N1088;
  assign N636 = N1064 & N1089;
  assign N635 = N1064 & N1090;
  assign N634 = N1064 & N1091;
  assign N633 = N1064 & N1092;
  assign N632 = N1064 & N1093;
  assign N631 = N1064 & N1094;
  assign N630 = N1065 & N1079;
  assign N629 = N1065 & N1080;
  assign N628 = N1065 & N1081;
  assign N627 = N1065 & N1082;
  assign N626 = N1065 & N1083;
  assign N625 = N1065 & N1084;
  assign N624 = N1065 & N1085;
  assign N623 = N1065 & N1086;
  assign N622 = N1065 & N1087;
  assign N621 = N1065 & N1088;
  assign N620 = N1065 & N1089;
  assign N619 = N1065 & N1090;
  assign N618 = N1065 & N1091;
  assign N617 = N1065 & N1092;
  assign N616 = N1065 & N1093;
  assign N615 = N1065 & N1094;
  assign N614 = N1066 & N1079;
  assign N613 = N1066 & N1080;
  assign N612 = N1066 & N1081;
  assign N611 = N1066 & N1082;
  assign N610 = N1066 & N1083;
  assign N609 = N1066 & N1084;
  assign N608 = N1066 & N1085;
  assign N607 = N1066 & N1086;
  assign N606 = N1066 & N1087;
  assign N605 = N1066 & N1088;
  assign N604 = N1066 & N1089;
  assign N603 = N1066 & N1090;
  assign N602 = N1066 & N1091;
  assign N601 = N1066 & N1092;
  assign N600 = N1066 & N1093;
  assign N599 = N1066 & N1094;
  assign N598 = N1067 & N1079;
  assign N597 = N1067 & N1080;
  assign N596 = N1067 & N1081;
  assign N595 = N1067 & N1082;
  assign N594 = N1067 & N1083;
  assign N593 = N1067 & N1084;
  assign N592 = N1067 & N1085;
  assign N591 = N1067 & N1086;
  assign N590 = N1067 & N1087;
  assign N589 = N1067 & N1088;
  assign N588 = N1067 & N1089;
  assign N587 = N1067 & N1090;
  assign N586 = N1067 & N1091;
  assign N585 = N1067 & N1092;
  assign N584 = N1067 & N1093;
  assign N583 = N1067 & N1094;
  assign N582 = N1068 & N1079;
  assign N581 = N1068 & N1080;
  assign N580 = N1068 & N1081;
  assign N579 = N1068 & N1082;
  assign N578 = N1068 & N1083;
  assign N577 = N1068 & N1084;
  assign N576 = N1068 & N1085;
  assign N575 = N1068 & N1086;
  assign N574 = N1068 & N1087;
  assign N573 = N1068 & N1088;
  assign N572 = N1068 & N1089;
  assign N571 = N1068 & N1090;
  assign N570 = N1068 & N1091;
  assign N569 = N1068 & N1092;
  assign N568 = N1068 & N1093;
  assign N567 = N1068 & N1094;
  assign N566 = N1069 & N1079;
  assign N565 = N1069 & N1080;
  assign N564 = N1069 & N1081;
  assign N563 = N1069 & N1082;
  assign N562 = N1069 & N1083;
  assign N561 = N1069 & N1084;
  assign N560 = N1069 & N1085;
  assign N559 = N1069 & N1086;
  assign N558 = N1069 & N1087;
  assign N557 = N1069 & N1088;
  assign N556 = N1069 & N1089;
  assign N555 = N1069 & N1090;
  assign N554 = N1069 & N1091;
  assign N553 = N1069 & N1092;
  assign N552 = N1069 & N1093;
  assign N551 = N1069 & N1094;
  assign N550 = N1070 & N1079;
  assign N549 = N1070 & N1080;
  assign N548 = N1070 & N1081;
  assign N547 = N1070 & N1082;
  assign N546 = N1070 & N1083;
  assign N545 = N1070 & N1084;
  assign N544 = N1070 & N1085;
  assign N543 = N1070 & N1086;
  assign N542 = N1070 & N1087;
  assign N541 = N1070 & N1088;
  assign N540 = N1070 & N1089;
  assign N539 = N1070 & N1090;
  assign N538 = N1070 & N1091;
  assign N537 = N1070 & N1092;
  assign N536 = N1070 & N1093;
  assign N535 = N1070 & N1094;
  assign { N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791 } = (N16)? { N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             (N534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N533;
  assign read_en = v_i & N1095;
  assign N1095 = ~w_i;
  assign N17 = ~addr_r[0];
  assign N18 = ~addr_r[1];
  assign N19 = N17 & N18;
  assign N20 = N17 & addr_r[1];
  assign N21 = addr_r[0] & N18;
  assign N22 = addr_r[0] & addr_r[1];
  assign N23 = ~addr_r[2];
  assign N24 = N19 & N23;
  assign N25 = N19 & addr_r[2];
  assign N26 = N21 & N23;
  assign N27 = N21 & addr_r[2];
  assign N28 = N20 & N23;
  assign N29 = N20 & addr_r[2];
  assign N30 = N22 & N23;
  assign N31 = N22 & addr_r[2];
  assign N32 = ~addr_r[3];
  assign N33 = N24 & N32;
  assign N34 = N24 & addr_r[3];
  assign N35 = N26 & N32;
  assign N36 = N26 & addr_r[3];
  assign N37 = N28 & N32;
  assign N38 = N28 & addr_r[3];
  assign N39 = N30 & N32;
  assign N40 = N30 & addr_r[3];
  assign N41 = N25 & N32;
  assign N42 = N25 & addr_r[3];
  assign N43 = N27 & N32;
  assign N44 = N27 & addr_r[3];
  assign N45 = N29 & N32;
  assign N46 = N29 & addr_r[3];
  assign N47 = N31 & N32;
  assign N48 = N31 & addr_r[3];
  assign N49 = ~addr_r[4];
  assign N50 = N33 & N49;
  assign N51 = N33 & addr_r[4];
  assign N52 = N35 & N49;
  assign N53 = N35 & addr_r[4];
  assign N54 = N37 & N49;
  assign N55 = N37 & addr_r[4];
  assign N56 = N39 & N49;
  assign N57 = N39 & addr_r[4];
  assign N58 = N41 & N49;
  assign N59 = N41 & addr_r[4];
  assign N60 = N43 & N49;
  assign N61 = N43 & addr_r[4];
  assign N62 = N45 & N49;
  assign N63 = N45 & addr_r[4];
  assign N64 = N47 & N49;
  assign N65 = N47 & addr_r[4];
  assign N66 = N34 & N49;
  assign N67 = N34 & addr_r[4];
  assign N68 = N36 & N49;
  assign N69 = N36 & addr_r[4];
  assign N70 = N38 & N49;
  assign N71 = N38 & addr_r[4];
  assign N72 = N40 & N49;
  assign N73 = N40 & addr_r[4];
  assign N74 = N42 & N49;
  assign N75 = N42 & addr_r[4];
  assign N76 = N44 & N49;
  assign N77 = N44 & addr_r[4];
  assign N78 = N46 & N49;
  assign N79 = N46 & addr_r[4];
  assign N80 = N48 & N49;
  assign N81 = N48 & addr_r[4];
  assign N82 = ~addr_r[5];
  assign N83 = N50 & N82;
  assign N84 = N50 & addr_r[5];
  assign N85 = N52 & N82;
  assign N86 = N52 & addr_r[5];
  assign N87 = N54 & N82;
  assign N88 = N54 & addr_r[5];
  assign N89 = N56 & N82;
  assign N90 = N56 & addr_r[5];
  assign N91 = N58 & N82;
  assign N92 = N58 & addr_r[5];
  assign N93 = N60 & N82;
  assign N94 = N60 & addr_r[5];
  assign N95 = N62 & N82;
  assign N96 = N62 & addr_r[5];
  assign N97 = N64 & N82;
  assign N98 = N64 & addr_r[5];
  assign N99 = N66 & N82;
  assign N100 = N66 & addr_r[5];
  assign N101 = N68 & N82;
  assign N102 = N68 & addr_r[5];
  assign N103 = N70 & N82;
  assign N104 = N70 & addr_r[5];
  assign N105 = N72 & N82;
  assign N106 = N72 & addr_r[5];
  assign N107 = N74 & N82;
  assign N108 = N74 & addr_r[5];
  assign N109 = N76 & N82;
  assign N110 = N76 & addr_r[5];
  assign N111 = N78 & N82;
  assign N112 = N78 & addr_r[5];
  assign N113 = N80 & N82;
  assign N114 = N80 & addr_r[5];
  assign N115 = N51 & N82;
  assign N116 = N51 & addr_r[5];
  assign N117 = N53 & N82;
  assign N118 = N53 & addr_r[5];
  assign N119 = N55 & N82;
  assign N120 = N55 & addr_r[5];
  assign N121 = N57 & N82;
  assign N122 = N57 & addr_r[5];
  assign N123 = N59 & N82;
  assign N124 = N59 & addr_r[5];
  assign N125 = N61 & N82;
  assign N126 = N61 & addr_r[5];
  assign N127 = N63 & N82;
  assign N128 = N63 & addr_r[5];
  assign N129 = N65 & N82;
  assign N130 = N65 & addr_r[5];
  assign N131 = N67 & N82;
  assign N132 = N67 & addr_r[5];
  assign N133 = N69 & N82;
  assign N134 = N69 & addr_r[5];
  assign N135 = N71 & N82;
  assign N136 = N71 & addr_r[5];
  assign N137 = N73 & N82;
  assign N138 = N73 & addr_r[5];
  assign N139 = N75 & N82;
  assign N140 = N75 & addr_r[5];
  assign N141 = N77 & N82;
  assign N142 = N77 & addr_r[5];
  assign N143 = N79 & N82;
  assign N144 = N79 & addr_r[5];
  assign N145 = N81 & N82;
  assign N146 = N81 & addr_r[5];
  assign N147 = ~addr_r[6];
  assign N148 = N83 & N147;
  assign N149 = N83 & addr_r[6];
  assign N150 = N85 & N147;
  assign N151 = N85 & addr_r[6];
  assign N152 = N87 & N147;
  assign N153 = N87 & addr_r[6];
  assign N154 = N89 & N147;
  assign N155 = N89 & addr_r[6];
  assign N156 = N91 & N147;
  assign N157 = N91 & addr_r[6];
  assign N158 = N93 & N147;
  assign N159 = N93 & addr_r[6];
  assign N160 = N95 & N147;
  assign N161 = N95 & addr_r[6];
  assign N162 = N97 & N147;
  assign N163 = N97 & addr_r[6];
  assign N164 = N99 & N147;
  assign N165 = N99 & addr_r[6];
  assign N166 = N101 & N147;
  assign N167 = N101 & addr_r[6];
  assign N168 = N103 & N147;
  assign N169 = N103 & addr_r[6];
  assign N170 = N105 & N147;
  assign N171 = N105 & addr_r[6];
  assign N172 = N107 & N147;
  assign N173 = N107 & addr_r[6];
  assign N174 = N109 & N147;
  assign N175 = N109 & addr_r[6];
  assign N176 = N111 & N147;
  assign N177 = N111 & addr_r[6];
  assign N178 = N113 & N147;
  assign N179 = N113 & addr_r[6];
  assign N180 = N115 & N147;
  assign N181 = N115 & addr_r[6];
  assign N182 = N117 & N147;
  assign N183 = N117 & addr_r[6];
  assign N184 = N119 & N147;
  assign N185 = N119 & addr_r[6];
  assign N186 = N121 & N147;
  assign N187 = N121 & addr_r[6];
  assign N188 = N123 & N147;
  assign N189 = N123 & addr_r[6];
  assign N190 = N125 & N147;
  assign N191 = N125 & addr_r[6];
  assign N192 = N127 & N147;
  assign N193 = N127 & addr_r[6];
  assign N194 = N129 & N147;
  assign N195 = N129 & addr_r[6];
  assign N196 = N131 & N147;
  assign N197 = N131 & addr_r[6];
  assign N198 = N133 & N147;
  assign N199 = N133 & addr_r[6];
  assign N200 = N135 & N147;
  assign N201 = N135 & addr_r[6];
  assign N202 = N137 & N147;
  assign N203 = N137 & addr_r[6];
  assign N204 = N139 & N147;
  assign N205 = N139 & addr_r[6];
  assign N206 = N141 & N147;
  assign N207 = N141 & addr_r[6];
  assign N208 = N143 & N147;
  assign N209 = N143 & addr_r[6];
  assign N210 = N145 & N147;
  assign N211 = N145 & addr_r[6];
  assign N212 = N84 & N147;
  assign N213 = N84 & addr_r[6];
  assign N214 = N86 & N147;
  assign N215 = N86 & addr_r[6];
  assign N216 = N88 & N147;
  assign N217 = N88 & addr_r[6];
  assign N218 = N90 & N147;
  assign N219 = N90 & addr_r[6];
  assign N220 = N92 & N147;
  assign N221 = N92 & addr_r[6];
  assign N222 = N94 & N147;
  assign N223 = N94 & addr_r[6];
  assign N224 = N96 & N147;
  assign N225 = N96 & addr_r[6];
  assign N226 = N98 & N147;
  assign N227 = N98 & addr_r[6];
  assign N228 = N100 & N147;
  assign N229 = N100 & addr_r[6];
  assign N230 = N102 & N147;
  assign N231 = N102 & addr_r[6];
  assign N232 = N104 & N147;
  assign N233 = N104 & addr_r[6];
  assign N234 = N106 & N147;
  assign N235 = N106 & addr_r[6];
  assign N236 = N108 & N147;
  assign N237 = N108 & addr_r[6];
  assign N238 = N110 & N147;
  assign N239 = N110 & addr_r[6];
  assign N240 = N112 & N147;
  assign N241 = N112 & addr_r[6];
  assign N242 = N114 & N147;
  assign N243 = N114 & addr_r[6];
  assign N244 = N116 & N147;
  assign N245 = N116 & addr_r[6];
  assign N246 = N118 & N147;
  assign N247 = N118 & addr_r[6];
  assign N248 = N120 & N147;
  assign N249 = N120 & addr_r[6];
  assign N250 = N122 & N147;
  assign N251 = N122 & addr_r[6];
  assign N252 = N124 & N147;
  assign N253 = N124 & addr_r[6];
  assign N254 = N126 & N147;
  assign N255 = N126 & addr_r[6];
  assign N256 = N128 & N147;
  assign N257 = N128 & addr_r[6];
  assign N258 = N130 & N147;
  assign N259 = N130 & addr_r[6];
  assign N260 = N132 & N147;
  assign N261 = N132 & addr_r[6];
  assign N262 = N134 & N147;
  assign N263 = N134 & addr_r[6];
  assign N264 = N136 & N147;
  assign N265 = N136 & addr_r[6];
  assign N266 = N138 & N147;
  assign N267 = N138 & addr_r[6];
  assign N268 = N140 & N147;
  assign N269 = N140 & addr_r[6];
  assign N270 = N142 & N147;
  assign N271 = N142 & addr_r[6];
  assign N272 = N144 & N147;
  assign N273 = N144 & addr_r[6];
  assign N274 = N146 & N147;
  assign N275 = N146 & addr_r[6];
  assign N276 = ~addr_r[7];
  assign N277 = N148 & N276;
  assign N278 = N148 & addr_r[7];
  assign N279 = N150 & N276;
  assign N280 = N150 & addr_r[7];
  assign N281 = N152 & N276;
  assign N282 = N152 & addr_r[7];
  assign N283 = N154 & N276;
  assign N284 = N154 & addr_r[7];
  assign N285 = N156 & N276;
  assign N286 = N156 & addr_r[7];
  assign N287 = N158 & N276;
  assign N288 = N158 & addr_r[7];
  assign N289 = N160 & N276;
  assign N290 = N160 & addr_r[7];
  assign N291 = N162 & N276;
  assign N292 = N162 & addr_r[7];
  assign N293 = N164 & N276;
  assign N294 = N164 & addr_r[7];
  assign N295 = N166 & N276;
  assign N296 = N166 & addr_r[7];
  assign N297 = N168 & N276;
  assign N298 = N168 & addr_r[7];
  assign N299 = N170 & N276;
  assign N300 = N170 & addr_r[7];
  assign N301 = N172 & N276;
  assign N302 = N172 & addr_r[7];
  assign N303 = N174 & N276;
  assign N304 = N174 & addr_r[7];
  assign N305 = N176 & N276;
  assign N306 = N176 & addr_r[7];
  assign N307 = N178 & N276;
  assign N308 = N178 & addr_r[7];
  assign N309 = N180 & N276;
  assign N310 = N180 & addr_r[7];
  assign N311 = N182 & N276;
  assign N312 = N182 & addr_r[7];
  assign N313 = N184 & N276;
  assign N314 = N184 & addr_r[7];
  assign N315 = N186 & N276;
  assign N316 = N186 & addr_r[7];
  assign N317 = N188 & N276;
  assign N318 = N188 & addr_r[7];
  assign N319 = N190 & N276;
  assign N320 = N190 & addr_r[7];
  assign N321 = N192 & N276;
  assign N322 = N192 & addr_r[7];
  assign N323 = N194 & N276;
  assign N324 = N194 & addr_r[7];
  assign N325 = N196 & N276;
  assign N326 = N196 & addr_r[7];
  assign N327 = N198 & N276;
  assign N328 = N198 & addr_r[7];
  assign N329 = N200 & N276;
  assign N330 = N200 & addr_r[7];
  assign N331 = N202 & N276;
  assign N332 = N202 & addr_r[7];
  assign N333 = N204 & N276;
  assign N334 = N204 & addr_r[7];
  assign N335 = N206 & N276;
  assign N336 = N206 & addr_r[7];
  assign N337 = N208 & N276;
  assign N338 = N208 & addr_r[7];
  assign N339 = N210 & N276;
  assign N340 = N210 & addr_r[7];
  assign N341 = N212 & N276;
  assign N342 = N212 & addr_r[7];
  assign N343 = N214 & N276;
  assign N344 = N214 & addr_r[7];
  assign N345 = N216 & N276;
  assign N346 = N216 & addr_r[7];
  assign N347 = N218 & N276;
  assign N348 = N218 & addr_r[7];
  assign N349 = N220 & N276;
  assign N350 = N220 & addr_r[7];
  assign N351 = N222 & N276;
  assign N352 = N222 & addr_r[7];
  assign N353 = N224 & N276;
  assign N354 = N224 & addr_r[7];
  assign N355 = N226 & N276;
  assign N356 = N226 & addr_r[7];
  assign N357 = N228 & N276;
  assign N358 = N228 & addr_r[7];
  assign N359 = N230 & N276;
  assign N360 = N230 & addr_r[7];
  assign N361 = N232 & N276;
  assign N362 = N232 & addr_r[7];
  assign N363 = N234 & N276;
  assign N364 = N234 & addr_r[7];
  assign N365 = N236 & N276;
  assign N366 = N236 & addr_r[7];
  assign N367 = N238 & N276;
  assign N368 = N238 & addr_r[7];
  assign N369 = N240 & N276;
  assign N370 = N240 & addr_r[7];
  assign N371 = N242 & N276;
  assign N372 = N242 & addr_r[7];
  assign N373 = N244 & N276;
  assign N374 = N244 & addr_r[7];
  assign N375 = N246 & N276;
  assign N376 = N246 & addr_r[7];
  assign N377 = N248 & N276;
  assign N378 = N248 & addr_r[7];
  assign N379 = N250 & N276;
  assign N380 = N250 & addr_r[7];
  assign N381 = N252 & N276;
  assign N382 = N252 & addr_r[7];
  assign N383 = N254 & N276;
  assign N384 = N254 & addr_r[7];
  assign N385 = N256 & N276;
  assign N386 = N256 & addr_r[7];
  assign N387 = N258 & N276;
  assign N388 = N258 & addr_r[7];
  assign N389 = N260 & N276;
  assign N390 = N260 & addr_r[7];
  assign N391 = N262 & N276;
  assign N392 = N262 & addr_r[7];
  assign N393 = N264 & N276;
  assign N394 = N264 & addr_r[7];
  assign N395 = N266 & N276;
  assign N396 = N266 & addr_r[7];
  assign N397 = N268 & N276;
  assign N398 = N268 & addr_r[7];
  assign N399 = N270 & N276;
  assign N400 = N270 & addr_r[7];
  assign N401 = N272 & N276;
  assign N402 = N272 & addr_r[7];
  assign N403 = N274 & N276;
  assign N404 = N274 & addr_r[7];
  assign N405 = N149 & N276;
  assign N406 = N149 & addr_r[7];
  assign N407 = N151 & N276;
  assign N408 = N151 & addr_r[7];
  assign N409 = N153 & N276;
  assign N410 = N153 & addr_r[7];
  assign N411 = N155 & N276;
  assign N412 = N155 & addr_r[7];
  assign N413 = N157 & N276;
  assign N414 = N157 & addr_r[7];
  assign N415 = N159 & N276;
  assign N416 = N159 & addr_r[7];
  assign N417 = N161 & N276;
  assign N418 = N161 & addr_r[7];
  assign N419 = N163 & N276;
  assign N420 = N163 & addr_r[7];
  assign N421 = N165 & N276;
  assign N422 = N165 & addr_r[7];
  assign N423 = N167 & N276;
  assign N424 = N167 & addr_r[7];
  assign N425 = N169 & N276;
  assign N426 = N169 & addr_r[7];
  assign N427 = N171 & N276;
  assign N428 = N171 & addr_r[7];
  assign N429 = N173 & N276;
  assign N430 = N173 & addr_r[7];
  assign N431 = N175 & N276;
  assign N432 = N175 & addr_r[7];
  assign N433 = N177 & N276;
  assign N434 = N177 & addr_r[7];
  assign N435 = N179 & N276;
  assign N436 = N179 & addr_r[7];
  assign N437 = N181 & N276;
  assign N438 = N181 & addr_r[7];
  assign N439 = N183 & N276;
  assign N440 = N183 & addr_r[7];
  assign N441 = N185 & N276;
  assign N442 = N185 & addr_r[7];
  assign N443 = N187 & N276;
  assign N444 = N187 & addr_r[7];
  assign N445 = N189 & N276;
  assign N446 = N189 & addr_r[7];
  assign N447 = N191 & N276;
  assign N448 = N191 & addr_r[7];
  assign N449 = N193 & N276;
  assign N450 = N193 & addr_r[7];
  assign N451 = N195 & N276;
  assign N452 = N195 & addr_r[7];
  assign N453 = N197 & N276;
  assign N454 = N197 & addr_r[7];
  assign N455 = N199 & N276;
  assign N456 = N199 & addr_r[7];
  assign N457 = N201 & N276;
  assign N458 = N201 & addr_r[7];
  assign N459 = N203 & N276;
  assign N460 = N203 & addr_r[7];
  assign N461 = N205 & N276;
  assign N462 = N205 & addr_r[7];
  assign N463 = N207 & N276;
  assign N464 = N207 & addr_r[7];
  assign N465 = N209 & N276;
  assign N466 = N209 & addr_r[7];
  assign N467 = N211 & N276;
  assign N468 = N211 & addr_r[7];
  assign N469 = N213 & N276;
  assign N470 = N213 & addr_r[7];
  assign N471 = N215 & N276;
  assign N472 = N215 & addr_r[7];
  assign N473 = N217 & N276;
  assign N474 = N217 & addr_r[7];
  assign N475 = N219 & N276;
  assign N476 = N219 & addr_r[7];
  assign N477 = N221 & N276;
  assign N478 = N221 & addr_r[7];
  assign N479 = N223 & N276;
  assign N480 = N223 & addr_r[7];
  assign N481 = N225 & N276;
  assign N482 = N225 & addr_r[7];
  assign N483 = N227 & N276;
  assign N484 = N227 & addr_r[7];
  assign N485 = N229 & N276;
  assign N486 = N229 & addr_r[7];
  assign N487 = N231 & N276;
  assign N488 = N231 & addr_r[7];
  assign N489 = N233 & N276;
  assign N490 = N233 & addr_r[7];
  assign N491 = N235 & N276;
  assign N492 = N235 & addr_r[7];
  assign N493 = N237 & N276;
  assign N494 = N237 & addr_r[7];
  assign N495 = N239 & N276;
  assign N496 = N239 & addr_r[7];
  assign N497 = N241 & N276;
  assign N498 = N241 & addr_r[7];
  assign N499 = N243 & N276;
  assign N500 = N243 & addr_r[7];
  assign N501 = N245 & N276;
  assign N502 = N245 & addr_r[7];
  assign N503 = N247 & N276;
  assign N504 = N247 & addr_r[7];
  assign N505 = N249 & N276;
  assign N506 = N249 & addr_r[7];
  assign N507 = N251 & N276;
  assign N508 = N251 & addr_r[7];
  assign N509 = N253 & N276;
  assign N510 = N253 & addr_r[7];
  assign N511 = N255 & N276;
  assign N512 = N255 & addr_r[7];
  assign N513 = N257 & N276;
  assign N514 = N257 & addr_r[7];
  assign N515 = N259 & N276;
  assign N516 = N259 & addr_r[7];
  assign N517 = N261 & N276;
  assign N518 = N261 & addr_r[7];
  assign N519 = N263 & N276;
  assign N520 = N263 & addr_r[7];
  assign N521 = N265 & N276;
  assign N522 = N265 & addr_r[7];
  assign N523 = N267 & N276;
  assign N524 = N267 & addr_r[7];
  assign N525 = N269 & N276;
  assign N526 = N269 & addr_r[7];
  assign N527 = N271 & N276;
  assign N528 = N271 & addr_r[7];
  assign N529 = N273 & N276;
  assign N530 = N273 & addr_r[7];
  assign N531 = N275 & N276;
  assign N532 = N275 & addr_r[7];
  assign N533 = v_i & w_i;
  assign N534 = ~N533;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { addr_r[7:0] } <= { addr_i[7:0] };
    end 
    if(N1046) begin
      { mem[2047:2040] } <= { data_i[7:0] };
    end 
    if(N1045) begin
      { mem[2039:2032] } <= { data_i[7:0] };
    end 
    if(N1044) begin
      { mem[2031:2024] } <= { data_i[7:0] };
    end 
    if(N1043) begin
      { mem[2023:2016] } <= { data_i[7:0] };
    end 
    if(N1042) begin
      { mem[2015:2008] } <= { data_i[7:0] };
    end 
    if(N1041) begin
      { mem[2007:2000] } <= { data_i[7:0] };
    end 
    if(N1040) begin
      { mem[1999:1992] } <= { data_i[7:0] };
    end 
    if(N1039) begin
      { mem[1991:1984] } <= { data_i[7:0] };
    end 
    if(N1038) begin
      { mem[1983:1976] } <= { data_i[7:0] };
    end 
    if(N1037) begin
      { mem[1975:1968] } <= { data_i[7:0] };
    end 
    if(N1036) begin
      { mem[1967:1960] } <= { data_i[7:0] };
    end 
    if(N1035) begin
      { mem[1959:1952] } <= { data_i[7:0] };
    end 
    if(N1034) begin
      { mem[1951:1944] } <= { data_i[7:0] };
    end 
    if(N1033) begin
      { mem[1943:1936] } <= { data_i[7:0] };
    end 
    if(N1032) begin
      { mem[1935:1928] } <= { data_i[7:0] };
    end 
    if(N1031) begin
      { mem[1927:1920] } <= { data_i[7:0] };
    end 
    if(N1030) begin
      { mem[1919:1912] } <= { data_i[7:0] };
    end 
    if(N1029) begin
      { mem[1911:1904] } <= { data_i[7:0] };
    end 
    if(N1028) begin
      { mem[1903:1896] } <= { data_i[7:0] };
    end 
    if(N1027) begin
      { mem[1895:1888] } <= { data_i[7:0] };
    end 
    if(N1026) begin
      { mem[1887:1880] } <= { data_i[7:0] };
    end 
    if(N1025) begin
      { mem[1879:1872] } <= { data_i[7:0] };
    end 
    if(N1024) begin
      { mem[1871:1864] } <= { data_i[7:0] };
    end 
    if(N1023) begin
      { mem[1863:1856] } <= { data_i[7:0] };
    end 
    if(N1022) begin
      { mem[1855:1848] } <= { data_i[7:0] };
    end 
    if(N1021) begin
      { mem[1847:1840] } <= { data_i[7:0] };
    end 
    if(N1020) begin
      { mem[1839:1832] } <= { data_i[7:0] };
    end 
    if(N1019) begin
      { mem[1831:1824] } <= { data_i[7:0] };
    end 
    if(N1018) begin
      { mem[1823:1816] } <= { data_i[7:0] };
    end 
    if(N1017) begin
      { mem[1815:1808] } <= { data_i[7:0] };
    end 
    if(N1016) begin
      { mem[1807:1800] } <= { data_i[7:0] };
    end 
    if(N1015) begin
      { mem[1799:1792] } <= { data_i[7:0] };
    end 
    if(N1014) begin
      { mem[1791:1784] } <= { data_i[7:0] };
    end 
    if(N1013) begin
      { mem[1783:1776] } <= { data_i[7:0] };
    end 
    if(N1012) begin
      { mem[1775:1768] } <= { data_i[7:0] };
    end 
    if(N1011) begin
      { mem[1767:1760] } <= { data_i[7:0] };
    end 
    if(N1010) begin
      { mem[1759:1752] } <= { data_i[7:0] };
    end 
    if(N1009) begin
      { mem[1751:1744] } <= { data_i[7:0] };
    end 
    if(N1008) begin
      { mem[1743:1736] } <= { data_i[7:0] };
    end 
    if(N1007) begin
      { mem[1735:1728] } <= { data_i[7:0] };
    end 
    if(N1006) begin
      { mem[1727:1720] } <= { data_i[7:0] };
    end 
    if(N1005) begin
      { mem[1719:1712] } <= { data_i[7:0] };
    end 
    if(N1004) begin
      { mem[1711:1704] } <= { data_i[7:0] };
    end 
    if(N1003) begin
      { mem[1703:1696] } <= { data_i[7:0] };
    end 
    if(N1002) begin
      { mem[1695:1688] } <= { data_i[7:0] };
    end 
    if(N1001) begin
      { mem[1687:1680] } <= { data_i[7:0] };
    end 
    if(N1000) begin
      { mem[1679:1672] } <= { data_i[7:0] };
    end 
    if(N999) begin
      { mem[1671:1664] } <= { data_i[7:0] };
    end 
    if(N998) begin
      { mem[1663:1656] } <= { data_i[7:0] };
    end 
    if(N997) begin
      { mem[1655:1648] } <= { data_i[7:0] };
    end 
    if(N996) begin
      { mem[1647:1640] } <= { data_i[7:0] };
    end 
    if(N995) begin
      { mem[1639:1632] } <= { data_i[7:0] };
    end 
    if(N994) begin
      { mem[1631:1624] } <= { data_i[7:0] };
    end 
    if(N993) begin
      { mem[1623:1616] } <= { data_i[7:0] };
    end 
    if(N992) begin
      { mem[1615:1608] } <= { data_i[7:0] };
    end 
    if(N991) begin
      { mem[1607:1600] } <= { data_i[7:0] };
    end 
    if(N990) begin
      { mem[1599:1592] } <= { data_i[7:0] };
    end 
    if(N989) begin
      { mem[1591:1584] } <= { data_i[7:0] };
    end 
    if(N988) begin
      { mem[1583:1576] } <= { data_i[7:0] };
    end 
    if(N987) begin
      { mem[1575:1568] } <= { data_i[7:0] };
    end 
    if(N986) begin
      { mem[1567:1560] } <= { data_i[7:0] };
    end 
    if(N985) begin
      { mem[1559:1552] } <= { data_i[7:0] };
    end 
    if(N984) begin
      { mem[1551:1544] } <= { data_i[7:0] };
    end 
    if(N983) begin
      { mem[1543:1536] } <= { data_i[7:0] };
    end 
    if(N982) begin
      { mem[1535:1528] } <= { data_i[7:0] };
    end 
    if(N981) begin
      { mem[1527:1520] } <= { data_i[7:0] };
    end 
    if(N980) begin
      { mem[1519:1512] } <= { data_i[7:0] };
    end 
    if(N979) begin
      { mem[1511:1504] } <= { data_i[7:0] };
    end 
    if(N978) begin
      { mem[1503:1496] } <= { data_i[7:0] };
    end 
    if(N977) begin
      { mem[1495:1488] } <= { data_i[7:0] };
    end 
    if(N976) begin
      { mem[1487:1480] } <= { data_i[7:0] };
    end 
    if(N975) begin
      { mem[1479:1472] } <= { data_i[7:0] };
    end 
    if(N974) begin
      { mem[1471:1464] } <= { data_i[7:0] };
    end 
    if(N973) begin
      { mem[1463:1456] } <= { data_i[7:0] };
    end 
    if(N972) begin
      { mem[1455:1448] } <= { data_i[7:0] };
    end 
    if(N971) begin
      { mem[1447:1440] } <= { data_i[7:0] };
    end 
    if(N970) begin
      { mem[1439:1432] } <= { data_i[7:0] };
    end 
    if(N969) begin
      { mem[1431:1424] } <= { data_i[7:0] };
    end 
    if(N968) begin
      { mem[1423:1416] } <= { data_i[7:0] };
    end 
    if(N967) begin
      { mem[1415:1408] } <= { data_i[7:0] };
    end 
    if(N966) begin
      { mem[1407:1400] } <= { data_i[7:0] };
    end 
    if(N965) begin
      { mem[1399:1392] } <= { data_i[7:0] };
    end 
    if(N964) begin
      { mem[1391:1384] } <= { data_i[7:0] };
    end 
    if(N963) begin
      { mem[1383:1376] } <= { data_i[7:0] };
    end 
    if(N962) begin
      { mem[1375:1368] } <= { data_i[7:0] };
    end 
    if(N961) begin
      { mem[1367:1360] } <= { data_i[7:0] };
    end 
    if(N960) begin
      { mem[1359:1352] } <= { data_i[7:0] };
    end 
    if(N959) begin
      { mem[1351:1344] } <= { data_i[7:0] };
    end 
    if(N958) begin
      { mem[1343:1336] } <= { data_i[7:0] };
    end 
    if(N957) begin
      { mem[1335:1328] } <= { data_i[7:0] };
    end 
    if(N956) begin
      { mem[1327:1320] } <= { data_i[7:0] };
    end 
    if(N955) begin
      { mem[1319:1312] } <= { data_i[7:0] };
    end 
    if(N954) begin
      { mem[1311:1304] } <= { data_i[7:0] };
    end 
    if(N953) begin
      { mem[1303:1296] } <= { data_i[7:0] };
    end 
    if(N952) begin
      { mem[1295:1288] } <= { data_i[7:0] };
    end 
    if(N951) begin
      { mem[1287:1280] } <= { data_i[7:0] };
    end 
    if(N950) begin
      { mem[1279:1272] } <= { data_i[7:0] };
    end 
    if(N949) begin
      { mem[1271:1264] } <= { data_i[7:0] };
    end 
    if(N948) begin
      { mem[1263:1256] } <= { data_i[7:0] };
    end 
    if(N947) begin
      { mem[1255:1248] } <= { data_i[7:0] };
    end 
    if(N946) begin
      { mem[1247:1240] } <= { data_i[7:0] };
    end 
    if(N945) begin
      { mem[1239:1232] } <= { data_i[7:0] };
    end 
    if(N944) begin
      { mem[1231:1224] } <= { data_i[7:0] };
    end 
    if(N943) begin
      { mem[1223:1216] } <= { data_i[7:0] };
    end 
    if(N942) begin
      { mem[1215:1208] } <= { data_i[7:0] };
    end 
    if(N941) begin
      { mem[1207:1200] } <= { data_i[7:0] };
    end 
    if(N940) begin
      { mem[1199:1192] } <= { data_i[7:0] };
    end 
    if(N939) begin
      { mem[1191:1184] } <= { data_i[7:0] };
    end 
    if(N938) begin
      { mem[1183:1176] } <= { data_i[7:0] };
    end 
    if(N937) begin
      { mem[1175:1168] } <= { data_i[7:0] };
    end 
    if(N936) begin
      { mem[1167:1160] } <= { data_i[7:0] };
    end 
    if(N935) begin
      { mem[1159:1152] } <= { data_i[7:0] };
    end 
    if(N934) begin
      { mem[1151:1144] } <= { data_i[7:0] };
    end 
    if(N933) begin
      { mem[1143:1136] } <= { data_i[7:0] };
    end 
    if(N932) begin
      { mem[1135:1128] } <= { data_i[7:0] };
    end 
    if(N931) begin
      { mem[1127:1120] } <= { data_i[7:0] };
    end 
    if(N930) begin
      { mem[1119:1112] } <= { data_i[7:0] };
    end 
    if(N929) begin
      { mem[1111:1104] } <= { data_i[7:0] };
    end 
    if(N928) begin
      { mem[1103:1096] } <= { data_i[7:0] };
    end 
    if(N927) begin
      { mem[1095:1088] } <= { data_i[7:0] };
    end 
    if(N926) begin
      { mem[1087:1080] } <= { data_i[7:0] };
    end 
    if(N925) begin
      { mem[1079:1072] } <= { data_i[7:0] };
    end 
    if(N924) begin
      { mem[1071:1064] } <= { data_i[7:0] };
    end 
    if(N923) begin
      { mem[1063:1056] } <= { data_i[7:0] };
    end 
    if(N922) begin
      { mem[1055:1048] } <= { data_i[7:0] };
    end 
    if(N921) begin
      { mem[1047:1040] } <= { data_i[7:0] };
    end 
    if(N920) begin
      { mem[1039:1032] } <= { data_i[7:0] };
    end 
    if(N919) begin
      { mem[1031:1024] } <= { data_i[7:0] };
    end 
    if(N918) begin
      { mem[1023:1016] } <= { data_i[7:0] };
    end 
    if(N917) begin
      { mem[1015:1008] } <= { data_i[7:0] };
    end 
    if(N916) begin
      { mem[1007:1000] } <= { data_i[7:0] };
    end 
    if(N915) begin
      { mem[999:992] } <= { data_i[7:0] };
    end 
    if(N914) begin
      { mem[991:984] } <= { data_i[7:0] };
    end 
    if(N913) begin
      { mem[983:976] } <= { data_i[7:0] };
    end 
    if(N912) begin
      { mem[975:968] } <= { data_i[7:0] };
    end 
    if(N911) begin
      { mem[967:960] } <= { data_i[7:0] };
    end 
    if(N910) begin
      { mem[959:952] } <= { data_i[7:0] };
    end 
    if(N909) begin
      { mem[951:944] } <= { data_i[7:0] };
    end 
    if(N908) begin
      { mem[943:936] } <= { data_i[7:0] };
    end 
    if(N907) begin
      { mem[935:928] } <= { data_i[7:0] };
    end 
    if(N906) begin
      { mem[927:920] } <= { data_i[7:0] };
    end 
    if(N905) begin
      { mem[919:912] } <= { data_i[7:0] };
    end 
    if(N904) begin
      { mem[911:904] } <= { data_i[7:0] };
    end 
    if(N903) begin
      { mem[903:896] } <= { data_i[7:0] };
    end 
    if(N902) begin
      { mem[895:888] } <= { data_i[7:0] };
    end 
    if(N901) begin
      { mem[887:880] } <= { data_i[7:0] };
    end 
    if(N900) begin
      { mem[879:872] } <= { data_i[7:0] };
    end 
    if(N899) begin
      { mem[871:864] } <= { data_i[7:0] };
    end 
    if(N898) begin
      { mem[863:856] } <= { data_i[7:0] };
    end 
    if(N897) begin
      { mem[855:848] } <= { data_i[7:0] };
    end 
    if(N896) begin
      { mem[847:840] } <= { data_i[7:0] };
    end 
    if(N895) begin
      { mem[839:832] } <= { data_i[7:0] };
    end 
    if(N894) begin
      { mem[831:824] } <= { data_i[7:0] };
    end 
    if(N893) begin
      { mem[823:816] } <= { data_i[7:0] };
    end 
    if(N892) begin
      { mem[815:808] } <= { data_i[7:0] };
    end 
    if(N891) begin
      { mem[807:800] } <= { data_i[7:0] };
    end 
    if(N890) begin
      { mem[799:792] } <= { data_i[7:0] };
    end 
    if(N889) begin
      { mem[791:784] } <= { data_i[7:0] };
    end 
    if(N888) begin
      { mem[783:776] } <= { data_i[7:0] };
    end 
    if(N887) begin
      { mem[775:768] } <= { data_i[7:0] };
    end 
    if(N886) begin
      { mem[767:760] } <= { data_i[7:0] };
    end 
    if(N885) begin
      { mem[759:752] } <= { data_i[7:0] };
    end 
    if(N884) begin
      { mem[751:744] } <= { data_i[7:0] };
    end 
    if(N883) begin
      { mem[743:736] } <= { data_i[7:0] };
    end 
    if(N882) begin
      { mem[735:728] } <= { data_i[7:0] };
    end 
    if(N881) begin
      { mem[727:720] } <= { data_i[7:0] };
    end 
    if(N880) begin
      { mem[719:712] } <= { data_i[7:0] };
    end 
    if(N879) begin
      { mem[711:704] } <= { data_i[7:0] };
    end 
    if(N878) begin
      { mem[703:696] } <= { data_i[7:0] };
    end 
    if(N877) begin
      { mem[695:688] } <= { data_i[7:0] };
    end 
    if(N876) begin
      { mem[687:680] } <= { data_i[7:0] };
    end 
    if(N875) begin
      { mem[679:672] } <= { data_i[7:0] };
    end 
    if(N874) begin
      { mem[671:664] } <= { data_i[7:0] };
    end 
    if(N873) begin
      { mem[663:656] } <= { data_i[7:0] };
    end 
    if(N872) begin
      { mem[655:648] } <= { data_i[7:0] };
    end 
    if(N871) begin
      { mem[647:640] } <= { data_i[7:0] };
    end 
    if(N870) begin
      { mem[639:632] } <= { data_i[7:0] };
    end 
    if(N869) begin
      { mem[631:624] } <= { data_i[7:0] };
    end 
    if(N868) begin
      { mem[623:616] } <= { data_i[7:0] };
    end 
    if(N867) begin
      { mem[615:608] } <= { data_i[7:0] };
    end 
    if(N866) begin
      { mem[607:600] } <= { data_i[7:0] };
    end 
    if(N865) begin
      { mem[599:592] } <= { data_i[7:0] };
    end 
    if(N864) begin
      { mem[591:584] } <= { data_i[7:0] };
    end 
    if(N863) begin
      { mem[583:576] } <= { data_i[7:0] };
    end 
    if(N862) begin
      { mem[575:568] } <= { data_i[7:0] };
    end 
    if(N861) begin
      { mem[567:560] } <= { data_i[7:0] };
    end 
    if(N860) begin
      { mem[559:552] } <= { data_i[7:0] };
    end 
    if(N859) begin
      { mem[551:544] } <= { data_i[7:0] };
    end 
    if(N858) begin
      { mem[543:536] } <= { data_i[7:0] };
    end 
    if(N857) begin
      { mem[535:528] } <= { data_i[7:0] };
    end 
    if(N856) begin
      { mem[527:520] } <= { data_i[7:0] };
    end 
    if(N855) begin
      { mem[519:512] } <= { data_i[7:0] };
    end 
    if(N854) begin
      { mem[511:504] } <= { data_i[7:0] };
    end 
    if(N853) begin
      { mem[503:496] } <= { data_i[7:0] };
    end 
    if(N852) begin
      { mem[495:488] } <= { data_i[7:0] };
    end 
    if(N851) begin
      { mem[487:480] } <= { data_i[7:0] };
    end 
    if(N850) begin
      { mem[479:472] } <= { data_i[7:0] };
    end 
    if(N849) begin
      { mem[471:464] } <= { data_i[7:0] };
    end 
    if(N848) begin
      { mem[463:456] } <= { data_i[7:0] };
    end 
    if(N847) begin
      { mem[455:448] } <= { data_i[7:0] };
    end 
    if(N846) begin
      { mem[447:440] } <= { data_i[7:0] };
    end 
    if(N845) begin
      { mem[439:432] } <= { data_i[7:0] };
    end 
    if(N844) begin
      { mem[431:424] } <= { data_i[7:0] };
    end 
    if(N843) begin
      { mem[423:416] } <= { data_i[7:0] };
    end 
    if(N842) begin
      { mem[415:408] } <= { data_i[7:0] };
    end 
    if(N841) begin
      { mem[407:400] } <= { data_i[7:0] };
    end 
    if(N840) begin
      { mem[399:392] } <= { data_i[7:0] };
    end 
    if(N839) begin
      { mem[391:384] } <= { data_i[7:0] };
    end 
    if(N838) begin
      { mem[383:376] } <= { data_i[7:0] };
    end 
    if(N837) begin
      { mem[375:368] } <= { data_i[7:0] };
    end 
    if(N836) begin
      { mem[367:360] } <= { data_i[7:0] };
    end 
    if(N835) begin
      { mem[359:352] } <= { data_i[7:0] };
    end 
    if(N834) begin
      { mem[351:344] } <= { data_i[7:0] };
    end 
    if(N833) begin
      { mem[343:336] } <= { data_i[7:0] };
    end 
    if(N832) begin
      { mem[335:328] } <= { data_i[7:0] };
    end 
    if(N831) begin
      { mem[327:320] } <= { data_i[7:0] };
    end 
    if(N830) begin
      { mem[319:312] } <= { data_i[7:0] };
    end 
    if(N829) begin
      { mem[311:304] } <= { data_i[7:0] };
    end 
    if(N828) begin
      { mem[303:296] } <= { data_i[7:0] };
    end 
    if(N827) begin
      { mem[295:288] } <= { data_i[7:0] };
    end 
    if(N826) begin
      { mem[287:280] } <= { data_i[7:0] };
    end 
    if(N825) begin
      { mem[279:272] } <= { data_i[7:0] };
    end 
    if(N824) begin
      { mem[271:264] } <= { data_i[7:0] };
    end 
    if(N823) begin
      { mem[263:256] } <= { data_i[7:0] };
    end 
    if(N822) begin
      { mem[255:248] } <= { data_i[7:0] };
    end 
    if(N821) begin
      { mem[247:240] } <= { data_i[7:0] };
    end 
    if(N820) begin
      { mem[239:232] } <= { data_i[7:0] };
    end 
    if(N819) begin
      { mem[231:224] } <= { data_i[7:0] };
    end 
    if(N818) begin
      { mem[223:216] } <= { data_i[7:0] };
    end 
    if(N817) begin
      { mem[215:208] } <= { data_i[7:0] };
    end 
    if(N816) begin
      { mem[207:200] } <= { data_i[7:0] };
    end 
    if(N815) begin
      { mem[199:192] } <= { data_i[7:0] };
    end 
    if(N814) begin
      { mem[191:184] } <= { data_i[7:0] };
    end 
    if(N813) begin
      { mem[183:176] } <= { data_i[7:0] };
    end 
    if(N812) begin
      { mem[175:168] } <= { data_i[7:0] };
    end 
    if(N811) begin
      { mem[167:160] } <= { data_i[7:0] };
    end 
    if(N810) begin
      { mem[159:152] } <= { data_i[7:0] };
    end 
    if(N809) begin
      { mem[151:144] } <= { data_i[7:0] };
    end 
    if(N808) begin
      { mem[143:136] } <= { data_i[7:0] };
    end 
    if(N807) begin
      { mem[135:128] } <= { data_i[7:0] };
    end 
    if(N806) begin
      { mem[127:120] } <= { data_i[7:0] };
    end 
    if(N805) begin
      { mem[119:112] } <= { data_i[7:0] };
    end 
    if(N804) begin
      { mem[111:104] } <= { data_i[7:0] };
    end 
    if(N803) begin
      { mem[103:96] } <= { data_i[7:0] };
    end 
    if(N802) begin
      { mem[95:88] } <= { data_i[7:0] };
    end 
    if(N801) begin
      { mem[87:80] } <= { data_i[7:0] };
    end 
    if(N800) begin
      { mem[79:72] } <= { data_i[7:0] };
    end 
    if(N799) begin
      { mem[71:64] } <= { data_i[7:0] };
    end 
    if(N798) begin
      { mem[63:56] } <= { data_i[7:0] };
    end 
    if(N797) begin
      { mem[55:48] } <= { data_i[7:0] };
    end 
    if(N796) begin
      { mem[47:40] } <= { data_i[7:0] };
    end 
    if(N795) begin
      { mem[39:32] } <= { data_i[7:0] };
    end 
    if(N794) begin
      { mem[31:24] } <= { data_i[7:0] };
    end 
    if(N793) begin
      { mem[23:16] } <= { data_i[7:0] };
    end 
    if(N792) begin
      { mem[15:8] } <= { data_i[7:0] };
    end 
    if(N791) begin
      { mem[7:0] } <= { data_i[7:0] };
    end 
  end


endmodule



module bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [7:0] addr_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [7:0] data_o;

  bsg_mem_1rw_sync_synth_width_p8_els_p256_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .v_i(v_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_synth_els_p256_latch_last_read_p1_data_width_p64
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [7:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;
  wire N0,N1,n_0_net__0_,n_1_net_,N2,N3,n_2_net__0_,n_3_net_,N4,n_4_net__0_,n_5_net_,
  N5,n_6_net__0_,n_7_net_,N6,n_8_net__0_,n_9_net_,N7,n_10_net__0_,n_11_net_,N8,
  n_12_net__0_,n_13_net_,N9,n_14_net__0_,n_15_net_,N10;

  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_0__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[7:0]),
    .addr_i(addr_i),
    .v_i(n_0_net__0_),
    .w_i(n_1_net_),
    .data_o(data_o[7:0])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_1__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[15:8]),
    .addr_i(addr_i),
    .v_i(n_2_net__0_),
    .w_i(n_3_net_),
    .data_o(data_o[15:8])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_2__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[23:16]),
    .addr_i(addr_i),
    .v_i(n_4_net__0_),
    .w_i(n_5_net_),
    .data_o(data_o[23:16])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_3__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[31:24]),
    .addr_i(addr_i),
    .v_i(n_6_net__0_),
    .w_i(n_7_net_),
    .data_o(data_o[31:24])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_4__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[39:32]),
    .addr_i(addr_i),
    .v_i(n_8_net__0_),
    .w_i(n_9_net_),
    .data_o(data_o[39:32])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_5__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[47:40]),
    .addr_i(addr_i),
    .v_i(n_10_net__0_),
    .w_i(n_11_net_),
    .data_o(data_o[47:40])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_6__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[55:48]),
    .addr_i(addr_i),
    .v_i(n_12_net__0_),
    .w_i(n_13_net_),
    .data_o(data_o[55:48])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8
  bk_7__mem_1rw_sync
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[63:56]),
    .addr_i(addr_i),
    .v_i(n_14_net__0_),
    .w_i(n_15_net_),
    .data_o(data_o[63:56])
  );

  assign N3 = (N0)? write_mask_i[0] : 
              (N1)? 1'b1 : 1'b0;
  assign N0 = w_i;
  assign N1 = N2;
  assign N4 = (N0)? write_mask_i[1] : 
              (N1)? 1'b1 : 1'b0;
  assign N5 = (N0)? write_mask_i[2] : 
              (N1)? 1'b1 : 1'b0;
  assign N6 = (N0)? write_mask_i[3] : 
              (N1)? 1'b1 : 1'b0;
  assign N7 = (N0)? write_mask_i[4] : 
              (N1)? 1'b1 : 1'b0;
  assign N8 = (N0)? write_mask_i[5] : 
              (N1)? 1'b1 : 1'b0;
  assign N9 = (N0)? write_mask_i[6] : 
              (N1)? 1'b1 : 1'b0;
  assign N10 = (N0)? write_mask_i[7] : 
               (N1)? 1'b1 : 1'b0;
  assign n_1_net_ = w_i & write_mask_i[0];
  assign N2 = ~w_i;
  assign n_0_net__0_ = v_i & N3;
  assign n_3_net_ = w_i & write_mask_i[1];
  assign n_2_net__0_ = v_i & N4;
  assign n_5_net_ = w_i & write_mask_i[2];
  assign n_4_net__0_ = v_i & N5;
  assign n_7_net_ = w_i & write_mask_i[3];
  assign n_6_net__0_ = v_i & N6;
  assign n_9_net_ = w_i & write_mask_i[4];
  assign n_8_net__0_ = v_i & N7;
  assign n_11_net_ = w_i & write_mask_i[5];
  assign n_10_net__0_ = v_i & N8;
  assign n_13_net_ = w_i & write_mask_i[6];
  assign n_12_net__0_ = v_i & N9;
  assign n_15_net_ = w_i & write_mask_i[7];
  assign n_14_net__0_ = v_i & N10;

endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p256_data_width_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [7:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  bsg_mem_1rw_sync_mask_write_byte_synth_els_p256_latch_last_read_p1_data_width_p64
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_width_p2_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [1:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[0] = i[0] | 1'b0;
  assign o[1] = i[1] | i[0];

endmodule



module bsg_priority_encode_one_hot_out_width_p2_lo_to_hi_p1
(
  i,
  o
);

  input [1:0] i;
  output [1:0] o;
  wire [1:0] o;
  wire N0;
  wire [1:1] scan_lo;

  bsg_scan_width_p2_or_p1_lo_to_hi_p1
  genblk1_scan
  (
    .i(i),
    .o({ scan_lo[1:1], o[0:0] })
  );

  assign o[1] = scan_lo[1] & N0;
  assign N0 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_priority_encode_width_p2_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  wire [1:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p2_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p2_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o[0]),
    .v_o(v_o)
  );


endmodule



module bsg_dff_en_width_p3_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  input en_i;
  reg [2:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[2:0] } <= { data_i[2:0] };
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p3
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  input en_i;
  wire [2:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p3_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p3_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [2:0] data_i;
  input [5:0] addr_i;
  input [2:0] w_mask_i;
  output [2:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [2:0] data_o,data_out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,read_en,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,llr_read_en_r,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621;
  reg [5:0] addr_r;
  reg [191:0] mem;
  assign data_out[2] = (N78)? mem[2] : 
                       (N80)? mem[5] : 
                       (N82)? mem[8] : 
                       (N84)? mem[11] : 
                       (N86)? mem[14] : 
                       (N88)? mem[17] : 
                       (N90)? mem[20] : 
                       (N92)? mem[23] : 
                       (N94)? mem[26] : 
                       (N96)? mem[29] : 
                       (N98)? mem[32] : 
                       (N100)? mem[35] : 
                       (N102)? mem[38] : 
                       (N104)? mem[41] : 
                       (N106)? mem[44] : 
                       (N108)? mem[47] : 
                       (N110)? mem[50] : 
                       (N112)? mem[53] : 
                       (N114)? mem[56] : 
                       (N116)? mem[59] : 
                       (N118)? mem[62] : 
                       (N120)? mem[65] : 
                       (N122)? mem[68] : 
                       (N124)? mem[71] : 
                       (N126)? mem[74] : 
                       (N128)? mem[77] : 
                       (N130)? mem[80] : 
                       (N132)? mem[83] : 
                       (N134)? mem[86] : 
                       (N136)? mem[89] : 
                       (N138)? mem[92] : 
                       (N140)? mem[95] : 
                       (N79)? mem[98] : 
                       (N81)? mem[101] : 
                       (N83)? mem[104] : 
                       (N85)? mem[107] : 
                       (N87)? mem[110] : 
                       (N89)? mem[113] : 
                       (N91)? mem[116] : 
                       (N93)? mem[119] : 
                       (N95)? mem[122] : 
                       (N97)? mem[125] : 
                       (N99)? mem[128] : 
                       (N101)? mem[131] : 
                       (N103)? mem[134] : 
                       (N105)? mem[137] : 
                       (N107)? mem[140] : 
                       (N109)? mem[143] : 
                       (N111)? mem[146] : 
                       (N113)? mem[149] : 
                       (N115)? mem[152] : 
                       (N117)? mem[155] : 
                       (N119)? mem[158] : 
                       (N121)? mem[161] : 
                       (N123)? mem[164] : 
                       (N125)? mem[167] : 
                       (N127)? mem[170] : 
                       (N129)? mem[173] : 
                       (N131)? mem[176] : 
                       (N133)? mem[179] : 
                       (N135)? mem[182] : 
                       (N137)? mem[185] : 
                       (N139)? mem[188] : 
                       (N141)? mem[191] : 1'b0;
  assign data_out[1] = (N78)? mem[1] : 
                       (N80)? mem[4] : 
                       (N82)? mem[7] : 
                       (N84)? mem[10] : 
                       (N86)? mem[13] : 
                       (N88)? mem[16] : 
                       (N90)? mem[19] : 
                       (N92)? mem[22] : 
                       (N94)? mem[25] : 
                       (N96)? mem[28] : 
                       (N98)? mem[31] : 
                       (N100)? mem[34] : 
                       (N102)? mem[37] : 
                       (N104)? mem[40] : 
                       (N106)? mem[43] : 
                       (N108)? mem[46] : 
                       (N110)? mem[49] : 
                       (N112)? mem[52] : 
                       (N114)? mem[55] : 
                       (N116)? mem[58] : 
                       (N118)? mem[61] : 
                       (N120)? mem[64] : 
                       (N122)? mem[67] : 
                       (N124)? mem[70] : 
                       (N126)? mem[73] : 
                       (N128)? mem[76] : 
                       (N130)? mem[79] : 
                       (N132)? mem[82] : 
                       (N134)? mem[85] : 
                       (N136)? mem[88] : 
                       (N138)? mem[91] : 
                       (N140)? mem[94] : 
                       (N79)? mem[97] : 
                       (N81)? mem[100] : 
                       (N83)? mem[103] : 
                       (N85)? mem[106] : 
                       (N87)? mem[109] : 
                       (N89)? mem[112] : 
                       (N91)? mem[115] : 
                       (N93)? mem[118] : 
                       (N95)? mem[121] : 
                       (N97)? mem[124] : 
                       (N99)? mem[127] : 
                       (N101)? mem[130] : 
                       (N103)? mem[133] : 
                       (N105)? mem[136] : 
                       (N107)? mem[139] : 
                       (N109)? mem[142] : 
                       (N111)? mem[145] : 
                       (N113)? mem[148] : 
                       (N115)? mem[151] : 
                       (N117)? mem[154] : 
                       (N119)? mem[157] : 
                       (N121)? mem[160] : 
                       (N123)? mem[163] : 
                       (N125)? mem[166] : 
                       (N127)? mem[169] : 
                       (N129)? mem[172] : 
                       (N131)? mem[175] : 
                       (N133)? mem[178] : 
                       (N135)? mem[181] : 
                       (N137)? mem[184] : 
                       (N139)? mem[187] : 
                       (N141)? mem[190] : 1'b0;
  assign data_out[0] = (N78)? mem[0] : 
                       (N80)? mem[3] : 
                       (N82)? mem[6] : 
                       (N84)? mem[9] : 
                       (N86)? mem[12] : 
                       (N88)? mem[15] : 
                       (N90)? mem[18] : 
                       (N92)? mem[21] : 
                       (N94)? mem[24] : 
                       (N96)? mem[27] : 
                       (N98)? mem[30] : 
                       (N100)? mem[33] : 
                       (N102)? mem[36] : 
                       (N104)? mem[39] : 
                       (N106)? mem[42] : 
                       (N108)? mem[45] : 
                       (N110)? mem[48] : 
                       (N112)? mem[51] : 
                       (N114)? mem[54] : 
                       (N116)? mem[57] : 
                       (N118)? mem[60] : 
                       (N120)? mem[63] : 
                       (N122)? mem[66] : 
                       (N124)? mem[69] : 
                       (N126)? mem[72] : 
                       (N128)? mem[75] : 
                       (N130)? mem[78] : 
                       (N132)? mem[81] : 
                       (N134)? mem[84] : 
                       (N136)? mem[87] : 
                       (N138)? mem[90] : 
                       (N140)? mem[93] : 
                       (N79)? mem[96] : 
                       (N81)? mem[99] : 
                       (N83)? mem[102] : 
                       (N85)? mem[105] : 
                       (N87)? mem[108] : 
                       (N89)? mem[111] : 
                       (N91)? mem[114] : 
                       (N93)? mem[117] : 
                       (N95)? mem[120] : 
                       (N97)? mem[123] : 
                       (N99)? mem[126] : 
                       (N101)? mem[129] : 
                       (N103)? mem[132] : 
                       (N105)? mem[135] : 
                       (N107)? mem[138] : 
                       (N109)? mem[141] : 
                       (N111)? mem[144] : 
                       (N113)? mem[147] : 
                       (N115)? mem[150] : 
                       (N117)? mem[153] : 
                       (N119)? mem[156] : 
                       (N121)? mem[159] : 
                       (N123)? mem[162] : 
                       (N125)? mem[165] : 
                       (N127)? mem[168] : 
                       (N129)? mem[171] : 
                       (N131)? mem[174] : 
                       (N133)? mem[177] : 
                       (N135)? mem[180] : 
                       (N137)? mem[183] : 
                       (N139)? mem[186] : 
                       (N141)? mem[189] : 1'b0;

  bsg_dff_width_p1
  llr_read_en_dff
  (
    .clk_i(clk_i),
    .data_i(read_en),
    .data_o(llr_read_en_r)
  );


  bsg_dff_en_bypass_width_p3
  llr_dff_bypass
  (
    .clk_i(clk_i),
    .en_i(llr_read_en_r),
    .data_i(data_out),
    .data_o(data_o)
  );

  assign N595 = ~addr_i[5];
  assign N596 = addr_i[3] & addr_i[4];
  assign N597 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N598 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N599 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N600 = addr_i[5] & N596;
  assign N601 = addr_i[5] & N597;
  assign N602 = addr_i[5] & N598;
  assign N603 = addr_i[5] & N599;
  assign N604 = N595 & N596;
  assign N605 = N595 & N597;
  assign N606 = N595 & N598;
  assign N607 = N595 & N599;
  assign N608 = ~addr_i[2];
  assign N609 = addr_i[0] & addr_i[1];
  assign N610 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N611 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N612 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N613 = addr_i[2] & N609;
  assign N614 = addr_i[2] & N610;
  assign N615 = addr_i[2] & N611;
  assign N616 = addr_i[2] & N612;
  assign N617 = N608 & N609;
  assign N618 = N608 & N610;
  assign N619 = N608 & N611;
  assign N620 = N608 & N612;
  assign N338 = N600 & N613;
  assign N337 = N600 & N614;
  assign N336 = N600 & N615;
  assign N335 = N600 & N616;
  assign N334 = N600 & N617;
  assign N333 = N600 & N618;
  assign N332 = N600 & N619;
  assign N331 = N600 & N620;
  assign N330 = N601 & N613;
  assign N329 = N601 & N614;
  assign N328 = N601 & N615;
  assign N327 = N601 & N616;
  assign N326 = N601 & N617;
  assign N325 = N601 & N618;
  assign N324 = N601 & N619;
  assign N323 = N601 & N620;
  assign N322 = N602 & N613;
  assign N321 = N602 & N614;
  assign N320 = N602 & N615;
  assign N319 = N602 & N616;
  assign N318 = N602 & N617;
  assign N317 = N602 & N618;
  assign N316 = N602 & N619;
  assign N315 = N602 & N620;
  assign N314 = N603 & N613;
  assign N313 = N603 & N614;
  assign N312 = N603 & N615;
  assign N311 = N603 & N616;
  assign N310 = N603 & N617;
  assign N309 = N603 & N618;
  assign N308 = N603 & N619;
  assign N307 = N603 & N620;
  assign N306 = N604 & N613;
  assign N305 = N604 & N614;
  assign N304 = N604 & N615;
  assign N303 = N604 & N616;
  assign N302 = N604 & N617;
  assign N301 = N604 & N618;
  assign N300 = N604 & N619;
  assign N299 = N604 & N620;
  assign N298 = N605 & N613;
  assign N297 = N605 & N614;
  assign N296 = N605 & N615;
  assign N295 = N605 & N616;
  assign N294 = N605 & N617;
  assign N293 = N605 & N618;
  assign N292 = N605 & N619;
  assign N291 = N605 & N620;
  assign N290 = N606 & N613;
  assign N289 = N606 & N614;
  assign N288 = N606 & N615;
  assign N287 = N606 & N616;
  assign N286 = N606 & N617;
  assign N285 = N606 & N618;
  assign N284 = N606 & N619;
  assign N283 = N606 & N620;
  assign N282 = N607 & N613;
  assign N281 = N607 & N614;
  assign N280 = N607 & N615;
  assign N279 = N607 & N616;
  assign N278 = N607 & N617;
  assign N277 = N607 & N618;
  assign N276 = N607 & N619;
  assign N275 = N607 & N620;
  assign { N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145 } = (N8)? { N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N144)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210 } = (N9)? { N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N209)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339 } = (N10)? { N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N274)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403 } = (N11)? { N402, N273, N208, N401, N272, N207, N400, N271, N206, N399, N270, N205, N398, N269, N204, N397, N268, N203, N396, N267, N202, N395, N266, N201, N394, N265, N200, N393, N264, N199, N392, N263, N198, N391, N262, N197, N390, N261, N196, N389, N260, N195, N388, N259, N194, N387, N258, N193, N386, N257, N192, N385, N256, N191, N384, N255, N190, N383, N254, N189, N382, N253, N188, N381, N252, N187, N380, N251, N186, N379, N250, N185, N378, N249, N184, N377, N248, N183, N376, N247, N182, N375, N246, N181, N374, N245, N180, N373, N244, N179, N372, N243, N178, N371, N242, N177, N370, N241, N176, N369, N240, N175, N368, N239, N174, N367, N238, N173, N366, N237, N172, N365, N236, N171, N364, N235, N170, N363, N234, N169, N362, N233, N168, N361, N232, N167, N360, N231, N166, N359, N230, N165, N358, N229, N164, N357, N228, N163, N356, N227, N162, N355, N226, N161, N354, N225, N160, N353, N224, N159, N352, N223, N158, N351, N222, N157, N350, N221, N156, N349, N220, N155, N348, N219, N154, N347, N218, N153, N346, N217, N152, N345, N216, N151, N344, N215, N150, N343, N214, N149, N342, N213, N148, N341, N212, N147, N340, N211, N146, N339, N210, N145 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N143)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = N142;
  assign read_en = v_i & N621;
  assign N621 = ~w_i;
  assign N12 = ~addr_r[0];
  assign N13 = ~addr_r[1];
  assign N14 = N12 & N13;
  assign N15 = N12 & addr_r[1];
  assign N16 = addr_r[0] & N13;
  assign N17 = addr_r[0] & addr_r[1];
  assign N18 = ~addr_r[2];
  assign N19 = N14 & N18;
  assign N20 = N14 & addr_r[2];
  assign N21 = N16 & N18;
  assign N22 = N16 & addr_r[2];
  assign N23 = N15 & N18;
  assign N24 = N15 & addr_r[2];
  assign N25 = N17 & N18;
  assign N26 = N17 & addr_r[2];
  assign N27 = ~addr_r[3];
  assign N28 = N19 & N27;
  assign N29 = N19 & addr_r[3];
  assign N30 = N21 & N27;
  assign N31 = N21 & addr_r[3];
  assign N32 = N23 & N27;
  assign N33 = N23 & addr_r[3];
  assign N34 = N25 & N27;
  assign N35 = N25 & addr_r[3];
  assign N36 = N20 & N27;
  assign N37 = N20 & addr_r[3];
  assign N38 = N22 & N27;
  assign N39 = N22 & addr_r[3];
  assign N40 = N24 & N27;
  assign N41 = N24 & addr_r[3];
  assign N42 = N26 & N27;
  assign N43 = N26 & addr_r[3];
  assign N44 = ~addr_r[4];
  assign N45 = N28 & N44;
  assign N46 = N28 & addr_r[4];
  assign N47 = N30 & N44;
  assign N48 = N30 & addr_r[4];
  assign N49 = N32 & N44;
  assign N50 = N32 & addr_r[4];
  assign N51 = N34 & N44;
  assign N52 = N34 & addr_r[4];
  assign N53 = N36 & N44;
  assign N54 = N36 & addr_r[4];
  assign N55 = N38 & N44;
  assign N56 = N38 & addr_r[4];
  assign N57 = N40 & N44;
  assign N58 = N40 & addr_r[4];
  assign N59 = N42 & N44;
  assign N60 = N42 & addr_r[4];
  assign N61 = N29 & N44;
  assign N62 = N29 & addr_r[4];
  assign N63 = N31 & N44;
  assign N64 = N31 & addr_r[4];
  assign N65 = N33 & N44;
  assign N66 = N33 & addr_r[4];
  assign N67 = N35 & N44;
  assign N68 = N35 & addr_r[4];
  assign N69 = N37 & N44;
  assign N70 = N37 & addr_r[4];
  assign N71 = N39 & N44;
  assign N72 = N39 & addr_r[4];
  assign N73 = N41 & N44;
  assign N74 = N41 & addr_r[4];
  assign N75 = N43 & N44;
  assign N76 = N43 & addr_r[4];
  assign N77 = ~addr_r[5];
  assign N78 = N45 & N77;
  assign N79 = N45 & addr_r[5];
  assign N80 = N47 & N77;
  assign N81 = N47 & addr_r[5];
  assign N82 = N49 & N77;
  assign N83 = N49 & addr_r[5];
  assign N84 = N51 & N77;
  assign N85 = N51 & addr_r[5];
  assign N86 = N53 & N77;
  assign N87 = N53 & addr_r[5];
  assign N88 = N55 & N77;
  assign N89 = N55 & addr_r[5];
  assign N90 = N57 & N77;
  assign N91 = N57 & addr_r[5];
  assign N92 = N59 & N77;
  assign N93 = N59 & addr_r[5];
  assign N94 = N61 & N77;
  assign N95 = N61 & addr_r[5];
  assign N96 = N63 & N77;
  assign N97 = N63 & addr_r[5];
  assign N98 = N65 & N77;
  assign N99 = N65 & addr_r[5];
  assign N100 = N67 & N77;
  assign N101 = N67 & addr_r[5];
  assign N102 = N69 & N77;
  assign N103 = N69 & addr_r[5];
  assign N104 = N71 & N77;
  assign N105 = N71 & addr_r[5];
  assign N106 = N73 & N77;
  assign N107 = N73 & addr_r[5];
  assign N108 = N75 & N77;
  assign N109 = N75 & addr_r[5];
  assign N110 = N46 & N77;
  assign N111 = N46 & addr_r[5];
  assign N112 = N48 & N77;
  assign N113 = N48 & addr_r[5];
  assign N114 = N50 & N77;
  assign N115 = N50 & addr_r[5];
  assign N116 = N52 & N77;
  assign N117 = N52 & addr_r[5];
  assign N118 = N54 & N77;
  assign N119 = N54 & addr_r[5];
  assign N120 = N56 & N77;
  assign N121 = N56 & addr_r[5];
  assign N122 = N58 & N77;
  assign N123 = N58 & addr_r[5];
  assign N124 = N60 & N77;
  assign N125 = N60 & addr_r[5];
  assign N126 = N62 & N77;
  assign N127 = N62 & addr_r[5];
  assign N128 = N64 & N77;
  assign N129 = N64 & addr_r[5];
  assign N130 = N66 & N77;
  assign N131 = N66 & addr_r[5];
  assign N132 = N68 & N77;
  assign N133 = N68 & addr_r[5];
  assign N134 = N70 & N77;
  assign N135 = N70 & addr_r[5];
  assign N136 = N72 & N77;
  assign N137 = N72 & addr_r[5];
  assign N138 = N74 & N77;
  assign N139 = N74 & addr_r[5];
  assign N140 = N76 & N77;
  assign N141 = N76 & addr_r[5];
  assign N142 = v_i & w_i;
  assign N143 = ~N142;
  assign N144 = ~w_mask_i[0];
  assign N209 = ~w_mask_i[1];
  assign N274 = ~w_mask_i[2];

  always @(posedge clk_i) begin
    if(1'b1) begin
      { addr_r[5:0] } <= { addr_i[5:0] };
    end 
    if(N594) begin
      { mem[191:191] } <= { data_i[2:2] };
    end 
    if(N593) begin
      { mem[190:190] } <= { data_i[1:1] };
    end 
    if(N592) begin
      { mem[189:189] } <= { data_i[0:0] };
    end 
    if(N591) begin
      { mem[188:188] } <= { data_i[2:2] };
    end 
    if(N590) begin
      { mem[187:187] } <= { data_i[1:1] };
    end 
    if(N589) begin
      { mem[186:186] } <= { data_i[0:0] };
    end 
    if(N588) begin
      { mem[185:185] } <= { data_i[2:2] };
    end 
    if(N587) begin
      { mem[184:184] } <= { data_i[1:1] };
    end 
    if(N586) begin
      { mem[183:183] } <= { data_i[0:0] };
    end 
    if(N585) begin
      { mem[182:182] } <= { data_i[2:2] };
    end 
    if(N584) begin
      { mem[181:181] } <= { data_i[1:1] };
    end 
    if(N583) begin
      { mem[180:180] } <= { data_i[0:0] };
    end 
    if(N582) begin
      { mem[179:179] } <= { data_i[2:2] };
    end 
    if(N581) begin
      { mem[178:178] } <= { data_i[1:1] };
    end 
    if(N580) begin
      { mem[177:177] } <= { data_i[0:0] };
    end 
    if(N579) begin
      { mem[176:176] } <= { data_i[2:2] };
    end 
    if(N578) begin
      { mem[175:175] } <= { data_i[1:1] };
    end 
    if(N577) begin
      { mem[174:174] } <= { data_i[0:0] };
    end 
    if(N576) begin
      { mem[173:173] } <= { data_i[2:2] };
    end 
    if(N575) begin
      { mem[172:172] } <= { data_i[1:1] };
    end 
    if(N574) begin
      { mem[171:171] } <= { data_i[0:0] };
    end 
    if(N573) begin
      { mem[170:170] } <= { data_i[2:2] };
    end 
    if(N572) begin
      { mem[169:169] } <= { data_i[1:1] };
    end 
    if(N571) begin
      { mem[168:168] } <= { data_i[0:0] };
    end 
    if(N570) begin
      { mem[167:167] } <= { data_i[2:2] };
    end 
    if(N569) begin
      { mem[166:166] } <= { data_i[1:1] };
    end 
    if(N568) begin
      { mem[165:165] } <= { data_i[0:0] };
    end 
    if(N567) begin
      { mem[164:164] } <= { data_i[2:2] };
    end 
    if(N566) begin
      { mem[163:163] } <= { data_i[1:1] };
    end 
    if(N565) begin
      { mem[162:162] } <= { data_i[0:0] };
    end 
    if(N564) begin
      { mem[161:161] } <= { data_i[2:2] };
    end 
    if(N563) begin
      { mem[160:160] } <= { data_i[1:1] };
    end 
    if(N562) begin
      { mem[159:159] } <= { data_i[0:0] };
    end 
    if(N561) begin
      { mem[158:158] } <= { data_i[2:2] };
    end 
    if(N560) begin
      { mem[157:157] } <= { data_i[1:1] };
    end 
    if(N559) begin
      { mem[156:156] } <= { data_i[0:0] };
    end 
    if(N558) begin
      { mem[155:155] } <= { data_i[2:2] };
    end 
    if(N557) begin
      { mem[154:154] } <= { data_i[1:1] };
    end 
    if(N556) begin
      { mem[153:153] } <= { data_i[0:0] };
    end 
    if(N555) begin
      { mem[152:152] } <= { data_i[2:2] };
    end 
    if(N554) begin
      { mem[151:151] } <= { data_i[1:1] };
    end 
    if(N553) begin
      { mem[150:150] } <= { data_i[0:0] };
    end 
    if(N552) begin
      { mem[149:149] } <= { data_i[2:2] };
    end 
    if(N551) begin
      { mem[148:148] } <= { data_i[1:1] };
    end 
    if(N550) begin
      { mem[147:147] } <= { data_i[0:0] };
    end 
    if(N549) begin
      { mem[146:146] } <= { data_i[2:2] };
    end 
    if(N548) begin
      { mem[145:145] } <= { data_i[1:1] };
    end 
    if(N547) begin
      { mem[144:144] } <= { data_i[0:0] };
    end 
    if(N546) begin
      { mem[143:143] } <= { data_i[2:2] };
    end 
    if(N545) begin
      { mem[142:142] } <= { data_i[1:1] };
    end 
    if(N544) begin
      { mem[141:141] } <= { data_i[0:0] };
    end 
    if(N543) begin
      { mem[140:140] } <= { data_i[2:2] };
    end 
    if(N542) begin
      { mem[139:139] } <= { data_i[1:1] };
    end 
    if(N541) begin
      { mem[138:138] } <= { data_i[0:0] };
    end 
    if(N540) begin
      { mem[137:137] } <= { data_i[2:2] };
    end 
    if(N539) begin
      { mem[136:136] } <= { data_i[1:1] };
    end 
    if(N538) begin
      { mem[135:135] } <= { data_i[0:0] };
    end 
    if(N537) begin
      { mem[134:134] } <= { data_i[2:2] };
    end 
    if(N536) begin
      { mem[133:133] } <= { data_i[1:1] };
    end 
    if(N535) begin
      { mem[132:132] } <= { data_i[0:0] };
    end 
    if(N534) begin
      { mem[131:131] } <= { data_i[2:2] };
    end 
    if(N533) begin
      { mem[130:130] } <= { data_i[1:1] };
    end 
    if(N532) begin
      { mem[129:129] } <= { data_i[0:0] };
    end 
    if(N531) begin
      { mem[128:128] } <= { data_i[2:2] };
    end 
    if(N530) begin
      { mem[127:127] } <= { data_i[1:1] };
    end 
    if(N529) begin
      { mem[126:126] } <= { data_i[0:0] };
    end 
    if(N528) begin
      { mem[125:125] } <= { data_i[2:2] };
    end 
    if(N527) begin
      { mem[124:124] } <= { data_i[1:1] };
    end 
    if(N526) begin
      { mem[123:123] } <= { data_i[0:0] };
    end 
    if(N525) begin
      { mem[122:122] } <= { data_i[2:2] };
    end 
    if(N524) begin
      { mem[121:121] } <= { data_i[1:1] };
    end 
    if(N523) begin
      { mem[120:120] } <= { data_i[0:0] };
    end 
    if(N522) begin
      { mem[119:119] } <= { data_i[2:2] };
    end 
    if(N521) begin
      { mem[118:118] } <= { data_i[1:1] };
    end 
    if(N520) begin
      { mem[117:117] } <= { data_i[0:0] };
    end 
    if(N519) begin
      { mem[116:116] } <= { data_i[2:2] };
    end 
    if(N518) begin
      { mem[115:115] } <= { data_i[1:1] };
    end 
    if(N517) begin
      { mem[114:114] } <= { data_i[0:0] };
    end 
    if(N516) begin
      { mem[113:113] } <= { data_i[2:2] };
    end 
    if(N515) begin
      { mem[112:112] } <= { data_i[1:1] };
    end 
    if(N514) begin
      { mem[111:111] } <= { data_i[0:0] };
    end 
    if(N513) begin
      { mem[110:110] } <= { data_i[2:2] };
    end 
    if(N512) begin
      { mem[109:109] } <= { data_i[1:1] };
    end 
    if(N511) begin
      { mem[108:108] } <= { data_i[0:0] };
    end 
    if(N510) begin
      { mem[107:107] } <= { data_i[2:2] };
    end 
    if(N509) begin
      { mem[106:106] } <= { data_i[1:1] };
    end 
    if(N508) begin
      { mem[105:105] } <= { data_i[0:0] };
    end 
    if(N507) begin
      { mem[104:104] } <= { data_i[2:2] };
    end 
    if(N506) begin
      { mem[103:103] } <= { data_i[1:1] };
    end 
    if(N505) begin
      { mem[102:102] } <= { data_i[0:0] };
    end 
    if(N504) begin
      { mem[101:101] } <= { data_i[2:2] };
    end 
    if(N503) begin
      { mem[100:100] } <= { data_i[1:1] };
    end 
    if(N502) begin
      { mem[99:99] } <= { data_i[0:0] };
    end 
    if(N501) begin
      { mem[98:98] } <= { data_i[2:2] };
    end 
    if(N500) begin
      { mem[97:97] } <= { data_i[1:1] };
    end 
    if(N499) begin
      { mem[96:96] } <= { data_i[0:0] };
    end 
    if(N498) begin
      { mem[95:95] } <= { data_i[2:2] };
    end 
    if(N497) begin
      { mem[94:94] } <= { data_i[1:1] };
    end 
    if(N496) begin
      { mem[93:93] } <= { data_i[0:0] };
    end 
    if(N495) begin
      { mem[92:92] } <= { data_i[2:2] };
    end 
    if(N494) begin
      { mem[91:91] } <= { data_i[1:1] };
    end 
    if(N493) begin
      { mem[90:90] } <= { data_i[0:0] };
    end 
    if(N492) begin
      { mem[89:89] } <= { data_i[2:2] };
    end 
    if(N491) begin
      { mem[88:88] } <= { data_i[1:1] };
    end 
    if(N490) begin
      { mem[87:87] } <= { data_i[0:0] };
    end 
    if(N489) begin
      { mem[86:86] } <= { data_i[2:2] };
    end 
    if(N488) begin
      { mem[85:85] } <= { data_i[1:1] };
    end 
    if(N487) begin
      { mem[84:84] } <= { data_i[0:0] };
    end 
    if(N486) begin
      { mem[83:83] } <= { data_i[2:2] };
    end 
    if(N485) begin
      { mem[82:82] } <= { data_i[1:1] };
    end 
    if(N484) begin
      { mem[81:81] } <= { data_i[0:0] };
    end 
    if(N483) begin
      { mem[80:80] } <= { data_i[2:2] };
    end 
    if(N482) begin
      { mem[79:79] } <= { data_i[1:1] };
    end 
    if(N481) begin
      { mem[78:78] } <= { data_i[0:0] };
    end 
    if(N480) begin
      { mem[77:77] } <= { data_i[2:2] };
    end 
    if(N479) begin
      { mem[76:76] } <= { data_i[1:1] };
    end 
    if(N478) begin
      { mem[75:75] } <= { data_i[0:0] };
    end 
    if(N477) begin
      { mem[74:74] } <= { data_i[2:2] };
    end 
    if(N476) begin
      { mem[73:73] } <= { data_i[1:1] };
    end 
    if(N475) begin
      { mem[72:72] } <= { data_i[0:0] };
    end 
    if(N474) begin
      { mem[71:71] } <= { data_i[2:2] };
    end 
    if(N473) begin
      { mem[70:70] } <= { data_i[1:1] };
    end 
    if(N472) begin
      { mem[69:69] } <= { data_i[0:0] };
    end 
    if(N471) begin
      { mem[68:68] } <= { data_i[2:2] };
    end 
    if(N470) begin
      { mem[67:67] } <= { data_i[1:1] };
    end 
    if(N469) begin
      { mem[66:66] } <= { data_i[0:0] };
    end 
    if(N468) begin
      { mem[65:65] } <= { data_i[2:2] };
    end 
    if(N467) begin
      { mem[64:64] } <= { data_i[1:1] };
    end 
    if(N466) begin
      { mem[63:63] } <= { data_i[0:0] };
    end 
    if(N465) begin
      { mem[62:62] } <= { data_i[2:2] };
    end 
    if(N464) begin
      { mem[61:61] } <= { data_i[1:1] };
    end 
    if(N463) begin
      { mem[60:60] } <= { data_i[0:0] };
    end 
    if(N462) begin
      { mem[59:59] } <= { data_i[2:2] };
    end 
    if(N461) begin
      { mem[58:58] } <= { data_i[1:1] };
    end 
    if(N460) begin
      { mem[57:57] } <= { data_i[0:0] };
    end 
    if(N459) begin
      { mem[56:56] } <= { data_i[2:2] };
    end 
    if(N458) begin
      { mem[55:55] } <= { data_i[1:1] };
    end 
    if(N457) begin
      { mem[54:54] } <= { data_i[0:0] };
    end 
    if(N456) begin
      { mem[53:53] } <= { data_i[2:2] };
    end 
    if(N455) begin
      { mem[52:52] } <= { data_i[1:1] };
    end 
    if(N454) begin
      { mem[51:51] } <= { data_i[0:0] };
    end 
    if(N453) begin
      { mem[50:50] } <= { data_i[2:2] };
    end 
    if(N452) begin
      { mem[49:49] } <= { data_i[1:1] };
    end 
    if(N451) begin
      { mem[48:48] } <= { data_i[0:0] };
    end 
    if(N450) begin
      { mem[47:47] } <= { data_i[2:2] };
    end 
    if(N449) begin
      { mem[46:46] } <= { data_i[1:1] };
    end 
    if(N448) begin
      { mem[45:45] } <= { data_i[0:0] };
    end 
    if(N447) begin
      { mem[44:44] } <= { data_i[2:2] };
    end 
    if(N446) begin
      { mem[43:43] } <= { data_i[1:1] };
    end 
    if(N445) begin
      { mem[42:42] } <= { data_i[0:0] };
    end 
    if(N444) begin
      { mem[41:41] } <= { data_i[2:2] };
    end 
    if(N443) begin
      { mem[40:40] } <= { data_i[1:1] };
    end 
    if(N442) begin
      { mem[39:39] } <= { data_i[0:0] };
    end 
    if(N441) begin
      { mem[38:38] } <= { data_i[2:2] };
    end 
    if(N440) begin
      { mem[37:37] } <= { data_i[1:1] };
    end 
    if(N439) begin
      { mem[36:36] } <= { data_i[0:0] };
    end 
    if(N438) begin
      { mem[35:35] } <= { data_i[2:2] };
    end 
    if(N437) begin
      { mem[34:34] } <= { data_i[1:1] };
    end 
    if(N436) begin
      { mem[33:33] } <= { data_i[0:0] };
    end 
    if(N435) begin
      { mem[32:32] } <= { data_i[2:2] };
    end 
    if(N434) begin
      { mem[31:31] } <= { data_i[1:1] };
    end 
    if(N433) begin
      { mem[30:30] } <= { data_i[0:0] };
    end 
    if(N432) begin
      { mem[29:29] } <= { data_i[2:2] };
    end 
    if(N431) begin
      { mem[28:28] } <= { data_i[1:1] };
    end 
    if(N430) begin
      { mem[27:27] } <= { data_i[0:0] };
    end 
    if(N429) begin
      { mem[26:26] } <= { data_i[2:2] };
    end 
    if(N428) begin
      { mem[25:25] } <= { data_i[1:1] };
    end 
    if(N427) begin
      { mem[24:24] } <= { data_i[0:0] };
    end 
    if(N426) begin
      { mem[23:23] } <= { data_i[2:2] };
    end 
    if(N425) begin
      { mem[22:22] } <= { data_i[1:1] };
    end 
    if(N424) begin
      { mem[21:21] } <= { data_i[0:0] };
    end 
    if(N423) begin
      { mem[20:20] } <= { data_i[2:2] };
    end 
    if(N422) begin
      { mem[19:19] } <= { data_i[1:1] };
    end 
    if(N421) begin
      { mem[18:18] } <= { data_i[0:0] };
    end 
    if(N420) begin
      { mem[17:17] } <= { data_i[2:2] };
    end 
    if(N419) begin
      { mem[16:16] } <= { data_i[1:1] };
    end 
    if(N418) begin
      { mem[15:15] } <= { data_i[0:0] };
    end 
    if(N417) begin
      { mem[14:14] } <= { data_i[2:2] };
    end 
    if(N416) begin
      { mem[13:13] } <= { data_i[1:1] };
    end 
    if(N415) begin
      { mem[12:12] } <= { data_i[0:0] };
    end 
    if(N414) begin
      { mem[11:11] } <= { data_i[2:2] };
    end 
    if(N413) begin
      { mem[10:10] } <= { data_i[1:1] };
    end 
    if(N412) begin
      { mem[9:9] } <= { data_i[0:0] };
    end 
    if(N411) begin
      { mem[8:8] } <= { data_i[2:2] };
    end 
    if(N410) begin
      { mem[7:7] } <= { data_i[1:1] };
    end 
    if(N409) begin
      { mem[6:6] } <= { data_i[0:0] };
    end 
    if(N408) begin
      { mem[5:5] } <= { data_i[2:2] };
    end 
    if(N407) begin
      { mem[4:4] } <= { data_i[1:1] };
    end 
    if(N406) begin
      { mem[3:3] } <= { data_i[0:0] };
    end 
    if(N405) begin
      { mem[2:2] } <= { data_i[2:2] };
    end 
    if(N404) begin
      { mem[1:1] } <= { data_i[1:1] };
    end 
    if(N403) begin
      { mem[0:0] } <= { data_i[0:0] };
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p3_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [2:0] data_i;
  input [5:0] addr_i;
  input [2:0] w_mask_i;
  output [2:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [2:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p3_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_lru_pseudo_tree_encode_ways_p2
(
  lru_i,
  way_id_o
);

  input [0:0] lru_i;
  output [0:0] way_id_o;
  wire [0:0] way_id_o;
  assign way_id_o[0] = lru_i[0];

endmodule



module bsg_lru_pseudo_tree_decode_ways_p2
(
  way_id_i,
  data_o,
  mask_o
);

  input [0:0] way_id_i;
  output [0:0] data_o;
  output [0:0] mask_o;
  wire [0:0] data_o,mask_o;
  wire N0;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[0];

endmodule



module bsg_decode_num_out_p2
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bsg_cache_miss_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p2
(
  clk_i,
  reset_i,
  miss_v_i,
  decode_v_i,
  addr_v_i,
  tag_v_i,
  valid_v_i,
  lock_v_i,
  tag_hit_way_id_i,
  tag_hit_found_i,
  sbuf_empty_i,
  dma_cmd_o,
  dma_way_o,
  dma_addr_o,
  dma_done_i,
  stat_info_i,
  stat_mem_v_o,
  stat_mem_w_o,
  stat_mem_addr_o,
  stat_mem_data_o,
  stat_mem_w_mask_o,
  tag_mem_v_o,
  tag_mem_w_o,
  tag_mem_addr_o,
  tag_mem_data_o,
  tag_mem_w_mask_o,
  done_o,
  recover_o,
  chosen_way_o,
  ack_i
);

  input [15:0] decode_v_i;
  input [27:0] addr_v_i;
  input [35:0] tag_v_i;
  input [1:0] valid_v_i;
  input [1:0] lock_v_i;
  input [0:0] tag_hit_way_id_i;
  output [3:0] dma_cmd_o;
  output [0:0] dma_way_o;
  output [27:0] dma_addr_o;
  input [2:0] stat_info_i;
  output [5:0] stat_mem_addr_o;
  output [2:0] stat_mem_data_o;
  output [2:0] stat_mem_w_mask_o;
  output [5:0] tag_mem_addr_o;
  output [39:0] tag_mem_data_o;
  output [39:0] tag_mem_w_mask_o;
  output [0:0] chosen_way_o;
  input clk_i;
  input reset_i;
  input miss_v_i;
  input tag_hit_found_i;
  input sbuf_empty_i;
  input dma_done_i;
  input ack_i;
  output stat_mem_v_o;
  output stat_mem_w_o;
  output tag_mem_v_o;
  output tag_mem_w_o;
  output done_o;
  output recover_o;
  wire [3:0] dma_cmd_o,miss_state_n;
  wire [27:0] dma_addr_o;
  wire [5:0] stat_mem_addr_o,tag_mem_addr_o;
  wire [2:0] stat_mem_data_o,stat_mem_w_mask_o;
  wire [39:0] tag_mem_data_o,tag_mem_w_mask_o;
  wire [0:0] chosen_way_o,invalid_way_id,lru_way_id,chosen_way_lru_data,chosen_way_lru_mask,
  backup_lru_way_id;
  wire stat_mem_v_o,stat_mem_w_o,tag_mem_v_o,tag_mem_w_o,done_o,recover_o,N0,N1,N2,N3,
  N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,n_0_net__1_,
  n_0_net__0_,invalid_exist,goto_flush_op,goto_lock_op,n_2_net__1_,n_2_net__0_,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,
  N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159;
  wire [1:0] chosen_way_decode;
  reg [0:0] dma_way_o;
  reg [3:0] miss_state_r;
  assign dma_addr_o[0] = 1'b0;
  assign dma_addr_o[1] = 1'b0;
  assign tag_mem_addr_o[5] = addr_v_i[9];
  assign stat_mem_addr_o[5] = addr_v_i[9];
  assign tag_mem_addr_o[4] = addr_v_i[8];
  assign stat_mem_addr_o[4] = addr_v_i[8];
  assign tag_mem_addr_o[3] = addr_v_i[7];
  assign stat_mem_addr_o[3] = addr_v_i[7];
  assign tag_mem_addr_o[2] = addr_v_i[6];
  assign stat_mem_addr_o[2] = addr_v_i[6];
  assign tag_mem_addr_o[1] = addr_v_i[5];
  assign stat_mem_addr_o[1] = addr_v_i[5];
  assign tag_mem_addr_o[0] = addr_v_i[4];
  assign stat_mem_addr_o[0] = addr_v_i[4];
  assign dma_cmd_o[0] = tag_mem_data_o[39];
  assign tag_mem_data_o[19] = tag_mem_data_o[39];

  bsg_priority_encode_width_p2_lo_to_hi_p1
  invalid_way_pe
  (
    .i({ n_0_net__1_, n_0_net__0_ }),
    .addr_o(invalid_way_id[0]),
    .v_o(invalid_exist)
  );


  bsg_lru_pseudo_tree_encode_ways_p2
  lru_encode
  (
    .lru_i(stat_info_i[0]),
    .way_id_o(lru_way_id[0])
  );


  bsg_lru_pseudo_tree_decode_ways_p2
  chosen_way_lru_decode
  (
    .way_id_i(chosen_way_o[0]),
    .data_o(chosen_way_lru_data[0]),
    .mask_o(chosen_way_lru_mask[0])
  );


  bsg_priority_encode_width_p2_lo_to_hi_p1
  backup_lru_pe
  (
    .i({ n_2_net__1_, n_2_net__0_ }),
    .addr_o(backup_lru_way_id[0])
  );


  bsg_decode_num_out_p2
  chosen_way_demux
  (
    .i(chosen_way_o[0]),
    .o(chosen_way_decode)
  );

  assign N25 = N21 & N22;
  assign N26 = N23 & N24;
  assign N27 = N25 & N26;
  assign N28 = miss_state_r[3] | N22;
  assign N29 = miss_state_r[1] | miss_state_r[0];
  assign N30 = N28 | N29;
  assign N32 = miss_state_r[3] | miss_state_r[2];
  assign N33 = miss_state_r[1] | N24;
  assign N34 = N32 | N33;
  assign N36 = miss_state_r[3] | miss_state_r[2];
  assign N37 = N23 | miss_state_r[0];
  assign N38 = N36 | N37;
  assign N40 = miss_state_r[3] | miss_state_r[2];
  assign N41 = N23 | N24;
  assign N42 = N40 | N41;
  assign N44 = miss_state_r[3] | N22;
  assign N45 = miss_state_r[1] | N24;
  assign N46 = N44 | N45;
  assign N48 = miss_state_r[3] | N22;
  assign N49 = N23 | miss_state_r[0];
  assign N50 = N48 | N49;
  assign N52 = miss_state_r[3] | N22;
  assign N53 = N23 | N24;
  assign N54 = N52 | N53;
  assign N56 = N21 | miss_state_r[2];
  assign N57 = miss_state_r[1] | miss_state_r[0];
  assign N58 = N56 | N57;
  assign N60 = miss_state_r[3] & miss_state_r[0];
  assign N61 = miss_state_r[3] & miss_state_r[1];
  assign N62 = miss_state_r[3] & miss_state_r[2];
  assign N74 = (N73)? lock_v_i[0] : 
               (N0)? lock_v_i[1] : 1'b0;
  assign N0 = lru_way_id[0];
  assign N79 = (N78)? stat_info_i[1] : 
               (N1)? stat_info_i[2] : 1'b0;
  assign N1 = N77;
  assign N80 = (N78)? valid_v_i[0] : 
               (N1)? valid_v_i[1] : 1'b0;
  assign N92 = (N91)? stat_info_i[1] : 
               (N2)? stat_info_i[2] : 1'b0;
  assign N2 = N86;
  assign N93 = (N91)? valid_v_i[0] : 
               (N2)? valid_v_i[1] : 1'b0;
  assign N97 = (N96)? tag_v_i[17] : 
               (N3)? tag_v_i[35] : 1'b0;
  assign N3 = dma_way_o[0];
  assign N98 = (N96)? tag_v_i[16] : 
               (N3)? tag_v_i[34] : 1'b0;
  assign N99 = (N96)? tag_v_i[15] : 
               (N3)? tag_v_i[33] : 1'b0;
  assign N100 = (N96)? tag_v_i[14] : 
                (N3)? tag_v_i[32] : 1'b0;
  assign N101 = (N96)? tag_v_i[13] : 
                (N3)? tag_v_i[31] : 1'b0;
  assign N102 = (N96)? tag_v_i[12] : 
                (N3)? tag_v_i[30] : 1'b0;
  assign N103 = (N96)? tag_v_i[11] : 
                (N3)? tag_v_i[29] : 1'b0;
  assign N104 = (N96)? tag_v_i[10] : 
                (N3)? tag_v_i[28] : 1'b0;
  assign N105 = (N96)? tag_v_i[9] : 
                (N3)? tag_v_i[27] : 1'b0;
  assign N106 = (N96)? tag_v_i[8] : 
                (N3)? tag_v_i[26] : 1'b0;
  assign N107 = (N96)? tag_v_i[7] : 
                (N3)? tag_v_i[25] : 1'b0;
  assign N108 = (N96)? tag_v_i[6] : 
                (N3)? tag_v_i[24] : 1'b0;
  assign N109 = (N96)? tag_v_i[5] : 
                (N3)? tag_v_i[23] : 1'b0;
  assign N110 = (N96)? tag_v_i[4] : 
                (N3)? tag_v_i[22] : 1'b0;
  assign N111 = (N96)? tag_v_i[3] : 
                (N3)? tag_v_i[21] : 1'b0;
  assign N112 = (N96)? tag_v_i[2] : 
                (N3)? tag_v_i[20] : 1'b0;
  assign N113 = (N96)? tag_v_i[1] : 
                (N3)? tag_v_i[19] : 1'b0;
  assign N114 = (N96)? tag_v_i[0] : 
                (N3)? tag_v_i[18] : 1'b0;
  assign N116 = (N96)? tag_v_i[17] : 
                (N3)? tag_v_i[35] : 1'b0;
  assign N117 = (N96)? tag_v_i[16] : 
                (N3)? tag_v_i[34] : 1'b0;
  assign N118 = (N96)? tag_v_i[15] : 
                (N3)? tag_v_i[33] : 1'b0;
  assign N119 = (N96)? tag_v_i[14] : 
                (N3)? tag_v_i[32] : 1'b0;
  assign N120 = (N96)? tag_v_i[13] : 
                (N3)? tag_v_i[31] : 1'b0;
  assign N121 = (N96)? tag_v_i[12] : 
                (N3)? tag_v_i[30] : 1'b0;
  assign N122 = (N96)? tag_v_i[11] : 
                (N3)? tag_v_i[29] : 1'b0;
  assign N123 = (N96)? tag_v_i[10] : 
                (N3)? tag_v_i[28] : 1'b0;
  assign N124 = (N96)? tag_v_i[9] : 
                (N3)? tag_v_i[27] : 1'b0;
  assign N125 = (N96)? tag_v_i[8] : 
                (N3)? tag_v_i[26] : 1'b0;
  assign N126 = (N96)? tag_v_i[7] : 
                (N3)? tag_v_i[25] : 1'b0;
  assign N127 = (N96)? tag_v_i[6] : 
                (N3)? tag_v_i[24] : 1'b0;
  assign N128 = (N96)? tag_v_i[5] : 
                (N3)? tag_v_i[23] : 1'b0;
  assign N129 = (N96)? tag_v_i[4] : 
                (N3)? tag_v_i[22] : 1'b0;
  assign N130 = (N96)? tag_v_i[3] : 
                (N3)? tag_v_i[21] : 1'b0;
  assign N131 = (N96)? tag_v_i[2] : 
                (N3)? tag_v_i[20] : 1'b0;
  assign N132 = (N96)? tag_v_i[1] : 
                (N3)? tag_v_i[19] : 1'b0;
  assign N133 = (N96)? tag_v_i[0] : 
                (N3)? tag_v_i[18] : 1'b0;
  assign { N69, N68, N67 } = (N4)? { 1'b0, 1'b0, 1'b1 } : 
                             (N142)? { 1'b0, 1'b1, 1'b0 } : 
                             (N66)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N4 = goto_flush_op;
  assign { N72, N71, N70 } = (N5)? { N69, N68, N67 } : 
                             (N6)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = miss_v_i;
  assign N6 = N64;
  assign N77 = (N7)? invalid_way_id[0] : 
               (N144)? backup_lru_way_id[0] : 
               (N76)? lru_way_id[0] : 1'b0;
  assign N7 = invalid_exist;
  assign N82 = ~N81;
  assign { N84, N83 } = (N8)? { N82, N81 } : 
                        (N9)? { 1'b1, 1'b0 } : 1'b0;
  assign N8 = dma_done_i;
  assign N9 = N115;
  assign N86 = (N10)? addr_v_i[10] : 
               (N85)? tag_hit_way_id_i[0] : 1'b0;
  assign N10 = decode_v_i[8];
  assign N95 = ~N94;
  assign N135 = (N8)? N134 : 
                (N9)? 1'b1 : 1'b0;
  assign stat_mem_v_o = (N11)? miss_v_i : 
                        (N12)? dma_done_i : 
                        (N13)? 1'b1 : 
                        (N14)? 1'b0 : 
                        (N15)? 1'b0 : 
                        (N16)? 1'b0 : 
                        (N17)? 1'b0 : 
                        (N18)? 1'b0 : 
                        (N19)? 1'b0 : 
                        (N20)? 1'b0 : 1'b0;
  assign N11 = N27;
  assign N12 = tag_mem_data_o[39];
  assign N13 = N35;
  assign N14 = N39;
  assign N15 = dma_cmd_o[1];
  assign N16 = N47;
  assign N17 = N51;
  assign N18 = N55;
  assign N19 = N59;
  assign N20 = N63;
  assign miss_state_n = (N11)? { 1'b0, N72, N71, N70 } : 
                        (N12)? { 1'b0, N84, dma_done_i, N83 } : 
                        (N13)? { 1'b0, N95, 1'b1, 1'b1 } : 
                        (N14)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                        (N15)? { 1'b0, dma_done_i, N115, 1'b1 } : 
                        (N16)? { 1'b0, 1'b1, dma_done_i, N135 } : 
                        (N17)? { 1'b0, 1'b1, 1'b1, dma_done_i } : 
                        (N18)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                        (N19)? { N136, 1'b0, 1'b0, 1'b0 } : 
                        (N20)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign chosen_way_o[0] = (N11)? dma_way_o[0] : 
                           (N12)? N77 : 
                           (N13)? N86 : 
                           (N14)? tag_hit_way_id_i[0] : 
                           (N15)? dma_way_o[0] : 
                           (N16)? dma_way_o[0] : 
                           (N17)? dma_way_o[0] : 
                           (N18)? dma_way_o[0] : 
                           (N19)? dma_way_o[0] : 
                           (N20)? dma_way_o[0] : 1'b0;
  assign dma_cmd_o[2] = (N17)? sbuf_empty_i : 
                        (N139)? 1'b0 : 1'b0;
  assign dma_cmd_o[3] = (N16)? sbuf_empty_i : 
                        (N140)? 1'b0 : 1'b0;
  assign dma_addr_o[3:2] = (N17)? addr_v_i[3:2] : 
                           (N139)? { 1'b0, 1'b0 } : 1'b0;
  assign dma_addr_o[27:4] = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N12)? addr_v_i[27:4] : 
                            (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N15)? { N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, addr_v_i[9:4] } : 
                            (N16)? { N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, addr_v_i[9:4] } : 
                            (N17)? addr_v_i[27:4] : 
                            (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_o = (N11)? 1'b0 : 
                        (N12)? dma_done_i : 
                        (N13)? 1'b1 : 
                        (N14)? 1'b0 : 
                        (N15)? 1'b0 : 
                        (N16)? 1'b0 : 
                        (N17)? 1'b0 : 
                        (N18)? 1'b0 : 
                        (N19)? 1'b0 : 
                        (N20)? 1'b0 : 1'b0;
  assign stat_mem_data_o = (N11)? { 1'b0, 1'b0, 1'b0 } : 
                           (N12)? { decode_v_i[10:10], decode_v_i[10:10], chosen_way_lru_data[0:0] } : 
                           (N13)? { 1'b0, 1'b0, 1'b0 } : 
                           (N14)? { 1'b0, 1'b0, 1'b0 } : 
                           (N15)? { 1'b0, 1'b0, 1'b0 } : 
                           (N16)? { 1'b0, 1'b0, 1'b0 } : 
                           (N17)? { 1'b0, 1'b0, 1'b0 } : 
                           (N18)? { 1'b0, 1'b0, 1'b0 } : 
                           (N19)? { 1'b0, 1'b0, 1'b0 } : 
                           (N20)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_mask_o = (N11)? { 1'b0, 1'b0, 1'b0 } : 
                             (N12)? { chosen_way_decode, chosen_way_lru_mask[0:0] } : 
                             (N13)? { chosen_way_decode, 1'b0 } : 
                             (N14)? { 1'b0, 1'b0, 1'b0 } : 
                             (N15)? { 1'b0, 1'b0, 1'b0 } : 
                             (N16)? { 1'b0, 1'b0, 1'b0 } : 
                             (N17)? { 1'b0, 1'b0, 1'b0 } : 
                             (N18)? { 1'b0, 1'b0, 1'b0 } : 
                             (N19)? { 1'b0, 1'b0, 1'b0 } : 
                             (N20)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_v_o = (N11)? 1'b0 : 
                       (N12)? dma_done_i : 
                       (N13)? 1'b1 : 
                       (N14)? 1'b1 : 
                       (N15)? 1'b0 : 
                       (N16)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N20)? 1'b0 : 1'b0;
  assign tag_mem_w_o = (N11)? 1'b0 : 
                       (N12)? dma_done_i : 
                       (N13)? 1'b1 : 
                       (N14)? 1'b1 : 
                       (N15)? 1'b0 : 
                       (N16)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N20)? 1'b0 : 1'b0;
  assign { tag_mem_w_mask_o[37:20], tag_mem_w_mask_o[17:0] } = (N12)? { chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode, chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                                                               (N138)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { tag_mem_w_mask_o[39:38], tag_mem_w_mask_o[19:18] } = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N12)? { chosen_way_decode[1:1], chosen_way_decode, chosen_way_decode[0:0] } : 
                                                                (N13)? { N89, N90, N87, N88 } : 
                                                                (N14)? { 1'b0, chosen_way_decode[1:1], 1'b0, chosen_way_decode[0:0] } : 
                                                                (N15)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N16)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N17)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N18)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N19)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N20)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { tag_mem_data_o[37:20], tag_mem_data_o[17:0] } = (N12)? { addr_v_i[27:10], addr_v_i[27:10] } : 
                                                           (N138)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { tag_mem_data_o[38:38], tag_mem_data_o[18:18] } = (N11)? { 1'b0, 1'b0 } : 
                                                            (N12)? { decode_v_i[2:2], decode_v_i[2:2] } : 
                                                            (N13)? { 1'b0, 1'b0 } : 
                                                            (N14)? { decode_v_i[2:2], decode_v_i[2:2] } : 
                                                            (N15)? { 1'b0, 1'b0 } : 
                                                            (N16)? { 1'b0, 1'b0 } : 
                                                            (N17)? { 1'b0, 1'b0 } : 
                                                            (N18)? { 1'b0, 1'b0 } : 
                                                            (N19)? { 1'b0, 1'b0 } : 
                                                            (N20)? { 1'b0, 1'b0 } : 1'b0;
  assign recover_o = (N11)? 1'b0 : 
                     (N12)? 1'b0 : 
                     (N13)? 1'b0 : 
                     (N14)? 1'b0 : 
                     (N15)? 1'b0 : 
                     (N16)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N18)? 1'b1 : 
                     (N19)? 1'b0 : 
                     (N20)? 1'b0 : 1'b0;
  assign done_o = (N11)? 1'b0 : 
                  (N12)? 1'b0 : 
                  (N13)? 1'b0 : 
                  (N14)? 1'b0 : 
                  (N15)? 1'b0 : 
                  (N16)? 1'b0 : 
                  (N17)? 1'b0 : 
                  (N18)? 1'b0 : 
                  (N19)? 1'b1 : 
                  (N20)? 1'b0 : 1'b0;
  assign n_0_net__1_ = N145 & N146;
  assign N145 = ~valid_v_i[1];
  assign N146 = ~lock_v_i[1];
  assign n_0_net__0_ = N147 & N148;
  assign N147 = ~valid_v_i[0];
  assign N148 = ~lock_v_i[0];
  assign goto_flush_op = N150 | decode_v_i[4];
  assign N150 = N149 | decode_v_i[5];
  assign N149 = decode_v_i[8] | decode_v_i[3];
  assign goto_lock_op = decode_v_i[1] | N151;
  assign N151 = decode_v_i[2] & tag_hit_found_i;
  assign n_2_net__1_ = ~lock_v_i[1];
  assign n_2_net__0_ = ~lock_v_i[0];
  assign N21 = ~miss_state_r[3];
  assign N22 = ~miss_state_r[2];
  assign N23 = ~miss_state_r[1];
  assign N24 = ~miss_state_r[0];
  assign N31 = ~N30;
  assign N35 = ~N34;
  assign N39 = ~N38;
  assign N43 = ~N42;
  assign N47 = ~N46;
  assign N51 = ~N50;
  assign N55 = ~N54;
  assign N59 = ~N58;
  assign N63 = N60 | N152;
  assign N152 = N61 | N62;
  assign tag_mem_data_o[39] = N31;
  assign dma_cmd_o[1] = N43;
  assign N64 = ~miss_v_i;
  assign N65 = goto_lock_op | goto_flush_op;
  assign N66 = ~N65;
  assign N73 = ~lru_way_id[0];
  assign N75 = N74 | invalid_exist;
  assign N76 = ~N75;
  assign N78 = ~N77;
  assign N81 = N79 & N80;
  assign N85 = ~decode_v_i[8];
  assign N87 = N153 & chosen_way_decode[0];
  assign N153 = decode_v_i[3] | decode_v_i[4];
  assign N88 = N154 & chosen_way_decode[0];
  assign N154 = decode_v_i[3] | decode_v_i[4];
  assign N89 = N155 & chosen_way_decode[1];
  assign N155 = decode_v_i[3] | decode_v_i[4];
  assign N90 = N156 & chosen_way_decode[1];
  assign N156 = decode_v_i[3] | decode_v_i[4];
  assign N91 = ~N86;
  assign N94 = N158 & N93;
  assign N158 = N157 & N92;
  assign N157 = ~decode_v_i[3];
  assign N96 = ~dma_way_o[0];
  assign N115 = ~dma_done_i;
  assign N134 = N159 | decode_v_i[5];
  assign N159 = decode_v_i[8] | decode_v_i[4];
  assign N136 = ~ack_i;
  assign N137 = ~tag_mem_data_o[39];
  assign N138 = N137;
  assign N139 = N50;
  assign N140 = N46;
  assign N141 = ~goto_flush_op;
  assign N142 = goto_lock_op & N141;
  assign N143 = ~invalid_exist;
  assign N144 = N74 & N143;

  always @(posedge clk_i) begin
    if(reset_i) begin
      { dma_way_o[0:0] } <= { 1'b0 };
      { miss_state_r[3:0] } <= { 1'b0, 1'b0, 1'b0, 1'b0 };
    end else if(1'b1) begin
      { dma_way_o[0:0] } <= { chosen_way_o[0:0] };
      { miss_state_r[3:0] } <= { miss_state_n[3:0] };
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p4
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [2:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  reg [2:0] count_o;
  assign { N8, N7, N6 } = { N14, N13, N12 } + up_i;
  assign { N11, N10, N9 } = (N0)? { 1'b0, 1'b0, 1'b0 } : 
                            (N1)? { N8, N7, N6 } : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign { N14, N13, N12 } = count_o * N4;
  assign N2 = ~reset_i;
  assign N3 = N2;
  assign N4 = ~clear_i;
  assign N5 = N3 & N4;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { count_o[2:0] } <= { N11, N10, N9 };
    end 
  end


endmodule



module bsg_circular_ptr_slots_p4_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] n_o,genblk1_genblk1_ptr_r_p1;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  reg [1:0] o;
  assign genblk1_genblk1_ptr_r_p1 = o + 1'b1;
  assign { N6, N5 } = (N0)? { 1'b0, 1'b0 } : 
                      (N1)? n_o : 1'b0;
  assign N0 = reset_i;
  assign N1 = N4;
  assign n_o = (N2)? genblk1_genblk1_ptr_r_p1 : 
               (N3)? o : 1'b0;
  assign N2 = add_i[0];
  assign N3 = N7;
  assign N4 = ~reset_i;
  assign N7 = ~add_i[0];

  always @(posedge clk) begin
    if(1'b1) begin
      { o[1:0] } <= { N6, N5 };
    end 
  end


endmodule



module bsg_fifo_tracker_els_p4
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,equal_ptrs,SYNOPSYS_UNCONNECTED_1,
  SYNOPSYS_UNCONNECTED_2;
  reg deq_r,enq_r;

  bsg_circular_ptr_slots_p4_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p4_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N5 = (N0)? 1'b1 : 
              (N9)? 1'b1 : 
              (N4)? 1'b0 : 1'b0;
  assign N0 = N2;
  assign N6 = (N0)? 1'b0 : 
              (N9)? enq_i : 1'b0;
  assign N7 = (N0)? 1'b1 : 
              (N9)? deq_i : 1'b0;
  assign N1 = enq_i | deq_i;
  assign N2 = reset_i;
  assign N3 = N1 | N2;
  assign N4 = ~N3;
  assign N8 = ~N2;
  assign N9 = N1 & N8;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(N5) begin
      deq_r <= N7;
      enq_r <= N6;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p4_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;
  reg [127:0] mem;
  assign r_data_o[31] = (N8)? mem[31] : 
                        (N10)? mem[63] : 
                        (N9)? mem[95] : 
                        (N11)? mem[127] : 1'b0;
  assign r_data_o[30] = (N8)? mem[30] : 
                        (N10)? mem[62] : 
                        (N9)? mem[94] : 
                        (N11)? mem[126] : 1'b0;
  assign r_data_o[29] = (N8)? mem[29] : 
                        (N10)? mem[61] : 
                        (N9)? mem[93] : 
                        (N11)? mem[125] : 1'b0;
  assign r_data_o[28] = (N8)? mem[28] : 
                        (N10)? mem[60] : 
                        (N9)? mem[92] : 
                        (N11)? mem[124] : 1'b0;
  assign r_data_o[27] = (N8)? mem[27] : 
                        (N10)? mem[59] : 
                        (N9)? mem[91] : 
                        (N11)? mem[123] : 1'b0;
  assign r_data_o[26] = (N8)? mem[26] : 
                        (N10)? mem[58] : 
                        (N9)? mem[90] : 
                        (N11)? mem[122] : 1'b0;
  assign r_data_o[25] = (N8)? mem[25] : 
                        (N10)? mem[57] : 
                        (N9)? mem[89] : 
                        (N11)? mem[121] : 1'b0;
  assign r_data_o[24] = (N8)? mem[24] : 
                        (N10)? mem[56] : 
                        (N9)? mem[88] : 
                        (N11)? mem[120] : 1'b0;
  assign r_data_o[23] = (N8)? mem[23] : 
                        (N10)? mem[55] : 
                        (N9)? mem[87] : 
                        (N11)? mem[119] : 1'b0;
  assign r_data_o[22] = (N8)? mem[22] : 
                        (N10)? mem[54] : 
                        (N9)? mem[86] : 
                        (N11)? mem[118] : 1'b0;
  assign r_data_o[21] = (N8)? mem[21] : 
                        (N10)? mem[53] : 
                        (N9)? mem[85] : 
                        (N11)? mem[117] : 1'b0;
  assign r_data_o[20] = (N8)? mem[20] : 
                        (N10)? mem[52] : 
                        (N9)? mem[84] : 
                        (N11)? mem[116] : 1'b0;
  assign r_data_o[19] = (N8)? mem[19] : 
                        (N10)? mem[51] : 
                        (N9)? mem[83] : 
                        (N11)? mem[115] : 1'b0;
  assign r_data_o[18] = (N8)? mem[18] : 
                        (N10)? mem[50] : 
                        (N9)? mem[82] : 
                        (N11)? mem[114] : 1'b0;
  assign r_data_o[17] = (N8)? mem[17] : 
                        (N10)? mem[49] : 
                        (N9)? mem[81] : 
                        (N11)? mem[113] : 1'b0;
  assign r_data_o[16] = (N8)? mem[16] : 
                        (N10)? mem[48] : 
                        (N9)? mem[80] : 
                        (N11)? mem[112] : 1'b0;
  assign r_data_o[15] = (N8)? mem[15] : 
                        (N10)? mem[47] : 
                        (N9)? mem[79] : 
                        (N11)? mem[111] : 1'b0;
  assign r_data_o[14] = (N8)? mem[14] : 
                        (N10)? mem[46] : 
                        (N9)? mem[78] : 
                        (N11)? mem[110] : 1'b0;
  assign r_data_o[13] = (N8)? mem[13] : 
                        (N10)? mem[45] : 
                        (N9)? mem[77] : 
                        (N11)? mem[109] : 1'b0;
  assign r_data_o[12] = (N8)? mem[12] : 
                        (N10)? mem[44] : 
                        (N9)? mem[76] : 
                        (N11)? mem[108] : 1'b0;
  assign r_data_o[11] = (N8)? mem[11] : 
                        (N10)? mem[43] : 
                        (N9)? mem[75] : 
                        (N11)? mem[107] : 1'b0;
  assign r_data_o[10] = (N8)? mem[10] : 
                        (N10)? mem[42] : 
                        (N9)? mem[74] : 
                        (N11)? mem[106] : 1'b0;
  assign r_data_o[9] = (N8)? mem[9] : 
                       (N10)? mem[41] : 
                       (N9)? mem[73] : 
                       (N11)? mem[105] : 1'b0;
  assign r_data_o[8] = (N8)? mem[8] : 
                       (N10)? mem[40] : 
                       (N9)? mem[72] : 
                       (N11)? mem[104] : 1'b0;
  assign r_data_o[7] = (N8)? mem[7] : 
                       (N10)? mem[39] : 
                       (N9)? mem[71] : 
                       (N11)? mem[103] : 1'b0;
  assign r_data_o[6] = (N8)? mem[6] : 
                       (N10)? mem[38] : 
                       (N9)? mem[70] : 
                       (N11)? mem[102] : 1'b0;
  assign r_data_o[5] = (N8)? mem[5] : 
                       (N10)? mem[37] : 
                       (N9)? mem[69] : 
                       (N11)? mem[101] : 1'b0;
  assign r_data_o[4] = (N8)? mem[4] : 
                       (N10)? mem[36] : 
                       (N9)? mem[68] : 
                       (N11)? mem[100] : 1'b0;
  assign r_data_o[3] = (N8)? mem[3] : 
                       (N10)? mem[35] : 
                       (N9)? mem[67] : 
                       (N11)? mem[99] : 1'b0;
  assign r_data_o[2] = (N8)? mem[2] : 
                       (N10)? mem[34] : 
                       (N9)? mem[66] : 
                       (N11)? mem[98] : 1'b0;
  assign r_data_o[1] = (N8)? mem[1] : 
                       (N10)? mem[33] : 
                       (N9)? mem[65] : 
                       (N11)? mem[97] : 1'b0;
  assign r_data_o[0] = (N8)? mem[0] : 
                       (N10)? mem[32] : 
                       (N9)? mem[64] : 
                       (N11)? mem[96] : 1'b0;
  assign N16 = w_addr_i[0] & w_addr_i[1];
  assign N15 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N14 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N13 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign { N20, N19, N18, N17 } = (N4)? { N16, N15, N14, N13 } : 
                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = w_v_i;
  assign N5 = N12;
  assign N6 = ~r_addr_i[0];
  assign N7 = ~r_addr_i[1];
  assign N8 = N6 & N7;
  assign N9 = N6 & r_addr_i[1];
  assign N10 = r_addr_i[0] & N7;
  assign N11 = r_addr_i[0] & r_addr_i[1];
  assign N12 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N20) begin
      { mem[127:96] } <= { w_data_i[31:0] };
    end 
    if(N19) begin
      { mem[95:64] } <= { w_data_i[31:0] };
    end 
    if(N18) begin
      { mem[63:32] } <= { w_data_i[31:0] };
    end 
    if(N17) begin
      { mem[31:0] } <= { w_data_i[31:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p4_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p4_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p32_els_p4_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enque,full,empty,SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p4
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p32_els_p4_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_o;
  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p32_els_p4
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p32_els_p4_ready_THEN_valid_p0
  unhardened_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [63:0] mem;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[62] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[61] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[60] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[59] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[58] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[57] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[56] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[55] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[45] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[44] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[43] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[42] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[41] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[40] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[39] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[38] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[37] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[36] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[35] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[34] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[33] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[63:32] } <= { w_data_i[31:0] };
    end 
    if(N7) begin
      { mem[31:0] } <= { w_data_i[31:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bsg_mux_width_p32_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [0:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[63] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[62] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[61] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[60] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[59] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[58] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[57] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[56] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[55] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[54] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[53] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[52] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[51] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[50] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[49] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[48] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[47] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[46] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[45] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[44] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[43] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[42] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[41] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[40] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[39] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[38] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[37] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[36] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[35] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[34] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[33] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[32] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_cache_dma_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p2_debug_p0
(
  clk_i,
  reset_i,
  dma_cmd_i,
  dma_way_i,
  dma_addr_i,
  done_o,
  snoop_word_o,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  data_mem_v_o,
  data_mem_w_o,
  data_mem_addr_o,
  data_mem_w_mask_o,
  data_mem_data_o,
  data_mem_data_i,
  dma_evict_o
);

  input [3:0] dma_cmd_i;
  input [0:0] dma_way_i;
  input [27:0] dma_addr_i;
  output [31:0] snoop_word_o;
  output [28:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  output [7:0] data_mem_addr_o;
  output [7:0] data_mem_w_mask_o;
  output [63:0] data_mem_data_o;
  input [63:0] data_mem_data_i;
  input clk_i;
  input reset_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output done_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output data_mem_v_o;
  output data_mem_w_o;
  output dma_evict_o;
  wire [28:0] dma_pkt_o;
  wire [31:0] dma_data_o,out_fifo_data_li;
  wire [7:0] data_mem_addr_o,data_mem_w_mask_o;
  wire [63:0] data_mem_data_o;
  wire done_o,dma_pkt_v_o,dma_data_ready_o,dma_data_v_o,data_mem_v_o,data_mem_w_o,
  dma_evict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,counter_clear,counter_up,in_fifo_v_lo,
  in_fifo_yumi_li,out_fifo_v_li,out_fifo_ready_lo,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,snoop_word_we,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76;
  wire [2:2] counter_r;
  wire [1:0] dma_state_n;
  reg [31:0] snoop_word_o;
  reg [1:0] dma_state_r;
  assign dma_pkt_o[0] = 1'b0;
  assign dma_pkt_o[1] = 1'b0;
  assign dma_pkt_o[2] = 1'b0;
  assign dma_pkt_o[3] = 1'b0;
  assign dma_pkt_o[27] = dma_addr_i[27];
  assign dma_pkt_o[26] = dma_addr_i[26];
  assign dma_pkt_o[25] = dma_addr_i[25];
  assign dma_pkt_o[24] = dma_addr_i[24];
  assign dma_pkt_o[23] = dma_addr_i[23];
  assign dma_pkt_o[22] = dma_addr_i[22];
  assign dma_pkt_o[21] = dma_addr_i[21];
  assign dma_pkt_o[20] = dma_addr_i[20];
  assign dma_pkt_o[19] = dma_addr_i[19];
  assign dma_pkt_o[18] = dma_addr_i[18];
  assign dma_pkt_o[17] = dma_addr_i[17];
  assign dma_pkt_o[16] = dma_addr_i[16];
  assign dma_pkt_o[15] = dma_addr_i[15];
  assign dma_pkt_o[14] = dma_addr_i[14];
  assign dma_pkt_o[13] = dma_addr_i[13];
  assign dma_pkt_o[12] = dma_addr_i[12];
  assign dma_pkt_o[11] = dma_addr_i[11];
  assign dma_pkt_o[10] = dma_addr_i[10];
  assign dma_pkt_o[9] = dma_addr_i[9];
  assign data_mem_addr_o[7] = dma_addr_i[9];
  assign dma_pkt_o[8] = dma_addr_i[8];
  assign data_mem_addr_o[6] = dma_addr_i[8];
  assign dma_pkt_o[7] = dma_addr_i[7];
  assign data_mem_addr_o[5] = dma_addr_i[7];
  assign dma_pkt_o[6] = dma_addr_i[6];
  assign data_mem_addr_o[4] = dma_addr_i[6];
  assign dma_pkt_o[5] = dma_addr_i[5];
  assign data_mem_addr_o[3] = dma_addr_i[5];
  assign dma_pkt_o[4] = dma_addr_i[4];
  assign data_mem_addr_o[2] = dma_addr_i[4];
  assign data_mem_w_mask_o[4] = data_mem_w_mask_o[7];
  assign data_mem_w_mask_o[5] = data_mem_w_mask_o[7];
  assign data_mem_w_mask_o[6] = data_mem_w_mask_o[7];
  assign data_mem_w_mask_o[0] = data_mem_w_mask_o[3];
  assign data_mem_w_mask_o[1] = data_mem_w_mask_o[3];
  assign data_mem_w_mask_o[2] = data_mem_w_mask_o[3];
  assign data_mem_data_o[31] = data_mem_data_o[63];
  assign data_mem_data_o[30] = data_mem_data_o[62];
  assign data_mem_data_o[29] = data_mem_data_o[61];
  assign data_mem_data_o[28] = data_mem_data_o[60];
  assign data_mem_data_o[27] = data_mem_data_o[59];
  assign data_mem_data_o[26] = data_mem_data_o[58];
  assign data_mem_data_o[25] = data_mem_data_o[57];
  assign data_mem_data_o[24] = data_mem_data_o[56];
  assign data_mem_data_o[23] = data_mem_data_o[55];
  assign data_mem_data_o[22] = data_mem_data_o[54];
  assign data_mem_data_o[21] = data_mem_data_o[53];
  assign data_mem_data_o[20] = data_mem_data_o[52];
  assign data_mem_data_o[19] = data_mem_data_o[51];
  assign data_mem_data_o[18] = data_mem_data_o[50];
  assign data_mem_data_o[17] = data_mem_data_o[49];
  assign data_mem_data_o[16] = data_mem_data_o[48];
  assign data_mem_data_o[15] = data_mem_data_o[47];
  assign data_mem_data_o[14] = data_mem_data_o[46];
  assign data_mem_data_o[13] = data_mem_data_o[45];
  assign data_mem_data_o[12] = data_mem_data_o[44];
  assign data_mem_data_o[11] = data_mem_data_o[43];
  assign data_mem_data_o[10] = data_mem_data_o[42];
  assign data_mem_data_o[9] = data_mem_data_o[41];
  assign data_mem_data_o[8] = data_mem_data_o[40];
  assign data_mem_data_o[7] = data_mem_data_o[39];
  assign data_mem_data_o[6] = data_mem_data_o[38];
  assign data_mem_data_o[5] = data_mem_data_o[37];
  assign data_mem_data_o[4] = data_mem_data_o[36];
  assign data_mem_data_o[3] = data_mem_data_o[35];
  assign data_mem_data_o[2] = data_mem_data_o[34];
  assign data_mem_data_o[1] = data_mem_data_o[33];
  assign data_mem_data_o[0] = data_mem_data_o[32];

  bsg_counter_clear_up_max_val_p4
  dma_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(counter_clear),
    .up_i(counter_up),
    .count_o({ counter_r[2:2], data_mem_addr_o[1:0] })
  );


  bsg_fifo_1r1w_small_width_p32_els_p4
  in_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(dma_data_v_i),
    .ready_o(dma_data_ready_o),
    .data_i(dma_data_i),
    .v_o(in_fifo_v_lo),
    .data_o(data_mem_data_o[63:32]),
    .yumi_i(in_fifo_yumi_li)
  );


  bsg_two_fifo_width_p32
  out_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(out_fifo_ready_lo),
    .data_i(out_fifo_data_li),
    .v_i(out_fifo_v_li),
    .v_o(dma_data_v_o),
    .data_o(dma_data_o),
    .yumi_i(dma_data_yumi_i)
  );


  bsg_decode_num_out_p2
  dma_way_demux
  (
    .i(dma_way_i[0]),
    .o({ data_mem_w_mask_o[7:7], data_mem_w_mask_o[3:3] })
  );


  bsg_mux_width_p32_els_p2
  write_data_mux
  (
    .data_i(data_mem_data_i),
    .sel_i(dma_way_i[0]),
    .data_o(out_fifo_data_li)
  );

  assign N12 = N11 & N64;
  assign N13 = dma_state_r[1] | N64;
  assign N15 = N11 | dma_state_r[0];
  assign N17 = dma_state_r[1] & dma_state_r[0];
  assign N18 = dma_cmd_i[1] | N35;
  assign N19 = N21 | N18;
  assign N21 = dma_cmd_i[3] | dma_cmd_i[2];
  assign N22 = N34 | dma_cmd_i[0];
  assign N23 = N21 | N22;
  assign N25 = dma_cmd_i[3] | N33;
  assign N26 = N25 | N29;
  assign N28 = N32 | dma_cmd_i[2];
  assign N29 = dma_cmd_i[1] | dma_cmd_i[0];
  assign N30 = N28 | N29;
  assign N36 = N32 & N33;
  assign N37 = N34 & N35;
  assign N38 = N36 & N37;
  assign N60 = dma_addr_i[3:2] == data_mem_addr_o[1:0];
  assign N64 = ~dma_state_r[0];
  assign N65 = N64 | dma_state_r[1];
  assign N66 = ~N65;
  assign N67 = ~counter_r[2];
  assign N68 = data_mem_addr_o[1] | N67;
  assign N69 = data_mem_addr_o[0] | N68;
  assign N70 = ~N69;
  assign N71 = ~data_mem_addr_o[1];
  assign N72 = ~data_mem_addr_o[0];
  assign N73 = N71 | counter_r[2];
  assign N74 = N72 | N73;
  assign N75 = ~N74;
  assign N44 = (N0)? 1'b1 : 
               (N1)? 1'b1 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N0 = N20;
  assign N1 = N24;
  assign N2 = N27;
  assign N3 = N31;
  assign N4 = N38;
  assign N45 = (N0)? 1'b0 : 
               (N1)? 1'b1 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N46 = (N0)? dma_pkt_yumi_i : 
               (N1)? dma_pkt_yumi_i : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N47 = (N0)? 1'b0 : 
               (N1)? 1'b0 : 
               (N2)? 1'b1 : 
               (N3)? 1'b1 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N48 = (N0)? 1'b0 : 
               (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b1 : 
               (N4)? 1'b0 : 
               (N43)? 1'b0 : 1'b0;
  assign N50 = ~N49;
  assign N55 = ~N54;
  assign counter_clear = (N5)? N47 : 
                         (N6)? N52 : 
                         (N7)? N57 : 
                         (N8)? 1'b0 : 1'b0;
  assign N5 = N12;
  assign N6 = N14;
  assign N7 = N16;
  assign N8 = N17;
  assign counter_up = (N5)? N48 : 
                      (N6)? N51 : 
                      (N7)? N56 : 
                      (N8)? 1'b0 : 1'b0;
  assign data_mem_v_o = (N5)? N48 : 
                        (N6)? in_fifo_v_lo : 
                        (N7)? N58 : 
                        (N8)? 1'b0 : 1'b0;
  assign dma_pkt_v_o = (N5)? N44 : 
                       (N6)? 1'b0 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b0 : 1'b0;
  assign dma_pkt_o[28] = (N5)? N45 : 
                         (N6)? 1'b0 : 
                         (N7)? 1'b0 : 
                         (N8)? 1'b0 : 1'b0;
  assign done_o = (N5)? N46 : 
                  (N6)? N53 : 
                  (N7)? N59 : 
                  (N8)? 1'b0 : 1'b0;
  assign dma_state_n = (N5)? { N31, N27 } : 
                       (N6)? { 1'b0, N50 } : 
                       (N7)? { N55, 1'b0 } : 
                       (N8)? { 1'b0, 1'b0 } : 1'b0;
  assign data_mem_w_o = (N5)? 1'b0 : 
                        (N6)? in_fifo_v_lo : 
                        (N7)? 1'b0 : 
                        (N8)? 1'b0 : 1'b0;
  assign in_fifo_yumi_li = (N5)? 1'b0 : 
                           (N6)? in_fifo_v_lo : 
                           (N7)? 1'b0 : 
                           (N8)? 1'b0 : 1'b0;
  assign out_fifo_v_li = (N5)? 1'b0 : 
                         (N6)? 1'b0 : 
                         (N7)? 1'b1 : 
                         (N8)? 1'b0 : 1'b0;
  assign dma_evict_o = (N5)? 1'b0 : 
                       (N6)? 1'b0 : 
                       (N7)? 1'b1 : 
                       (N8)? 1'b0 : 1'b0;
  assign N63 = (N9)? 1'b0 : 
               (N10)? snoop_word_we : 1'b0;
  assign N9 = N62;
  assign N10 = N61;
  assign N11 = ~dma_state_r[1];
  assign N14 = ~N13;
  assign N16 = ~N15;
  assign N20 = ~N19;
  assign N24 = ~N23;
  assign N27 = ~N26;
  assign N31 = ~N30;
  assign N32 = ~dma_cmd_i[3];
  assign N33 = ~dma_cmd_i[2];
  assign N34 = ~dma_cmd_i[1];
  assign N35 = ~dma_cmd_i[0];
  assign N39 = N24 | N20;
  assign N40 = N27 | N39;
  assign N41 = N31 | N40;
  assign N42 = N38 | N41;
  assign N43 = ~N42;
  assign N49 = N75 & in_fifo_v_lo;
  assign N51 = in_fifo_v_lo & N74;
  assign N52 = in_fifo_v_lo & N75;
  assign N53 = N75 & in_fifo_v_lo;
  assign N54 = N70 & out_fifo_ready_lo;
  assign N56 = out_fifo_ready_lo & N69;
  assign N57 = out_fifo_ready_lo & N70;
  assign N58 = out_fifo_ready_lo & N69;
  assign N59 = N70 & out_fifo_ready_lo;
  assign snoop_word_we = N76 & in_fifo_v_lo;
  assign N76 = N66 & N60;
  assign N61 = ~reset_i;
  assign N62 = reset_i;

  always @(posedge clk_i) begin
    if(N63) begin
      { snoop_word_o[31:0] } <= { data_mem_data_o[63:32] };
    end 
    if(reset_i) begin
      { dma_state_r[1:0] } <= { 1'b0, 1'b0 };
    end else if(1'b1) begin
      { dma_state_r[1:0] } <= { dma_state_n[1:0] };
    end 
  end


endmodule



module bsg_cache_sbuf_queue_width_p65
(
  clk_i,
  data_i,
  el0_en_i,
  el1_en_i,
  mux0_sel_i,
  mux1_sel_i,
  el0_snoop_o,
  el1_snoop_o,
  data_o
);

  input [64:0] data_i;
  output [64:0] el0_snoop_o;
  output [64:0] el1_snoop_o;
  output [64:0] data_o;
  input clk_i;
  input el0_en_i;
  input el1_en_i;
  input mux0_sel_i;
  input mux1_sel_i;
  wire [64:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70;
  reg [64:0] el0_snoop_o,el1_snoop_o;
  assign { N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 } = (N0)? el0_snoop_o : 
                                                                                                                                                                                                                                                                                                                                              (N1)? data_i : 1'b0;
  assign N0 = mux0_sel_i;
  assign N1 = N4;
  assign data_o = (N2)? el1_snoop_o : 
                  (N3)? data_i : 1'b0;
  assign N2 = mux1_sel_i;
  assign N3 = N70;
  assign N4 = ~mux0_sel_i;
  assign N70 = ~mux1_sel_i;

  always @(posedge clk_i) begin
    if(el0_en_i) begin
      { el0_snoop_o[64:0] } <= { data_i[64:0] };
    end 
    if(el1_en_i) begin
      { el1_snoop_o[64:0] } <= { N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 };
    end 
  end


endmodule



module bsg_mux_segmented_segments_p4_segment_width_p8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [31:0] data0_i;
  input [31:0] data1_i;
  input [3:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  assign data_o[7:0] = (N0)? data1_i[7:0] : 
                       (N4)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] : 
                        (N5)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] : 
                         (N6)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] : 
                         (N7)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign N4 = ~sel_i[0];
  assign N5 = ~sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = ~sel_i[3];

endmodule



module bsg_cache_sbuf_data_width_p32_addr_width_p28_ways_p2
(
  clk_i,
  reset_i,
  sbuf_entry_i,
  v_i,
  sbuf_entry_o,
  v_o,
  yumi_i,
  empty_o,
  bypass_addr_i,
  bypass_v_i,
  bypass_data_o,
  bypass_mask_o
);

  input [64:0] sbuf_entry_i;
  output [64:0] sbuf_entry_o;
  input [27:0] bypass_addr_i;
  output [31:0] bypass_data_o;
  output [3:0] bypass_mask_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input bypass_v_i;
  output v_o;
  output empty_o;
  wire [64:0] sbuf_entry_o,el0,el1;
  wire v_o,empty_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,el0_valid,el1_valid,
  el0_enable,N14,el1_enable,mux0_sel,mux1_sel,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,tag_hit0_n,tag_hit1_n,tag_hit2_n,n_2_net__3_,n_2_net__2_,n_2_net__1_,
  n_2_net__0_,n_4_net__3_,n_4_net__2_,n_4_net__1_,n_4_net__0_,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83;
  wire [3:3] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  wire [3:0] bypass_mask_n;
  wire [31:0] el0or1_data,bypass_data_n;
  reg [1:0] num_els_r;
  reg [31:0] bypass_data_o;
  reg [3:0] bypass_mask_o;
  assign N8 = N6 & N7;
  assign N9 = num_els_r[1] | N7;
  assign N11 = N6 | num_els_r[0];
  assign N13 = num_els_r[1] & num_els_r[0];

  bsg_cache_sbuf_queue_width_p65
  sbq
  (
    .clk_i(clk_i),
    .data_i(sbuf_entry_i),
    .el0_en_i(el0_enable),
    .el1_en_i(el1_enable),
    .mux0_sel_i(mux0_sel),
    .mux1_sel_i(mux1_sel),
    .el0_snoop_o(el0),
    .el1_snoop_o(el1),
    .data_o(sbuf_entry_o)
  );

  assign tag_hit0_n = bypass_addr_i[27:2] == el0[64:39];
  assign tag_hit1_n = bypass_addr_i[27:2] == el1[64:39];
  assign tag_hit2_n = bypass_addr_i[27:2] == sbuf_entry_i[64:39];

  bsg_mux_segmented_segments_p4_segment_width_p8
  mux_segmented_merge0
  (
    .data0_i(el1[36:5]),
    .data1_i(el0[36:5]),
    .sel_i({ n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_segments_p4_segment_width_p8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(sbuf_entry_i[36:5]),
    .sel_i({ n_4_net__3_, n_4_net__2_, n_4_net__1_, n_4_net__0_ }),
    .data_o(bypass_data_n)
  );

  assign { N20, N19 } = num_els_r + v_i;
  assign { N23, N22 } = { N20, N19 } - N21;
  assign v_o = (N0)? v_i : 
               (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N8;
  assign N1 = N10;
  assign N2 = N12;
  assign N3 = N13;
  assign empty_o = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 1'b0;
  assign el0_valid = (N0)? 1'b0 : 
                     (N1)? 1'b0 : 
                     (N2)? 1'b1 : 
                     (N3)? 1'b0 : 1'b0;
  assign el1_valid = (N0)? 1'b0 : 
                     (N1)? 1'b1 : 
                     (N2)? 1'b1 : 
                     (N3)? 1'b0 : 1'b0;
  assign el0_enable = (N0)? 1'b0 : 
                      (N1)? N15 : 
                      (N2)? N17 : 
                      (N3)? 1'b0 : 1'b0;
  assign el1_enable = (N0)? N14 : 
                      (N1)? N16 : 
                      (N2)? yumi_i : 
                      (N3)? 1'b0 : 1'b0;
  assign mux0_sel = (N0)? 1'b0 : 
                    (N1)? 1'b0 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign mux1_sel = (N0)? 1'b0 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign { N25, N24 } = (N4)? { 1'b0, 1'b0 } : 
                        (N5)? { N23, N22 } : 1'b0;
  assign N4 = reset_i;
  assign N5 = N18;
  assign N28 = (N4)? 1'b1 : 
               (N66)? 1'b1 : 
               (N27)? 1'b0 : 1'b0;
  assign { N32, N31, N30, N29 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N66)? bypass_mask_n : 1'b0;
  assign { N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                              (N66)? bypass_data_n : 1'b0;
  assign N6 = ~num_els_r[1];
  assign N7 = ~num_els_r[0];
  assign N10 = ~N9;
  assign N12 = ~N11;
  assign N14 = v_i & N67;
  assign N67 = ~yumi_i;
  assign N15 = v_i & N67;
  assign N16 = v_i & yumi_i;
  assign N17 = v_i & yumi_i;
  assign N18 = ~reset_i;
  assign N21 = v_o & yumi_i;
  assign tag_hit0x4[3] = tag_hit0_n & el0_valid;
  assign tag_hit1x4[3] = tag_hit1_n & el1_valid;
  assign tag_hit2x4[3] = tag_hit2_n & v_i;
  assign bypass_mask_n[3] = N70 | N71;
  assign N70 = N68 | N69;
  assign N68 = tag_hit0x4[3] & el0[4];
  assign N69 = tag_hit1x4[3] & el1[4];
  assign N71 = tag_hit2x4[3] & sbuf_entry_i[4];
  assign bypass_mask_n[2] = N74 | N75;
  assign N74 = N72 | N73;
  assign N72 = tag_hit0x4[3] & el0[3];
  assign N73 = tag_hit1x4[3] & el1[3];
  assign N75 = tag_hit2x4[3] & sbuf_entry_i[3];
  assign bypass_mask_n[1] = N78 | N79;
  assign N78 = N76 | N77;
  assign N76 = tag_hit0x4[3] & el0[2];
  assign N77 = tag_hit1x4[3] & el1[2];
  assign N79 = tag_hit2x4[3] & sbuf_entry_i[2];
  assign bypass_mask_n[0] = N82 | N83;
  assign N82 = N80 | N81;
  assign N80 = tag_hit0x4[3] & el0[1];
  assign N81 = tag_hit1x4[3] & el1[1];
  assign N83 = tag_hit2x4[3] & sbuf_entry_i[1];
  assign n_2_net__3_ = tag_hit0x4[3] & el0[4];
  assign n_2_net__2_ = tag_hit0x4[3] & el0[3];
  assign n_2_net__1_ = tag_hit0x4[3] & el0[2];
  assign n_2_net__0_ = tag_hit0x4[3] & el0[1];
  assign n_4_net__3_ = tag_hit2x4[3] & sbuf_entry_i[4];
  assign n_4_net__2_ = tag_hit2x4[3] & sbuf_entry_i[3];
  assign n_4_net__1_ = tag_hit2x4[3] & sbuf_entry_i[2];
  assign n_4_net__0_ = tag_hit2x4[3] & sbuf_entry_i[1];
  assign N26 = bypass_v_i | reset_i;
  assign N27 = ~N26;
  assign N65 = ~reset_i;
  assign N66 = bypass_v_i & N65;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { num_els_r[1:0] } <= { N25, N24 };
    end 
    if(N28) begin
      { bypass_data_o[31:0] } <= { N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33 };
      { bypass_mask_o[3:0] } <= { N32, N31, N30, N29 };
    end 
  end


endmodule



module bsg_mux_width_p32_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [95:0] data_i;
  input [1:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[31] = (N2)? data_i[31] : 
                      (N3)? data_i[63] : 
                      (N4)? data_i[95] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[30] = (N2)? data_i[30] : 
                      (N3)? data_i[62] : 
                      (N4)? data_i[94] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N3)? data_i[61] : 
                      (N4)? data_i[93] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N3)? data_i[60] : 
                      (N4)? data_i[92] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N3)? data_i[59] : 
                      (N4)? data_i[91] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N3)? data_i[58] : 
                      (N4)? data_i[90] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N3)? data_i[57] : 
                      (N4)? data_i[89] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N3)? data_i[56] : 
                      (N4)? data_i[88] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N3)? data_i[55] : 
                      (N4)? data_i[87] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N3)? data_i[54] : 
                      (N4)? data_i[86] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N3)? data_i[53] : 
                      (N4)? data_i[85] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N3)? data_i[52] : 
                      (N4)? data_i[84] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N3)? data_i[51] : 
                      (N4)? data_i[83] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N3)? data_i[50] : 
                      (N4)? data_i[82] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N3)? data_i[49] : 
                      (N4)? data_i[81] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N3)? data_i[48] : 
                      (N4)? data_i[80] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N3)? data_i[47] : 
                      (N4)? data_i[79] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N3)? data_i[46] : 
                      (N4)? data_i[78] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N3)? data_i[45] : 
                      (N4)? data_i[77] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N3)? data_i[44] : 
                      (N4)? data_i[76] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N3)? data_i[43] : 
                      (N4)? data_i[75] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N3)? data_i[42] : 
                      (N4)? data_i[74] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N3)? data_i[41] : 
                     (N4)? data_i[73] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N3)? data_i[40] : 
                     (N4)? data_i[72] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N3)? data_i[39] : 
                     (N4)? data_i[71] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N3)? data_i[38] : 
                     (N4)? data_i[70] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N3)? data_i[37] : 
                     (N4)? data_i[69] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N3)? data_i[36] : 
                     (N4)? data_i[68] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[35] : 
                     (N4)? data_i[67] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[34] : 
                     (N4)? data_i[66] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[33] : 
                     (N4)? data_i[65] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[32] : 
                     (N4)? data_i[64] : 1'b0;

endmodule



module bsg_mux_width_p4_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [11:0] data_i;
  input [1:0] sel_i;
  output [3:0] data_o;
  wire [3:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[7] : 
                     (N4)? data_i[11] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[6] : 
                     (N4)? data_i[10] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[5] : 
                     (N4)? data_i[9] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[4] : 
                     (N4)? data_i[8] : 1'b0;

endmodule



module bsg_decode_num_out_p4
(
  i,
  o
);

  input [1:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_mux_width_p8_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [1:0] sel_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[15] : 
                     (N3)? data_i[23] : 
                     (N5)? data_i[31] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[14] : 
                     (N3)? data_i[22] : 
                     (N5)? data_i[30] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[13] : 
                     (N3)? data_i[21] : 
                     (N5)? data_i[29] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[12] : 
                     (N3)? data_i[20] : 
                     (N5)? data_i[28] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[11] : 
                     (N3)? data_i[19] : 
                     (N5)? data_i[27] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[10] : 
                     (N3)? data_i[18] : 
                     (N5)? data_i[26] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[9] : 
                     (N3)? data_i[17] : 
                     (N5)? data_i[25] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[8] : 
                     (N3)? data_i[16] : 
                     (N5)? data_i[24] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p16_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [0:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[31] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[30] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[29] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[28] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[27] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[26] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[25] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[24] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[23] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[22] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[21] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[20] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[19] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[18] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[17] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[16] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_cache
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [68:0] cache_pkt_i;
  output [31:0] data_o;
  output [28:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output ready_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output v_we_o;
  wire [31:0] data_o,dma_data_o,snoop_word_lo,bypass_data_lo,sbuf_data_in,ld_data_way_picked,
  bypass_data_masked,snoop_or_ld_data,expanded_mask_v,ld_data_masked,
  ld_data_final_lo;
  wire [28:0] dma_pkt_o;
  wire ready_o,v_o,dma_pkt_v_o,dma_data_ready_o,dma_data_v_o,v_we_o,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,
  N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,
  N121,N122,tag_mem_v_li,tag_mem_w_li,data_mem_v_li,data_mem_w_li,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  tag_hit_found,ld_st_miss,N255,N256,tagfl_hit,aflinv_hit,N257,N258,N259,N260,
  N261,N262,alock_miss,N263,N264,N265,N266,N267,aunlock_hit,miss_v,retval_op_v,
  stat_mem_v_li,stat_mem_w_li,sbuf_empty_li,dma_done_li,miss_stat_mem_v_lo,
  miss_stat_mem_w_lo,miss_tag_mem_v_lo,miss_tag_mem_w_lo,recover_lo,miss_done_lo,n_0_net_,
  dma_data_mem_v_lo,dma_data_mem_w_lo,dma_evict_lo,sbuf_entry_li_data__31_,
  sbuf_entry_li_data__30_,sbuf_entry_li_data__29_,sbuf_entry_li_data__28_,
  sbuf_entry_li_data__27_,sbuf_entry_li_data__26_,sbuf_entry_li_data__25_,sbuf_entry_li_data__24_,
  sbuf_entry_li_data__23_,sbuf_entry_li_data__22_,sbuf_entry_li_data__21_,
  sbuf_entry_li_data__20_,sbuf_entry_li_data__19_,sbuf_entry_li_data__18_,
  sbuf_entry_li_data__17_,sbuf_entry_li_data__16_,sbuf_entry_li_data__15_,sbuf_entry_li_data__14_,
  sbuf_entry_li_data__13_,sbuf_entry_li_data__12_,sbuf_entry_li_data__11_,
  sbuf_entry_li_data__10_,sbuf_entry_li_data__9_,sbuf_entry_li_data__8_,sbuf_entry_li_data__7_,
  sbuf_entry_li_data__6_,sbuf_entry_li_data__5_,sbuf_entry_li_data__4_,
  sbuf_entry_li_data__3_,sbuf_entry_li_data__2_,sbuf_entry_li_data__1_,
  sbuf_entry_li_data__0_,sbuf_entry_li_mask__3_,sbuf_entry_li_mask__2_,sbuf_entry_li_mask__1_,
  sbuf_entry_li_mask__0_,sbuf_entry_li_way_id__0_,sbuf_v_li,sbuf_v_lo,sbuf_yumi_li,
  bypass_v_li,sbuf_mask_in_mux_li_1__3_,sbuf_mask_in_mux_li_1__2_,
  sbuf_mask_in_mux_li_1__1_,sbuf_mask_in_mux_li_1__0_,sbuf_mask_in_mux_li_0__3_,sbuf_mask_in_mux_li_0__2_,
  sbuf_mask_in_mux_li_0__1_,sbuf_mask_in_mux_li_0__0_,N268,N269,N270,N271,N272,
  N273,ld_data_final_li_1__31_,ld_data_final_li_1__30_,ld_data_final_li_1__29_,
  ld_data_final_li_1__28_,ld_data_final_li_1__27_,ld_data_final_li_1__26_,
  ld_data_final_li_1__25_,ld_data_final_li_1__24_,ld_data_final_li_1__23_,
  ld_data_final_li_1__22_,ld_data_final_li_1__21_,ld_data_final_li_1__20_,ld_data_final_li_1__19_,
  ld_data_final_li_1__18_,ld_data_final_li_1__17_,ld_data_final_li_1__16_,
  ld_data_final_li_0__31_,ld_data_final_li_0__30_,ld_data_final_li_0__29_,
  ld_data_final_li_0__28_,ld_data_final_li_0__27_,ld_data_final_li_0__26_,ld_data_final_li_0__25_,
  ld_data_final_li_0__24_,ld_data_final_li_0__23_,ld_data_final_li_0__22_,
  ld_data_final_li_0__21_,ld_data_final_li_0__20_,ld_data_final_li_0__19_,
  ld_data_final_li_0__18_,ld_data_final_li_0__17_,ld_data_final_li_0__16_,ld_data_final_li_0__15_,
  ld_data_final_li_0__14_,ld_data_final_li_0__13_,ld_data_final_li_0__12_,
  ld_data_final_li_0__11_,ld_data_final_li_0__10_,ld_data_final_li_0__9_,ld_data_final_li_0__8_,
  N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
  N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,
  N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,
  N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,
  N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,tl_ready,N349,N350,
  tagst_write_en,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,
  N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,
  N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,
  N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,
  N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,
  N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439;
  wire [15:0] decode,ld_data_sel_1__non_max_size_byte_sel;
  wire [5:0] tag_mem_addr_li,stat_mem_addr_li,miss_stat_mem_addr_lo,miss_tag_mem_addr_lo;
  wire [39:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo,miss_tag_mem_data_lo,
  miss_tag_mem_w_mask_lo;
  wire [7:0] data_mem_addr_li,data_mem_w_mask_li,dma_data_mem_addr_lo,dma_data_mem_w_mask_lo,
  sbuf_data_mem_w_mask,ld_data_sel_0__non_max_size_byte_sel;
  wire [63:0] data_mem_data_li,data_mem_data_lo,dma_data_mem_data_lo;
  wire [1:0] tag_hit_v,sbuf_way_decode,sbuf_in_sel_1__non_max_size_decode_lo,addr_way_decode;
  wire [0:0] tag_hit_way_id,dma_way_lo,chosen_way_lo,plru_decode_data_lo,plru_decode_mask_lo;
  wire [2:0] stat_mem_data_li,stat_mem_w_mask_li,stat_mem_data_lo,miss_stat_mem_data_lo,
  miss_stat_mem_w_mask_lo;
  wire [3:0] dma_cmd_lo,bypass_mask_lo,sbuf_mask_in,sbuf_in_sel_0__non_max_size_decode_lo;
  wire [27:0] dma_addr_lo;
  wire [64:0] sbuf_entry_lo;
  reg [31:0] data_tl_r,data_v_r;
  reg v_tl_r,v_v_r;
  reg [15:0] decode_tl_r,decode_v_r;
  reg [3:0] mask_tl_r,mask_v_r;
  reg [27:0] addr_tl_r,addr_v_r;
  reg [63:0] ld_data_v_r;
  reg [35:0] tag_v_r;
  reg [1:0] valid_v_r,lock_v_r;

  bsg_cache_pkt_decode_data_width_p32_addr_width_p28
  cache_pkt_decoder
  (
    .cache_pkt_i(cache_pkt_i),
    .decode_o(decode)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p40_els_p64_latch_last_read_p1
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(tag_mem_v_li),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p256_data_width_p64_latch_last_read_p1
  data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li),
    .data_i(data_mem_data_li),
    .write_mask_i(data_mem_w_mask_li),
    .data_o(data_mem_data_lo)
  );

  assign N253 = addr_v_r[27:10] == tag_v_r[17:0];
  assign N254 = addr_v_r[27:10] == tag_v_r[35:18];

  bsg_priority_encode_width_p2_lo_to_hi_p1
  tag_hit_pe
  (
    .i(tag_hit_v),
    .addr_o(tag_hit_way_id[0]),
    .v_o(tag_hit_found)
  );

  assign N256 = (N255)? valid_v_r[0] : 
                (N0)? valid_v_r[1] : 1'b0;
  assign N0 = addr_v_r[10];
  assign N260 = (N259)? lock_v_r[0] : 
                (N1)? lock_v_r[1] : 1'b0;
  assign N1 = tag_hit_way_id[0];
  assign N266 = (N265)? lock_v_r[0] : 
                (N1)? lock_v_r[1] : 1'b0;

  bsg_mem_1rw_sync_mask_write_bit_width_p3_els_p64_latch_last_read_p1
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(stat_mem_v_li),
    .w_mask_i(stat_mem_w_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_data_lo)
  );


  bsg_cache_miss_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p2
  miss
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .miss_v_i(miss_v),
    .decode_v_i(decode_v_r),
    .addr_v_i(addr_v_r),
    .tag_v_i(tag_v_r),
    .valid_v_i(valid_v_r),
    .lock_v_i(lock_v_r),
    .tag_hit_way_id_i(tag_hit_way_id[0]),
    .tag_hit_found_i(tag_hit_found),
    .sbuf_empty_i(sbuf_empty_li),
    .dma_cmd_o(dma_cmd_lo),
    .dma_way_o(dma_way_lo[0]),
    .dma_addr_o(dma_addr_lo),
    .dma_done_i(dma_done_li),
    .stat_info_i(stat_mem_data_lo),
    .stat_mem_v_o(miss_stat_mem_v_lo),
    .stat_mem_w_o(miss_stat_mem_w_lo),
    .stat_mem_addr_o(miss_stat_mem_addr_lo),
    .stat_mem_data_o(miss_stat_mem_data_lo),
    .stat_mem_w_mask_o(miss_stat_mem_w_mask_lo),
    .tag_mem_v_o(miss_tag_mem_v_lo),
    .tag_mem_w_o(miss_tag_mem_w_lo),
    .tag_mem_addr_o(miss_tag_mem_addr_lo),
    .tag_mem_data_o(miss_tag_mem_data_lo),
    .tag_mem_w_mask_o(miss_tag_mem_w_mask_lo),
    .done_o(miss_done_lo),
    .recover_o(recover_lo),
    .chosen_way_o(chosen_way_lo[0]),
    .ack_i(n_0_net_)
  );


  bsg_cache_dma_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p2_debug_p0
  dma
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .dma_cmd_i(dma_cmd_lo),
    .dma_way_i(dma_way_lo[0]),
    .dma_addr_i(dma_addr_lo),
    .done_o(dma_done_li),
    .snoop_word_o(snoop_word_lo),
    .dma_pkt_o(dma_pkt_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_i(dma_data_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_ready_o(dma_data_ready_o),
    .dma_data_o(dma_data_o),
    .dma_data_v_o(dma_data_v_o),
    .dma_data_yumi_i(dma_data_yumi_i),
    .data_mem_v_o(dma_data_mem_v_lo),
    .data_mem_w_o(dma_data_mem_w_lo),
    .data_mem_addr_o(dma_data_mem_addr_lo),
    .data_mem_w_mask_o(dma_data_mem_w_mask_lo),
    .data_mem_data_o(dma_data_mem_data_lo),
    .data_mem_data_i(data_mem_data_lo),
    .dma_evict_o(dma_evict_lo)
  );


  bsg_cache_sbuf_data_width_p32_addr_width_p28_ways_p2
  sbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .sbuf_entry_i({ addr_v_r, sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_, sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_, sbuf_entry_li_way_id__0_ }),
    .v_i(sbuf_v_li),
    .sbuf_entry_o(sbuf_entry_lo),
    .v_o(sbuf_v_lo),
    .yumi_i(sbuf_yumi_li),
    .empty_o(sbuf_empty_li),
    .bypass_addr_i(addr_tl_r),
    .bypass_v_i(bypass_v_li),
    .bypass_data_o(bypass_data_lo),
    .bypass_mask_o(bypass_mask_lo)
  );


  bsg_decode_num_out_p2
  sbuf_way_demux
  (
    .i(sbuf_entry_lo[0]),
    .o(sbuf_way_decode)
  );


  bsg_mux_width_p32_els_p3
  sbuf_data_in_mux
  (
    .data_i({ data_v_r, data_v_r[15:0], data_v_r[15:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0] }),
    .sel_i(decode_v_r[15:14]),
    .data_o(sbuf_data_in)
  );


  bsg_mux_width_p4_els_p3
  sbuf_mask_in_mux
  (
    .data_i({ 1'b1, 1'b1, 1'b1, 1'b1, sbuf_mask_in_mux_li_1__3_, sbuf_mask_in_mux_li_1__2_, sbuf_mask_in_mux_li_1__1_, sbuf_mask_in_mux_li_1__0_, sbuf_mask_in_mux_li_0__3_, sbuf_mask_in_mux_li_0__2_, sbuf_mask_in_mux_li_0__1_, sbuf_mask_in_mux_li_0__0_ }),
    .sel_i(decode_v_r[15:14]),
    .data_o(sbuf_mask_in)
  );


  bsg_decode_num_out_p4
  sbuf_in_sel_0__non_max_size_dec
  (
    .i(addr_v_r[1:0]),
    .o(sbuf_in_sel_0__non_max_size_decode_lo)
  );


  bsg_expand_bitmask
  sbuf_in_sel_0__non_max_size_exp
  (
    .i(sbuf_in_sel_0__non_max_size_decode_lo),
    .o({ sbuf_mask_in_mux_li_0__3_, sbuf_mask_in_mux_li_0__2_, sbuf_mask_in_mux_li_0__1_, sbuf_mask_in_mux_li_0__0_ })
  );


  bsg_decode_num_out_p2
  sbuf_in_sel_1__non_max_size_dec
  (
    .i(addr_v_r[1]),
    .o(sbuf_in_sel_1__non_max_size_decode_lo)
  );


  bsg_expand_bitmask
  sbuf_in_sel_1__non_max_size_exp
  (
    .i(sbuf_in_sel_1__non_max_size_decode_lo),
    .o({ sbuf_mask_in_mux_li_1__3_, sbuf_mask_in_mux_li_1__2_, sbuf_mask_in_mux_li_1__1_, sbuf_mask_in_mux_li_1__0_ })
  );


  bsg_mux_width_p32_els_p2
  ld_data_mux
  (
    .data_i(ld_data_v_r),
    .sel_i(tag_hit_way_id[0]),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_segmented_segments_p4_segment_width_p8
  bypass_mux_segmented
  (
    .data0_i(ld_data_way_picked),
    .data1_i(bypass_data_lo),
    .sel_i(bypass_mask_lo),
    .data_o(bypass_data_masked)
  );


  bsg_expand_bitmask
  mask_v_expand
  (
    .i(mask_v_r),
    .o(expanded_mask_v)
  );


  bsg_mux_width_p8_els_p4
  ld_data_sel_0__non_max_size_byte_mux
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[1:0]),
    .data_o(ld_data_sel_0__non_max_size_byte_sel)
  );


  bsg_mux_width_p16_els_p2
  ld_data_sel_1__non_max_size_byte_mux
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[1]),
    .data_o(ld_data_sel_1__non_max_size_byte_sel)
  );


  bsg_mux_width_p32_els_p3
  ld_data_size_mux
  (
    .data_i({ snoop_or_ld_data, ld_data_final_li_1__31_, ld_data_final_li_1__30_, ld_data_final_li_1__29_, ld_data_final_li_1__28_, ld_data_final_li_1__27_, ld_data_final_li_1__26_, ld_data_final_li_1__25_, ld_data_final_li_1__24_, ld_data_final_li_1__23_, ld_data_final_li_1__22_, ld_data_final_li_1__21_, ld_data_final_li_1__20_, ld_data_final_li_1__19_, ld_data_final_li_1__18_, ld_data_final_li_1__17_, ld_data_final_li_1__16_, ld_data_sel_1__non_max_size_byte_sel, ld_data_final_li_0__31_, ld_data_final_li_0__30_, ld_data_final_li_0__29_, ld_data_final_li_0__28_, ld_data_final_li_0__27_, ld_data_final_li_0__26_, ld_data_final_li_0__25_, ld_data_final_li_0__24_, ld_data_final_li_0__23_, ld_data_final_li_0__22_, ld_data_final_li_0__21_, ld_data_final_li_0__20_, ld_data_final_li_0__19_, ld_data_final_li_0__18_, ld_data_final_li_0__17_, ld_data_final_li_0__16_, ld_data_final_li_0__15_, ld_data_final_li_0__14_, ld_data_final_li_0__13_, ld_data_final_li_0__12_, ld_data_final_li_0__11_, ld_data_final_li_0__10_, ld_data_final_li_0__9_, ld_data_final_li_0__8_, ld_data_sel_0__non_max_size_byte_sel }),
    .sel_i(decode_v_r[15:14]),
    .data_o(ld_data_final_lo)
  );

  assign N282 = (N281)? lock_v_r[0] : 
                (N0)? lock_v_r[1] : 1'b0;
  assign N284 = (N283)? valid_v_r[0] : 
                (N0)? valid_v_r[1] : 1'b0;
  assign N286 = (N285)? tag_v_r[17] : 
                (N0)? tag_v_r[35] : 1'b0;
  assign N287 = (N285)? tag_v_r[16] : 
                (N0)? tag_v_r[34] : 1'b0;
  assign N288 = (N285)? tag_v_r[15] : 
                (N0)? tag_v_r[33] : 1'b0;
  assign N289 = (N285)? tag_v_r[14] : 
                (N0)? tag_v_r[32] : 1'b0;
  assign N290 = (N285)? tag_v_r[13] : 
                (N0)? tag_v_r[31] : 1'b0;
  assign N291 = (N285)? tag_v_r[12] : 
                (N0)? tag_v_r[30] : 1'b0;
  assign N292 = (N285)? tag_v_r[11] : 
                (N0)? tag_v_r[29] : 1'b0;
  assign N293 = (N285)? tag_v_r[10] : 
                (N0)? tag_v_r[28] : 1'b0;
  assign N294 = (N285)? tag_v_r[9] : 
                (N0)? tag_v_r[27] : 1'b0;
  assign N295 = (N285)? tag_v_r[8] : 
                (N0)? tag_v_r[26] : 1'b0;
  assign N296 = (N285)? tag_v_r[7] : 
                (N0)? tag_v_r[25] : 1'b0;
  assign N297 = (N285)? tag_v_r[6] : 
                (N0)? tag_v_r[24] : 1'b0;
  assign N298 = (N285)? tag_v_r[5] : 
                (N0)? tag_v_r[23] : 1'b0;
  assign N299 = (N285)? tag_v_r[4] : 
                (N0)? tag_v_r[22] : 1'b0;
  assign N300 = (N285)? tag_v_r[3] : 
                (N0)? tag_v_r[21] : 1'b0;
  assign N301 = (N285)? tag_v_r[2] : 
                (N0)? tag_v_r[20] : 1'b0;
  assign N302 = (N285)? tag_v_r[1] : 
                (N0)? tag_v_r[19] : 1'b0;
  assign N303 = (N285)? tag_v_r[0] : 
                (N0)? tag_v_r[18] : 1'b0;

  bsg_decode_num_out_p2
  addr_way_demux
  (
    .i(cache_pkt_i[46]),
    .o(addr_way_decode)
  );


  bsg_lru_pseudo_tree_decode_ways_p2
  plru_decode
  (
    .way_id_i(tag_hit_way_id[0]),
    .data_o(plru_decode_data_lo[0]),
    .mask_o(plru_decode_mask_lo[0])
  );

  assign N38 = (N2)? 1'b1 : 
               (N122)? 1'b1 : 
               (N37)? 1'b0 : 1'b0;
  assign N2 = N35;
  assign N39 = (N2)? 1'b0 : 
               (N122)? v_i : 1'b0;
  assign N40 = (N2)? 1'b1 : 
               (N122)? v_i : 
               (N37)? 1'b0 : 1'b0;
  assign { N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                              (N122)? decode : 1'b0;
  assign { N60, N59, N58, N57 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N122)? cache_pkt_i[3:0] : 1'b0;
  assign { N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                          (N122)? cache_pkt_i[63:36] : 1'b0;
  assign { N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                   (N122)? cache_pkt_i[35:4] : 1'b0;
  assign N126 = (N3)? 1'b1 : 
                (N252)? 1'b1 : 
                (N125)? 1'b0 : 1'b0;
  assign N3 = N123;
  assign N127 = (N3)? 1'b0 : 
                (N252)? v_tl_r : 1'b0;
  assign { N132, N128 } = (N3)? { 1'b1, 1'b1 } : 
                          (N252)? { v_tl_r, v_tl_r } : 
                          (N125)? { 1'b0, 1'b0 } : 1'b0;
  assign { N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N131, N130, N129 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                      (N252)? { tag_mem_data_lo[37:20], tag_mem_data_lo[17:0] } : 1'b0;
  assign { N169, N168, N167, N166 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N252)? mask_tl_r : 1'b0;
  assign { N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                              (N252)? decode_tl_r : 1'b0;
  assign { N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                      (N252)? addr_tl_r : 1'b0;
  assign { N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N252)? data_tl_r : 1'b0;
  assign { N247, N246 } = (N3)? { 1'b0, 1'b0 } : 
                          (N252)? { tag_mem_data_lo[39:39], tag_mem_data_lo[19:19] } : 1'b0;
  assign { N249, N248 } = (N3)? { 1'b0, 1'b0 } : 
                          (N252)? { tag_mem_data_lo[38:38], tag_mem_data_lo[18:18] } : 1'b0;
  assign N250 = (N3)? 1'b0 : 
                (N252)? v_tl_r : 
                (N125)? 1'b0 : 1'b0;
  assign N262 = (N4)? N261 : 
                (N5)? 1'b1 : 1'b0;
  assign N4 = N258;
  assign N5 = N257;
  assign N267 = (N6)? N266 : 
                (N7)? 1'b0 : 1'b0;
  assign N6 = N264;
  assign N7 = N263;
  assign { sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_ } = (N8)? data_v_r : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N269)? sbuf_data_in : 1'b0;
  assign N8 = N268;
  assign { sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_ } = (N9)? mask_v_r : 
                                                                                                              (N271)? sbuf_mask_in : 1'b0;
  assign N9 = N270;
  assign snoop_or_ld_data = (N10)? snoop_word_lo : 
                            (N11)? bypass_data_masked : 1'b0;
  assign N10 = N273;
  assign N11 = N272;
  assign { N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304 } = (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N282, N284 } : 
                                                                                                                                                                                                              (N337)? { 1'b0, 1'b0, 1'b0, 1'b0, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, addr_v_r[9:4], 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N340)? ld_data_masked : 
                                                                                                                                                                                                              (N280)? ld_data_final_lo : 1'b0;
  assign N12 = N275;
  assign data_o = (N13)? { N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304 } : 
                  (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = retval_op_v;
  assign N14 = N274;
  assign N343 = (N15)? miss_done_lo : 
                (N16)? 1'b1 : 1'b0;
  assign N15 = N342;
  assign N16 = N341;
  assign v_we_o = (N17)? N345 : 
                  (N18)? 1'b1 : 1'b0;
  assign N17 = v_v_r;
  assign N18 = N344;
  assign tl_ready = (N19)? N348 : 
                    (N20)? 1'b1 : 1'b0;
  assign N19 = N347;
  assign N20 = N346;
  assign ready_o = (N21)? N350 : 
                   (N22)? tl_ready : 1'b0;
  assign N21 = v_tl_r;
  assign N22 = N349;
  assign tag_mem_w_li = (N23)? miss_tag_mem_w_lo : 
                        (N24)? tagst_write_en : 1'b0;
  assign N23 = N352;
  assign N24 = N351;
  assign { N362, N361, N360, N359, N358, N357 } = (N25)? addr_tl_r[9:4] : 
                                                  (N364)? miss_tag_mem_addr_lo : 
                                                  (N356)? cache_pkt_i[45:40] : 1'b0;
  assign N25 = recover_lo;
  assign tag_mem_addr_li = (N26)? { N362, N361, N360, N359, N358, N357 } : 
                           (N27)? cache_pkt_i[45:40] : 1'b0;
  assign N26 = N354;
  assign N27 = N353;
  assign tag_mem_data_li = (N26)? miss_tag_mem_data_lo : 
                           (N27)? { cache_pkt_i[35:34], cache_pkt_i[21:4], cache_pkt_i[35:34], cache_pkt_i[21:4] } : 1'b0;
  assign tag_mem_w_mask_li = (N26)? miss_tag_mem_w_mask_lo : 
                             (N27)? { addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode, addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0] } : 1'b0;
  assign data_mem_data_li = (N28)? dma_data_mem_data_lo : 
                            (N29)? { sbuf_entry_lo[36:5], sbuf_entry_lo[36:5] } : 1'b0;
  assign N28 = dma_data_mem_w_lo;
  assign N29 = N365;
  assign data_mem_addr_li = (N25)? addr_tl_r[9:2] : 
                            (N370)? dma_data_mem_addr_lo : 
                            (N373)? cache_pkt_i[45:38] : 
                            (N369)? sbuf_entry_lo[46:39] : 1'b0;
  assign data_mem_w_mask_li = (N28)? dma_data_mem_w_mask_lo : 
                              (N29)? sbuf_data_mem_w_mask : 1'b0;
  assign { N384, N383, N382 } = (N30)? { 1'b0, 1'b0, 1'b0 } : 
                                (N379)? { decode_v_r[10:10], decode_v_r[10:10], plru_decode_data_lo[0:0] } : 1'b0;
  assign N30 = N378;
  assign { N387, N386, N385 } = (N30)? { 1'b1, 1'b1, 1'b1 } : 
                                (N379)? { N380, N381, plru_decode_mask_lo[0:0] } : 1'b0;
  assign stat_mem_v_li = (N31)? miss_stat_mem_v_lo : 
                         (N32)? N376 : 1'b0;
  assign N31 = N375;
  assign N32 = N374;
  assign stat_mem_w_li = (N31)? miss_stat_mem_w_lo : 
                         (N32)? N377 : 1'b0;
  assign stat_mem_addr_li = (N31)? miss_stat_mem_addr_lo : 
                            (N32)? addr_v_r[9:4] : 1'b0;
  assign stat_mem_data_li = (N31)? miss_stat_mem_data_lo : 
                            (N32)? { N384, N383, N382 } : 1'b0;
  assign stat_mem_w_mask_li = (N31)? miss_stat_mem_w_mask_lo : 
                              (N32)? { N387, N386, N385 } : 1'b0;
  assign sbuf_entry_li_way_id__0_ = (N33)? chosen_way_lo[0] : 
                                    (N34)? tag_hit_way_id[0] : 1'b0;
  assign N33 = N389;
  assign N34 = N388;
  assign N35 = reset_i;
  assign N36 = ready_o | N35;
  assign N37 = ~N36;
  assign N121 = ~N35;
  assign N122 = ready_o & N121;
  assign N123 = reset_i;
  assign N124 = v_we_o | N123;
  assign N125 = ~N124;
  assign N251 = ~N123;
  assign N252 = v_we_o & N251;
  assign tag_hit_v[0] = N253 & valid_v_r[0];
  assign tag_hit_v[1] = N254 & valid_v_r[1];
  assign ld_st_miss = N390 & N391;
  assign N390 = ~tag_hit_found;
  assign N391 = decode_v_r[11] | decode_v_r[10];
  assign N255 = ~addr_v_r[10];
  assign tagfl_hit = decode_v_r[8] & N256;
  assign aflinv_hit = N393 & tag_hit_found;
  assign N393 = N392 | decode_v_r[3];
  assign N392 = decode_v_r[5] | decode_v_r[4];
  assign N257 = ~tag_hit_found;
  assign N258 = tag_hit_found;
  assign N259 = ~tag_hit_way_id[0];
  assign N261 = ~N260;
  assign alock_miss = decode_v_r[2] & N262;
  assign N263 = ~tag_hit_found;
  assign N264 = tag_hit_found;
  assign N265 = ~tag_hit_way_id[0];
  assign aunlock_hit = decode_v_r[1] & N267;
  assign miss_v = N395 & N399;
  assign N395 = N394 & v_v_r;
  assign N394 = ~decode_v_r[9];
  assign N399 = N398 | aunlock_hit;
  assign N398 = N397 | alock_miss;
  assign N397 = N396 | aflinv_hit;
  assign N396 = ld_st_miss | tagfl_hit;
  assign retval_op_v = N400 | decode_v_r[6];
  assign N400 = decode_v_r[11] | decode_v_r[7];
  assign n_0_net_ = v_o & yumi_i;
  assign sbuf_data_mem_w_mask[3] = sbuf_way_decode[0] & sbuf_entry_lo[4];
  assign sbuf_data_mem_w_mask[2] = sbuf_way_decode[0] & sbuf_entry_lo[3];
  assign sbuf_data_mem_w_mask[1] = sbuf_way_decode[0] & sbuf_entry_lo[2];
  assign sbuf_data_mem_w_mask[0] = sbuf_way_decode[0] & sbuf_entry_lo[1];
  assign sbuf_data_mem_w_mask[7] = sbuf_way_decode[1] & sbuf_entry_lo[4];
  assign sbuf_data_mem_w_mask[6] = sbuf_way_decode[1] & sbuf_entry_lo[3];
  assign sbuf_data_mem_w_mask[5] = sbuf_way_decode[1] & sbuf_entry_lo[2];
  assign sbuf_data_mem_w_mask[4] = sbuf_way_decode[1] & sbuf_entry_lo[1];
  assign N268 = decode_v_r[12];
  assign N269 = ~N268;
  assign N270 = decode_v_r[12];
  assign N271 = ~N270;
  assign N272 = ~miss_v;
  assign N273 = miss_v;
  assign ld_data_masked[31] = snoop_or_ld_data[31] & expanded_mask_v[31];
  assign ld_data_masked[30] = snoop_or_ld_data[30] & expanded_mask_v[30];
  assign ld_data_masked[29] = snoop_or_ld_data[29] & expanded_mask_v[29];
  assign ld_data_masked[28] = snoop_or_ld_data[28] & expanded_mask_v[28];
  assign ld_data_masked[27] = snoop_or_ld_data[27] & expanded_mask_v[27];
  assign ld_data_masked[26] = snoop_or_ld_data[26] & expanded_mask_v[26];
  assign ld_data_masked[25] = snoop_or_ld_data[25] & expanded_mask_v[25];
  assign ld_data_masked[24] = snoop_or_ld_data[24] & expanded_mask_v[24];
  assign ld_data_masked[23] = snoop_or_ld_data[23] & expanded_mask_v[23];
  assign ld_data_masked[22] = snoop_or_ld_data[22] & expanded_mask_v[22];
  assign ld_data_masked[21] = snoop_or_ld_data[21] & expanded_mask_v[21];
  assign ld_data_masked[20] = snoop_or_ld_data[20] & expanded_mask_v[20];
  assign ld_data_masked[19] = snoop_or_ld_data[19] & expanded_mask_v[19];
  assign ld_data_masked[18] = snoop_or_ld_data[18] & expanded_mask_v[18];
  assign ld_data_masked[17] = snoop_or_ld_data[17] & expanded_mask_v[17];
  assign ld_data_masked[16] = snoop_or_ld_data[16] & expanded_mask_v[16];
  assign ld_data_masked[15] = snoop_or_ld_data[15] & expanded_mask_v[15];
  assign ld_data_masked[14] = snoop_or_ld_data[14] & expanded_mask_v[14];
  assign ld_data_masked[13] = snoop_or_ld_data[13] & expanded_mask_v[13];
  assign ld_data_masked[12] = snoop_or_ld_data[12] & expanded_mask_v[12];
  assign ld_data_masked[11] = snoop_or_ld_data[11] & expanded_mask_v[11];
  assign ld_data_masked[10] = snoop_or_ld_data[10] & expanded_mask_v[10];
  assign ld_data_masked[9] = snoop_or_ld_data[9] & expanded_mask_v[9];
  assign ld_data_masked[8] = snoop_or_ld_data[8] & expanded_mask_v[8];
  assign ld_data_masked[7] = snoop_or_ld_data[7] & expanded_mask_v[7];
  assign ld_data_masked[6] = snoop_or_ld_data[6] & expanded_mask_v[6];
  assign ld_data_masked[5] = snoop_or_ld_data[5] & expanded_mask_v[5];
  assign ld_data_masked[4] = snoop_or_ld_data[4] & expanded_mask_v[4];
  assign ld_data_masked[3] = snoop_or_ld_data[3] & expanded_mask_v[3];
  assign ld_data_masked[2] = snoop_or_ld_data[2] & expanded_mask_v[2];
  assign ld_data_masked[1] = snoop_or_ld_data[1] & expanded_mask_v[1];
  assign ld_data_masked[0] = snoop_or_ld_data[0] & expanded_mask_v[0];
  assign ld_data_final_li_0__31_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__30_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__29_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__28_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__27_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__26_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__25_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__24_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__23_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__22_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__21_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__20_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__19_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__18_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__17_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__16_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__15_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__14_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__13_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__12_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__11_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__10_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__9_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_0__8_ = decode_v_r[13] & ld_data_sel_0__non_max_size_byte_sel[7];
  assign ld_data_final_li_1__31_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__30_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__29_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__28_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__27_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__26_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__25_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__24_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__23_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__22_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__21_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__20_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__19_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__18_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__17_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign ld_data_final_li_1__16_ = decode_v_r[13] & ld_data_sel_1__non_max_size_byte_sel[15];
  assign N274 = ~retval_op_v;
  assign N275 = decode_v_r[7];
  assign N276 = decode_v_r[6];
  assign N277 = decode_v_r[12];
  assign N278 = N276 | N275;
  assign N279 = N277 | N278;
  assign N280 = ~N279;
  assign N281 = ~addr_v_r[10];
  assign N283 = ~addr_v_r[10];
  assign N285 = ~addr_v_r[10];
  assign N336 = ~N275;
  assign N337 = N276 & N336;
  assign N338 = ~N276;
  assign N339 = N336 & N338;
  assign N340 = N277 & N339;
  assign N341 = ~miss_v;
  assign N342 = miss_v;
  assign v_o = v_v_r & N343;
  assign N344 = ~v_v_r;
  assign N345 = v_o & yumi_i;
  assign N346 = ~miss_v;
  assign N347 = miss_v;
  assign N348 = N408 & N409;
  assign N408 = N406 & N407;
  assign N406 = N404 & N405;
  assign N404 = N402 & N403;
  assign N402 = ~N401;
  assign N401 = decode[9] & v_i;
  assign N403 = ~miss_tag_mem_v_lo;
  assign N405 = ~dma_data_mem_v_lo;
  assign N407 = ~recover_lo;
  assign N409 = ~dma_evict_lo;
  assign N349 = ~v_tl_r;
  assign N350 = v_we_o & tl_ready;
  assign tagst_write_en = N410 & v_i;
  assign N410 = decode[9] & ready_o;
  assign tag_mem_v_li = N416 | N418;
  assign N416 = N415 | miss_tag_mem_v_lo;
  assign N415 = N412 | N414;
  assign N412 = N411 & v_i;
  assign N411 = decode[0] & ready_o;
  assign N414 = N413 & v_tl_r;
  assign N413 = recover_lo & decode_tl_r[0];
  assign N418 = N417 & v_i;
  assign N417 = decode[9] & ready_o;
  assign N351 = ~miss_v;
  assign N352 = miss_v;
  assign N353 = ~miss_v;
  assign N354 = miss_v;
  assign N355 = miss_tag_mem_v_lo | recover_lo;
  assign N356 = ~N355;
  assign N363 = ~recover_lo;
  assign N364 = miss_tag_mem_v_lo & N363;
  assign data_mem_v_li = N424 | N425;
  assign N424 = N423 | dma_data_mem_v_lo;
  assign N423 = N420 | N422;
  assign N420 = N419 & ready_o;
  assign N419 = v_i & decode[11];
  assign N422 = N421 & decode_tl_r[11];
  assign N421 = v_tl_r & recover_lo;
  assign N425 = sbuf_v_lo & sbuf_yumi_li;
  assign data_mem_w_li = dma_data_mem_w_lo | N426;
  assign N426 = sbuf_v_lo & sbuf_yumi_li;
  assign N365 = ~dma_data_mem_w_lo;
  assign N366 = N427 & ready_o;
  assign N427 = decode[11] & v_i;
  assign N367 = dma_data_mem_v_lo | recover_lo;
  assign N368 = N366 | N367;
  assign N369 = ~N368;
  assign N370 = dma_data_mem_v_lo & N363;
  assign N371 = ~dma_data_mem_v_lo;
  assign N372 = N363 & N371;
  assign N373 = N366 & N372;
  assign N374 = ~miss_v;
  assign N375 = miss_v;
  assign N376 = N430 & yumi_i;
  assign N430 = N429 & v_o;
  assign N429 = N428 | decode_v_r[9];
  assign N428 = decode_v_r[10] | decode_v_r[11];
  assign N377 = N433 & yumi_i;
  assign N433 = N432 & v_o;
  assign N432 = N431 | decode_v_r[9];
  assign N431 = decode_v_r[10] | decode_v_r[11];
  assign N378 = decode_v_r[9];
  assign N379 = ~N378;
  assign N380 = decode_v_r[10] & tag_hit_v[1];
  assign N381 = decode_v_r[10] & tag_hit_v[0];
  assign sbuf_v_li = N434 & yumi_i;
  assign N434 = decode_v_r[10] & v_o;
  assign N388 = ~miss_v;
  assign N389 = miss_v;
  assign sbuf_yumi_li = N438 & N405;
  assign N438 = sbuf_v_lo & N437;
  assign N437 = ~N436;
  assign N436 = N435 & ready_o;
  assign N435 = decode[11] & v_i;
  assign bypass_v_li = N439 & v_we_o;
  assign N439 = decode_tl_r[11] & v_tl_r;

  always @(posedge clk_i) begin
    if(N40) begin
      { data_tl_r[31:0] } <= { N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89 };
      { decode_tl_r[15:0] } <= { N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41 };
      { mask_tl_r[3:0] } <= { N60, N59, N58, N57 };
      { addr_tl_r[27:0] } <= { N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61 };
    end 
    if(N38) begin
      v_tl_r <= N39;
    end 
    if(N250) begin
      { ld_data_v_r[63:0] } <= { data_mem_data_lo[63:0] };
    end 
    if(N126) begin
      v_v_r <= N127;
    end 
    if(N132) begin
      { tag_v_r[35:3] } <= { N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133 };
      { mask_v_r[0:0] } <= { N166 };
      { lock_v_r[1:0] } <= { N249, N248 };
    end 
    if(N128) begin
      { tag_v_r[2:0] } <= { N131, N130, N129 };
      { mask_v_r[3:1] } <= { N169, N168, N167 };
      { decode_v_r[15:0] } <= { N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170 };
      { addr_v_r[27:0] } <= { N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186 };
      { data_v_r[31:0] } <= { N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214 };
      { valid_v_r[1:0] } <= { N247, N246 };
    end 
  end


endmodule

