

module top
(
  clk_i,
  reset_i,
  calibration_done_i,
  channel_active_i,
  in_v_i,
  in_data_i,
  in_yumi_o,
  in_v_o,
  in_data_o,
  in_yumi_i,
  out_me_v_i,
  out_me_data_i,
  out_me_ready_o,
  out_me_v_o,
  out_me_data_o,
  out_me_ready_i
);

  input [15:0] channel_active_i;
  input [15:0] in_v_i;
  input [511:0] in_data_i;
  output [15:0] in_yumi_o;
  output [15:0] in_v_o;
  output [511:0] in_data_o;
  input [15:0] in_yumi_i;
  input [15:0] out_me_v_i;
  input [511:0] out_me_data_i;
  output [15:0] out_me_ready_o;
  output [15:0] out_me_v_o;
  output [511:0] out_me_data_o;
  input [15:0] out_me_ready_i;
  input clk_i;
  input reset_i;
  input calibration_done_i;

  bsg_sbox
  wrapper
  (
    .channel_active_i(channel_active_i),
    .in_v_i(in_v_i),
    .in_data_i(in_data_i),
    .in_yumi_o(in_yumi_o),
    .in_v_o(in_v_o),
    .in_data_o(in_data_o),
    .in_yumi_i(in_yumi_i),
    .out_me_v_i(out_me_v_i),
    .out_me_data_i(out_me_data_i),
    .out_me_ready_o(out_me_ready_o),
    .out_me_v_o(out_me_v_o),
    .out_me_data_o(out_me_data_o),
    .out_me_ready_i(out_me_ready_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .calibration_done_i(calibration_done_i)
  );


endmodule



module bsg_scatter_gather_vec_size_lp16
(
  vec_i,
  fwd_o,
  fwd_datapath_o,
  bk_o,
  bk_datapath_o
);

  input [15:0] vec_i;
  output [63:0] fwd_o;
  output [63:0] fwd_datapath_o;
  output [63:0] bk_o;
  output [63:0] bk_datapath_o;
  wire [63:0] fwd_o,fwd_datapath_o,bk_o,bk_datapath_o;

endmodule



module bsg_sbox
(
  clk_i,
  reset_i,
  calibration_done_i,
  channel_active_i,
  in_v_i,
  in_data_i,
  in_yumi_o,
  in_v_o,
  in_data_o,
  in_yumi_i,
  out_me_v_i,
  out_me_data_i,
  out_me_ready_o,
  out_me_v_o,
  out_me_data_o,
  out_me_ready_i
);

  input [15:0] channel_active_i;
  input [15:0] in_v_i;
  input [511:0] in_data_i;
  output [15:0] in_yumi_o;
  output [15:0] in_v_o;
  output [511:0] in_data_o;
  input [15:0] in_yumi_i;
  input [15:0] out_me_v_i;
  input [511:0] out_me_data_i;
  output [15:0] out_me_ready_o;
  output [15:0] out_me_v_o;
  output [511:0] out_me_data_o;
  input [15:0] out_me_ready_i;
  input clk_i;
  input reset_i;
  input calibration_done_i;
  wire [15:0] in_yumi_o,in_v_o,out_me_ready_o,out_me_v_o;
  wire [511:0] in_data_o,out_me_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,in_data_i_15__31_,in_data_i_15__30_,in_data_i_15__29_,
  in_data_i_15__28_,in_data_i_15__27_,in_data_i_15__26_,in_data_i_15__25_,
  in_data_i_15__24_,in_data_i_15__23_,in_data_i_15__22_,in_data_i_15__21_,in_data_i_15__20_,
  in_data_i_15__19_,in_data_i_15__18_,in_data_i_15__17_,in_data_i_15__16_,
  in_data_i_15__15_,in_data_i_15__14_,in_data_i_15__13_,in_data_i_15__12_,in_data_i_15__11_,
  in_data_i_15__10_,in_data_i_15__9_,in_data_i_15__8_,in_data_i_15__7_,
  in_data_i_15__6_,in_data_i_15__5_,in_data_i_15__4_,in_data_i_15__3_,in_data_i_15__2_,
  in_data_i_15__1_,in_data_i_15__0_,out_me_data_i_0__31_,out_me_data_i_0__30_,
  out_me_data_i_0__29_,out_me_data_i_0__28_,out_me_data_i_0__27_,out_me_data_i_0__26_,
  out_me_data_i_0__25_,out_me_data_i_0__24_,out_me_data_i_0__23_,out_me_data_i_0__22_,
  out_me_data_i_0__21_,out_me_data_i_0__20_,out_me_data_i_0__19_,out_me_data_i_0__18_,
  out_me_data_i_0__17_,out_me_data_i_0__16_,out_me_data_i_0__15_,
  out_me_data_i_0__14_,out_me_data_i_0__13_,out_me_data_i_0__12_,out_me_data_i_0__11_,
  out_me_data_i_0__10_,out_me_data_i_0__9_,out_me_data_i_0__8_,out_me_data_i_0__7_,
  out_me_data_i_0__6_,out_me_data_i_0__5_,out_me_data_i_0__4_,out_me_data_i_0__3_,
  out_me_data_i_0__2_,out_me_data_i_0__1_,out_me_data_i_0__0_,fwd_dpath_sel_r_56,
  fwd_dpath_sel_r_53,fwd_dpath_sel_r_52,fwd_dpath_sel_r_49,fwd_dpath_sel_r_48,
  fwd_dpath_sel_r_46,fwd_dpath_sel_r_45,fwd_dpath_sel_r_44,fwd_dpath_sel_r_42,fwd_dpath_sel_r_41,
  fwd_dpath_sel_r_40,fwd_dpath_sel_r_38,fwd_dpath_sel_r_37,fwd_dpath_sel_r_36,
  bk_dpath_sel_r_30,bk_dpath_sel_r_29,bk_dpath_sel_r_28,bk_dpath_sel_r_26,
  bk_dpath_sel_r_25,bk_dpath_sel_r_24,bk_dpath_sel_r_22,bk_dpath_sel_r_21,bk_dpath_sel_r_20,
  bk_dpath_sel_r_18,bk_dpath_sel_r_17,bk_dpath_sel_r_16,bk_dpath_sel_r_13,
  bk_dpath_sel_r_12,bk_dpath_sel_r_9,bk_dpath_sel_r_8,bk_dpath_sel_r_4,N538,N539,N540,N541,
  N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__15_ ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__14_ ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__13_ ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__12_ ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__11_ ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__10_ ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__9_ ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__8_ ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__7_ ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__6_ ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__5_ ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__4_ ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__3_ ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__2_ ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__1_ ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__0_ ,
  N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,
  N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,
  N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,
  N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,
  N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,
  N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,
  N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,
  N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,
  N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__15_ ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__14_ ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__13_ ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__12_ ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__11_ ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__10_ ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__9_ ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__8_ ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__7_ ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__6_ ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__5_ ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__4_ ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__3_ ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__2_ ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__1_ ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__0_ ,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,
  N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,
  N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,
  N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,
  N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,
  N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,
  N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,
  N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__15_ ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__14_ ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__13_ ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__12_ ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__11_ ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__10_ ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__9_ ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__8_ ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__7_ ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__6_ ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__5_ ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__4_ ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__3_ ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__2_ ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__1_ ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__0_ ,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__15_ ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__14_ ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__13_ ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__12_ ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__11_ ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__10_ ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__9_ ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__8_ ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__7_ ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__6_ ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__5_ ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__4_ ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__3_ ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__2_ ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__1_ ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__0_ ,
  N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,
  N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,
  N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,
  N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,
  N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,
  N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,
  N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,
  N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,
  N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__15_ ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__14_ ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__13_ ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__12_ ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__11_ ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__10_ ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__9_ ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__8_ ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__7_ ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__6_ ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__5_ ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__4_ ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__3_ ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__2_ ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__1_ ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__0_ ,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,
  N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,
  N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,
  N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,
  N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,
  N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,
  N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
  N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,
  N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,
  N1187,N1188,N1189,N1190,N1191,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__15_ ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__14_ ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__13_ ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__12_ ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__11_ ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__10_ ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__9_ ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__8_ ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__7_ ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__6_ ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__5_ ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__4_ ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__3_ ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__2_ ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__1_ ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__0_ ,N1192,N1193,N1194,N1195,
  N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,
  N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,
  N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,
  N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,
  N1316,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__15_ ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__14_ ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__13_ ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__12_ ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__11_ ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__10_ ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__9_ ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__8_ ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__7_ ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__6_ ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__5_ ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__4_ ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__3_ ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__2_ ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__1_ ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__0_ ,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__15_ ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__14_ ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__13_ ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__12_ ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__11_ ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__10_ ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__9_ ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__8_ ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__7_ ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__6_ ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__5_ ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__4_ ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__3_ ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__2_ ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__1_ ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__0_ ,
  N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,
  N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,
  N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,
  N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,
  N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,
  N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,
  N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,
  N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
  N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,
  N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__15_ ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__14_ ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__13_ ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__12_ ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__11_ ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__10_ ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__9_ ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__8_ ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__7_ ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__6_ ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__5_ ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__4_ ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__3_ ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__2_ ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__1_ ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__0_ ,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,
  N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,
  N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,
  N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,
  N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,
  N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,
  N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__15_ ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__14_ ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__13_ ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__12_ ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__11_ ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__10_ ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__9_ ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__8_ ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__7_ ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__6_ ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__5_ ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__4_ ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__3_ ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__2_ ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__1_ ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__0_ ,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,
  N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,
  N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,
  N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,
  N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,
  N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,
  N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,
  N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,
  N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,
  N1822,N1823,N1824,N1825,N1826,N1827,N1828,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__15_ ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__14_ ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__13_ ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__12_ ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__11_ ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__10_ ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__9_ ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__8_ ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__7_ ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__6_ ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__5_ ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__4_ ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__3_ ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__2_ ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__1_ ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__0_ ,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,
  N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,
  N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,
  N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,
  N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,
  N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,
  N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
  N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,
  N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,
  N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__15_ ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__14_ ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__13_ ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__12_ ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__11_ ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__10_ ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__9_ ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__8_ ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__7_ ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__6_ ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__5_ ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__4_ ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__3_ ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__2_ ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__1_ ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__0_ ,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,
  N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,
  N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,
  N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,
  N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,
  N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,
  N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,
  N2044,N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,
  N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,
  N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__15_ ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__14_ ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__13_ ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__12_ ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__11_ ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__10_ ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__9_ ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__8_ ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__7_ ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__6_ ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__5_ ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__4_ ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__3_ ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__2_ ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__1_ ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__0_ ,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,
  N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,
  N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,
  N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,
  N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,
  N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,
  N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,
  N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,
  N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,
  N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__15_ ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__14_ ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__13_ ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__12_ ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__11_ ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__10_ ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__9_ ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__8_ ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__7_ ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__6_ ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__5_ ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__4_ ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__3_ ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__2_ ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__1_ ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__0_ ,N2205,N2206,N2207,N2208,N2209,N2210,N2211,
  N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,N2225,
  N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,
  N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,
  N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,N2265,
  N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,
  N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,N2291,
  N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,N2305,
  N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
  N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__15_ ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__14_ ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__13_ ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__12_ ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__11_ ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__10_ ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__9_ ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__8_ ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__7_ ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__6_ ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__5_ ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__4_ ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__3_ ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__2_ ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__1_ ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__0_ ,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,
  N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,
  N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,
  N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,
  N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,
  N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,
  N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,
  N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,
  N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,
  N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,N2451,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__15_ ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__14_ ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__13_ ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__12_ ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__11_ ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__10_ ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__9_ ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__8_ ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__7_ ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__6_ ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__5_ ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__4_ ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__3_ ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__2_ ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__1_ ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__0_ ,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,
  N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,
  N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,
  N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,
  N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,
  N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,
  N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,
  N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,
  N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,
  N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,
  N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,
  N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,
  N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,
  N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,
  N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,
  N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,
  N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,
  N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,
  N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,
  N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,
  N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,
  N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,
  N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,
  N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,
  N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,
  N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,
  N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,
  N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,
  N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,
  N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,
  N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,
  N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,
  N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,
  N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
  N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,
  N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,
  N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,
  N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,
  N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,
  N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,
  N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,
  N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,
  N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,
  N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,
  N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,
  N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055;
  wire [63:0] fwd_sel,fwd_dpath_sel,bk_sel,bk_dpath_sel,fwd_sel_r,bk_sel_r;
  wire [34:0] fwd_dpath_sel_r;
  wire [63:32] bk_dpath_sel_r;
  reg fwd_sel_r_63_sv2v_reg,fwd_sel_r_62_sv2v_reg,fwd_sel_r_61_sv2v_reg,
  fwd_sel_r_60_sv2v_reg,fwd_sel_r_59_sv2v_reg,fwd_sel_r_58_sv2v_reg,fwd_sel_r_57_sv2v_reg,
  fwd_sel_r_56_sv2v_reg,fwd_sel_r_55_sv2v_reg,fwd_sel_r_54_sv2v_reg,
  fwd_sel_r_53_sv2v_reg,fwd_sel_r_52_sv2v_reg,fwd_sel_r_51_sv2v_reg,fwd_sel_r_50_sv2v_reg,
  fwd_sel_r_49_sv2v_reg,fwd_sel_r_48_sv2v_reg,fwd_sel_r_47_sv2v_reg,fwd_sel_r_46_sv2v_reg,
  fwd_sel_r_45_sv2v_reg,fwd_sel_r_44_sv2v_reg,fwd_sel_r_43_sv2v_reg,
  fwd_sel_r_42_sv2v_reg,fwd_sel_r_41_sv2v_reg,fwd_sel_r_40_sv2v_reg,fwd_sel_r_39_sv2v_reg,
  fwd_sel_r_38_sv2v_reg,fwd_sel_r_37_sv2v_reg,fwd_sel_r_36_sv2v_reg,fwd_sel_r_35_sv2v_reg,
  fwd_sel_r_34_sv2v_reg,fwd_sel_r_33_sv2v_reg,fwd_sel_r_32_sv2v_reg,
  fwd_sel_r_31_sv2v_reg,fwd_sel_r_30_sv2v_reg,fwd_sel_r_29_sv2v_reg,fwd_sel_r_28_sv2v_reg,
  fwd_sel_r_27_sv2v_reg,fwd_sel_r_26_sv2v_reg,fwd_sel_r_25_sv2v_reg,fwd_sel_r_24_sv2v_reg,
  fwd_sel_r_23_sv2v_reg,fwd_sel_r_22_sv2v_reg,fwd_sel_r_21_sv2v_reg,
  fwd_sel_r_20_sv2v_reg,fwd_sel_r_19_sv2v_reg,fwd_sel_r_18_sv2v_reg,fwd_sel_r_17_sv2v_reg,
  fwd_sel_r_16_sv2v_reg,fwd_sel_r_15_sv2v_reg,fwd_sel_r_14_sv2v_reg,
  fwd_sel_r_13_sv2v_reg,fwd_sel_r_12_sv2v_reg,fwd_sel_r_11_sv2v_reg,fwd_sel_r_10_sv2v_reg,
  fwd_sel_r_9_sv2v_reg,fwd_sel_r_8_sv2v_reg,fwd_sel_r_7_sv2v_reg,fwd_sel_r_6_sv2v_reg,
  fwd_sel_r_5_sv2v_reg,fwd_sel_r_4_sv2v_reg,fwd_sel_r_3_sv2v_reg,fwd_sel_r_2_sv2v_reg,
  fwd_sel_r_1_sv2v_reg,fwd_sel_r_0_sv2v_reg,fwd_dpath_sel_r_56_sv2v_reg,
  fwd_dpath_sel_r_53_sv2v_reg,fwd_dpath_sel_r_52_sv2v_reg,fwd_dpath_sel_r_49_sv2v_reg,
  fwd_dpath_sel_r_48_sv2v_reg,fwd_dpath_sel_r_46_sv2v_reg,fwd_dpath_sel_r_45_sv2v_reg,
  fwd_dpath_sel_r_44_sv2v_reg,fwd_dpath_sel_r_42_sv2v_reg,fwd_dpath_sel_r_41_sv2v_reg,
  fwd_dpath_sel_r_40_sv2v_reg,fwd_dpath_sel_r_38_sv2v_reg,
  fwd_dpath_sel_r_37_sv2v_reg,fwd_dpath_sel_r_36_sv2v_reg,fwd_dpath_sel_r_34_sv2v_reg,
  fwd_dpath_sel_r_33_sv2v_reg,fwd_dpath_sel_r_32_sv2v_reg,fwd_dpath_sel_r_31_sv2v_reg,
  fwd_dpath_sel_r_30_sv2v_reg,fwd_dpath_sel_r_29_sv2v_reg,fwd_dpath_sel_r_28_sv2v_reg,
  fwd_dpath_sel_r_27_sv2v_reg,fwd_dpath_sel_r_26_sv2v_reg,fwd_dpath_sel_r_25_sv2v_reg,
  fwd_dpath_sel_r_24_sv2v_reg,fwd_dpath_sel_r_23_sv2v_reg,fwd_dpath_sel_r_22_sv2v_reg,
  fwd_dpath_sel_r_21_sv2v_reg,fwd_dpath_sel_r_20_sv2v_reg,fwd_dpath_sel_r_19_sv2v_reg,
  fwd_dpath_sel_r_18_sv2v_reg,fwd_dpath_sel_r_17_sv2v_reg,
  fwd_dpath_sel_r_16_sv2v_reg,fwd_dpath_sel_r_15_sv2v_reg,fwd_dpath_sel_r_14_sv2v_reg,
  fwd_dpath_sel_r_13_sv2v_reg,fwd_dpath_sel_r_12_sv2v_reg,fwd_dpath_sel_r_11_sv2v_reg,
  fwd_dpath_sel_r_10_sv2v_reg,fwd_dpath_sel_r_9_sv2v_reg,fwd_dpath_sel_r_8_sv2v_reg,
  fwd_dpath_sel_r_7_sv2v_reg,fwd_dpath_sel_r_6_sv2v_reg,fwd_dpath_sel_r_5_sv2v_reg,
  fwd_dpath_sel_r_4_sv2v_reg,fwd_dpath_sel_r_3_sv2v_reg,fwd_dpath_sel_r_2_sv2v_reg,
  fwd_dpath_sel_r_1_sv2v_reg,fwd_dpath_sel_r_0_sv2v_reg,bk_sel_r_63_sv2v_reg,
  bk_sel_r_62_sv2v_reg,bk_sel_r_61_sv2v_reg,bk_sel_r_60_sv2v_reg,bk_sel_r_59_sv2v_reg,
  bk_sel_r_58_sv2v_reg,bk_sel_r_57_sv2v_reg,bk_sel_r_56_sv2v_reg,bk_sel_r_55_sv2v_reg,
  bk_sel_r_54_sv2v_reg,bk_sel_r_53_sv2v_reg,bk_sel_r_52_sv2v_reg,bk_sel_r_51_sv2v_reg,
  bk_sel_r_50_sv2v_reg,bk_sel_r_49_sv2v_reg,bk_sel_r_48_sv2v_reg,bk_sel_r_47_sv2v_reg,
  bk_sel_r_46_sv2v_reg,bk_sel_r_45_sv2v_reg,bk_sel_r_44_sv2v_reg,
  bk_sel_r_43_sv2v_reg,bk_sel_r_42_sv2v_reg,bk_sel_r_41_sv2v_reg,bk_sel_r_40_sv2v_reg,
  bk_sel_r_39_sv2v_reg,bk_sel_r_38_sv2v_reg,bk_sel_r_37_sv2v_reg,bk_sel_r_36_sv2v_reg,
  bk_sel_r_35_sv2v_reg,bk_sel_r_34_sv2v_reg,bk_sel_r_33_sv2v_reg,bk_sel_r_32_sv2v_reg,
  bk_sel_r_31_sv2v_reg,bk_sel_r_30_sv2v_reg,bk_sel_r_29_sv2v_reg,bk_sel_r_28_sv2v_reg,
  bk_sel_r_27_sv2v_reg,bk_sel_r_26_sv2v_reg,bk_sel_r_25_sv2v_reg,bk_sel_r_24_sv2v_reg,
  bk_sel_r_23_sv2v_reg,bk_sel_r_22_sv2v_reg,bk_sel_r_21_sv2v_reg,
  bk_sel_r_20_sv2v_reg,bk_sel_r_19_sv2v_reg,bk_sel_r_18_sv2v_reg,bk_sel_r_17_sv2v_reg,
  bk_sel_r_16_sv2v_reg,bk_sel_r_15_sv2v_reg,bk_sel_r_14_sv2v_reg,bk_sel_r_13_sv2v_reg,
  bk_sel_r_12_sv2v_reg,bk_sel_r_11_sv2v_reg,bk_sel_r_10_sv2v_reg,bk_sel_r_9_sv2v_reg,
  bk_sel_r_8_sv2v_reg,bk_sel_r_7_sv2v_reg,bk_sel_r_6_sv2v_reg,bk_sel_r_5_sv2v_reg,
  bk_sel_r_4_sv2v_reg,bk_sel_r_3_sv2v_reg,bk_sel_r_2_sv2v_reg,bk_sel_r_1_sv2v_reg,
  bk_sel_r_0_sv2v_reg,bk_dpath_sel_r_63_sv2v_reg,bk_dpath_sel_r_62_sv2v_reg,
  bk_dpath_sel_r_61_sv2v_reg,bk_dpath_sel_r_60_sv2v_reg,bk_dpath_sel_r_59_sv2v_reg,
  bk_dpath_sel_r_58_sv2v_reg,bk_dpath_sel_r_57_sv2v_reg,bk_dpath_sel_r_56_sv2v_reg,
  bk_dpath_sel_r_55_sv2v_reg,bk_dpath_sel_r_54_sv2v_reg,bk_dpath_sel_r_53_sv2v_reg,
  bk_dpath_sel_r_52_sv2v_reg,bk_dpath_sel_r_51_sv2v_reg,bk_dpath_sel_r_50_sv2v_reg,
  bk_dpath_sel_r_49_sv2v_reg,bk_dpath_sel_r_48_sv2v_reg,bk_dpath_sel_r_47_sv2v_reg,
  bk_dpath_sel_r_46_sv2v_reg,bk_dpath_sel_r_45_sv2v_reg,bk_dpath_sel_r_44_sv2v_reg,
  bk_dpath_sel_r_43_sv2v_reg,bk_dpath_sel_r_42_sv2v_reg,bk_dpath_sel_r_41_sv2v_reg,
  bk_dpath_sel_r_40_sv2v_reg,bk_dpath_sel_r_39_sv2v_reg,bk_dpath_sel_r_38_sv2v_reg,
  bk_dpath_sel_r_37_sv2v_reg,bk_dpath_sel_r_36_sv2v_reg,bk_dpath_sel_r_35_sv2v_reg,
  bk_dpath_sel_r_34_sv2v_reg,bk_dpath_sel_r_33_sv2v_reg,bk_dpath_sel_r_32_sv2v_reg,
  bk_dpath_sel_r_30_sv2v_reg,bk_dpath_sel_r_29_sv2v_reg,bk_dpath_sel_r_28_sv2v_reg,
  bk_dpath_sel_r_26_sv2v_reg,bk_dpath_sel_r_25_sv2v_reg,bk_dpath_sel_r_24_sv2v_reg,
  bk_dpath_sel_r_22_sv2v_reg,bk_dpath_sel_r_21_sv2v_reg,
  bk_dpath_sel_r_20_sv2v_reg,bk_dpath_sel_r_18_sv2v_reg,bk_dpath_sel_r_17_sv2v_reg,
  bk_dpath_sel_r_16_sv2v_reg,bk_dpath_sel_r_13_sv2v_reg,bk_dpath_sel_r_12_sv2v_reg,
  bk_dpath_sel_r_9_sv2v_reg,bk_dpath_sel_r_8_sv2v_reg,bk_dpath_sel_r_4_sv2v_reg,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__15__sv2v_reg ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__14__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__13__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__12__sv2v_reg ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__11__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__10__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__9__sv2v_reg ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__8__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__7__sv2v_reg ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__6__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__5__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__4__sv2v_reg ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__3__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__2__sv2v_reg ,
  \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__1__sv2v_reg ,\sbox_0_.fi1hot.fwd_sel_one_hot_r_0__0__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__15__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__14__sv2v_reg ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__13__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__12__sv2v_reg ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__11__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__10__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__9__sv2v_reg ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__8__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__7__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__6__sv2v_reg ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__5__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__4__sv2v_reg ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__3__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__2__sv2v_reg ,
  \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__1__sv2v_reg ,\sbox_1_.fi1hot.fwd_sel_one_hot_r_1__0__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__15__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__14__sv2v_reg ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__13__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__12__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__11__sv2v_reg ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__10__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__9__sv2v_reg ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__8__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__7__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__6__sv2v_reg ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__5__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__4__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__3__sv2v_reg ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__2__sv2v_reg ,
  \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__1__sv2v_reg ,\sbox_2_.fi1hot.fwd_sel_one_hot_r_2__0__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__15__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__14__sv2v_reg ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__13__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__12__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__11__sv2v_reg ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__10__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__9__sv2v_reg ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__8__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__7__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__6__sv2v_reg ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__5__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__4__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__3__sv2v_reg ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__2__sv2v_reg ,
  \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__1__sv2v_reg ,\sbox_3_.fi1hot.fwd_sel_one_hot_r_3__0__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__15__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__14__sv2v_reg ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__13__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__12__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__11__sv2v_reg ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__10__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__9__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__8__sv2v_reg ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__7__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__6__sv2v_reg ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__5__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__4__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__3__sv2v_reg ,\sbox_4_.fi1hot.fwd_sel_one_hot_r_4__2__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__1__sv2v_reg ,
  \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__0__sv2v_reg ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__15__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__14__sv2v_reg ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__13__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__12__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__11__sv2v_reg ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__10__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__9__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__8__sv2v_reg ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__7__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__6__sv2v_reg ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__5__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__4__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__3__sv2v_reg ,\sbox_5_.fi1hot.fwd_sel_one_hot_r_5__2__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__1__sv2v_reg ,
  \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__0__sv2v_reg ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__15__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__14__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__13__sv2v_reg ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__12__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__11__sv2v_reg ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__10__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__9__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__8__sv2v_reg ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__7__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__6__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__5__sv2v_reg ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__4__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__3__sv2v_reg ,\sbox_6_.fi1hot.fwd_sel_one_hot_r_6__2__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__1__sv2v_reg ,
  \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__0__sv2v_reg ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__15__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__14__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__13__sv2v_reg ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__12__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__11__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__10__sv2v_reg ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__9__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__8__sv2v_reg ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__7__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__6__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__5__sv2v_reg ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__4__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__3__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__2__sv2v_reg ,\sbox_7_.fi1hot.fwd_sel_one_hot_r_7__1__sv2v_reg ,
  \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__0__sv2v_reg ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__15__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__14__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__13__sv2v_reg ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__12__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__11__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__10__sv2v_reg ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__9__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__8__sv2v_reg ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__7__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__6__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__5__sv2v_reg ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__4__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__3__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__2__sv2v_reg ,\sbox_8_.fi1hot.fwd_sel_one_hot_r_8__1__sv2v_reg ,
  \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__0__sv2v_reg ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__15__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__14__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__13__sv2v_reg ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__12__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__11__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__10__sv2v_reg ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__9__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__8__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__7__sv2v_reg ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__6__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__5__sv2v_reg ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__4__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__3__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__2__sv2v_reg ,\sbox_9_.fi1hot.fwd_sel_one_hot_r_9__1__sv2v_reg ,
  \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__0__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__15__sv2v_reg ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__14__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__13__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__12__sv2v_reg ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__11__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__10__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__9__sv2v_reg ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__8__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__7__sv2v_reg ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__6__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__5__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__4__sv2v_reg ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__3__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__2__sv2v_reg ,
  \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__1__sv2v_reg ,\sbox_10_.fi1hot.fwd_sel_one_hot_r_10__0__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__15__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__14__sv2v_reg ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__13__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__12__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__11__sv2v_reg ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__10__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__9__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__8__sv2v_reg ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__7__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__6__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__5__sv2v_reg ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__4__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__3__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__2__sv2v_reg ,\sbox_11_.fi1hot.fwd_sel_one_hot_r_11__1__sv2v_reg ,
  \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__0__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__15__sv2v_reg ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__14__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__13__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__12__sv2v_reg ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__11__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__10__sv2v_reg ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__9__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__8__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__7__sv2v_reg ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__6__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__5__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__4__sv2v_reg ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__3__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__2__sv2v_reg ,
  \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__1__sv2v_reg ,\sbox_12_.fi1hot.fwd_sel_one_hot_r_12__0__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__15__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__14__sv2v_reg ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__13__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__12__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__11__sv2v_reg ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__10__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__9__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__8__sv2v_reg ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__7__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__6__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__5__sv2v_reg ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__4__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__3__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__2__sv2v_reg ,\sbox_13_.fi1hot.fwd_sel_one_hot_r_13__1__sv2v_reg ,
  \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__0__sv2v_reg ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__15__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__14__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__13__sv2v_reg ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__12__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__11__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__10__sv2v_reg ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__9__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__8__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__7__sv2v_reg ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__6__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__5__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__4__sv2v_reg ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__3__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__2__sv2v_reg ,
  \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__1__sv2v_reg ,\sbox_14_.fi1hot.fwd_sel_one_hot_r_14__0__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__15__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__14__sv2v_reg ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__13__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__12__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__11__sv2v_reg ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__10__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__9__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__8__sv2v_reg ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__7__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__6__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__5__sv2v_reg ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__4__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__3__sv2v_reg ,\sbox_15_.fi1hot.fwd_sel_one_hot_r_15__2__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__1__sv2v_reg ,
  \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__0__sv2v_reg ;
  assign fwd_sel_r[63] = fwd_sel_r_63_sv2v_reg;
  assign fwd_sel_r[62] = fwd_sel_r_62_sv2v_reg;
  assign fwd_sel_r[61] = fwd_sel_r_61_sv2v_reg;
  assign fwd_sel_r[60] = fwd_sel_r_60_sv2v_reg;
  assign fwd_sel_r[59] = fwd_sel_r_59_sv2v_reg;
  assign fwd_sel_r[58] = fwd_sel_r_58_sv2v_reg;
  assign fwd_sel_r[57] = fwd_sel_r_57_sv2v_reg;
  assign fwd_sel_r[56] = fwd_sel_r_56_sv2v_reg;
  assign fwd_sel_r[55] = fwd_sel_r_55_sv2v_reg;
  assign fwd_sel_r[54] = fwd_sel_r_54_sv2v_reg;
  assign fwd_sel_r[53] = fwd_sel_r_53_sv2v_reg;
  assign fwd_sel_r[52] = fwd_sel_r_52_sv2v_reg;
  assign fwd_sel_r[51] = fwd_sel_r_51_sv2v_reg;
  assign fwd_sel_r[50] = fwd_sel_r_50_sv2v_reg;
  assign fwd_sel_r[49] = fwd_sel_r_49_sv2v_reg;
  assign fwd_sel_r[48] = fwd_sel_r_48_sv2v_reg;
  assign fwd_sel_r[47] = fwd_sel_r_47_sv2v_reg;
  assign fwd_sel_r[46] = fwd_sel_r_46_sv2v_reg;
  assign fwd_sel_r[45] = fwd_sel_r_45_sv2v_reg;
  assign fwd_sel_r[44] = fwd_sel_r_44_sv2v_reg;
  assign fwd_sel_r[43] = fwd_sel_r_43_sv2v_reg;
  assign fwd_sel_r[42] = fwd_sel_r_42_sv2v_reg;
  assign fwd_sel_r[41] = fwd_sel_r_41_sv2v_reg;
  assign fwd_sel_r[40] = fwd_sel_r_40_sv2v_reg;
  assign fwd_sel_r[39] = fwd_sel_r_39_sv2v_reg;
  assign fwd_sel_r[38] = fwd_sel_r_38_sv2v_reg;
  assign fwd_sel_r[37] = fwd_sel_r_37_sv2v_reg;
  assign fwd_sel_r[36] = fwd_sel_r_36_sv2v_reg;
  assign fwd_sel_r[35] = fwd_sel_r_35_sv2v_reg;
  assign fwd_sel_r[34] = fwd_sel_r_34_sv2v_reg;
  assign fwd_sel_r[33] = fwd_sel_r_33_sv2v_reg;
  assign fwd_sel_r[32] = fwd_sel_r_32_sv2v_reg;
  assign fwd_sel_r[31] = fwd_sel_r_31_sv2v_reg;
  assign fwd_sel_r[30] = fwd_sel_r_30_sv2v_reg;
  assign fwd_sel_r[29] = fwd_sel_r_29_sv2v_reg;
  assign fwd_sel_r[28] = fwd_sel_r_28_sv2v_reg;
  assign fwd_sel_r[27] = fwd_sel_r_27_sv2v_reg;
  assign fwd_sel_r[26] = fwd_sel_r_26_sv2v_reg;
  assign fwd_sel_r[25] = fwd_sel_r_25_sv2v_reg;
  assign fwd_sel_r[24] = fwd_sel_r_24_sv2v_reg;
  assign fwd_sel_r[23] = fwd_sel_r_23_sv2v_reg;
  assign fwd_sel_r[22] = fwd_sel_r_22_sv2v_reg;
  assign fwd_sel_r[21] = fwd_sel_r_21_sv2v_reg;
  assign fwd_sel_r[20] = fwd_sel_r_20_sv2v_reg;
  assign fwd_sel_r[19] = fwd_sel_r_19_sv2v_reg;
  assign fwd_sel_r[18] = fwd_sel_r_18_sv2v_reg;
  assign fwd_sel_r[17] = fwd_sel_r_17_sv2v_reg;
  assign fwd_sel_r[16] = fwd_sel_r_16_sv2v_reg;
  assign fwd_sel_r[15] = fwd_sel_r_15_sv2v_reg;
  assign fwd_sel_r[14] = fwd_sel_r_14_sv2v_reg;
  assign fwd_sel_r[13] = fwd_sel_r_13_sv2v_reg;
  assign fwd_sel_r[12] = fwd_sel_r_12_sv2v_reg;
  assign fwd_sel_r[11] = fwd_sel_r_11_sv2v_reg;
  assign fwd_sel_r[10] = fwd_sel_r_10_sv2v_reg;
  assign fwd_sel_r[9] = fwd_sel_r_9_sv2v_reg;
  assign fwd_sel_r[8] = fwd_sel_r_8_sv2v_reg;
  assign fwd_sel_r[7] = fwd_sel_r_7_sv2v_reg;
  assign fwd_sel_r[6] = fwd_sel_r_6_sv2v_reg;
  assign fwd_sel_r[5] = fwd_sel_r_5_sv2v_reg;
  assign fwd_sel_r[4] = fwd_sel_r_4_sv2v_reg;
  assign fwd_sel_r[3] = fwd_sel_r_3_sv2v_reg;
  assign fwd_sel_r[2] = fwd_sel_r_2_sv2v_reg;
  assign fwd_sel_r[1] = fwd_sel_r_1_sv2v_reg;
  assign fwd_sel_r[0] = fwd_sel_r_0_sv2v_reg;
  assign fwd_dpath_sel_r_56 = fwd_dpath_sel_r_56_sv2v_reg;
  assign fwd_dpath_sel_r_53 = fwd_dpath_sel_r_53_sv2v_reg;
  assign fwd_dpath_sel_r_52 = fwd_dpath_sel_r_52_sv2v_reg;
  assign fwd_dpath_sel_r_49 = fwd_dpath_sel_r_49_sv2v_reg;
  assign fwd_dpath_sel_r_48 = fwd_dpath_sel_r_48_sv2v_reg;
  assign fwd_dpath_sel_r_46 = fwd_dpath_sel_r_46_sv2v_reg;
  assign fwd_dpath_sel_r_45 = fwd_dpath_sel_r_45_sv2v_reg;
  assign fwd_dpath_sel_r_44 = fwd_dpath_sel_r_44_sv2v_reg;
  assign fwd_dpath_sel_r_42 = fwd_dpath_sel_r_42_sv2v_reg;
  assign fwd_dpath_sel_r_41 = fwd_dpath_sel_r_41_sv2v_reg;
  assign fwd_dpath_sel_r_40 = fwd_dpath_sel_r_40_sv2v_reg;
  assign fwd_dpath_sel_r_38 = fwd_dpath_sel_r_38_sv2v_reg;
  assign fwd_dpath_sel_r_37 = fwd_dpath_sel_r_37_sv2v_reg;
  assign fwd_dpath_sel_r_36 = fwd_dpath_sel_r_36_sv2v_reg;
  assign fwd_dpath_sel_r[34] = fwd_dpath_sel_r_34_sv2v_reg;
  assign fwd_dpath_sel_r[33] = fwd_dpath_sel_r_33_sv2v_reg;
  assign fwd_dpath_sel_r[32] = fwd_dpath_sel_r_32_sv2v_reg;
  assign fwd_dpath_sel_r[31] = fwd_dpath_sel_r_31_sv2v_reg;
  assign fwd_dpath_sel_r[30] = fwd_dpath_sel_r_30_sv2v_reg;
  assign fwd_dpath_sel_r[29] = fwd_dpath_sel_r_29_sv2v_reg;
  assign fwd_dpath_sel_r[28] = fwd_dpath_sel_r_28_sv2v_reg;
  assign fwd_dpath_sel_r[27] = fwd_dpath_sel_r_27_sv2v_reg;
  assign fwd_dpath_sel_r[26] = fwd_dpath_sel_r_26_sv2v_reg;
  assign fwd_dpath_sel_r[25] = fwd_dpath_sel_r_25_sv2v_reg;
  assign fwd_dpath_sel_r[24] = fwd_dpath_sel_r_24_sv2v_reg;
  assign fwd_dpath_sel_r[23] = fwd_dpath_sel_r_23_sv2v_reg;
  assign fwd_dpath_sel_r[22] = fwd_dpath_sel_r_22_sv2v_reg;
  assign fwd_dpath_sel_r[21] = fwd_dpath_sel_r_21_sv2v_reg;
  assign fwd_dpath_sel_r[20] = fwd_dpath_sel_r_20_sv2v_reg;
  assign fwd_dpath_sel_r[19] = fwd_dpath_sel_r_19_sv2v_reg;
  assign fwd_dpath_sel_r[18] = fwd_dpath_sel_r_18_sv2v_reg;
  assign fwd_dpath_sel_r[17] = fwd_dpath_sel_r_17_sv2v_reg;
  assign fwd_dpath_sel_r[16] = fwd_dpath_sel_r_16_sv2v_reg;
  assign fwd_dpath_sel_r[15] = fwd_dpath_sel_r_15_sv2v_reg;
  assign fwd_dpath_sel_r[14] = fwd_dpath_sel_r_14_sv2v_reg;
  assign fwd_dpath_sel_r[13] = fwd_dpath_sel_r_13_sv2v_reg;
  assign fwd_dpath_sel_r[12] = fwd_dpath_sel_r_12_sv2v_reg;
  assign fwd_dpath_sel_r[11] = fwd_dpath_sel_r_11_sv2v_reg;
  assign fwd_dpath_sel_r[10] = fwd_dpath_sel_r_10_sv2v_reg;
  assign fwd_dpath_sel_r[9] = fwd_dpath_sel_r_9_sv2v_reg;
  assign fwd_dpath_sel_r[8] = fwd_dpath_sel_r_8_sv2v_reg;
  assign fwd_dpath_sel_r[7] = fwd_dpath_sel_r_7_sv2v_reg;
  assign fwd_dpath_sel_r[6] = fwd_dpath_sel_r_6_sv2v_reg;
  assign fwd_dpath_sel_r[5] = fwd_dpath_sel_r_5_sv2v_reg;
  assign fwd_dpath_sel_r[4] = fwd_dpath_sel_r_4_sv2v_reg;
  assign fwd_dpath_sel_r[3] = fwd_dpath_sel_r_3_sv2v_reg;
  assign fwd_dpath_sel_r[2] = fwd_dpath_sel_r_2_sv2v_reg;
  assign fwd_dpath_sel_r[1] = fwd_dpath_sel_r_1_sv2v_reg;
  assign fwd_dpath_sel_r[0] = fwd_dpath_sel_r_0_sv2v_reg;
  assign bk_sel_r[63] = bk_sel_r_63_sv2v_reg;
  assign bk_sel_r[62] = bk_sel_r_62_sv2v_reg;
  assign bk_sel_r[61] = bk_sel_r_61_sv2v_reg;
  assign bk_sel_r[60] = bk_sel_r_60_sv2v_reg;
  assign bk_sel_r[59] = bk_sel_r_59_sv2v_reg;
  assign bk_sel_r[58] = bk_sel_r_58_sv2v_reg;
  assign bk_sel_r[57] = bk_sel_r_57_sv2v_reg;
  assign bk_sel_r[56] = bk_sel_r_56_sv2v_reg;
  assign bk_sel_r[55] = bk_sel_r_55_sv2v_reg;
  assign bk_sel_r[54] = bk_sel_r_54_sv2v_reg;
  assign bk_sel_r[53] = bk_sel_r_53_sv2v_reg;
  assign bk_sel_r[52] = bk_sel_r_52_sv2v_reg;
  assign bk_sel_r[51] = bk_sel_r_51_sv2v_reg;
  assign bk_sel_r[50] = bk_sel_r_50_sv2v_reg;
  assign bk_sel_r[49] = bk_sel_r_49_sv2v_reg;
  assign bk_sel_r[48] = bk_sel_r_48_sv2v_reg;
  assign bk_sel_r[47] = bk_sel_r_47_sv2v_reg;
  assign bk_sel_r[46] = bk_sel_r_46_sv2v_reg;
  assign bk_sel_r[45] = bk_sel_r_45_sv2v_reg;
  assign bk_sel_r[44] = bk_sel_r_44_sv2v_reg;
  assign bk_sel_r[43] = bk_sel_r_43_sv2v_reg;
  assign bk_sel_r[42] = bk_sel_r_42_sv2v_reg;
  assign bk_sel_r[41] = bk_sel_r_41_sv2v_reg;
  assign bk_sel_r[40] = bk_sel_r_40_sv2v_reg;
  assign bk_sel_r[39] = bk_sel_r_39_sv2v_reg;
  assign bk_sel_r[38] = bk_sel_r_38_sv2v_reg;
  assign bk_sel_r[37] = bk_sel_r_37_sv2v_reg;
  assign bk_sel_r[36] = bk_sel_r_36_sv2v_reg;
  assign bk_sel_r[35] = bk_sel_r_35_sv2v_reg;
  assign bk_sel_r[34] = bk_sel_r_34_sv2v_reg;
  assign bk_sel_r[33] = bk_sel_r_33_sv2v_reg;
  assign bk_sel_r[32] = bk_sel_r_32_sv2v_reg;
  assign bk_sel_r[31] = bk_sel_r_31_sv2v_reg;
  assign bk_sel_r[30] = bk_sel_r_30_sv2v_reg;
  assign bk_sel_r[29] = bk_sel_r_29_sv2v_reg;
  assign bk_sel_r[28] = bk_sel_r_28_sv2v_reg;
  assign bk_sel_r[27] = bk_sel_r_27_sv2v_reg;
  assign bk_sel_r[26] = bk_sel_r_26_sv2v_reg;
  assign bk_sel_r[25] = bk_sel_r_25_sv2v_reg;
  assign bk_sel_r[24] = bk_sel_r_24_sv2v_reg;
  assign bk_sel_r[23] = bk_sel_r_23_sv2v_reg;
  assign bk_sel_r[22] = bk_sel_r_22_sv2v_reg;
  assign bk_sel_r[21] = bk_sel_r_21_sv2v_reg;
  assign bk_sel_r[20] = bk_sel_r_20_sv2v_reg;
  assign bk_sel_r[19] = bk_sel_r_19_sv2v_reg;
  assign bk_sel_r[18] = bk_sel_r_18_sv2v_reg;
  assign bk_sel_r[17] = bk_sel_r_17_sv2v_reg;
  assign bk_sel_r[16] = bk_sel_r_16_sv2v_reg;
  assign bk_sel_r[15] = bk_sel_r_15_sv2v_reg;
  assign bk_sel_r[14] = bk_sel_r_14_sv2v_reg;
  assign bk_sel_r[13] = bk_sel_r_13_sv2v_reg;
  assign bk_sel_r[12] = bk_sel_r_12_sv2v_reg;
  assign bk_sel_r[11] = bk_sel_r_11_sv2v_reg;
  assign bk_sel_r[10] = bk_sel_r_10_sv2v_reg;
  assign bk_sel_r[9] = bk_sel_r_9_sv2v_reg;
  assign bk_sel_r[8] = bk_sel_r_8_sv2v_reg;
  assign bk_sel_r[7] = bk_sel_r_7_sv2v_reg;
  assign bk_sel_r[6] = bk_sel_r_6_sv2v_reg;
  assign bk_sel_r[5] = bk_sel_r_5_sv2v_reg;
  assign bk_sel_r[4] = bk_sel_r_4_sv2v_reg;
  assign bk_sel_r[3] = bk_sel_r_3_sv2v_reg;
  assign bk_sel_r[2] = bk_sel_r_2_sv2v_reg;
  assign bk_sel_r[1] = bk_sel_r_1_sv2v_reg;
  assign bk_sel_r[0] = bk_sel_r_0_sv2v_reg;
  assign bk_dpath_sel_r[63] = bk_dpath_sel_r_63_sv2v_reg;
  assign bk_dpath_sel_r[62] = bk_dpath_sel_r_62_sv2v_reg;
  assign bk_dpath_sel_r[61] = bk_dpath_sel_r_61_sv2v_reg;
  assign bk_dpath_sel_r[60] = bk_dpath_sel_r_60_sv2v_reg;
  assign bk_dpath_sel_r[59] = bk_dpath_sel_r_59_sv2v_reg;
  assign bk_dpath_sel_r[58] = bk_dpath_sel_r_58_sv2v_reg;
  assign bk_dpath_sel_r[57] = bk_dpath_sel_r_57_sv2v_reg;
  assign bk_dpath_sel_r[56] = bk_dpath_sel_r_56_sv2v_reg;
  assign bk_dpath_sel_r[55] = bk_dpath_sel_r_55_sv2v_reg;
  assign bk_dpath_sel_r[54] = bk_dpath_sel_r_54_sv2v_reg;
  assign bk_dpath_sel_r[53] = bk_dpath_sel_r_53_sv2v_reg;
  assign bk_dpath_sel_r[52] = bk_dpath_sel_r_52_sv2v_reg;
  assign bk_dpath_sel_r[51] = bk_dpath_sel_r_51_sv2v_reg;
  assign bk_dpath_sel_r[50] = bk_dpath_sel_r_50_sv2v_reg;
  assign bk_dpath_sel_r[49] = bk_dpath_sel_r_49_sv2v_reg;
  assign bk_dpath_sel_r[48] = bk_dpath_sel_r_48_sv2v_reg;
  assign bk_dpath_sel_r[47] = bk_dpath_sel_r_47_sv2v_reg;
  assign bk_dpath_sel_r[46] = bk_dpath_sel_r_46_sv2v_reg;
  assign bk_dpath_sel_r[45] = bk_dpath_sel_r_45_sv2v_reg;
  assign bk_dpath_sel_r[44] = bk_dpath_sel_r_44_sv2v_reg;
  assign bk_dpath_sel_r[43] = bk_dpath_sel_r_43_sv2v_reg;
  assign bk_dpath_sel_r[42] = bk_dpath_sel_r_42_sv2v_reg;
  assign bk_dpath_sel_r[41] = bk_dpath_sel_r_41_sv2v_reg;
  assign bk_dpath_sel_r[40] = bk_dpath_sel_r_40_sv2v_reg;
  assign bk_dpath_sel_r[39] = bk_dpath_sel_r_39_sv2v_reg;
  assign bk_dpath_sel_r[38] = bk_dpath_sel_r_38_sv2v_reg;
  assign bk_dpath_sel_r[37] = bk_dpath_sel_r_37_sv2v_reg;
  assign bk_dpath_sel_r[36] = bk_dpath_sel_r_36_sv2v_reg;
  assign bk_dpath_sel_r[35] = bk_dpath_sel_r_35_sv2v_reg;
  assign bk_dpath_sel_r[34] = bk_dpath_sel_r_34_sv2v_reg;
  assign bk_dpath_sel_r[33] = bk_dpath_sel_r_33_sv2v_reg;
  assign bk_dpath_sel_r[32] = bk_dpath_sel_r_32_sv2v_reg;
  assign bk_dpath_sel_r_30 = bk_dpath_sel_r_30_sv2v_reg;
  assign bk_dpath_sel_r_29 = bk_dpath_sel_r_29_sv2v_reg;
  assign bk_dpath_sel_r_28 = bk_dpath_sel_r_28_sv2v_reg;
  assign bk_dpath_sel_r_26 = bk_dpath_sel_r_26_sv2v_reg;
  assign bk_dpath_sel_r_25 = bk_dpath_sel_r_25_sv2v_reg;
  assign bk_dpath_sel_r_24 = bk_dpath_sel_r_24_sv2v_reg;
  assign bk_dpath_sel_r_22 = bk_dpath_sel_r_22_sv2v_reg;
  assign bk_dpath_sel_r_21 = bk_dpath_sel_r_21_sv2v_reg;
  assign bk_dpath_sel_r_20 = bk_dpath_sel_r_20_sv2v_reg;
  assign bk_dpath_sel_r_18 = bk_dpath_sel_r_18_sv2v_reg;
  assign bk_dpath_sel_r_17 = bk_dpath_sel_r_17_sv2v_reg;
  assign bk_dpath_sel_r_16 = bk_dpath_sel_r_16_sv2v_reg;
  assign bk_dpath_sel_r_13 = bk_dpath_sel_r_13_sv2v_reg;
  assign bk_dpath_sel_r_12 = bk_dpath_sel_r_12_sv2v_reg;
  assign bk_dpath_sel_r_9 = bk_dpath_sel_r_9_sv2v_reg;
  assign bk_dpath_sel_r_8 = bk_dpath_sel_r_8_sv2v_reg;
  assign bk_dpath_sel_r_4 = bk_dpath_sel_r_4_sv2v_reg;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__15_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__15__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__14_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__14__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__13_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__13__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__12_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__12__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__11_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__11__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__10_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__10__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__9_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__9__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__8_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__8__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__7_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__7__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__6_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__6__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__5_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__5__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__4_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__4__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__3_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__3__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__2_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__2__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__1_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__1__sv2v_reg ;
  assign \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__0_  = \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__0__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__15_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__15__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__14_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__14__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__13_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__13__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__12_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__12__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__11_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__11__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__10_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__10__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__9_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__9__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__8_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__8__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__7_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__7__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__6_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__6__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__5_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__5__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__4_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__4__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__3_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__3__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__2_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__2__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__1_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__1__sv2v_reg ;
  assign \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__0_  = \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__0__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__15_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__15__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__14_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__14__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__13_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__13__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__12_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__12__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__11_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__11__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__10_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__10__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__9_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__9__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__8_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__8__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__7_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__7__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__6_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__6__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__5_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__5__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__4_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__4__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__3_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__3__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__2_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__2__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__1_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__1__sv2v_reg ;
  assign \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__0_  = \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__0__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__15_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__15__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__14_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__14__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__13_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__13__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__12_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__12__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__11_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__11__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__10_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__10__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__9_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__9__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__8_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__8__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__7_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__7__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__6_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__6__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__5_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__5__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__4_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__4__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__3_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__3__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__2_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__2__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__1_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__1__sv2v_reg ;
  assign \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__0_  = \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__0__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__15_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__15__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__14_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__14__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__13_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__13__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__12_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__12__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__11_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__11__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__10_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__10__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__9_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__9__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__8_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__8__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__7_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__7__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__6_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__6__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__5_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__5__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__4_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__4__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__3_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__3__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__2_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__2__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__1_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__1__sv2v_reg ;
  assign \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__0_  = \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__0__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__15_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__15__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__14_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__14__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__13_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__13__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__12_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__12__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__11_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__11__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__10_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__10__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__9_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__9__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__8_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__8__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__7_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__7__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__6_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__6__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__5_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__5__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__4_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__4__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__3_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__3__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__2_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__2__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__1_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__1__sv2v_reg ;
  assign \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__0_  = \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__0__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__15_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__15__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__14_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__14__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__13_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__13__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__12_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__12__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__11_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__11__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__10_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__10__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__9_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__9__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__8_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__8__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__7_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__7__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__6_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__6__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__5_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__5__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__4_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__4__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__3_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__3__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__2_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__2__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__1_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__1__sv2v_reg ;
  assign \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__0_  = \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__0__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__15_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__15__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__14_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__14__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__13_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__13__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__12_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__12__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__11_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__11__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__10_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__10__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__9_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__9__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__8_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__8__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__7_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__7__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__6_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__6__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__5_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__5__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__4_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__4__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__3_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__3__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__2_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__2__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__1_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__1__sv2v_reg ;
  assign \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__0_  = \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__0__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__15_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__15__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__14_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__14__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__13_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__13__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__12_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__12__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__11_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__11__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__10_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__10__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__9_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__9__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__8_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__8__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__7_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__7__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__6_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__6__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__5_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__5__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__4_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__4__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__3_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__3__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__2_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__2__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__1_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__1__sv2v_reg ;
  assign \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__0_  = \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__0__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__15_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__15__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__14_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__14__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__13_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__13__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__12_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__12__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__11_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__11__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__10_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__10__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__9_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__9__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__8_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__8__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__7_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__7__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__6_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__6__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__5_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__5__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__4_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__4__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__3_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__3__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__2_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__2__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__1_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__1__sv2v_reg ;
  assign \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__0_  = \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__0__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__15_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__15__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__14_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__14__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__13_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__13__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__12_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__12__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__11_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__11__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__10_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__10__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__9_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__9__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__8_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__8__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__7_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__7__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__6_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__6__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__5_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__5__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__4_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__4__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__3_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__3__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__2_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__2__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__1_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__1__sv2v_reg ;
  assign \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__0_  = \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__0__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__15_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__15__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__14_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__14__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__13_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__13__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__12_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__12__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__11_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__11__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__10_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__10__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__9_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__9__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__8_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__8__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__7_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__7__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__6_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__6__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__5_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__5__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__4_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__4__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__3_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__3__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__2_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__2__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__1_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__1__sv2v_reg ;
  assign \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__0_  = \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__0__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__15_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__15__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__14_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__14__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__13_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__13__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__12_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__12__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__11_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__11__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__10_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__10__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__9_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__9__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__8_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__8__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__7_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__7__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__6_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__6__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__5_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__5__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__4_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__4__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__3_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__3__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__2_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__2__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__1_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__1__sv2v_reg ;
  assign \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__0_  = \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__0__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__15_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__15__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__14_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__14__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__13_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__13__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__12_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__12__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__11_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__11__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__10_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__10__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__9_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__9__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__8_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__8__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__7_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__7__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__6_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__6__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__5_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__5__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__4_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__4__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__3_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__3__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__2_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__2__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__1_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__1__sv2v_reg ;
  assign \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__0_  = \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__0__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__15_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__15__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__14_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__14__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__13_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__13__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__12_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__12__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__11_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__11__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__10_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__10__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__9_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__9__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__8_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__8__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__7_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__7__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__6_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__6__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__5_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__5__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__4_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__4__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__3_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__3__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__2_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__2__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__1_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__1__sv2v_reg ;
  assign \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__0_  = \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__0__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__15_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__15__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__14_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__14__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__13_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__13__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__12_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__12__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__11_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__11__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__10_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__10__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__9_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__9__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__8_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__8__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__7_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__7__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__6_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__6__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__5_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__5__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__4_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__4__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__3_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__3__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__2_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__2__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__1_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__1__sv2v_reg ;
  assign \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__0_  = \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__0__sv2v_reg ;
  assign in_data_i_15__31_ = in_data_i[511];
  assign in_data_o[511] = in_data_i_15__31_;
  assign in_data_i_15__30_ = in_data_i[510];
  assign in_data_o[510] = in_data_i_15__30_;
  assign in_data_i_15__29_ = in_data_i[509];
  assign in_data_o[509] = in_data_i_15__29_;
  assign in_data_i_15__28_ = in_data_i[508];
  assign in_data_o[508] = in_data_i_15__28_;
  assign in_data_i_15__27_ = in_data_i[507];
  assign in_data_o[507] = in_data_i_15__27_;
  assign in_data_i_15__26_ = in_data_i[506];
  assign in_data_o[506] = in_data_i_15__26_;
  assign in_data_i_15__25_ = in_data_i[505];
  assign in_data_o[505] = in_data_i_15__25_;
  assign in_data_i_15__24_ = in_data_i[504];
  assign in_data_o[504] = in_data_i_15__24_;
  assign in_data_i_15__23_ = in_data_i[503];
  assign in_data_o[503] = in_data_i_15__23_;
  assign in_data_i_15__22_ = in_data_i[502];
  assign in_data_o[502] = in_data_i_15__22_;
  assign in_data_i_15__21_ = in_data_i[501];
  assign in_data_o[501] = in_data_i_15__21_;
  assign in_data_i_15__20_ = in_data_i[500];
  assign in_data_o[500] = in_data_i_15__20_;
  assign in_data_i_15__19_ = in_data_i[499];
  assign in_data_o[499] = in_data_i_15__19_;
  assign in_data_i_15__18_ = in_data_i[498];
  assign in_data_o[498] = in_data_i_15__18_;
  assign in_data_i_15__17_ = in_data_i[497];
  assign in_data_o[497] = in_data_i_15__17_;
  assign in_data_i_15__16_ = in_data_i[496];
  assign in_data_o[496] = in_data_i_15__16_;
  assign in_data_i_15__15_ = in_data_i[495];
  assign in_data_o[495] = in_data_i_15__15_;
  assign in_data_i_15__14_ = in_data_i[494];
  assign in_data_o[494] = in_data_i_15__14_;
  assign in_data_i_15__13_ = in_data_i[493];
  assign in_data_o[493] = in_data_i_15__13_;
  assign in_data_i_15__12_ = in_data_i[492];
  assign in_data_o[492] = in_data_i_15__12_;
  assign in_data_i_15__11_ = in_data_i[491];
  assign in_data_o[491] = in_data_i_15__11_;
  assign in_data_i_15__10_ = in_data_i[490];
  assign in_data_o[490] = in_data_i_15__10_;
  assign in_data_i_15__9_ = in_data_i[489];
  assign in_data_o[489] = in_data_i_15__9_;
  assign in_data_i_15__8_ = in_data_i[488];
  assign in_data_o[488] = in_data_i_15__8_;
  assign in_data_i_15__7_ = in_data_i[487];
  assign in_data_o[487] = in_data_i_15__7_;
  assign in_data_i_15__6_ = in_data_i[486];
  assign in_data_o[486] = in_data_i_15__6_;
  assign in_data_i_15__5_ = in_data_i[485];
  assign in_data_o[485] = in_data_i_15__5_;
  assign in_data_i_15__4_ = in_data_i[484];
  assign in_data_o[484] = in_data_i_15__4_;
  assign in_data_i_15__3_ = in_data_i[483];
  assign in_data_o[483] = in_data_i_15__3_;
  assign in_data_i_15__2_ = in_data_i[482];
  assign in_data_o[482] = in_data_i_15__2_;
  assign in_data_i_15__1_ = in_data_i[481];
  assign in_data_o[481] = in_data_i_15__1_;
  assign in_data_i_15__0_ = in_data_i[480];
  assign in_data_o[480] = in_data_i_15__0_;
  assign out_me_data_i_0__31_ = out_me_data_i[31];
  assign out_me_data_o[31] = out_me_data_i_0__31_;
  assign out_me_data_i_0__30_ = out_me_data_i[30];
  assign out_me_data_o[30] = out_me_data_i_0__30_;
  assign out_me_data_i_0__29_ = out_me_data_i[29];
  assign out_me_data_o[29] = out_me_data_i_0__29_;
  assign out_me_data_i_0__28_ = out_me_data_i[28];
  assign out_me_data_o[28] = out_me_data_i_0__28_;
  assign out_me_data_i_0__27_ = out_me_data_i[27];
  assign out_me_data_o[27] = out_me_data_i_0__27_;
  assign out_me_data_i_0__26_ = out_me_data_i[26];
  assign out_me_data_o[26] = out_me_data_i_0__26_;
  assign out_me_data_i_0__25_ = out_me_data_i[25];
  assign out_me_data_o[25] = out_me_data_i_0__25_;
  assign out_me_data_i_0__24_ = out_me_data_i[24];
  assign out_me_data_o[24] = out_me_data_i_0__24_;
  assign out_me_data_i_0__23_ = out_me_data_i[23];
  assign out_me_data_o[23] = out_me_data_i_0__23_;
  assign out_me_data_i_0__22_ = out_me_data_i[22];
  assign out_me_data_o[22] = out_me_data_i_0__22_;
  assign out_me_data_i_0__21_ = out_me_data_i[21];
  assign out_me_data_o[21] = out_me_data_i_0__21_;
  assign out_me_data_i_0__20_ = out_me_data_i[20];
  assign out_me_data_o[20] = out_me_data_i_0__20_;
  assign out_me_data_i_0__19_ = out_me_data_i[19];
  assign out_me_data_o[19] = out_me_data_i_0__19_;
  assign out_me_data_i_0__18_ = out_me_data_i[18];
  assign out_me_data_o[18] = out_me_data_i_0__18_;
  assign out_me_data_i_0__17_ = out_me_data_i[17];
  assign out_me_data_o[17] = out_me_data_i_0__17_;
  assign out_me_data_i_0__16_ = out_me_data_i[16];
  assign out_me_data_o[16] = out_me_data_i_0__16_;
  assign out_me_data_i_0__15_ = out_me_data_i[15];
  assign out_me_data_o[15] = out_me_data_i_0__15_;
  assign out_me_data_i_0__14_ = out_me_data_i[14];
  assign out_me_data_o[14] = out_me_data_i_0__14_;
  assign out_me_data_i_0__13_ = out_me_data_i[13];
  assign out_me_data_o[13] = out_me_data_i_0__13_;
  assign out_me_data_i_0__12_ = out_me_data_i[12];
  assign out_me_data_o[12] = out_me_data_i_0__12_;
  assign out_me_data_i_0__11_ = out_me_data_i[11];
  assign out_me_data_o[11] = out_me_data_i_0__11_;
  assign out_me_data_i_0__10_ = out_me_data_i[10];
  assign out_me_data_o[10] = out_me_data_i_0__10_;
  assign out_me_data_i_0__9_ = out_me_data_i[9];
  assign out_me_data_o[9] = out_me_data_i_0__9_;
  assign out_me_data_i_0__8_ = out_me_data_i[8];
  assign out_me_data_o[8] = out_me_data_i_0__8_;
  assign out_me_data_i_0__7_ = out_me_data_i[7];
  assign out_me_data_o[7] = out_me_data_i_0__7_;
  assign out_me_data_i_0__6_ = out_me_data_i[6];
  assign out_me_data_o[6] = out_me_data_i_0__6_;
  assign out_me_data_i_0__5_ = out_me_data_i[5];
  assign out_me_data_o[5] = out_me_data_i_0__5_;
  assign out_me_data_i_0__4_ = out_me_data_i[4];
  assign out_me_data_o[4] = out_me_data_i_0__4_;
  assign out_me_data_i_0__3_ = out_me_data_i[3];
  assign out_me_data_o[3] = out_me_data_i_0__3_;
  assign out_me_data_i_0__2_ = out_me_data_i[2];
  assign out_me_data_o[2] = out_me_data_i_0__2_;
  assign out_me_data_i_0__1_ = out_me_data_i[1];
  assign out_me_data_o[1] = out_me_data_i_0__1_;
  assign out_me_data_i_0__0_ = out_me_data_i[0];
  assign out_me_data_o[0] = out_me_data_i_0__0_;

  bsg_scatter_gather_vec_size_lp16
  bsg
  (
    .vec_i(channel_active_i),
    .fwd_o(fwd_sel),
    .fwd_datapath_o(fwd_dpath_sel),
    .bk_o(bk_sel),
    .bk_datapath_o(bk_dpath_sel)
  );

  assign in_yumi_o[0] = (N570)? in_yumi_i[0] : 
                        (N572)? in_yumi_i[1] : 
                        (N574)? in_yumi_i[2] : 
                        (N576)? in_yumi_i[3] : 
                        (N578)? in_yumi_i[4] : 
                        (N580)? in_yumi_i[5] : 
                        (N582)? in_yumi_i[6] : 
                        (N584)? in_yumi_i[7] : 
                        (N571)? in_yumi_i[8] : 
                        (N573)? in_yumi_i[9] : 
                        (N575)? in_yumi_i[10] : 
                        (N577)? in_yumi_i[11] : 
                        (N579)? in_yumi_i[12] : 
                        (N581)? in_yumi_i[13] : 
                        (N583)? in_yumi_i[14] : 
                        (N585)? in_yumi_i[15] : 1'b0;
  assign in_data_o[31] = (N602)? in_data_i[31] : 
                         (N604)? in_data_i[63] : 
                         (N606)? in_data_i[95] : 
                         (N608)? in_data_i[127] : 
                         (N610)? in_data_i[159] : 
                         (N612)? in_data_i[191] : 
                         (N614)? in_data_i[223] : 
                         (N616)? in_data_i[255] : 
                         (N603)? in_data_i[287] : 
                         (N605)? in_data_i[319] : 
                         (N607)? in_data_i[351] : 
                         (N609)? in_data_i[383] : 
                         (N611)? in_data_i[415] : 
                         (N613)? in_data_i[447] : 
                         (N615)? in_data_i[479] : 
                         (N617)? in_data_i_15__31_ : 1'b0;
  assign in_data_o[30] = (N602)? in_data_i[30] : 
                         (N604)? in_data_i[62] : 
                         (N606)? in_data_i[94] : 
                         (N608)? in_data_i[126] : 
                         (N610)? in_data_i[158] : 
                         (N612)? in_data_i[190] : 
                         (N614)? in_data_i[222] : 
                         (N616)? in_data_i[254] : 
                         (N603)? in_data_i[286] : 
                         (N605)? in_data_i[318] : 
                         (N607)? in_data_i[350] : 
                         (N609)? in_data_i[382] : 
                         (N611)? in_data_i[414] : 
                         (N613)? in_data_i[446] : 
                         (N615)? in_data_i[478] : 
                         (N617)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[29] = (N602)? in_data_i[29] : 
                         (N604)? in_data_i[61] : 
                         (N606)? in_data_i[93] : 
                         (N608)? in_data_i[125] : 
                         (N610)? in_data_i[157] : 
                         (N612)? in_data_i[189] : 
                         (N614)? in_data_i[221] : 
                         (N616)? in_data_i[253] : 
                         (N603)? in_data_i[285] : 
                         (N605)? in_data_i[317] : 
                         (N607)? in_data_i[349] : 
                         (N609)? in_data_i[381] : 
                         (N611)? in_data_i[413] : 
                         (N613)? in_data_i[445] : 
                         (N615)? in_data_i[477] : 
                         (N617)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[28] = (N602)? in_data_i[28] : 
                         (N604)? in_data_i[60] : 
                         (N606)? in_data_i[92] : 
                         (N608)? in_data_i[124] : 
                         (N610)? in_data_i[156] : 
                         (N612)? in_data_i[188] : 
                         (N614)? in_data_i[220] : 
                         (N616)? in_data_i[252] : 
                         (N603)? in_data_i[284] : 
                         (N605)? in_data_i[316] : 
                         (N607)? in_data_i[348] : 
                         (N609)? in_data_i[380] : 
                         (N611)? in_data_i[412] : 
                         (N613)? in_data_i[444] : 
                         (N615)? in_data_i[476] : 
                         (N617)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[27] = (N602)? in_data_i[27] : 
                         (N604)? in_data_i[59] : 
                         (N606)? in_data_i[91] : 
                         (N608)? in_data_i[123] : 
                         (N610)? in_data_i[155] : 
                         (N612)? in_data_i[187] : 
                         (N614)? in_data_i[219] : 
                         (N616)? in_data_i[251] : 
                         (N603)? in_data_i[283] : 
                         (N605)? in_data_i[315] : 
                         (N607)? in_data_i[347] : 
                         (N609)? in_data_i[379] : 
                         (N611)? in_data_i[411] : 
                         (N613)? in_data_i[443] : 
                         (N615)? in_data_i[475] : 
                         (N617)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[26] = (N602)? in_data_i[26] : 
                         (N604)? in_data_i[58] : 
                         (N606)? in_data_i[90] : 
                         (N608)? in_data_i[122] : 
                         (N610)? in_data_i[154] : 
                         (N612)? in_data_i[186] : 
                         (N614)? in_data_i[218] : 
                         (N616)? in_data_i[250] : 
                         (N603)? in_data_i[282] : 
                         (N605)? in_data_i[314] : 
                         (N607)? in_data_i[346] : 
                         (N609)? in_data_i[378] : 
                         (N611)? in_data_i[410] : 
                         (N613)? in_data_i[442] : 
                         (N615)? in_data_i[474] : 
                         (N617)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[25] = (N602)? in_data_i[25] : 
                         (N604)? in_data_i[57] : 
                         (N606)? in_data_i[89] : 
                         (N608)? in_data_i[121] : 
                         (N610)? in_data_i[153] : 
                         (N612)? in_data_i[185] : 
                         (N614)? in_data_i[217] : 
                         (N616)? in_data_i[249] : 
                         (N603)? in_data_i[281] : 
                         (N605)? in_data_i[313] : 
                         (N607)? in_data_i[345] : 
                         (N609)? in_data_i[377] : 
                         (N611)? in_data_i[409] : 
                         (N613)? in_data_i[441] : 
                         (N615)? in_data_i[473] : 
                         (N617)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[24] = (N602)? in_data_i[24] : 
                         (N604)? in_data_i[56] : 
                         (N606)? in_data_i[88] : 
                         (N608)? in_data_i[120] : 
                         (N610)? in_data_i[152] : 
                         (N612)? in_data_i[184] : 
                         (N614)? in_data_i[216] : 
                         (N616)? in_data_i[248] : 
                         (N603)? in_data_i[280] : 
                         (N605)? in_data_i[312] : 
                         (N607)? in_data_i[344] : 
                         (N609)? in_data_i[376] : 
                         (N611)? in_data_i[408] : 
                         (N613)? in_data_i[440] : 
                         (N615)? in_data_i[472] : 
                         (N617)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[23] = (N602)? in_data_i[23] : 
                         (N604)? in_data_i[55] : 
                         (N606)? in_data_i[87] : 
                         (N608)? in_data_i[119] : 
                         (N610)? in_data_i[151] : 
                         (N612)? in_data_i[183] : 
                         (N614)? in_data_i[215] : 
                         (N616)? in_data_i[247] : 
                         (N603)? in_data_i[279] : 
                         (N605)? in_data_i[311] : 
                         (N607)? in_data_i[343] : 
                         (N609)? in_data_i[375] : 
                         (N611)? in_data_i[407] : 
                         (N613)? in_data_i[439] : 
                         (N615)? in_data_i[471] : 
                         (N617)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[22] = (N602)? in_data_i[22] : 
                         (N604)? in_data_i[54] : 
                         (N606)? in_data_i[86] : 
                         (N608)? in_data_i[118] : 
                         (N610)? in_data_i[150] : 
                         (N612)? in_data_i[182] : 
                         (N614)? in_data_i[214] : 
                         (N616)? in_data_i[246] : 
                         (N603)? in_data_i[278] : 
                         (N605)? in_data_i[310] : 
                         (N607)? in_data_i[342] : 
                         (N609)? in_data_i[374] : 
                         (N611)? in_data_i[406] : 
                         (N613)? in_data_i[438] : 
                         (N615)? in_data_i[470] : 
                         (N617)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[21] = (N602)? in_data_i[21] : 
                         (N604)? in_data_i[53] : 
                         (N606)? in_data_i[85] : 
                         (N608)? in_data_i[117] : 
                         (N610)? in_data_i[149] : 
                         (N612)? in_data_i[181] : 
                         (N614)? in_data_i[213] : 
                         (N616)? in_data_i[245] : 
                         (N603)? in_data_i[277] : 
                         (N605)? in_data_i[309] : 
                         (N607)? in_data_i[341] : 
                         (N609)? in_data_i[373] : 
                         (N611)? in_data_i[405] : 
                         (N613)? in_data_i[437] : 
                         (N615)? in_data_i[469] : 
                         (N617)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[20] = (N602)? in_data_i[20] : 
                         (N604)? in_data_i[52] : 
                         (N606)? in_data_i[84] : 
                         (N608)? in_data_i[116] : 
                         (N610)? in_data_i[148] : 
                         (N612)? in_data_i[180] : 
                         (N614)? in_data_i[212] : 
                         (N616)? in_data_i[244] : 
                         (N603)? in_data_i[276] : 
                         (N605)? in_data_i[308] : 
                         (N607)? in_data_i[340] : 
                         (N609)? in_data_i[372] : 
                         (N611)? in_data_i[404] : 
                         (N613)? in_data_i[436] : 
                         (N615)? in_data_i[468] : 
                         (N617)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[19] = (N602)? in_data_i[19] : 
                         (N604)? in_data_i[51] : 
                         (N606)? in_data_i[83] : 
                         (N608)? in_data_i[115] : 
                         (N610)? in_data_i[147] : 
                         (N612)? in_data_i[179] : 
                         (N614)? in_data_i[211] : 
                         (N616)? in_data_i[243] : 
                         (N603)? in_data_i[275] : 
                         (N605)? in_data_i[307] : 
                         (N607)? in_data_i[339] : 
                         (N609)? in_data_i[371] : 
                         (N611)? in_data_i[403] : 
                         (N613)? in_data_i[435] : 
                         (N615)? in_data_i[467] : 
                         (N617)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[18] = (N602)? in_data_i[18] : 
                         (N604)? in_data_i[50] : 
                         (N606)? in_data_i[82] : 
                         (N608)? in_data_i[114] : 
                         (N610)? in_data_i[146] : 
                         (N612)? in_data_i[178] : 
                         (N614)? in_data_i[210] : 
                         (N616)? in_data_i[242] : 
                         (N603)? in_data_i[274] : 
                         (N605)? in_data_i[306] : 
                         (N607)? in_data_i[338] : 
                         (N609)? in_data_i[370] : 
                         (N611)? in_data_i[402] : 
                         (N613)? in_data_i[434] : 
                         (N615)? in_data_i[466] : 
                         (N617)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[17] = (N602)? in_data_i[17] : 
                         (N604)? in_data_i[49] : 
                         (N606)? in_data_i[81] : 
                         (N608)? in_data_i[113] : 
                         (N610)? in_data_i[145] : 
                         (N612)? in_data_i[177] : 
                         (N614)? in_data_i[209] : 
                         (N616)? in_data_i[241] : 
                         (N603)? in_data_i[273] : 
                         (N605)? in_data_i[305] : 
                         (N607)? in_data_i[337] : 
                         (N609)? in_data_i[369] : 
                         (N611)? in_data_i[401] : 
                         (N613)? in_data_i[433] : 
                         (N615)? in_data_i[465] : 
                         (N617)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[16] = (N602)? in_data_i[16] : 
                         (N604)? in_data_i[48] : 
                         (N606)? in_data_i[80] : 
                         (N608)? in_data_i[112] : 
                         (N610)? in_data_i[144] : 
                         (N612)? in_data_i[176] : 
                         (N614)? in_data_i[208] : 
                         (N616)? in_data_i[240] : 
                         (N603)? in_data_i[272] : 
                         (N605)? in_data_i[304] : 
                         (N607)? in_data_i[336] : 
                         (N609)? in_data_i[368] : 
                         (N611)? in_data_i[400] : 
                         (N613)? in_data_i[432] : 
                         (N615)? in_data_i[464] : 
                         (N617)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[15] = (N602)? in_data_i[15] : 
                         (N604)? in_data_i[47] : 
                         (N606)? in_data_i[79] : 
                         (N608)? in_data_i[111] : 
                         (N610)? in_data_i[143] : 
                         (N612)? in_data_i[175] : 
                         (N614)? in_data_i[207] : 
                         (N616)? in_data_i[239] : 
                         (N603)? in_data_i[271] : 
                         (N605)? in_data_i[303] : 
                         (N607)? in_data_i[335] : 
                         (N609)? in_data_i[367] : 
                         (N611)? in_data_i[399] : 
                         (N613)? in_data_i[431] : 
                         (N615)? in_data_i[463] : 
                         (N617)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[14] = (N602)? in_data_i[14] : 
                         (N604)? in_data_i[46] : 
                         (N606)? in_data_i[78] : 
                         (N608)? in_data_i[110] : 
                         (N610)? in_data_i[142] : 
                         (N612)? in_data_i[174] : 
                         (N614)? in_data_i[206] : 
                         (N616)? in_data_i[238] : 
                         (N603)? in_data_i[270] : 
                         (N605)? in_data_i[302] : 
                         (N607)? in_data_i[334] : 
                         (N609)? in_data_i[366] : 
                         (N611)? in_data_i[398] : 
                         (N613)? in_data_i[430] : 
                         (N615)? in_data_i[462] : 
                         (N617)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[13] = (N602)? in_data_i[13] : 
                         (N604)? in_data_i[45] : 
                         (N606)? in_data_i[77] : 
                         (N608)? in_data_i[109] : 
                         (N610)? in_data_i[141] : 
                         (N612)? in_data_i[173] : 
                         (N614)? in_data_i[205] : 
                         (N616)? in_data_i[237] : 
                         (N603)? in_data_i[269] : 
                         (N605)? in_data_i[301] : 
                         (N607)? in_data_i[333] : 
                         (N609)? in_data_i[365] : 
                         (N611)? in_data_i[397] : 
                         (N613)? in_data_i[429] : 
                         (N615)? in_data_i[461] : 
                         (N617)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[12] = (N602)? in_data_i[12] : 
                         (N604)? in_data_i[44] : 
                         (N606)? in_data_i[76] : 
                         (N608)? in_data_i[108] : 
                         (N610)? in_data_i[140] : 
                         (N612)? in_data_i[172] : 
                         (N614)? in_data_i[204] : 
                         (N616)? in_data_i[236] : 
                         (N603)? in_data_i[268] : 
                         (N605)? in_data_i[300] : 
                         (N607)? in_data_i[332] : 
                         (N609)? in_data_i[364] : 
                         (N611)? in_data_i[396] : 
                         (N613)? in_data_i[428] : 
                         (N615)? in_data_i[460] : 
                         (N617)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[11] = (N602)? in_data_i[11] : 
                         (N604)? in_data_i[43] : 
                         (N606)? in_data_i[75] : 
                         (N608)? in_data_i[107] : 
                         (N610)? in_data_i[139] : 
                         (N612)? in_data_i[171] : 
                         (N614)? in_data_i[203] : 
                         (N616)? in_data_i[235] : 
                         (N603)? in_data_i[267] : 
                         (N605)? in_data_i[299] : 
                         (N607)? in_data_i[331] : 
                         (N609)? in_data_i[363] : 
                         (N611)? in_data_i[395] : 
                         (N613)? in_data_i[427] : 
                         (N615)? in_data_i[459] : 
                         (N617)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[10] = (N602)? in_data_i[10] : 
                         (N604)? in_data_i[42] : 
                         (N606)? in_data_i[74] : 
                         (N608)? in_data_i[106] : 
                         (N610)? in_data_i[138] : 
                         (N612)? in_data_i[170] : 
                         (N614)? in_data_i[202] : 
                         (N616)? in_data_i[234] : 
                         (N603)? in_data_i[266] : 
                         (N605)? in_data_i[298] : 
                         (N607)? in_data_i[330] : 
                         (N609)? in_data_i[362] : 
                         (N611)? in_data_i[394] : 
                         (N613)? in_data_i[426] : 
                         (N615)? in_data_i[458] : 
                         (N617)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[9] = (N602)? in_data_i[9] : 
                        (N604)? in_data_i[41] : 
                        (N606)? in_data_i[73] : 
                        (N608)? in_data_i[105] : 
                        (N610)? in_data_i[137] : 
                        (N612)? in_data_i[169] : 
                        (N614)? in_data_i[201] : 
                        (N616)? in_data_i[233] : 
                        (N603)? in_data_i[265] : 
                        (N605)? in_data_i[297] : 
                        (N607)? in_data_i[329] : 
                        (N609)? in_data_i[361] : 
                        (N611)? in_data_i[393] : 
                        (N613)? in_data_i[425] : 
                        (N615)? in_data_i[457] : 
                        (N617)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[8] = (N602)? in_data_i[8] : 
                        (N604)? in_data_i[40] : 
                        (N606)? in_data_i[72] : 
                        (N608)? in_data_i[104] : 
                        (N610)? in_data_i[136] : 
                        (N612)? in_data_i[168] : 
                        (N614)? in_data_i[200] : 
                        (N616)? in_data_i[232] : 
                        (N603)? in_data_i[264] : 
                        (N605)? in_data_i[296] : 
                        (N607)? in_data_i[328] : 
                        (N609)? in_data_i[360] : 
                        (N611)? in_data_i[392] : 
                        (N613)? in_data_i[424] : 
                        (N615)? in_data_i[456] : 
                        (N617)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[7] = (N602)? in_data_i[7] : 
                        (N604)? in_data_i[39] : 
                        (N606)? in_data_i[71] : 
                        (N608)? in_data_i[103] : 
                        (N610)? in_data_i[135] : 
                        (N612)? in_data_i[167] : 
                        (N614)? in_data_i[199] : 
                        (N616)? in_data_i[231] : 
                        (N603)? in_data_i[263] : 
                        (N605)? in_data_i[295] : 
                        (N607)? in_data_i[327] : 
                        (N609)? in_data_i[359] : 
                        (N611)? in_data_i[391] : 
                        (N613)? in_data_i[423] : 
                        (N615)? in_data_i[455] : 
                        (N617)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[6] = (N602)? in_data_i[6] : 
                        (N604)? in_data_i[38] : 
                        (N606)? in_data_i[70] : 
                        (N608)? in_data_i[102] : 
                        (N610)? in_data_i[134] : 
                        (N612)? in_data_i[166] : 
                        (N614)? in_data_i[198] : 
                        (N616)? in_data_i[230] : 
                        (N603)? in_data_i[262] : 
                        (N605)? in_data_i[294] : 
                        (N607)? in_data_i[326] : 
                        (N609)? in_data_i[358] : 
                        (N611)? in_data_i[390] : 
                        (N613)? in_data_i[422] : 
                        (N615)? in_data_i[454] : 
                        (N617)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[5] = (N602)? in_data_i[5] : 
                        (N604)? in_data_i[37] : 
                        (N606)? in_data_i[69] : 
                        (N608)? in_data_i[101] : 
                        (N610)? in_data_i[133] : 
                        (N612)? in_data_i[165] : 
                        (N614)? in_data_i[197] : 
                        (N616)? in_data_i[229] : 
                        (N603)? in_data_i[261] : 
                        (N605)? in_data_i[293] : 
                        (N607)? in_data_i[325] : 
                        (N609)? in_data_i[357] : 
                        (N611)? in_data_i[389] : 
                        (N613)? in_data_i[421] : 
                        (N615)? in_data_i[453] : 
                        (N617)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[4] = (N602)? in_data_i[4] : 
                        (N604)? in_data_i[36] : 
                        (N606)? in_data_i[68] : 
                        (N608)? in_data_i[100] : 
                        (N610)? in_data_i[132] : 
                        (N612)? in_data_i[164] : 
                        (N614)? in_data_i[196] : 
                        (N616)? in_data_i[228] : 
                        (N603)? in_data_i[260] : 
                        (N605)? in_data_i[292] : 
                        (N607)? in_data_i[324] : 
                        (N609)? in_data_i[356] : 
                        (N611)? in_data_i[388] : 
                        (N613)? in_data_i[420] : 
                        (N615)? in_data_i[452] : 
                        (N617)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[3] = (N602)? in_data_i[3] : 
                        (N604)? in_data_i[35] : 
                        (N606)? in_data_i[67] : 
                        (N608)? in_data_i[99] : 
                        (N610)? in_data_i[131] : 
                        (N612)? in_data_i[163] : 
                        (N614)? in_data_i[195] : 
                        (N616)? in_data_i[227] : 
                        (N603)? in_data_i[259] : 
                        (N605)? in_data_i[291] : 
                        (N607)? in_data_i[323] : 
                        (N609)? in_data_i[355] : 
                        (N611)? in_data_i[387] : 
                        (N613)? in_data_i[419] : 
                        (N615)? in_data_i[451] : 
                        (N617)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[2] = (N602)? in_data_i[2] : 
                        (N604)? in_data_i[34] : 
                        (N606)? in_data_i[66] : 
                        (N608)? in_data_i[98] : 
                        (N610)? in_data_i[130] : 
                        (N612)? in_data_i[162] : 
                        (N614)? in_data_i[194] : 
                        (N616)? in_data_i[226] : 
                        (N603)? in_data_i[258] : 
                        (N605)? in_data_i[290] : 
                        (N607)? in_data_i[322] : 
                        (N609)? in_data_i[354] : 
                        (N611)? in_data_i[386] : 
                        (N613)? in_data_i[418] : 
                        (N615)? in_data_i[450] : 
                        (N617)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[1] = (N602)? in_data_i[1] : 
                        (N604)? in_data_i[33] : 
                        (N606)? in_data_i[65] : 
                        (N608)? in_data_i[97] : 
                        (N610)? in_data_i[129] : 
                        (N612)? in_data_i[161] : 
                        (N614)? in_data_i[193] : 
                        (N616)? in_data_i[225] : 
                        (N603)? in_data_i[257] : 
                        (N605)? in_data_i[289] : 
                        (N607)? in_data_i[321] : 
                        (N609)? in_data_i[353] : 
                        (N611)? in_data_i[385] : 
                        (N613)? in_data_i[417] : 
                        (N615)? in_data_i[449] : 
                        (N617)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[0] = (N602)? in_data_i[0] : 
                        (N604)? in_data_i[32] : 
                        (N606)? in_data_i[64] : 
                        (N608)? in_data_i[96] : 
                        (N610)? in_data_i[128] : 
                        (N612)? in_data_i[160] : 
                        (N614)? in_data_i[192] : 
                        (N616)? in_data_i[224] : 
                        (N603)? in_data_i[256] : 
                        (N605)? in_data_i[288] : 
                        (N607)? in_data_i[320] : 
                        (N609)? in_data_i[352] : 
                        (N611)? in_data_i[384] : 
                        (N613)? in_data_i[416] : 
                        (N615)? in_data_i[448] : 
                        (N617)? in_data_i_15__0_ : 1'b0;
  assign out_me_v_o[0] = (N630)? out_me_v_i[0] : 
                         (N632)? out_me_v_i[1] : 
                         (N634)? out_me_v_i[2] : 
                         (N636)? out_me_v_i[3] : 
                         (N638)? out_me_v_i[4] : 
                         (N640)? out_me_v_i[5] : 
                         (N642)? out_me_v_i[6] : 
                         (N644)? out_me_v_i[7] : 
                         (N631)? out_me_v_i[8] : 
                         (N633)? out_me_v_i[9] : 
                         (N635)? out_me_v_i[10] : 
                         (N637)? out_me_v_i[11] : 
                         (N639)? out_me_v_i[12] : 
                         (N641)? out_me_v_i[13] : 
                         (N643)? out_me_v_i[14] : 
                         (N645)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[0] = (N662)? out_me_ready_i[0] : 
                             (N664)? out_me_ready_i[1] : 
                             (N666)? out_me_ready_i[2] : 
                             (N668)? out_me_ready_i[3] : 
                             (N670)? out_me_ready_i[4] : 
                             (N672)? out_me_ready_i[5] : 
                             (N674)? out_me_ready_i[6] : 
                             (N676)? out_me_ready_i[7] : 
                             (N663)? out_me_ready_i[8] : 
                             (N665)? out_me_ready_i[9] : 
                             (N667)? out_me_ready_i[10] : 
                             (N669)? out_me_ready_i[11] : 
                             (N671)? out_me_ready_i[12] : 
                             (N673)? out_me_ready_i[13] : 
                             (N675)? out_me_ready_i[14] : 
                             (N677)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[1] = (N710)? in_yumi_i[0] : 
                        (N712)? in_yumi_i[1] : 
                        (N714)? in_yumi_i[2] : 
                        (N716)? in_yumi_i[3] : 
                        (N718)? in_yumi_i[4] : 
                        (N720)? in_yumi_i[5] : 
                        (N722)? in_yumi_i[6] : 
                        (N724)? in_yumi_i[7] : 
                        (N711)? in_yumi_i[8] : 
                        (N713)? in_yumi_i[9] : 
                        (N715)? in_yumi_i[10] : 
                        (N717)? in_yumi_i[11] : 
                        (N719)? in_yumi_i[12] : 
                        (N721)? in_yumi_i[13] : 
                        (N723)? in_yumi_i[14] : 
                        (N725)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[1] = (N753)? out_me_v_i[0] : 
                         (N755)? out_me_v_i[1] : 
                         (N757)? out_me_v_i[2] : 
                         (N759)? out_me_v_i[3] : 
                         (N761)? out_me_v_i[4] : 
                         (N763)? out_me_v_i[5] : 
                         (N765)? out_me_v_i[6] : 
                         (N767)? out_me_v_i[7] : 
                         (N754)? out_me_v_i[8] : 
                         (N756)? out_me_v_i[9] : 
                         (N758)? out_me_v_i[10] : 
                         (N760)? out_me_v_i[11] : 
                         (N762)? out_me_v_i[12] : 
                         (N764)? out_me_v_i[13] : 
                         (N766)? out_me_v_i[14] : 
                         (N768)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[1] = (N785)? out_me_ready_i[0] : 
                             (N787)? out_me_ready_i[1] : 
                             (N789)? out_me_ready_i[2] : 
                             (N791)? out_me_ready_i[3] : 
                             (N793)? out_me_ready_i[4] : 
                             (N795)? out_me_ready_i[5] : 
                             (N797)? out_me_ready_i[6] : 
                             (N799)? out_me_ready_i[7] : 
                             (N786)? out_me_ready_i[8] : 
                             (N788)? out_me_ready_i[9] : 
                             (N790)? out_me_ready_i[10] : 
                             (N792)? out_me_ready_i[11] : 
                             (N794)? out_me_ready_i[12] : 
                             (N796)? out_me_ready_i[13] : 
                             (N798)? out_me_ready_i[14] : 
                             (N800)? out_me_ready_i[15] : 1'b0;
  assign out_me_data_o[63] = (N801)? out_me_data_i_0__31_ : 
                             (N0)? out_me_data_i[63] : 1'b0;
  assign N0 = bk_dpath_sel_r_4;
  assign out_me_data_o[62] = (N801)? out_me_data_i_0__30_ : 
                             (N0)? out_me_data_i[62] : 1'b0;
  assign out_me_data_o[61] = (N801)? out_me_data_i_0__29_ : 
                             (N0)? out_me_data_i[61] : 1'b0;
  assign out_me_data_o[60] = (N801)? out_me_data_i_0__28_ : 
                             (N0)? out_me_data_i[60] : 1'b0;
  assign out_me_data_o[59] = (N801)? out_me_data_i_0__27_ : 
                             (N0)? out_me_data_i[59] : 1'b0;
  assign out_me_data_o[58] = (N801)? out_me_data_i_0__26_ : 
                             (N0)? out_me_data_i[58] : 1'b0;
  assign out_me_data_o[57] = (N801)? out_me_data_i_0__25_ : 
                             (N0)? out_me_data_i[57] : 1'b0;
  assign out_me_data_o[56] = (N801)? out_me_data_i_0__24_ : 
                             (N0)? out_me_data_i[56] : 1'b0;
  assign out_me_data_o[55] = (N801)? out_me_data_i_0__23_ : 
                             (N0)? out_me_data_i[55] : 1'b0;
  assign out_me_data_o[54] = (N801)? out_me_data_i_0__22_ : 
                             (N0)? out_me_data_i[54] : 1'b0;
  assign out_me_data_o[53] = (N801)? out_me_data_i_0__21_ : 
                             (N0)? out_me_data_i[53] : 1'b0;
  assign out_me_data_o[52] = (N801)? out_me_data_i_0__20_ : 
                             (N0)? out_me_data_i[52] : 1'b0;
  assign out_me_data_o[51] = (N801)? out_me_data_i_0__19_ : 
                             (N0)? out_me_data_i[51] : 1'b0;
  assign out_me_data_o[50] = (N801)? out_me_data_i_0__18_ : 
                             (N0)? out_me_data_i[50] : 1'b0;
  assign out_me_data_o[49] = (N801)? out_me_data_i_0__17_ : 
                             (N0)? out_me_data_i[49] : 1'b0;
  assign out_me_data_o[48] = (N801)? out_me_data_i_0__16_ : 
                             (N0)? out_me_data_i[48] : 1'b0;
  assign out_me_data_o[47] = (N801)? out_me_data_i_0__15_ : 
                             (N0)? out_me_data_i[47] : 1'b0;
  assign out_me_data_o[46] = (N801)? out_me_data_i_0__14_ : 
                             (N0)? out_me_data_i[46] : 1'b0;
  assign out_me_data_o[45] = (N801)? out_me_data_i_0__13_ : 
                             (N0)? out_me_data_i[45] : 1'b0;
  assign out_me_data_o[44] = (N801)? out_me_data_i_0__12_ : 
                             (N0)? out_me_data_i[44] : 1'b0;
  assign out_me_data_o[43] = (N801)? out_me_data_i_0__11_ : 
                             (N0)? out_me_data_i[43] : 1'b0;
  assign out_me_data_o[42] = (N801)? out_me_data_i_0__10_ : 
                             (N0)? out_me_data_i[42] : 1'b0;
  assign out_me_data_o[41] = (N801)? out_me_data_i_0__9_ : 
                             (N0)? out_me_data_i[41] : 1'b0;
  assign out_me_data_o[40] = (N801)? out_me_data_i_0__8_ : 
                             (N0)? out_me_data_i[40] : 1'b0;
  assign out_me_data_o[39] = (N801)? out_me_data_i_0__7_ : 
                             (N0)? out_me_data_i[39] : 1'b0;
  assign out_me_data_o[38] = (N801)? out_me_data_i_0__6_ : 
                             (N0)? out_me_data_i[38] : 1'b0;
  assign out_me_data_o[37] = (N801)? out_me_data_i_0__5_ : 
                             (N0)? out_me_data_i[37] : 1'b0;
  assign out_me_data_o[36] = (N801)? out_me_data_i_0__4_ : 
                             (N0)? out_me_data_i[36] : 1'b0;
  assign out_me_data_o[35] = (N801)? out_me_data_i_0__3_ : 
                             (N0)? out_me_data_i[35] : 1'b0;
  assign out_me_data_o[34] = (N801)? out_me_data_i_0__2_ : 
                             (N0)? out_me_data_i[34] : 1'b0;
  assign out_me_data_o[33] = (N801)? out_me_data_i_0__1_ : 
                             (N0)? out_me_data_i[33] : 1'b0;
  assign out_me_data_o[32] = (N801)? out_me_data_i_0__0_ : 
                             (N0)? out_me_data_i[32] : 1'b0;
  assign in_yumi_o[2] = (N834)? in_yumi_i[0] : 
                        (N836)? in_yumi_i[1] : 
                        (N838)? in_yumi_i[2] : 
                        (N840)? in_yumi_i[3] : 
                        (N842)? in_yumi_i[4] : 
                        (N844)? in_yumi_i[5] : 
                        (N846)? in_yumi_i[6] : 
                        (N848)? in_yumi_i[7] : 
                        (N835)? in_yumi_i[8] : 
                        (N837)? in_yumi_i[9] : 
                        (N839)? in_yumi_i[10] : 
                        (N841)? in_yumi_i[11] : 
                        (N843)? in_yumi_i[12] : 
                        (N845)? in_yumi_i[13] : 
                        (N847)? in_yumi_i[14] : 
                        (N849)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[2] = (N876)? out_me_v_i[0] : 
                         (N878)? out_me_v_i[1] : 
                         (N880)? out_me_v_i[2] : 
                         (N882)? out_me_v_i[3] : 
                         (N884)? out_me_v_i[4] : 
                         (N886)? out_me_v_i[5] : 
                         (N888)? out_me_v_i[6] : 
                         (N890)? out_me_v_i[7] : 
                         (N877)? out_me_v_i[8] : 
                         (N879)? out_me_v_i[9] : 
                         (N881)? out_me_v_i[10] : 
                         (N883)? out_me_v_i[11] : 
                         (N885)? out_me_v_i[12] : 
                         (N887)? out_me_v_i[13] : 
                         (N889)? out_me_v_i[14] : 
                         (N891)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[2] = (N908)? out_me_ready_i[0] : 
                             (N910)? out_me_ready_i[1] : 
                             (N912)? out_me_ready_i[2] : 
                             (N914)? out_me_ready_i[3] : 
                             (N916)? out_me_ready_i[4] : 
                             (N918)? out_me_ready_i[5] : 
                             (N920)? out_me_ready_i[6] : 
                             (N922)? out_me_ready_i[7] : 
                             (N909)? out_me_ready_i[8] : 
                             (N911)? out_me_ready_i[9] : 
                             (N913)? out_me_ready_i[10] : 
                             (N915)? out_me_ready_i[11] : 
                             (N917)? out_me_ready_i[12] : 
                             (N919)? out_me_ready_i[13] : 
                             (N921)? out_me_ready_i[14] : 
                             (N923)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[3] = (N957)? in_yumi_i[0] : 
                        (N959)? in_yumi_i[1] : 
                        (N961)? in_yumi_i[2] : 
                        (N963)? in_yumi_i[3] : 
                        (N965)? in_yumi_i[4] : 
                        (N967)? in_yumi_i[5] : 
                        (N969)? in_yumi_i[6] : 
                        (N971)? in_yumi_i[7] : 
                        (N958)? in_yumi_i[8] : 
                        (N960)? in_yumi_i[9] : 
                        (N962)? in_yumi_i[10] : 
                        (N964)? in_yumi_i[11] : 
                        (N966)? in_yumi_i[12] : 
                        (N968)? in_yumi_i[13] : 
                        (N970)? in_yumi_i[14] : 
                        (N972)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[3] = (N998)? out_me_v_i[0] : 
                         (N1000)? out_me_v_i[1] : 
                         (N1002)? out_me_v_i[2] : 
                         (N1004)? out_me_v_i[3] : 
                         (N1006)? out_me_v_i[4] : 
                         (N1008)? out_me_v_i[5] : 
                         (N1010)? out_me_v_i[6] : 
                         (N1012)? out_me_v_i[7] : 
                         (N999)? out_me_v_i[8] : 
                         (N1001)? out_me_v_i[9] : 
                         (N1003)? out_me_v_i[10] : 
                         (N1005)? out_me_v_i[11] : 
                         (N1007)? out_me_v_i[12] : 
                         (N1009)? out_me_v_i[13] : 
                         (N1011)? out_me_v_i[14] : 
                         (N1013)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[3] = (N1030)? out_me_ready_i[0] : 
                             (N1032)? out_me_ready_i[1] : 
                             (N1034)? out_me_ready_i[2] : 
                             (N1036)? out_me_ready_i[3] : 
                             (N1038)? out_me_ready_i[4] : 
                             (N1040)? out_me_ready_i[5] : 
                             (N1042)? out_me_ready_i[6] : 
                             (N1044)? out_me_ready_i[7] : 
                             (N1031)? out_me_ready_i[8] : 
                             (N1033)? out_me_ready_i[9] : 
                             (N1035)? out_me_ready_i[10] : 
                             (N1037)? out_me_ready_i[11] : 
                             (N1039)? out_me_ready_i[12] : 
                             (N1041)? out_me_ready_i[13] : 
                             (N1043)? out_me_ready_i[14] : 
                             (N1045)? out_me_ready_i[15] : 1'b0;
  assign out_me_data_o[127] = (N1048)? out_me_data_i_0__31_ : 
                              (N1050)? out_me_data_i[63] : 
                              (N1049)? out_me_data_i[95] : 
                              (N1051)? out_me_data_i[127] : 1'b0;
  assign out_me_data_o[126] = (N1048)? out_me_data_i_0__30_ : 
                              (N1050)? out_me_data_i[62] : 
                              (N1049)? out_me_data_i[94] : 
                              (N1051)? out_me_data_i[126] : 1'b0;
  assign out_me_data_o[125] = (N1048)? out_me_data_i_0__29_ : 
                              (N1050)? out_me_data_i[61] : 
                              (N1049)? out_me_data_i[93] : 
                              (N1051)? out_me_data_i[125] : 1'b0;
  assign out_me_data_o[124] = (N1048)? out_me_data_i_0__28_ : 
                              (N1050)? out_me_data_i[60] : 
                              (N1049)? out_me_data_i[92] : 
                              (N1051)? out_me_data_i[124] : 1'b0;
  assign out_me_data_o[123] = (N1048)? out_me_data_i_0__27_ : 
                              (N1050)? out_me_data_i[59] : 
                              (N1049)? out_me_data_i[91] : 
                              (N1051)? out_me_data_i[123] : 1'b0;
  assign out_me_data_o[122] = (N1048)? out_me_data_i_0__26_ : 
                              (N1050)? out_me_data_i[58] : 
                              (N1049)? out_me_data_i[90] : 
                              (N1051)? out_me_data_i[122] : 1'b0;
  assign out_me_data_o[121] = (N1048)? out_me_data_i_0__25_ : 
                              (N1050)? out_me_data_i[57] : 
                              (N1049)? out_me_data_i[89] : 
                              (N1051)? out_me_data_i[121] : 1'b0;
  assign out_me_data_o[120] = (N1048)? out_me_data_i_0__24_ : 
                              (N1050)? out_me_data_i[56] : 
                              (N1049)? out_me_data_i[88] : 
                              (N1051)? out_me_data_i[120] : 1'b0;
  assign out_me_data_o[119] = (N1048)? out_me_data_i_0__23_ : 
                              (N1050)? out_me_data_i[55] : 
                              (N1049)? out_me_data_i[87] : 
                              (N1051)? out_me_data_i[119] : 1'b0;
  assign out_me_data_o[118] = (N1048)? out_me_data_i_0__22_ : 
                              (N1050)? out_me_data_i[54] : 
                              (N1049)? out_me_data_i[86] : 
                              (N1051)? out_me_data_i[118] : 1'b0;
  assign out_me_data_o[117] = (N1048)? out_me_data_i_0__21_ : 
                              (N1050)? out_me_data_i[53] : 
                              (N1049)? out_me_data_i[85] : 
                              (N1051)? out_me_data_i[117] : 1'b0;
  assign out_me_data_o[116] = (N1048)? out_me_data_i_0__20_ : 
                              (N1050)? out_me_data_i[52] : 
                              (N1049)? out_me_data_i[84] : 
                              (N1051)? out_me_data_i[116] : 1'b0;
  assign out_me_data_o[115] = (N1048)? out_me_data_i_0__19_ : 
                              (N1050)? out_me_data_i[51] : 
                              (N1049)? out_me_data_i[83] : 
                              (N1051)? out_me_data_i[115] : 1'b0;
  assign out_me_data_o[114] = (N1048)? out_me_data_i_0__18_ : 
                              (N1050)? out_me_data_i[50] : 
                              (N1049)? out_me_data_i[82] : 
                              (N1051)? out_me_data_i[114] : 1'b0;
  assign out_me_data_o[113] = (N1048)? out_me_data_i_0__17_ : 
                              (N1050)? out_me_data_i[49] : 
                              (N1049)? out_me_data_i[81] : 
                              (N1051)? out_me_data_i[113] : 1'b0;
  assign out_me_data_o[112] = (N1048)? out_me_data_i_0__16_ : 
                              (N1050)? out_me_data_i[48] : 
                              (N1049)? out_me_data_i[80] : 
                              (N1051)? out_me_data_i[112] : 1'b0;
  assign out_me_data_o[111] = (N1048)? out_me_data_i_0__15_ : 
                              (N1050)? out_me_data_i[47] : 
                              (N1049)? out_me_data_i[79] : 
                              (N1051)? out_me_data_i[111] : 1'b0;
  assign out_me_data_o[110] = (N1048)? out_me_data_i_0__14_ : 
                              (N1050)? out_me_data_i[46] : 
                              (N1049)? out_me_data_i[78] : 
                              (N1051)? out_me_data_i[110] : 1'b0;
  assign out_me_data_o[109] = (N1048)? out_me_data_i_0__13_ : 
                              (N1050)? out_me_data_i[45] : 
                              (N1049)? out_me_data_i[77] : 
                              (N1051)? out_me_data_i[109] : 1'b0;
  assign out_me_data_o[108] = (N1048)? out_me_data_i_0__12_ : 
                              (N1050)? out_me_data_i[44] : 
                              (N1049)? out_me_data_i[76] : 
                              (N1051)? out_me_data_i[108] : 1'b0;
  assign out_me_data_o[107] = (N1048)? out_me_data_i_0__11_ : 
                              (N1050)? out_me_data_i[43] : 
                              (N1049)? out_me_data_i[75] : 
                              (N1051)? out_me_data_i[107] : 1'b0;
  assign out_me_data_o[106] = (N1048)? out_me_data_i_0__10_ : 
                              (N1050)? out_me_data_i[42] : 
                              (N1049)? out_me_data_i[74] : 
                              (N1051)? out_me_data_i[106] : 1'b0;
  assign out_me_data_o[105] = (N1048)? out_me_data_i_0__9_ : 
                              (N1050)? out_me_data_i[41] : 
                              (N1049)? out_me_data_i[73] : 
                              (N1051)? out_me_data_i[105] : 1'b0;
  assign out_me_data_o[104] = (N1048)? out_me_data_i_0__8_ : 
                              (N1050)? out_me_data_i[40] : 
                              (N1049)? out_me_data_i[72] : 
                              (N1051)? out_me_data_i[104] : 1'b0;
  assign out_me_data_o[103] = (N1048)? out_me_data_i_0__7_ : 
                              (N1050)? out_me_data_i[39] : 
                              (N1049)? out_me_data_i[71] : 
                              (N1051)? out_me_data_i[103] : 1'b0;
  assign out_me_data_o[102] = (N1048)? out_me_data_i_0__6_ : 
                              (N1050)? out_me_data_i[38] : 
                              (N1049)? out_me_data_i[70] : 
                              (N1051)? out_me_data_i[102] : 1'b0;
  assign out_me_data_o[101] = (N1048)? out_me_data_i_0__5_ : 
                              (N1050)? out_me_data_i[37] : 
                              (N1049)? out_me_data_i[69] : 
                              (N1051)? out_me_data_i[101] : 1'b0;
  assign out_me_data_o[100] = (N1048)? out_me_data_i_0__4_ : 
                              (N1050)? out_me_data_i[36] : 
                              (N1049)? out_me_data_i[68] : 
                              (N1051)? out_me_data_i[100] : 1'b0;
  assign out_me_data_o[99] = (N1048)? out_me_data_i_0__3_ : 
                             (N1050)? out_me_data_i[35] : 
                             (N1049)? out_me_data_i[67] : 
                             (N1051)? out_me_data_i[99] : 1'b0;
  assign out_me_data_o[98] = (N1048)? out_me_data_i_0__2_ : 
                             (N1050)? out_me_data_i[34] : 
                             (N1049)? out_me_data_i[66] : 
                             (N1051)? out_me_data_i[98] : 1'b0;
  assign out_me_data_o[97] = (N1048)? out_me_data_i_0__1_ : 
                             (N1050)? out_me_data_i[33] : 
                             (N1049)? out_me_data_i[65] : 
                             (N1051)? out_me_data_i[97] : 1'b0;
  assign out_me_data_o[96] = (N1048)? out_me_data_i_0__0_ : 
                             (N1050)? out_me_data_i[32] : 
                             (N1049)? out_me_data_i[64] : 
                             (N1051)? out_me_data_i[96] : 1'b0;
  assign in_yumi_o[4] = (N1084)? in_yumi_i[0] : 
                        (N1086)? in_yumi_i[1] : 
                        (N1088)? in_yumi_i[2] : 
                        (N1090)? in_yumi_i[3] : 
                        (N1092)? in_yumi_i[4] : 
                        (N1094)? in_yumi_i[5] : 
                        (N1096)? in_yumi_i[6] : 
                        (N1098)? in_yumi_i[7] : 
                        (N1085)? in_yumi_i[8] : 
                        (N1087)? in_yumi_i[9] : 
                        (N1089)? in_yumi_i[10] : 
                        (N1091)? in_yumi_i[11] : 
                        (N1093)? in_yumi_i[12] : 
                        (N1095)? in_yumi_i[13] : 
                        (N1097)? in_yumi_i[14] : 
                        (N1099)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[4] = (N1124)? out_me_v_i[0] : 
                         (N1126)? out_me_v_i[1] : 
                         (N1128)? out_me_v_i[2] : 
                         (N1130)? out_me_v_i[3] : 
                         (N1132)? out_me_v_i[4] : 
                         (N1134)? out_me_v_i[5] : 
                         (N1136)? out_me_v_i[6] : 
                         (N1138)? out_me_v_i[7] : 
                         (N1125)? out_me_v_i[8] : 
                         (N1127)? out_me_v_i[9] : 
                         (N1129)? out_me_v_i[10] : 
                         (N1131)? out_me_v_i[11] : 
                         (N1133)? out_me_v_i[12] : 
                         (N1135)? out_me_v_i[13] : 
                         (N1137)? out_me_v_i[14] : 
                         (N1139)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[4] = (N1156)? out_me_ready_i[0] : 
                             (N1158)? out_me_ready_i[1] : 
                             (N1160)? out_me_ready_i[2] : 
                             (N1162)? out_me_ready_i[3] : 
                             (N1164)? out_me_ready_i[4] : 
                             (N1166)? out_me_ready_i[5] : 
                             (N1168)? out_me_ready_i[6] : 
                             (N1170)? out_me_ready_i[7] : 
                             (N1157)? out_me_ready_i[8] : 
                             (N1159)? out_me_ready_i[9] : 
                             (N1161)? out_me_ready_i[10] : 
                             (N1163)? out_me_ready_i[11] : 
                             (N1165)? out_me_ready_i[12] : 
                             (N1167)? out_me_ready_i[13] : 
                             (N1169)? out_me_ready_i[14] : 
                             (N1171)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[5] = (N1208)? in_yumi_i[0] : 
                        (N1210)? in_yumi_i[1] : 
                        (N1212)? in_yumi_i[2] : 
                        (N1214)? in_yumi_i[3] : 
                        (N1216)? in_yumi_i[4] : 
                        (N1218)? in_yumi_i[5] : 
                        (N1220)? in_yumi_i[6] : 
                        (N1222)? in_yumi_i[7] : 
                        (N1209)? in_yumi_i[8] : 
                        (N1211)? in_yumi_i[9] : 
                        (N1213)? in_yumi_i[10] : 
                        (N1215)? in_yumi_i[11] : 
                        (N1217)? in_yumi_i[12] : 
                        (N1219)? in_yumi_i[13] : 
                        (N1221)? in_yumi_i[14] : 
                        (N1223)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[5] = (N1247)? out_me_v_i[0] : 
                         (N1249)? out_me_v_i[1] : 
                         (N1251)? out_me_v_i[2] : 
                         (N1253)? out_me_v_i[3] : 
                         (N1255)? out_me_v_i[4] : 
                         (N1257)? out_me_v_i[5] : 
                         (N1259)? out_me_v_i[6] : 
                         (N1261)? out_me_v_i[7] : 
                         (N1248)? out_me_v_i[8] : 
                         (N1250)? out_me_v_i[9] : 
                         (N1252)? out_me_v_i[10] : 
                         (N1254)? out_me_v_i[11] : 
                         (N1256)? out_me_v_i[12] : 
                         (N1258)? out_me_v_i[13] : 
                         (N1260)? out_me_v_i[14] : 
                         (N1262)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[5] = (N1279)? out_me_ready_i[0] : 
                             (N1281)? out_me_ready_i[1] : 
                             (N1283)? out_me_ready_i[2] : 
                             (N1285)? out_me_ready_i[3] : 
                             (N1287)? out_me_ready_i[4] : 
                             (N1289)? out_me_ready_i[5] : 
                             (N1291)? out_me_ready_i[6] : 
                             (N1293)? out_me_ready_i[7] : 
                             (N1280)? out_me_ready_i[8] : 
                             (N1282)? out_me_ready_i[9] : 
                             (N1284)? out_me_ready_i[10] : 
                             (N1286)? out_me_ready_i[11] : 
                             (N1288)? out_me_ready_i[12] : 
                             (N1290)? out_me_ready_i[13] : 
                             (N1292)? out_me_ready_i[14] : 
                             (N1294)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[6] = (N1333)? in_yumi_i[0] : 
                        (N1335)? in_yumi_i[1] : 
                        (N1337)? in_yumi_i[2] : 
                        (N1339)? in_yumi_i[3] : 
                        (N1341)? in_yumi_i[4] : 
                        (N1343)? in_yumi_i[5] : 
                        (N1345)? in_yumi_i[6] : 
                        (N1347)? in_yumi_i[7] : 
                        (N1334)? in_yumi_i[8] : 
                        (N1336)? in_yumi_i[9] : 
                        (N1338)? in_yumi_i[10] : 
                        (N1340)? in_yumi_i[11] : 
                        (N1342)? in_yumi_i[12] : 
                        (N1344)? in_yumi_i[13] : 
                        (N1346)? in_yumi_i[14] : 
                        (N1348)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[6] = (N1371)? out_me_v_i[0] : 
                         (N1373)? out_me_v_i[1] : 
                         (N1375)? out_me_v_i[2] : 
                         (N1377)? out_me_v_i[3] : 
                         (N1379)? out_me_v_i[4] : 
                         (N1381)? out_me_v_i[5] : 
                         (N1383)? out_me_v_i[6] : 
                         (N1385)? out_me_v_i[7] : 
                         (N1372)? out_me_v_i[8] : 
                         (N1374)? out_me_v_i[9] : 
                         (N1376)? out_me_v_i[10] : 
                         (N1378)? out_me_v_i[11] : 
                         (N1380)? out_me_v_i[12] : 
                         (N1382)? out_me_v_i[13] : 
                         (N1384)? out_me_v_i[14] : 
                         (N1386)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[6] = (N1403)? out_me_ready_i[0] : 
                             (N1405)? out_me_ready_i[1] : 
                             (N1407)? out_me_ready_i[2] : 
                             (N1409)? out_me_ready_i[3] : 
                             (N1411)? out_me_ready_i[4] : 
                             (N1413)? out_me_ready_i[5] : 
                             (N1415)? out_me_ready_i[6] : 
                             (N1417)? out_me_ready_i[7] : 
                             (N1404)? out_me_ready_i[8] : 
                             (N1406)? out_me_ready_i[9] : 
                             (N1408)? out_me_ready_i[10] : 
                             (N1410)? out_me_ready_i[11] : 
                             (N1412)? out_me_ready_i[12] : 
                             (N1414)? out_me_ready_i[13] : 
                             (N1416)? out_me_ready_i[14] : 
                             (N1418)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[7] = (N1458)? in_yumi_i[0] : 
                        (N1460)? in_yumi_i[1] : 
                        (N1462)? in_yumi_i[2] : 
                        (N1464)? in_yumi_i[3] : 
                        (N1466)? in_yumi_i[4] : 
                        (N1468)? in_yumi_i[5] : 
                        (N1470)? in_yumi_i[6] : 
                        (N1472)? in_yumi_i[7] : 
                        (N1459)? in_yumi_i[8] : 
                        (N1461)? in_yumi_i[9] : 
                        (N1463)? in_yumi_i[10] : 
                        (N1465)? in_yumi_i[11] : 
                        (N1467)? in_yumi_i[12] : 
                        (N1469)? in_yumi_i[13] : 
                        (N1471)? in_yumi_i[14] : 
                        (N1473)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[7] = (N1494)? out_me_v_i[0] : 
                         (N1496)? out_me_v_i[1] : 
                         (N1498)? out_me_v_i[2] : 
                         (N1500)? out_me_v_i[3] : 
                         (N1502)? out_me_v_i[4] : 
                         (N1504)? out_me_v_i[5] : 
                         (N1506)? out_me_v_i[6] : 
                         (N1508)? out_me_v_i[7] : 
                         (N1495)? out_me_v_i[8] : 
                         (N1497)? out_me_v_i[9] : 
                         (N1499)? out_me_v_i[10] : 
                         (N1501)? out_me_v_i[11] : 
                         (N1503)? out_me_v_i[12] : 
                         (N1505)? out_me_v_i[13] : 
                         (N1507)? out_me_v_i[14] : 
                         (N1509)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[7] = (N1526)? out_me_ready_i[0] : 
                             (N1528)? out_me_ready_i[1] : 
                             (N1530)? out_me_ready_i[2] : 
                             (N1532)? out_me_ready_i[3] : 
                             (N1534)? out_me_ready_i[4] : 
                             (N1536)? out_me_ready_i[5] : 
                             (N1538)? out_me_ready_i[6] : 
                             (N1540)? out_me_ready_i[7] : 
                             (N1527)? out_me_ready_i[8] : 
                             (N1529)? out_me_ready_i[9] : 
                             (N1531)? out_me_ready_i[10] : 
                             (N1533)? out_me_ready_i[11] : 
                             (N1535)? out_me_ready_i[12] : 
                             (N1537)? out_me_ready_i[13] : 
                             (N1539)? out_me_ready_i[14] : 
                             (N1541)? out_me_ready_i[15] : 1'b0;
  assign out_me_data_o[255] = (N1549)? out_me_data_i_0__31_ : 
                              (N1551)? out_me_data_i[63] : 
                              (N1553)? out_me_data_i[95] : 
                              (N1555)? out_me_data_i[127] : 
                              (N1550)? out_me_data_i[159] : 
                              (N1552)? out_me_data_i[191] : 
                              (N1554)? out_me_data_i[223] : 
                              (N1556)? out_me_data_i[255] : 1'b0;
  assign out_me_data_o[254] = (N1549)? out_me_data_i_0__30_ : 
                              (N1551)? out_me_data_i[62] : 
                              (N1553)? out_me_data_i[94] : 
                              (N1555)? out_me_data_i[126] : 
                              (N1550)? out_me_data_i[158] : 
                              (N1552)? out_me_data_i[190] : 
                              (N1554)? out_me_data_i[222] : 
                              (N1556)? out_me_data_i[254] : 1'b0;
  assign out_me_data_o[253] = (N1549)? out_me_data_i_0__29_ : 
                              (N1551)? out_me_data_i[61] : 
                              (N1553)? out_me_data_i[93] : 
                              (N1555)? out_me_data_i[125] : 
                              (N1550)? out_me_data_i[157] : 
                              (N1552)? out_me_data_i[189] : 
                              (N1554)? out_me_data_i[221] : 
                              (N1556)? out_me_data_i[253] : 1'b0;
  assign out_me_data_o[252] = (N1549)? out_me_data_i_0__28_ : 
                              (N1551)? out_me_data_i[60] : 
                              (N1553)? out_me_data_i[92] : 
                              (N1555)? out_me_data_i[124] : 
                              (N1550)? out_me_data_i[156] : 
                              (N1552)? out_me_data_i[188] : 
                              (N1554)? out_me_data_i[220] : 
                              (N1556)? out_me_data_i[252] : 1'b0;
  assign out_me_data_o[251] = (N1549)? out_me_data_i_0__27_ : 
                              (N1551)? out_me_data_i[59] : 
                              (N1553)? out_me_data_i[91] : 
                              (N1555)? out_me_data_i[123] : 
                              (N1550)? out_me_data_i[155] : 
                              (N1552)? out_me_data_i[187] : 
                              (N1554)? out_me_data_i[219] : 
                              (N1556)? out_me_data_i[251] : 1'b0;
  assign out_me_data_o[250] = (N1549)? out_me_data_i_0__26_ : 
                              (N1551)? out_me_data_i[58] : 
                              (N1553)? out_me_data_i[90] : 
                              (N1555)? out_me_data_i[122] : 
                              (N1550)? out_me_data_i[154] : 
                              (N1552)? out_me_data_i[186] : 
                              (N1554)? out_me_data_i[218] : 
                              (N1556)? out_me_data_i[250] : 1'b0;
  assign out_me_data_o[249] = (N1549)? out_me_data_i_0__25_ : 
                              (N1551)? out_me_data_i[57] : 
                              (N1553)? out_me_data_i[89] : 
                              (N1555)? out_me_data_i[121] : 
                              (N1550)? out_me_data_i[153] : 
                              (N1552)? out_me_data_i[185] : 
                              (N1554)? out_me_data_i[217] : 
                              (N1556)? out_me_data_i[249] : 1'b0;
  assign out_me_data_o[248] = (N1549)? out_me_data_i_0__24_ : 
                              (N1551)? out_me_data_i[56] : 
                              (N1553)? out_me_data_i[88] : 
                              (N1555)? out_me_data_i[120] : 
                              (N1550)? out_me_data_i[152] : 
                              (N1552)? out_me_data_i[184] : 
                              (N1554)? out_me_data_i[216] : 
                              (N1556)? out_me_data_i[248] : 1'b0;
  assign out_me_data_o[247] = (N1549)? out_me_data_i_0__23_ : 
                              (N1551)? out_me_data_i[55] : 
                              (N1553)? out_me_data_i[87] : 
                              (N1555)? out_me_data_i[119] : 
                              (N1550)? out_me_data_i[151] : 
                              (N1552)? out_me_data_i[183] : 
                              (N1554)? out_me_data_i[215] : 
                              (N1556)? out_me_data_i[247] : 1'b0;
  assign out_me_data_o[246] = (N1549)? out_me_data_i_0__22_ : 
                              (N1551)? out_me_data_i[54] : 
                              (N1553)? out_me_data_i[86] : 
                              (N1555)? out_me_data_i[118] : 
                              (N1550)? out_me_data_i[150] : 
                              (N1552)? out_me_data_i[182] : 
                              (N1554)? out_me_data_i[214] : 
                              (N1556)? out_me_data_i[246] : 1'b0;
  assign out_me_data_o[245] = (N1549)? out_me_data_i_0__21_ : 
                              (N1551)? out_me_data_i[53] : 
                              (N1553)? out_me_data_i[85] : 
                              (N1555)? out_me_data_i[117] : 
                              (N1550)? out_me_data_i[149] : 
                              (N1552)? out_me_data_i[181] : 
                              (N1554)? out_me_data_i[213] : 
                              (N1556)? out_me_data_i[245] : 1'b0;
  assign out_me_data_o[244] = (N1549)? out_me_data_i_0__20_ : 
                              (N1551)? out_me_data_i[52] : 
                              (N1553)? out_me_data_i[84] : 
                              (N1555)? out_me_data_i[116] : 
                              (N1550)? out_me_data_i[148] : 
                              (N1552)? out_me_data_i[180] : 
                              (N1554)? out_me_data_i[212] : 
                              (N1556)? out_me_data_i[244] : 1'b0;
  assign out_me_data_o[243] = (N1549)? out_me_data_i_0__19_ : 
                              (N1551)? out_me_data_i[51] : 
                              (N1553)? out_me_data_i[83] : 
                              (N1555)? out_me_data_i[115] : 
                              (N1550)? out_me_data_i[147] : 
                              (N1552)? out_me_data_i[179] : 
                              (N1554)? out_me_data_i[211] : 
                              (N1556)? out_me_data_i[243] : 1'b0;
  assign out_me_data_o[242] = (N1549)? out_me_data_i_0__18_ : 
                              (N1551)? out_me_data_i[50] : 
                              (N1553)? out_me_data_i[82] : 
                              (N1555)? out_me_data_i[114] : 
                              (N1550)? out_me_data_i[146] : 
                              (N1552)? out_me_data_i[178] : 
                              (N1554)? out_me_data_i[210] : 
                              (N1556)? out_me_data_i[242] : 1'b0;
  assign out_me_data_o[241] = (N1549)? out_me_data_i_0__17_ : 
                              (N1551)? out_me_data_i[49] : 
                              (N1553)? out_me_data_i[81] : 
                              (N1555)? out_me_data_i[113] : 
                              (N1550)? out_me_data_i[145] : 
                              (N1552)? out_me_data_i[177] : 
                              (N1554)? out_me_data_i[209] : 
                              (N1556)? out_me_data_i[241] : 1'b0;
  assign out_me_data_o[240] = (N1549)? out_me_data_i_0__16_ : 
                              (N1551)? out_me_data_i[48] : 
                              (N1553)? out_me_data_i[80] : 
                              (N1555)? out_me_data_i[112] : 
                              (N1550)? out_me_data_i[144] : 
                              (N1552)? out_me_data_i[176] : 
                              (N1554)? out_me_data_i[208] : 
                              (N1556)? out_me_data_i[240] : 1'b0;
  assign out_me_data_o[239] = (N1549)? out_me_data_i_0__15_ : 
                              (N1551)? out_me_data_i[47] : 
                              (N1553)? out_me_data_i[79] : 
                              (N1555)? out_me_data_i[111] : 
                              (N1550)? out_me_data_i[143] : 
                              (N1552)? out_me_data_i[175] : 
                              (N1554)? out_me_data_i[207] : 
                              (N1556)? out_me_data_i[239] : 1'b0;
  assign out_me_data_o[238] = (N1549)? out_me_data_i_0__14_ : 
                              (N1551)? out_me_data_i[46] : 
                              (N1553)? out_me_data_i[78] : 
                              (N1555)? out_me_data_i[110] : 
                              (N1550)? out_me_data_i[142] : 
                              (N1552)? out_me_data_i[174] : 
                              (N1554)? out_me_data_i[206] : 
                              (N1556)? out_me_data_i[238] : 1'b0;
  assign out_me_data_o[237] = (N1549)? out_me_data_i_0__13_ : 
                              (N1551)? out_me_data_i[45] : 
                              (N1553)? out_me_data_i[77] : 
                              (N1555)? out_me_data_i[109] : 
                              (N1550)? out_me_data_i[141] : 
                              (N1552)? out_me_data_i[173] : 
                              (N1554)? out_me_data_i[205] : 
                              (N1556)? out_me_data_i[237] : 1'b0;
  assign out_me_data_o[236] = (N1549)? out_me_data_i_0__12_ : 
                              (N1551)? out_me_data_i[44] : 
                              (N1553)? out_me_data_i[76] : 
                              (N1555)? out_me_data_i[108] : 
                              (N1550)? out_me_data_i[140] : 
                              (N1552)? out_me_data_i[172] : 
                              (N1554)? out_me_data_i[204] : 
                              (N1556)? out_me_data_i[236] : 1'b0;
  assign out_me_data_o[235] = (N1549)? out_me_data_i_0__11_ : 
                              (N1551)? out_me_data_i[43] : 
                              (N1553)? out_me_data_i[75] : 
                              (N1555)? out_me_data_i[107] : 
                              (N1550)? out_me_data_i[139] : 
                              (N1552)? out_me_data_i[171] : 
                              (N1554)? out_me_data_i[203] : 
                              (N1556)? out_me_data_i[235] : 1'b0;
  assign out_me_data_o[234] = (N1549)? out_me_data_i_0__10_ : 
                              (N1551)? out_me_data_i[42] : 
                              (N1553)? out_me_data_i[74] : 
                              (N1555)? out_me_data_i[106] : 
                              (N1550)? out_me_data_i[138] : 
                              (N1552)? out_me_data_i[170] : 
                              (N1554)? out_me_data_i[202] : 
                              (N1556)? out_me_data_i[234] : 1'b0;
  assign out_me_data_o[233] = (N1549)? out_me_data_i_0__9_ : 
                              (N1551)? out_me_data_i[41] : 
                              (N1553)? out_me_data_i[73] : 
                              (N1555)? out_me_data_i[105] : 
                              (N1550)? out_me_data_i[137] : 
                              (N1552)? out_me_data_i[169] : 
                              (N1554)? out_me_data_i[201] : 
                              (N1556)? out_me_data_i[233] : 1'b0;
  assign out_me_data_o[232] = (N1549)? out_me_data_i_0__8_ : 
                              (N1551)? out_me_data_i[40] : 
                              (N1553)? out_me_data_i[72] : 
                              (N1555)? out_me_data_i[104] : 
                              (N1550)? out_me_data_i[136] : 
                              (N1552)? out_me_data_i[168] : 
                              (N1554)? out_me_data_i[200] : 
                              (N1556)? out_me_data_i[232] : 1'b0;
  assign out_me_data_o[231] = (N1549)? out_me_data_i_0__7_ : 
                              (N1551)? out_me_data_i[39] : 
                              (N1553)? out_me_data_i[71] : 
                              (N1555)? out_me_data_i[103] : 
                              (N1550)? out_me_data_i[135] : 
                              (N1552)? out_me_data_i[167] : 
                              (N1554)? out_me_data_i[199] : 
                              (N1556)? out_me_data_i[231] : 1'b0;
  assign out_me_data_o[230] = (N1549)? out_me_data_i_0__6_ : 
                              (N1551)? out_me_data_i[38] : 
                              (N1553)? out_me_data_i[70] : 
                              (N1555)? out_me_data_i[102] : 
                              (N1550)? out_me_data_i[134] : 
                              (N1552)? out_me_data_i[166] : 
                              (N1554)? out_me_data_i[198] : 
                              (N1556)? out_me_data_i[230] : 1'b0;
  assign out_me_data_o[229] = (N1549)? out_me_data_i_0__5_ : 
                              (N1551)? out_me_data_i[37] : 
                              (N1553)? out_me_data_i[69] : 
                              (N1555)? out_me_data_i[101] : 
                              (N1550)? out_me_data_i[133] : 
                              (N1552)? out_me_data_i[165] : 
                              (N1554)? out_me_data_i[197] : 
                              (N1556)? out_me_data_i[229] : 1'b0;
  assign out_me_data_o[228] = (N1549)? out_me_data_i_0__4_ : 
                              (N1551)? out_me_data_i[36] : 
                              (N1553)? out_me_data_i[68] : 
                              (N1555)? out_me_data_i[100] : 
                              (N1550)? out_me_data_i[132] : 
                              (N1552)? out_me_data_i[164] : 
                              (N1554)? out_me_data_i[196] : 
                              (N1556)? out_me_data_i[228] : 1'b0;
  assign out_me_data_o[227] = (N1549)? out_me_data_i_0__3_ : 
                              (N1551)? out_me_data_i[35] : 
                              (N1553)? out_me_data_i[67] : 
                              (N1555)? out_me_data_i[99] : 
                              (N1550)? out_me_data_i[131] : 
                              (N1552)? out_me_data_i[163] : 
                              (N1554)? out_me_data_i[195] : 
                              (N1556)? out_me_data_i[227] : 1'b0;
  assign out_me_data_o[226] = (N1549)? out_me_data_i_0__2_ : 
                              (N1551)? out_me_data_i[34] : 
                              (N1553)? out_me_data_i[66] : 
                              (N1555)? out_me_data_i[98] : 
                              (N1550)? out_me_data_i[130] : 
                              (N1552)? out_me_data_i[162] : 
                              (N1554)? out_me_data_i[194] : 
                              (N1556)? out_me_data_i[226] : 1'b0;
  assign out_me_data_o[225] = (N1549)? out_me_data_i_0__1_ : 
                              (N1551)? out_me_data_i[33] : 
                              (N1553)? out_me_data_i[65] : 
                              (N1555)? out_me_data_i[97] : 
                              (N1550)? out_me_data_i[129] : 
                              (N1552)? out_me_data_i[161] : 
                              (N1554)? out_me_data_i[193] : 
                              (N1556)? out_me_data_i[225] : 1'b0;
  assign out_me_data_o[224] = (N1549)? out_me_data_i_0__0_ : 
                              (N1551)? out_me_data_i[32] : 
                              (N1553)? out_me_data_i[64] : 
                              (N1555)? out_me_data_i[96] : 
                              (N1550)? out_me_data_i[128] : 
                              (N1552)? out_me_data_i[160] : 
                              (N1554)? out_me_data_i[192] : 
                              (N1556)? out_me_data_i[224] : 1'b0;
  assign in_yumi_o[8] = (N1589)? in_yumi_i[0] : 
                        (N1591)? in_yumi_i[1] : 
                        (N1593)? in_yumi_i[2] : 
                        (N1595)? in_yumi_i[3] : 
                        (N1597)? in_yumi_i[4] : 
                        (N1599)? in_yumi_i[5] : 
                        (N1601)? in_yumi_i[6] : 
                        (N1603)? in_yumi_i[7] : 
                        (N1590)? in_yumi_i[8] : 
                        (N1592)? in_yumi_i[9] : 
                        (N1594)? in_yumi_i[10] : 
                        (N1596)? in_yumi_i[11] : 
                        (N1598)? in_yumi_i[12] : 
                        (N1600)? in_yumi_i[13] : 
                        (N1602)? in_yumi_i[14] : 
                        (N1604)? in_yumi_i[15] : 1'b0;
  assign in_data_o[287] = (N1612)? in_data_i[287] : 
                          (N1614)? in_data_i[319] : 
                          (N1616)? in_data_i[351] : 
                          (N1618)? in_data_i[383] : 
                          (N1613)? in_data_i[415] : 
                          (N1615)? in_data_i[447] : 
                          (N1617)? in_data_i[479] : 
                          (N1619)? in_data_i_15__31_ : 1'b0;
  assign in_data_o[286] = (N1612)? in_data_i[286] : 
                          (N1614)? in_data_i[318] : 
                          (N1616)? in_data_i[350] : 
                          (N1618)? in_data_i[382] : 
                          (N1613)? in_data_i[414] : 
                          (N1615)? in_data_i[446] : 
                          (N1617)? in_data_i[478] : 
                          (N1619)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[285] = (N1612)? in_data_i[285] : 
                          (N1614)? in_data_i[317] : 
                          (N1616)? in_data_i[349] : 
                          (N1618)? in_data_i[381] : 
                          (N1613)? in_data_i[413] : 
                          (N1615)? in_data_i[445] : 
                          (N1617)? in_data_i[477] : 
                          (N1619)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[284] = (N1612)? in_data_i[284] : 
                          (N1614)? in_data_i[316] : 
                          (N1616)? in_data_i[348] : 
                          (N1618)? in_data_i[380] : 
                          (N1613)? in_data_i[412] : 
                          (N1615)? in_data_i[444] : 
                          (N1617)? in_data_i[476] : 
                          (N1619)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[283] = (N1612)? in_data_i[283] : 
                          (N1614)? in_data_i[315] : 
                          (N1616)? in_data_i[347] : 
                          (N1618)? in_data_i[379] : 
                          (N1613)? in_data_i[411] : 
                          (N1615)? in_data_i[443] : 
                          (N1617)? in_data_i[475] : 
                          (N1619)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[282] = (N1612)? in_data_i[282] : 
                          (N1614)? in_data_i[314] : 
                          (N1616)? in_data_i[346] : 
                          (N1618)? in_data_i[378] : 
                          (N1613)? in_data_i[410] : 
                          (N1615)? in_data_i[442] : 
                          (N1617)? in_data_i[474] : 
                          (N1619)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[281] = (N1612)? in_data_i[281] : 
                          (N1614)? in_data_i[313] : 
                          (N1616)? in_data_i[345] : 
                          (N1618)? in_data_i[377] : 
                          (N1613)? in_data_i[409] : 
                          (N1615)? in_data_i[441] : 
                          (N1617)? in_data_i[473] : 
                          (N1619)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[280] = (N1612)? in_data_i[280] : 
                          (N1614)? in_data_i[312] : 
                          (N1616)? in_data_i[344] : 
                          (N1618)? in_data_i[376] : 
                          (N1613)? in_data_i[408] : 
                          (N1615)? in_data_i[440] : 
                          (N1617)? in_data_i[472] : 
                          (N1619)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[279] = (N1612)? in_data_i[279] : 
                          (N1614)? in_data_i[311] : 
                          (N1616)? in_data_i[343] : 
                          (N1618)? in_data_i[375] : 
                          (N1613)? in_data_i[407] : 
                          (N1615)? in_data_i[439] : 
                          (N1617)? in_data_i[471] : 
                          (N1619)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[278] = (N1612)? in_data_i[278] : 
                          (N1614)? in_data_i[310] : 
                          (N1616)? in_data_i[342] : 
                          (N1618)? in_data_i[374] : 
                          (N1613)? in_data_i[406] : 
                          (N1615)? in_data_i[438] : 
                          (N1617)? in_data_i[470] : 
                          (N1619)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[277] = (N1612)? in_data_i[277] : 
                          (N1614)? in_data_i[309] : 
                          (N1616)? in_data_i[341] : 
                          (N1618)? in_data_i[373] : 
                          (N1613)? in_data_i[405] : 
                          (N1615)? in_data_i[437] : 
                          (N1617)? in_data_i[469] : 
                          (N1619)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[276] = (N1612)? in_data_i[276] : 
                          (N1614)? in_data_i[308] : 
                          (N1616)? in_data_i[340] : 
                          (N1618)? in_data_i[372] : 
                          (N1613)? in_data_i[404] : 
                          (N1615)? in_data_i[436] : 
                          (N1617)? in_data_i[468] : 
                          (N1619)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[275] = (N1612)? in_data_i[275] : 
                          (N1614)? in_data_i[307] : 
                          (N1616)? in_data_i[339] : 
                          (N1618)? in_data_i[371] : 
                          (N1613)? in_data_i[403] : 
                          (N1615)? in_data_i[435] : 
                          (N1617)? in_data_i[467] : 
                          (N1619)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[274] = (N1612)? in_data_i[274] : 
                          (N1614)? in_data_i[306] : 
                          (N1616)? in_data_i[338] : 
                          (N1618)? in_data_i[370] : 
                          (N1613)? in_data_i[402] : 
                          (N1615)? in_data_i[434] : 
                          (N1617)? in_data_i[466] : 
                          (N1619)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[273] = (N1612)? in_data_i[273] : 
                          (N1614)? in_data_i[305] : 
                          (N1616)? in_data_i[337] : 
                          (N1618)? in_data_i[369] : 
                          (N1613)? in_data_i[401] : 
                          (N1615)? in_data_i[433] : 
                          (N1617)? in_data_i[465] : 
                          (N1619)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[272] = (N1612)? in_data_i[272] : 
                          (N1614)? in_data_i[304] : 
                          (N1616)? in_data_i[336] : 
                          (N1618)? in_data_i[368] : 
                          (N1613)? in_data_i[400] : 
                          (N1615)? in_data_i[432] : 
                          (N1617)? in_data_i[464] : 
                          (N1619)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[271] = (N1612)? in_data_i[271] : 
                          (N1614)? in_data_i[303] : 
                          (N1616)? in_data_i[335] : 
                          (N1618)? in_data_i[367] : 
                          (N1613)? in_data_i[399] : 
                          (N1615)? in_data_i[431] : 
                          (N1617)? in_data_i[463] : 
                          (N1619)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[270] = (N1612)? in_data_i[270] : 
                          (N1614)? in_data_i[302] : 
                          (N1616)? in_data_i[334] : 
                          (N1618)? in_data_i[366] : 
                          (N1613)? in_data_i[398] : 
                          (N1615)? in_data_i[430] : 
                          (N1617)? in_data_i[462] : 
                          (N1619)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[269] = (N1612)? in_data_i[269] : 
                          (N1614)? in_data_i[301] : 
                          (N1616)? in_data_i[333] : 
                          (N1618)? in_data_i[365] : 
                          (N1613)? in_data_i[397] : 
                          (N1615)? in_data_i[429] : 
                          (N1617)? in_data_i[461] : 
                          (N1619)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[268] = (N1612)? in_data_i[268] : 
                          (N1614)? in_data_i[300] : 
                          (N1616)? in_data_i[332] : 
                          (N1618)? in_data_i[364] : 
                          (N1613)? in_data_i[396] : 
                          (N1615)? in_data_i[428] : 
                          (N1617)? in_data_i[460] : 
                          (N1619)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[267] = (N1612)? in_data_i[267] : 
                          (N1614)? in_data_i[299] : 
                          (N1616)? in_data_i[331] : 
                          (N1618)? in_data_i[363] : 
                          (N1613)? in_data_i[395] : 
                          (N1615)? in_data_i[427] : 
                          (N1617)? in_data_i[459] : 
                          (N1619)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[266] = (N1612)? in_data_i[266] : 
                          (N1614)? in_data_i[298] : 
                          (N1616)? in_data_i[330] : 
                          (N1618)? in_data_i[362] : 
                          (N1613)? in_data_i[394] : 
                          (N1615)? in_data_i[426] : 
                          (N1617)? in_data_i[458] : 
                          (N1619)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[265] = (N1612)? in_data_i[265] : 
                          (N1614)? in_data_i[297] : 
                          (N1616)? in_data_i[329] : 
                          (N1618)? in_data_i[361] : 
                          (N1613)? in_data_i[393] : 
                          (N1615)? in_data_i[425] : 
                          (N1617)? in_data_i[457] : 
                          (N1619)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[264] = (N1612)? in_data_i[264] : 
                          (N1614)? in_data_i[296] : 
                          (N1616)? in_data_i[328] : 
                          (N1618)? in_data_i[360] : 
                          (N1613)? in_data_i[392] : 
                          (N1615)? in_data_i[424] : 
                          (N1617)? in_data_i[456] : 
                          (N1619)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[263] = (N1612)? in_data_i[263] : 
                          (N1614)? in_data_i[295] : 
                          (N1616)? in_data_i[327] : 
                          (N1618)? in_data_i[359] : 
                          (N1613)? in_data_i[391] : 
                          (N1615)? in_data_i[423] : 
                          (N1617)? in_data_i[455] : 
                          (N1619)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[262] = (N1612)? in_data_i[262] : 
                          (N1614)? in_data_i[294] : 
                          (N1616)? in_data_i[326] : 
                          (N1618)? in_data_i[358] : 
                          (N1613)? in_data_i[390] : 
                          (N1615)? in_data_i[422] : 
                          (N1617)? in_data_i[454] : 
                          (N1619)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[261] = (N1612)? in_data_i[261] : 
                          (N1614)? in_data_i[293] : 
                          (N1616)? in_data_i[325] : 
                          (N1618)? in_data_i[357] : 
                          (N1613)? in_data_i[389] : 
                          (N1615)? in_data_i[421] : 
                          (N1617)? in_data_i[453] : 
                          (N1619)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[260] = (N1612)? in_data_i[260] : 
                          (N1614)? in_data_i[292] : 
                          (N1616)? in_data_i[324] : 
                          (N1618)? in_data_i[356] : 
                          (N1613)? in_data_i[388] : 
                          (N1615)? in_data_i[420] : 
                          (N1617)? in_data_i[452] : 
                          (N1619)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[259] = (N1612)? in_data_i[259] : 
                          (N1614)? in_data_i[291] : 
                          (N1616)? in_data_i[323] : 
                          (N1618)? in_data_i[355] : 
                          (N1613)? in_data_i[387] : 
                          (N1615)? in_data_i[419] : 
                          (N1617)? in_data_i[451] : 
                          (N1619)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[258] = (N1612)? in_data_i[258] : 
                          (N1614)? in_data_i[290] : 
                          (N1616)? in_data_i[322] : 
                          (N1618)? in_data_i[354] : 
                          (N1613)? in_data_i[386] : 
                          (N1615)? in_data_i[418] : 
                          (N1617)? in_data_i[450] : 
                          (N1619)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[257] = (N1612)? in_data_i[257] : 
                          (N1614)? in_data_i[289] : 
                          (N1616)? in_data_i[321] : 
                          (N1618)? in_data_i[353] : 
                          (N1613)? in_data_i[385] : 
                          (N1615)? in_data_i[417] : 
                          (N1617)? in_data_i[449] : 
                          (N1619)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[256] = (N1612)? in_data_i[256] : 
                          (N1614)? in_data_i[288] : 
                          (N1616)? in_data_i[320] : 
                          (N1618)? in_data_i[352] : 
                          (N1613)? in_data_i[384] : 
                          (N1615)? in_data_i[416] : 
                          (N1617)? in_data_i[448] : 
                          (N1619)? in_data_i_15__0_ : 1'b0;
  assign out_me_v_o[8] = (N1632)? out_me_v_i[0] : 
                         (N1634)? out_me_v_i[1] : 
                         (N1636)? out_me_v_i[2] : 
                         (N1638)? out_me_v_i[3] : 
                         (N1640)? out_me_v_i[4] : 
                         (N1642)? out_me_v_i[5] : 
                         (N1644)? out_me_v_i[6] : 
                         (N1646)? out_me_v_i[7] : 
                         (N1633)? out_me_v_i[8] : 
                         (N1635)? out_me_v_i[9] : 
                         (N1637)? out_me_v_i[10] : 
                         (N1639)? out_me_v_i[11] : 
                         (N1641)? out_me_v_i[12] : 
                         (N1643)? out_me_v_i[13] : 
                         (N1645)? out_me_v_i[14] : 
                         (N1647)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[8] = (N1664)? out_me_ready_i[0] : 
                             (N1666)? out_me_ready_i[1] : 
                             (N1668)? out_me_ready_i[2] : 
                             (N1670)? out_me_ready_i[3] : 
                             (N1672)? out_me_ready_i[4] : 
                             (N1674)? out_me_ready_i[5] : 
                             (N1676)? out_me_ready_i[6] : 
                             (N1678)? out_me_ready_i[7] : 
                             (N1665)? out_me_ready_i[8] : 
                             (N1667)? out_me_ready_i[9] : 
                             (N1669)? out_me_ready_i[10] : 
                             (N1671)? out_me_ready_i[11] : 
                             (N1673)? out_me_ready_i[12] : 
                             (N1675)? out_me_ready_i[13] : 
                             (N1677)? out_me_ready_i[14] : 
                             (N1679)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[9] = (N1720)? in_yumi_i[0] : 
                        (N1722)? in_yumi_i[1] : 
                        (N1724)? in_yumi_i[2] : 
                        (N1726)? in_yumi_i[3] : 
                        (N1728)? in_yumi_i[4] : 
                        (N1730)? in_yumi_i[5] : 
                        (N1732)? in_yumi_i[6] : 
                        (N1734)? in_yumi_i[7] : 
                        (N1721)? in_yumi_i[8] : 
                        (N1723)? in_yumi_i[9] : 
                        (N1725)? in_yumi_i[10] : 
                        (N1727)? in_yumi_i[11] : 
                        (N1729)? in_yumi_i[12] : 
                        (N1731)? in_yumi_i[13] : 
                        (N1733)? in_yumi_i[14] : 
                        (N1735)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[9] = (N1755)? out_me_v_i[0] : 
                         (N1757)? out_me_v_i[1] : 
                         (N1759)? out_me_v_i[2] : 
                         (N1761)? out_me_v_i[3] : 
                         (N1763)? out_me_v_i[4] : 
                         (N1765)? out_me_v_i[5] : 
                         (N1767)? out_me_v_i[6] : 
                         (N1769)? out_me_v_i[7] : 
                         (N1756)? out_me_v_i[8] : 
                         (N1758)? out_me_v_i[9] : 
                         (N1760)? out_me_v_i[10] : 
                         (N1762)? out_me_v_i[11] : 
                         (N1764)? out_me_v_i[12] : 
                         (N1766)? out_me_v_i[13] : 
                         (N1768)? out_me_v_i[14] : 
                         (N1770)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[9] = (N1787)? out_me_ready_i[0] : 
                             (N1789)? out_me_ready_i[1] : 
                             (N1791)? out_me_ready_i[2] : 
                             (N1793)? out_me_ready_i[3] : 
                             (N1795)? out_me_ready_i[4] : 
                             (N1797)? out_me_ready_i[5] : 
                             (N1799)? out_me_ready_i[6] : 
                             (N1801)? out_me_ready_i[7] : 
                             (N1788)? out_me_ready_i[8] : 
                             (N1790)? out_me_ready_i[9] : 
                             (N1792)? out_me_ready_i[10] : 
                             (N1794)? out_me_ready_i[11] : 
                             (N1796)? out_me_ready_i[12] : 
                             (N1798)? out_me_ready_i[13] : 
                             (N1800)? out_me_ready_i[14] : 
                             (N1802)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[10] = (N1845)? in_yumi_i[0] : 
                         (N1847)? in_yumi_i[1] : 
                         (N1849)? in_yumi_i[2] : 
                         (N1851)? in_yumi_i[3] : 
                         (N1853)? in_yumi_i[4] : 
                         (N1855)? in_yumi_i[5] : 
                         (N1857)? in_yumi_i[6] : 
                         (N1859)? in_yumi_i[7] : 
                         (N1846)? in_yumi_i[8] : 
                         (N1848)? in_yumi_i[9] : 
                         (N1850)? in_yumi_i[10] : 
                         (N1852)? in_yumi_i[11] : 
                         (N1854)? in_yumi_i[12] : 
                         (N1856)? in_yumi_i[13] : 
                         (N1858)? in_yumi_i[14] : 
                         (N1860)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[10] = (N1879)? out_me_v_i[0] : 
                          (N1881)? out_me_v_i[1] : 
                          (N1883)? out_me_v_i[2] : 
                          (N1885)? out_me_v_i[3] : 
                          (N1887)? out_me_v_i[4] : 
                          (N1889)? out_me_v_i[5] : 
                          (N1891)? out_me_v_i[6] : 
                          (N1893)? out_me_v_i[7] : 
                          (N1880)? out_me_v_i[8] : 
                          (N1882)? out_me_v_i[9] : 
                          (N1884)? out_me_v_i[10] : 
                          (N1886)? out_me_v_i[11] : 
                          (N1888)? out_me_v_i[12] : 
                          (N1890)? out_me_v_i[13] : 
                          (N1892)? out_me_v_i[14] : 
                          (N1894)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[10] = (N1911)? out_me_ready_i[0] : 
                              (N1913)? out_me_ready_i[1] : 
                              (N1915)? out_me_ready_i[2] : 
                              (N1917)? out_me_ready_i[3] : 
                              (N1919)? out_me_ready_i[4] : 
                              (N1921)? out_me_ready_i[5] : 
                              (N1923)? out_me_ready_i[6] : 
                              (N1925)? out_me_ready_i[7] : 
                              (N1912)? out_me_ready_i[8] : 
                              (N1914)? out_me_ready_i[9] : 
                              (N1916)? out_me_ready_i[10] : 
                              (N1918)? out_me_ready_i[11] : 
                              (N1920)? out_me_ready_i[12] : 
                              (N1922)? out_me_ready_i[13] : 
                              (N1924)? out_me_ready_i[14] : 
                              (N1926)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[11] = (N1970)? in_yumi_i[0] : 
                         (N1972)? in_yumi_i[1] : 
                         (N1974)? in_yumi_i[2] : 
                         (N1976)? in_yumi_i[3] : 
                         (N1978)? in_yumi_i[4] : 
                         (N1980)? in_yumi_i[5] : 
                         (N1982)? in_yumi_i[6] : 
                         (N1984)? in_yumi_i[7] : 
                         (N1971)? in_yumi_i[8] : 
                         (N1973)? in_yumi_i[9] : 
                         (N1975)? in_yumi_i[10] : 
                         (N1977)? in_yumi_i[11] : 
                         (N1979)? in_yumi_i[12] : 
                         (N1981)? in_yumi_i[13] : 
                         (N1983)? in_yumi_i[14] : 
                         (N1985)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[11] = (N2002)? out_me_v_i[0] : 
                          (N2004)? out_me_v_i[1] : 
                          (N2006)? out_me_v_i[2] : 
                          (N2008)? out_me_v_i[3] : 
                          (N2010)? out_me_v_i[4] : 
                          (N2012)? out_me_v_i[5] : 
                          (N2014)? out_me_v_i[6] : 
                          (N2016)? out_me_v_i[7] : 
                          (N2003)? out_me_v_i[8] : 
                          (N2005)? out_me_v_i[9] : 
                          (N2007)? out_me_v_i[10] : 
                          (N2009)? out_me_v_i[11] : 
                          (N2011)? out_me_v_i[12] : 
                          (N2013)? out_me_v_i[13] : 
                          (N2015)? out_me_v_i[14] : 
                          (N2017)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[11] = (N2034)? out_me_ready_i[0] : 
                              (N2036)? out_me_ready_i[1] : 
                              (N2038)? out_me_ready_i[2] : 
                              (N2040)? out_me_ready_i[3] : 
                              (N2042)? out_me_ready_i[4] : 
                              (N2044)? out_me_ready_i[5] : 
                              (N2046)? out_me_ready_i[6] : 
                              (N2048)? out_me_ready_i[7] : 
                              (N2035)? out_me_ready_i[8] : 
                              (N2037)? out_me_ready_i[9] : 
                              (N2039)? out_me_ready_i[10] : 
                              (N2041)? out_me_ready_i[11] : 
                              (N2043)? out_me_ready_i[12] : 
                              (N2045)? out_me_ready_i[13] : 
                              (N2047)? out_me_ready_i[14] : 
                              (N2049)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[12] = (N2094)? in_yumi_i[0] : 
                         (N2096)? in_yumi_i[1] : 
                         (N2098)? in_yumi_i[2] : 
                         (N2100)? in_yumi_i[3] : 
                         (N2102)? in_yumi_i[4] : 
                         (N2104)? in_yumi_i[5] : 
                         (N2106)? in_yumi_i[6] : 
                         (N2108)? in_yumi_i[7] : 
                         (N2095)? in_yumi_i[8] : 
                         (N2097)? in_yumi_i[9] : 
                         (N2099)? in_yumi_i[10] : 
                         (N2101)? in_yumi_i[11] : 
                         (N2103)? in_yumi_i[12] : 
                         (N2105)? in_yumi_i[13] : 
                         (N2107)? in_yumi_i[14] : 
                         (N2109)? in_yumi_i[15] : 1'b0;
  assign in_data_o[415] = (N2112)? in_data_i[415] : 
                          (N2114)? in_data_i[447] : 
                          (N2113)? in_data_i[479] : 
                          (N2115)? in_data_i_15__31_ : 1'b0;
  assign in_data_o[414] = (N2112)? in_data_i[414] : 
                          (N2114)? in_data_i[446] : 
                          (N2113)? in_data_i[478] : 
                          (N2115)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[413] = (N2112)? in_data_i[413] : 
                          (N2114)? in_data_i[445] : 
                          (N2113)? in_data_i[477] : 
                          (N2115)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[412] = (N2112)? in_data_i[412] : 
                          (N2114)? in_data_i[444] : 
                          (N2113)? in_data_i[476] : 
                          (N2115)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[411] = (N2112)? in_data_i[411] : 
                          (N2114)? in_data_i[443] : 
                          (N2113)? in_data_i[475] : 
                          (N2115)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[410] = (N2112)? in_data_i[410] : 
                          (N2114)? in_data_i[442] : 
                          (N2113)? in_data_i[474] : 
                          (N2115)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[409] = (N2112)? in_data_i[409] : 
                          (N2114)? in_data_i[441] : 
                          (N2113)? in_data_i[473] : 
                          (N2115)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[408] = (N2112)? in_data_i[408] : 
                          (N2114)? in_data_i[440] : 
                          (N2113)? in_data_i[472] : 
                          (N2115)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[407] = (N2112)? in_data_i[407] : 
                          (N2114)? in_data_i[439] : 
                          (N2113)? in_data_i[471] : 
                          (N2115)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[406] = (N2112)? in_data_i[406] : 
                          (N2114)? in_data_i[438] : 
                          (N2113)? in_data_i[470] : 
                          (N2115)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[405] = (N2112)? in_data_i[405] : 
                          (N2114)? in_data_i[437] : 
                          (N2113)? in_data_i[469] : 
                          (N2115)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[404] = (N2112)? in_data_i[404] : 
                          (N2114)? in_data_i[436] : 
                          (N2113)? in_data_i[468] : 
                          (N2115)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[403] = (N2112)? in_data_i[403] : 
                          (N2114)? in_data_i[435] : 
                          (N2113)? in_data_i[467] : 
                          (N2115)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[402] = (N2112)? in_data_i[402] : 
                          (N2114)? in_data_i[434] : 
                          (N2113)? in_data_i[466] : 
                          (N2115)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[401] = (N2112)? in_data_i[401] : 
                          (N2114)? in_data_i[433] : 
                          (N2113)? in_data_i[465] : 
                          (N2115)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[400] = (N2112)? in_data_i[400] : 
                          (N2114)? in_data_i[432] : 
                          (N2113)? in_data_i[464] : 
                          (N2115)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[399] = (N2112)? in_data_i[399] : 
                          (N2114)? in_data_i[431] : 
                          (N2113)? in_data_i[463] : 
                          (N2115)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[398] = (N2112)? in_data_i[398] : 
                          (N2114)? in_data_i[430] : 
                          (N2113)? in_data_i[462] : 
                          (N2115)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[397] = (N2112)? in_data_i[397] : 
                          (N2114)? in_data_i[429] : 
                          (N2113)? in_data_i[461] : 
                          (N2115)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[396] = (N2112)? in_data_i[396] : 
                          (N2114)? in_data_i[428] : 
                          (N2113)? in_data_i[460] : 
                          (N2115)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[395] = (N2112)? in_data_i[395] : 
                          (N2114)? in_data_i[427] : 
                          (N2113)? in_data_i[459] : 
                          (N2115)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[394] = (N2112)? in_data_i[394] : 
                          (N2114)? in_data_i[426] : 
                          (N2113)? in_data_i[458] : 
                          (N2115)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[393] = (N2112)? in_data_i[393] : 
                          (N2114)? in_data_i[425] : 
                          (N2113)? in_data_i[457] : 
                          (N2115)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[392] = (N2112)? in_data_i[392] : 
                          (N2114)? in_data_i[424] : 
                          (N2113)? in_data_i[456] : 
                          (N2115)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[391] = (N2112)? in_data_i[391] : 
                          (N2114)? in_data_i[423] : 
                          (N2113)? in_data_i[455] : 
                          (N2115)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[390] = (N2112)? in_data_i[390] : 
                          (N2114)? in_data_i[422] : 
                          (N2113)? in_data_i[454] : 
                          (N2115)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[389] = (N2112)? in_data_i[389] : 
                          (N2114)? in_data_i[421] : 
                          (N2113)? in_data_i[453] : 
                          (N2115)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[388] = (N2112)? in_data_i[388] : 
                          (N2114)? in_data_i[420] : 
                          (N2113)? in_data_i[452] : 
                          (N2115)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[387] = (N2112)? in_data_i[387] : 
                          (N2114)? in_data_i[419] : 
                          (N2113)? in_data_i[451] : 
                          (N2115)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[386] = (N2112)? in_data_i[386] : 
                          (N2114)? in_data_i[418] : 
                          (N2113)? in_data_i[450] : 
                          (N2115)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[385] = (N2112)? in_data_i[385] : 
                          (N2114)? in_data_i[417] : 
                          (N2113)? in_data_i[449] : 
                          (N2115)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[384] = (N2112)? in_data_i[384] : 
                          (N2114)? in_data_i[416] : 
                          (N2113)? in_data_i[448] : 
                          (N2115)? in_data_i_15__0_ : 1'b0;
  assign out_me_v_o[12] = (N2128)? out_me_v_i[0] : 
                          (N2130)? out_me_v_i[1] : 
                          (N2132)? out_me_v_i[2] : 
                          (N2134)? out_me_v_i[3] : 
                          (N2136)? out_me_v_i[4] : 
                          (N2138)? out_me_v_i[5] : 
                          (N2140)? out_me_v_i[6] : 
                          (N2142)? out_me_v_i[7] : 
                          (N2129)? out_me_v_i[8] : 
                          (N2131)? out_me_v_i[9] : 
                          (N2133)? out_me_v_i[10] : 
                          (N2135)? out_me_v_i[11] : 
                          (N2137)? out_me_v_i[12] : 
                          (N2139)? out_me_v_i[13] : 
                          (N2141)? out_me_v_i[14] : 
                          (N2143)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[12] = (N2160)? out_me_ready_i[0] : 
                              (N2162)? out_me_ready_i[1] : 
                              (N2164)? out_me_ready_i[2] : 
                              (N2166)? out_me_ready_i[3] : 
                              (N2168)? out_me_ready_i[4] : 
                              (N2170)? out_me_ready_i[5] : 
                              (N2172)? out_me_ready_i[6] : 
                              (N2174)? out_me_ready_i[7] : 
                              (N2161)? out_me_ready_i[8] : 
                              (N2163)? out_me_ready_i[9] : 
                              (N2165)? out_me_ready_i[10] : 
                              (N2167)? out_me_ready_i[11] : 
                              (N2169)? out_me_ready_i[12] : 
                              (N2171)? out_me_ready_i[13] : 
                              (N2173)? out_me_ready_i[14] : 
                              (N2175)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[13] = (N2221)? in_yumi_i[0] : 
                         (N2223)? in_yumi_i[1] : 
                         (N2225)? in_yumi_i[2] : 
                         (N2227)? in_yumi_i[3] : 
                         (N2229)? in_yumi_i[4] : 
                         (N2231)? in_yumi_i[5] : 
                         (N2233)? in_yumi_i[6] : 
                         (N2235)? in_yumi_i[7] : 
                         (N2222)? in_yumi_i[8] : 
                         (N2224)? in_yumi_i[9] : 
                         (N2226)? in_yumi_i[10] : 
                         (N2228)? in_yumi_i[11] : 
                         (N2230)? in_yumi_i[12] : 
                         (N2232)? in_yumi_i[13] : 
                         (N2234)? in_yumi_i[14] : 
                         (N2236)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[13] = (N2250)? out_me_v_i[0] : 
                          (N2252)? out_me_v_i[1] : 
                          (N2254)? out_me_v_i[2] : 
                          (N2256)? out_me_v_i[3] : 
                          (N2258)? out_me_v_i[4] : 
                          (N2260)? out_me_v_i[5] : 
                          (N2262)? out_me_v_i[6] : 
                          (N2264)? out_me_v_i[7] : 
                          (N2251)? out_me_v_i[8] : 
                          (N2253)? out_me_v_i[9] : 
                          (N2255)? out_me_v_i[10] : 
                          (N2257)? out_me_v_i[11] : 
                          (N2259)? out_me_v_i[12] : 
                          (N2261)? out_me_v_i[13] : 
                          (N2263)? out_me_v_i[14] : 
                          (N2265)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[13] = (N2282)? out_me_ready_i[0] : 
                              (N2284)? out_me_ready_i[1] : 
                              (N2286)? out_me_ready_i[2] : 
                              (N2288)? out_me_ready_i[3] : 
                              (N2290)? out_me_ready_i[4] : 
                              (N2292)? out_me_ready_i[5] : 
                              (N2294)? out_me_ready_i[6] : 
                              (N2296)? out_me_ready_i[7] : 
                              (N2283)? out_me_ready_i[8] : 
                              (N2285)? out_me_ready_i[9] : 
                              (N2287)? out_me_ready_i[10] : 
                              (N2289)? out_me_ready_i[11] : 
                              (N2291)? out_me_ready_i[12] : 
                              (N2293)? out_me_ready_i[13] : 
                              (N2295)? out_me_ready_i[14] : 
                              (N2297)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[14] = (N2344)? in_yumi_i[0] : 
                         (N2346)? in_yumi_i[1] : 
                         (N2348)? in_yumi_i[2] : 
                         (N2350)? in_yumi_i[3] : 
                         (N2352)? in_yumi_i[4] : 
                         (N2354)? in_yumi_i[5] : 
                         (N2356)? in_yumi_i[6] : 
                         (N2358)? in_yumi_i[7] : 
                         (N2345)? in_yumi_i[8] : 
                         (N2347)? in_yumi_i[9] : 
                         (N2349)? in_yumi_i[10] : 
                         (N2351)? in_yumi_i[11] : 
                         (N2353)? in_yumi_i[12] : 
                         (N2355)? in_yumi_i[13] : 
                         (N2357)? in_yumi_i[14] : 
                         (N2359)? in_yumi_i[15] : 1'b0;
  assign in_data_o[479] = (N2360)? in_data_i[479] : 
                          (N1)? in_data_i_15__31_ : 1'b0;
  assign N1 = fwd_dpath_sel_r_56;
  assign in_data_o[478] = (N2360)? in_data_i[478] : 
                          (N1)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[477] = (N2360)? in_data_i[477] : 
                          (N1)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[476] = (N2360)? in_data_i[476] : 
                          (N1)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[475] = (N2360)? in_data_i[475] : 
                          (N1)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[474] = (N2360)? in_data_i[474] : 
                          (N1)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[473] = (N2360)? in_data_i[473] : 
                          (N1)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[472] = (N2360)? in_data_i[472] : 
                          (N1)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[471] = (N2360)? in_data_i[471] : 
                          (N1)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[470] = (N2360)? in_data_i[470] : 
                          (N1)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[469] = (N2360)? in_data_i[469] : 
                          (N1)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[468] = (N2360)? in_data_i[468] : 
                          (N1)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[467] = (N2360)? in_data_i[467] : 
                          (N1)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[466] = (N2360)? in_data_i[466] : 
                          (N1)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[465] = (N2360)? in_data_i[465] : 
                          (N1)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[464] = (N2360)? in_data_i[464] : 
                          (N1)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[463] = (N2360)? in_data_i[463] : 
                          (N1)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[462] = (N2360)? in_data_i[462] : 
                          (N1)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[461] = (N2360)? in_data_i[461] : 
                          (N1)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[460] = (N2360)? in_data_i[460] : 
                          (N1)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[459] = (N2360)? in_data_i[459] : 
                          (N1)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[458] = (N2360)? in_data_i[458] : 
                          (N1)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[457] = (N2360)? in_data_i[457] : 
                          (N1)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[456] = (N2360)? in_data_i[456] : 
                          (N1)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[455] = (N2360)? in_data_i[455] : 
                          (N1)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[454] = (N2360)? in_data_i[454] : 
                          (N1)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[453] = (N2360)? in_data_i[453] : 
                          (N1)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[452] = (N2360)? in_data_i[452] : 
                          (N1)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[451] = (N2360)? in_data_i[451] : 
                          (N1)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[450] = (N2360)? in_data_i[450] : 
                          (N1)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[449] = (N2360)? in_data_i[449] : 
                          (N1)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[448] = (N2360)? in_data_i[448] : 
                          (N1)? in_data_i_15__0_ : 1'b0;
  assign out_me_v_o[14] = (N2373)? out_me_v_i[0] : 
                          (N2375)? out_me_v_i[1] : 
                          (N2377)? out_me_v_i[2] : 
                          (N2379)? out_me_v_i[3] : 
                          (N2381)? out_me_v_i[4] : 
                          (N2383)? out_me_v_i[5] : 
                          (N2385)? out_me_v_i[6] : 
                          (N2387)? out_me_v_i[7] : 
                          (N2374)? out_me_v_i[8] : 
                          (N2376)? out_me_v_i[9] : 
                          (N2378)? out_me_v_i[10] : 
                          (N2380)? out_me_v_i[11] : 
                          (N2382)? out_me_v_i[12] : 
                          (N2384)? out_me_v_i[13] : 
                          (N2386)? out_me_v_i[14] : 
                          (N2388)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[14] = (N2405)? out_me_ready_i[0] : 
                              (N2407)? out_me_ready_i[1] : 
                              (N2409)? out_me_ready_i[2] : 
                              (N2411)? out_me_ready_i[3] : 
                              (N2413)? out_me_ready_i[4] : 
                              (N2415)? out_me_ready_i[5] : 
                              (N2417)? out_me_ready_i[6] : 
                              (N2419)? out_me_ready_i[7] : 
                              (N2406)? out_me_ready_i[8] : 
                              (N2408)? out_me_ready_i[9] : 
                              (N2410)? out_me_ready_i[10] : 
                              (N2412)? out_me_ready_i[11] : 
                              (N2414)? out_me_ready_i[12] : 
                              (N2416)? out_me_ready_i[13] : 
                              (N2418)? out_me_ready_i[14] : 
                              (N2420)? out_me_ready_i[15] : 1'b0;
  assign in_yumi_o[15] = (N2468)? in_yumi_i[0] : 
                         (N2470)? in_yumi_i[1] : 
                         (N2472)? in_yumi_i[2] : 
                         (N2474)? in_yumi_i[3] : 
                         (N2476)? in_yumi_i[4] : 
                         (N2478)? in_yumi_i[5] : 
                         (N2480)? in_yumi_i[6] : 
                         (N2482)? in_yumi_i[7] : 
                         (N2469)? in_yumi_i[8] : 
                         (N2471)? in_yumi_i[9] : 
                         (N2473)? in_yumi_i[10] : 
                         (N2475)? in_yumi_i[11] : 
                         (N2477)? in_yumi_i[12] : 
                         (N2479)? in_yumi_i[13] : 
                         (N2481)? in_yumi_i[14] : 
                         (N2483)? in_yumi_i[15] : 1'b0;
  assign out_me_v_o[15] = (N2496)? out_me_v_i[0] : 
                          (N2498)? out_me_v_i[1] : 
                          (N2500)? out_me_v_i[2] : 
                          (N2502)? out_me_v_i[3] : 
                          (N2504)? out_me_v_i[4] : 
                          (N2506)? out_me_v_i[5] : 
                          (N2508)? out_me_v_i[6] : 
                          (N2510)? out_me_v_i[7] : 
                          (N2497)? out_me_v_i[8] : 
                          (N2499)? out_me_v_i[9] : 
                          (N2501)? out_me_v_i[10] : 
                          (N2503)? out_me_v_i[11] : 
                          (N2505)? out_me_v_i[12] : 
                          (N2507)? out_me_v_i[13] : 
                          (N2509)? out_me_v_i[14] : 
                          (N2511)? out_me_v_i[15] : 1'b0;
  assign out_me_ready_o[15] = (N2528)? out_me_ready_i[0] : 
                              (N2530)? out_me_ready_i[1] : 
                              (N2532)? out_me_ready_i[2] : 
                              (N2534)? out_me_ready_i[3] : 
                              (N2536)? out_me_ready_i[4] : 
                              (N2538)? out_me_ready_i[5] : 
                              (N2540)? out_me_ready_i[6] : 
                              (N2542)? out_me_ready_i[7] : 
                              (N2529)? out_me_ready_i[8] : 
                              (N2531)? out_me_ready_i[9] : 
                              (N2533)? out_me_ready_i[10] : 
                              (N2535)? out_me_ready_i[11] : 
                              (N2537)? out_me_ready_i[12] : 
                              (N2539)? out_me_ready_i[13] : 
                              (N2541)? out_me_ready_i[14] : 
                              (N2543)? out_me_ready_i[15] : 1'b0;
  assign out_me_data_o[511] = (N2560)? out_me_data_i_0__31_ : 
                              (N2562)? out_me_data_i[63] : 
                              (N2564)? out_me_data_i[95] : 
                              (N2566)? out_me_data_i[127] : 
                              (N2568)? out_me_data_i[159] : 
                              (N2570)? out_me_data_i[191] : 
                              (N2572)? out_me_data_i[223] : 
                              (N2574)? out_me_data_i[255] : 
                              (N2561)? out_me_data_i[287] : 
                              (N2563)? out_me_data_i[319] : 
                              (N2565)? out_me_data_i[351] : 
                              (N2567)? out_me_data_i[383] : 
                              (N2569)? out_me_data_i[415] : 
                              (N2571)? out_me_data_i[447] : 
                              (N2573)? out_me_data_i[479] : 
                              (N2575)? out_me_data_i[511] : 1'b0;
  assign out_me_data_o[510] = (N2560)? out_me_data_i_0__30_ : 
                              (N2562)? out_me_data_i[62] : 
                              (N2564)? out_me_data_i[94] : 
                              (N2566)? out_me_data_i[126] : 
                              (N2568)? out_me_data_i[158] : 
                              (N2570)? out_me_data_i[190] : 
                              (N2572)? out_me_data_i[222] : 
                              (N2574)? out_me_data_i[254] : 
                              (N2561)? out_me_data_i[286] : 
                              (N2563)? out_me_data_i[318] : 
                              (N2565)? out_me_data_i[350] : 
                              (N2567)? out_me_data_i[382] : 
                              (N2569)? out_me_data_i[414] : 
                              (N2571)? out_me_data_i[446] : 
                              (N2573)? out_me_data_i[478] : 
                              (N2575)? out_me_data_i[510] : 1'b0;
  assign out_me_data_o[509] = (N2560)? out_me_data_i_0__29_ : 
                              (N2562)? out_me_data_i[61] : 
                              (N2564)? out_me_data_i[93] : 
                              (N2566)? out_me_data_i[125] : 
                              (N2568)? out_me_data_i[157] : 
                              (N2570)? out_me_data_i[189] : 
                              (N2572)? out_me_data_i[221] : 
                              (N2574)? out_me_data_i[253] : 
                              (N2561)? out_me_data_i[285] : 
                              (N2563)? out_me_data_i[317] : 
                              (N2565)? out_me_data_i[349] : 
                              (N2567)? out_me_data_i[381] : 
                              (N2569)? out_me_data_i[413] : 
                              (N2571)? out_me_data_i[445] : 
                              (N2573)? out_me_data_i[477] : 
                              (N2575)? out_me_data_i[509] : 1'b0;
  assign out_me_data_o[508] = (N2560)? out_me_data_i_0__28_ : 
                              (N2562)? out_me_data_i[60] : 
                              (N2564)? out_me_data_i[92] : 
                              (N2566)? out_me_data_i[124] : 
                              (N2568)? out_me_data_i[156] : 
                              (N2570)? out_me_data_i[188] : 
                              (N2572)? out_me_data_i[220] : 
                              (N2574)? out_me_data_i[252] : 
                              (N2561)? out_me_data_i[284] : 
                              (N2563)? out_me_data_i[316] : 
                              (N2565)? out_me_data_i[348] : 
                              (N2567)? out_me_data_i[380] : 
                              (N2569)? out_me_data_i[412] : 
                              (N2571)? out_me_data_i[444] : 
                              (N2573)? out_me_data_i[476] : 
                              (N2575)? out_me_data_i[508] : 1'b0;
  assign out_me_data_o[507] = (N2560)? out_me_data_i_0__27_ : 
                              (N2562)? out_me_data_i[59] : 
                              (N2564)? out_me_data_i[91] : 
                              (N2566)? out_me_data_i[123] : 
                              (N2568)? out_me_data_i[155] : 
                              (N2570)? out_me_data_i[187] : 
                              (N2572)? out_me_data_i[219] : 
                              (N2574)? out_me_data_i[251] : 
                              (N2561)? out_me_data_i[283] : 
                              (N2563)? out_me_data_i[315] : 
                              (N2565)? out_me_data_i[347] : 
                              (N2567)? out_me_data_i[379] : 
                              (N2569)? out_me_data_i[411] : 
                              (N2571)? out_me_data_i[443] : 
                              (N2573)? out_me_data_i[475] : 
                              (N2575)? out_me_data_i[507] : 1'b0;
  assign out_me_data_o[506] = (N2560)? out_me_data_i_0__26_ : 
                              (N2562)? out_me_data_i[58] : 
                              (N2564)? out_me_data_i[90] : 
                              (N2566)? out_me_data_i[122] : 
                              (N2568)? out_me_data_i[154] : 
                              (N2570)? out_me_data_i[186] : 
                              (N2572)? out_me_data_i[218] : 
                              (N2574)? out_me_data_i[250] : 
                              (N2561)? out_me_data_i[282] : 
                              (N2563)? out_me_data_i[314] : 
                              (N2565)? out_me_data_i[346] : 
                              (N2567)? out_me_data_i[378] : 
                              (N2569)? out_me_data_i[410] : 
                              (N2571)? out_me_data_i[442] : 
                              (N2573)? out_me_data_i[474] : 
                              (N2575)? out_me_data_i[506] : 1'b0;
  assign out_me_data_o[505] = (N2560)? out_me_data_i_0__25_ : 
                              (N2562)? out_me_data_i[57] : 
                              (N2564)? out_me_data_i[89] : 
                              (N2566)? out_me_data_i[121] : 
                              (N2568)? out_me_data_i[153] : 
                              (N2570)? out_me_data_i[185] : 
                              (N2572)? out_me_data_i[217] : 
                              (N2574)? out_me_data_i[249] : 
                              (N2561)? out_me_data_i[281] : 
                              (N2563)? out_me_data_i[313] : 
                              (N2565)? out_me_data_i[345] : 
                              (N2567)? out_me_data_i[377] : 
                              (N2569)? out_me_data_i[409] : 
                              (N2571)? out_me_data_i[441] : 
                              (N2573)? out_me_data_i[473] : 
                              (N2575)? out_me_data_i[505] : 1'b0;
  assign out_me_data_o[504] = (N2560)? out_me_data_i_0__24_ : 
                              (N2562)? out_me_data_i[56] : 
                              (N2564)? out_me_data_i[88] : 
                              (N2566)? out_me_data_i[120] : 
                              (N2568)? out_me_data_i[152] : 
                              (N2570)? out_me_data_i[184] : 
                              (N2572)? out_me_data_i[216] : 
                              (N2574)? out_me_data_i[248] : 
                              (N2561)? out_me_data_i[280] : 
                              (N2563)? out_me_data_i[312] : 
                              (N2565)? out_me_data_i[344] : 
                              (N2567)? out_me_data_i[376] : 
                              (N2569)? out_me_data_i[408] : 
                              (N2571)? out_me_data_i[440] : 
                              (N2573)? out_me_data_i[472] : 
                              (N2575)? out_me_data_i[504] : 1'b0;
  assign out_me_data_o[503] = (N2560)? out_me_data_i_0__23_ : 
                              (N2562)? out_me_data_i[55] : 
                              (N2564)? out_me_data_i[87] : 
                              (N2566)? out_me_data_i[119] : 
                              (N2568)? out_me_data_i[151] : 
                              (N2570)? out_me_data_i[183] : 
                              (N2572)? out_me_data_i[215] : 
                              (N2574)? out_me_data_i[247] : 
                              (N2561)? out_me_data_i[279] : 
                              (N2563)? out_me_data_i[311] : 
                              (N2565)? out_me_data_i[343] : 
                              (N2567)? out_me_data_i[375] : 
                              (N2569)? out_me_data_i[407] : 
                              (N2571)? out_me_data_i[439] : 
                              (N2573)? out_me_data_i[471] : 
                              (N2575)? out_me_data_i[503] : 1'b0;
  assign out_me_data_o[502] = (N2560)? out_me_data_i_0__22_ : 
                              (N2562)? out_me_data_i[54] : 
                              (N2564)? out_me_data_i[86] : 
                              (N2566)? out_me_data_i[118] : 
                              (N2568)? out_me_data_i[150] : 
                              (N2570)? out_me_data_i[182] : 
                              (N2572)? out_me_data_i[214] : 
                              (N2574)? out_me_data_i[246] : 
                              (N2561)? out_me_data_i[278] : 
                              (N2563)? out_me_data_i[310] : 
                              (N2565)? out_me_data_i[342] : 
                              (N2567)? out_me_data_i[374] : 
                              (N2569)? out_me_data_i[406] : 
                              (N2571)? out_me_data_i[438] : 
                              (N2573)? out_me_data_i[470] : 
                              (N2575)? out_me_data_i[502] : 1'b0;
  assign out_me_data_o[501] = (N2560)? out_me_data_i_0__21_ : 
                              (N2562)? out_me_data_i[53] : 
                              (N2564)? out_me_data_i[85] : 
                              (N2566)? out_me_data_i[117] : 
                              (N2568)? out_me_data_i[149] : 
                              (N2570)? out_me_data_i[181] : 
                              (N2572)? out_me_data_i[213] : 
                              (N2574)? out_me_data_i[245] : 
                              (N2561)? out_me_data_i[277] : 
                              (N2563)? out_me_data_i[309] : 
                              (N2565)? out_me_data_i[341] : 
                              (N2567)? out_me_data_i[373] : 
                              (N2569)? out_me_data_i[405] : 
                              (N2571)? out_me_data_i[437] : 
                              (N2573)? out_me_data_i[469] : 
                              (N2575)? out_me_data_i[501] : 1'b0;
  assign out_me_data_o[500] = (N2560)? out_me_data_i_0__20_ : 
                              (N2562)? out_me_data_i[52] : 
                              (N2564)? out_me_data_i[84] : 
                              (N2566)? out_me_data_i[116] : 
                              (N2568)? out_me_data_i[148] : 
                              (N2570)? out_me_data_i[180] : 
                              (N2572)? out_me_data_i[212] : 
                              (N2574)? out_me_data_i[244] : 
                              (N2561)? out_me_data_i[276] : 
                              (N2563)? out_me_data_i[308] : 
                              (N2565)? out_me_data_i[340] : 
                              (N2567)? out_me_data_i[372] : 
                              (N2569)? out_me_data_i[404] : 
                              (N2571)? out_me_data_i[436] : 
                              (N2573)? out_me_data_i[468] : 
                              (N2575)? out_me_data_i[500] : 1'b0;
  assign out_me_data_o[499] = (N2560)? out_me_data_i_0__19_ : 
                              (N2562)? out_me_data_i[51] : 
                              (N2564)? out_me_data_i[83] : 
                              (N2566)? out_me_data_i[115] : 
                              (N2568)? out_me_data_i[147] : 
                              (N2570)? out_me_data_i[179] : 
                              (N2572)? out_me_data_i[211] : 
                              (N2574)? out_me_data_i[243] : 
                              (N2561)? out_me_data_i[275] : 
                              (N2563)? out_me_data_i[307] : 
                              (N2565)? out_me_data_i[339] : 
                              (N2567)? out_me_data_i[371] : 
                              (N2569)? out_me_data_i[403] : 
                              (N2571)? out_me_data_i[435] : 
                              (N2573)? out_me_data_i[467] : 
                              (N2575)? out_me_data_i[499] : 1'b0;
  assign out_me_data_o[498] = (N2560)? out_me_data_i_0__18_ : 
                              (N2562)? out_me_data_i[50] : 
                              (N2564)? out_me_data_i[82] : 
                              (N2566)? out_me_data_i[114] : 
                              (N2568)? out_me_data_i[146] : 
                              (N2570)? out_me_data_i[178] : 
                              (N2572)? out_me_data_i[210] : 
                              (N2574)? out_me_data_i[242] : 
                              (N2561)? out_me_data_i[274] : 
                              (N2563)? out_me_data_i[306] : 
                              (N2565)? out_me_data_i[338] : 
                              (N2567)? out_me_data_i[370] : 
                              (N2569)? out_me_data_i[402] : 
                              (N2571)? out_me_data_i[434] : 
                              (N2573)? out_me_data_i[466] : 
                              (N2575)? out_me_data_i[498] : 1'b0;
  assign out_me_data_o[497] = (N2560)? out_me_data_i_0__17_ : 
                              (N2562)? out_me_data_i[49] : 
                              (N2564)? out_me_data_i[81] : 
                              (N2566)? out_me_data_i[113] : 
                              (N2568)? out_me_data_i[145] : 
                              (N2570)? out_me_data_i[177] : 
                              (N2572)? out_me_data_i[209] : 
                              (N2574)? out_me_data_i[241] : 
                              (N2561)? out_me_data_i[273] : 
                              (N2563)? out_me_data_i[305] : 
                              (N2565)? out_me_data_i[337] : 
                              (N2567)? out_me_data_i[369] : 
                              (N2569)? out_me_data_i[401] : 
                              (N2571)? out_me_data_i[433] : 
                              (N2573)? out_me_data_i[465] : 
                              (N2575)? out_me_data_i[497] : 1'b0;
  assign out_me_data_o[496] = (N2560)? out_me_data_i_0__16_ : 
                              (N2562)? out_me_data_i[48] : 
                              (N2564)? out_me_data_i[80] : 
                              (N2566)? out_me_data_i[112] : 
                              (N2568)? out_me_data_i[144] : 
                              (N2570)? out_me_data_i[176] : 
                              (N2572)? out_me_data_i[208] : 
                              (N2574)? out_me_data_i[240] : 
                              (N2561)? out_me_data_i[272] : 
                              (N2563)? out_me_data_i[304] : 
                              (N2565)? out_me_data_i[336] : 
                              (N2567)? out_me_data_i[368] : 
                              (N2569)? out_me_data_i[400] : 
                              (N2571)? out_me_data_i[432] : 
                              (N2573)? out_me_data_i[464] : 
                              (N2575)? out_me_data_i[496] : 1'b0;
  assign out_me_data_o[495] = (N2560)? out_me_data_i_0__15_ : 
                              (N2562)? out_me_data_i[47] : 
                              (N2564)? out_me_data_i[79] : 
                              (N2566)? out_me_data_i[111] : 
                              (N2568)? out_me_data_i[143] : 
                              (N2570)? out_me_data_i[175] : 
                              (N2572)? out_me_data_i[207] : 
                              (N2574)? out_me_data_i[239] : 
                              (N2561)? out_me_data_i[271] : 
                              (N2563)? out_me_data_i[303] : 
                              (N2565)? out_me_data_i[335] : 
                              (N2567)? out_me_data_i[367] : 
                              (N2569)? out_me_data_i[399] : 
                              (N2571)? out_me_data_i[431] : 
                              (N2573)? out_me_data_i[463] : 
                              (N2575)? out_me_data_i[495] : 1'b0;
  assign out_me_data_o[494] = (N2560)? out_me_data_i_0__14_ : 
                              (N2562)? out_me_data_i[46] : 
                              (N2564)? out_me_data_i[78] : 
                              (N2566)? out_me_data_i[110] : 
                              (N2568)? out_me_data_i[142] : 
                              (N2570)? out_me_data_i[174] : 
                              (N2572)? out_me_data_i[206] : 
                              (N2574)? out_me_data_i[238] : 
                              (N2561)? out_me_data_i[270] : 
                              (N2563)? out_me_data_i[302] : 
                              (N2565)? out_me_data_i[334] : 
                              (N2567)? out_me_data_i[366] : 
                              (N2569)? out_me_data_i[398] : 
                              (N2571)? out_me_data_i[430] : 
                              (N2573)? out_me_data_i[462] : 
                              (N2575)? out_me_data_i[494] : 1'b0;
  assign out_me_data_o[493] = (N2560)? out_me_data_i_0__13_ : 
                              (N2562)? out_me_data_i[45] : 
                              (N2564)? out_me_data_i[77] : 
                              (N2566)? out_me_data_i[109] : 
                              (N2568)? out_me_data_i[141] : 
                              (N2570)? out_me_data_i[173] : 
                              (N2572)? out_me_data_i[205] : 
                              (N2574)? out_me_data_i[237] : 
                              (N2561)? out_me_data_i[269] : 
                              (N2563)? out_me_data_i[301] : 
                              (N2565)? out_me_data_i[333] : 
                              (N2567)? out_me_data_i[365] : 
                              (N2569)? out_me_data_i[397] : 
                              (N2571)? out_me_data_i[429] : 
                              (N2573)? out_me_data_i[461] : 
                              (N2575)? out_me_data_i[493] : 1'b0;
  assign out_me_data_o[492] = (N2560)? out_me_data_i_0__12_ : 
                              (N2562)? out_me_data_i[44] : 
                              (N2564)? out_me_data_i[76] : 
                              (N2566)? out_me_data_i[108] : 
                              (N2568)? out_me_data_i[140] : 
                              (N2570)? out_me_data_i[172] : 
                              (N2572)? out_me_data_i[204] : 
                              (N2574)? out_me_data_i[236] : 
                              (N2561)? out_me_data_i[268] : 
                              (N2563)? out_me_data_i[300] : 
                              (N2565)? out_me_data_i[332] : 
                              (N2567)? out_me_data_i[364] : 
                              (N2569)? out_me_data_i[396] : 
                              (N2571)? out_me_data_i[428] : 
                              (N2573)? out_me_data_i[460] : 
                              (N2575)? out_me_data_i[492] : 1'b0;
  assign out_me_data_o[491] = (N2560)? out_me_data_i_0__11_ : 
                              (N2562)? out_me_data_i[43] : 
                              (N2564)? out_me_data_i[75] : 
                              (N2566)? out_me_data_i[107] : 
                              (N2568)? out_me_data_i[139] : 
                              (N2570)? out_me_data_i[171] : 
                              (N2572)? out_me_data_i[203] : 
                              (N2574)? out_me_data_i[235] : 
                              (N2561)? out_me_data_i[267] : 
                              (N2563)? out_me_data_i[299] : 
                              (N2565)? out_me_data_i[331] : 
                              (N2567)? out_me_data_i[363] : 
                              (N2569)? out_me_data_i[395] : 
                              (N2571)? out_me_data_i[427] : 
                              (N2573)? out_me_data_i[459] : 
                              (N2575)? out_me_data_i[491] : 1'b0;
  assign out_me_data_o[490] = (N2560)? out_me_data_i_0__10_ : 
                              (N2562)? out_me_data_i[42] : 
                              (N2564)? out_me_data_i[74] : 
                              (N2566)? out_me_data_i[106] : 
                              (N2568)? out_me_data_i[138] : 
                              (N2570)? out_me_data_i[170] : 
                              (N2572)? out_me_data_i[202] : 
                              (N2574)? out_me_data_i[234] : 
                              (N2561)? out_me_data_i[266] : 
                              (N2563)? out_me_data_i[298] : 
                              (N2565)? out_me_data_i[330] : 
                              (N2567)? out_me_data_i[362] : 
                              (N2569)? out_me_data_i[394] : 
                              (N2571)? out_me_data_i[426] : 
                              (N2573)? out_me_data_i[458] : 
                              (N2575)? out_me_data_i[490] : 1'b0;
  assign out_me_data_o[489] = (N2560)? out_me_data_i_0__9_ : 
                              (N2562)? out_me_data_i[41] : 
                              (N2564)? out_me_data_i[73] : 
                              (N2566)? out_me_data_i[105] : 
                              (N2568)? out_me_data_i[137] : 
                              (N2570)? out_me_data_i[169] : 
                              (N2572)? out_me_data_i[201] : 
                              (N2574)? out_me_data_i[233] : 
                              (N2561)? out_me_data_i[265] : 
                              (N2563)? out_me_data_i[297] : 
                              (N2565)? out_me_data_i[329] : 
                              (N2567)? out_me_data_i[361] : 
                              (N2569)? out_me_data_i[393] : 
                              (N2571)? out_me_data_i[425] : 
                              (N2573)? out_me_data_i[457] : 
                              (N2575)? out_me_data_i[489] : 1'b0;
  assign out_me_data_o[488] = (N2560)? out_me_data_i_0__8_ : 
                              (N2562)? out_me_data_i[40] : 
                              (N2564)? out_me_data_i[72] : 
                              (N2566)? out_me_data_i[104] : 
                              (N2568)? out_me_data_i[136] : 
                              (N2570)? out_me_data_i[168] : 
                              (N2572)? out_me_data_i[200] : 
                              (N2574)? out_me_data_i[232] : 
                              (N2561)? out_me_data_i[264] : 
                              (N2563)? out_me_data_i[296] : 
                              (N2565)? out_me_data_i[328] : 
                              (N2567)? out_me_data_i[360] : 
                              (N2569)? out_me_data_i[392] : 
                              (N2571)? out_me_data_i[424] : 
                              (N2573)? out_me_data_i[456] : 
                              (N2575)? out_me_data_i[488] : 1'b0;
  assign out_me_data_o[487] = (N2560)? out_me_data_i_0__7_ : 
                              (N2562)? out_me_data_i[39] : 
                              (N2564)? out_me_data_i[71] : 
                              (N2566)? out_me_data_i[103] : 
                              (N2568)? out_me_data_i[135] : 
                              (N2570)? out_me_data_i[167] : 
                              (N2572)? out_me_data_i[199] : 
                              (N2574)? out_me_data_i[231] : 
                              (N2561)? out_me_data_i[263] : 
                              (N2563)? out_me_data_i[295] : 
                              (N2565)? out_me_data_i[327] : 
                              (N2567)? out_me_data_i[359] : 
                              (N2569)? out_me_data_i[391] : 
                              (N2571)? out_me_data_i[423] : 
                              (N2573)? out_me_data_i[455] : 
                              (N2575)? out_me_data_i[487] : 1'b0;
  assign out_me_data_o[486] = (N2560)? out_me_data_i_0__6_ : 
                              (N2562)? out_me_data_i[38] : 
                              (N2564)? out_me_data_i[70] : 
                              (N2566)? out_me_data_i[102] : 
                              (N2568)? out_me_data_i[134] : 
                              (N2570)? out_me_data_i[166] : 
                              (N2572)? out_me_data_i[198] : 
                              (N2574)? out_me_data_i[230] : 
                              (N2561)? out_me_data_i[262] : 
                              (N2563)? out_me_data_i[294] : 
                              (N2565)? out_me_data_i[326] : 
                              (N2567)? out_me_data_i[358] : 
                              (N2569)? out_me_data_i[390] : 
                              (N2571)? out_me_data_i[422] : 
                              (N2573)? out_me_data_i[454] : 
                              (N2575)? out_me_data_i[486] : 1'b0;
  assign out_me_data_o[485] = (N2560)? out_me_data_i_0__5_ : 
                              (N2562)? out_me_data_i[37] : 
                              (N2564)? out_me_data_i[69] : 
                              (N2566)? out_me_data_i[101] : 
                              (N2568)? out_me_data_i[133] : 
                              (N2570)? out_me_data_i[165] : 
                              (N2572)? out_me_data_i[197] : 
                              (N2574)? out_me_data_i[229] : 
                              (N2561)? out_me_data_i[261] : 
                              (N2563)? out_me_data_i[293] : 
                              (N2565)? out_me_data_i[325] : 
                              (N2567)? out_me_data_i[357] : 
                              (N2569)? out_me_data_i[389] : 
                              (N2571)? out_me_data_i[421] : 
                              (N2573)? out_me_data_i[453] : 
                              (N2575)? out_me_data_i[485] : 1'b0;
  assign out_me_data_o[484] = (N2560)? out_me_data_i_0__4_ : 
                              (N2562)? out_me_data_i[36] : 
                              (N2564)? out_me_data_i[68] : 
                              (N2566)? out_me_data_i[100] : 
                              (N2568)? out_me_data_i[132] : 
                              (N2570)? out_me_data_i[164] : 
                              (N2572)? out_me_data_i[196] : 
                              (N2574)? out_me_data_i[228] : 
                              (N2561)? out_me_data_i[260] : 
                              (N2563)? out_me_data_i[292] : 
                              (N2565)? out_me_data_i[324] : 
                              (N2567)? out_me_data_i[356] : 
                              (N2569)? out_me_data_i[388] : 
                              (N2571)? out_me_data_i[420] : 
                              (N2573)? out_me_data_i[452] : 
                              (N2575)? out_me_data_i[484] : 1'b0;
  assign out_me_data_o[483] = (N2560)? out_me_data_i_0__3_ : 
                              (N2562)? out_me_data_i[35] : 
                              (N2564)? out_me_data_i[67] : 
                              (N2566)? out_me_data_i[99] : 
                              (N2568)? out_me_data_i[131] : 
                              (N2570)? out_me_data_i[163] : 
                              (N2572)? out_me_data_i[195] : 
                              (N2574)? out_me_data_i[227] : 
                              (N2561)? out_me_data_i[259] : 
                              (N2563)? out_me_data_i[291] : 
                              (N2565)? out_me_data_i[323] : 
                              (N2567)? out_me_data_i[355] : 
                              (N2569)? out_me_data_i[387] : 
                              (N2571)? out_me_data_i[419] : 
                              (N2573)? out_me_data_i[451] : 
                              (N2575)? out_me_data_i[483] : 1'b0;
  assign out_me_data_o[482] = (N2560)? out_me_data_i_0__2_ : 
                              (N2562)? out_me_data_i[34] : 
                              (N2564)? out_me_data_i[66] : 
                              (N2566)? out_me_data_i[98] : 
                              (N2568)? out_me_data_i[130] : 
                              (N2570)? out_me_data_i[162] : 
                              (N2572)? out_me_data_i[194] : 
                              (N2574)? out_me_data_i[226] : 
                              (N2561)? out_me_data_i[258] : 
                              (N2563)? out_me_data_i[290] : 
                              (N2565)? out_me_data_i[322] : 
                              (N2567)? out_me_data_i[354] : 
                              (N2569)? out_me_data_i[386] : 
                              (N2571)? out_me_data_i[418] : 
                              (N2573)? out_me_data_i[450] : 
                              (N2575)? out_me_data_i[482] : 1'b0;
  assign out_me_data_o[481] = (N2560)? out_me_data_i_0__1_ : 
                              (N2562)? out_me_data_i[33] : 
                              (N2564)? out_me_data_i[65] : 
                              (N2566)? out_me_data_i[97] : 
                              (N2568)? out_me_data_i[129] : 
                              (N2570)? out_me_data_i[161] : 
                              (N2572)? out_me_data_i[193] : 
                              (N2574)? out_me_data_i[225] : 
                              (N2561)? out_me_data_i[257] : 
                              (N2563)? out_me_data_i[289] : 
                              (N2565)? out_me_data_i[321] : 
                              (N2567)? out_me_data_i[353] : 
                              (N2569)? out_me_data_i[385] : 
                              (N2571)? out_me_data_i[417] : 
                              (N2573)? out_me_data_i[449] : 
                              (N2575)? out_me_data_i[481] : 1'b0;
  assign out_me_data_o[480] = (N2560)? out_me_data_i_0__0_ : 
                              (N2562)? out_me_data_i[32] : 
                              (N2564)? out_me_data_i[64] : 
                              (N2566)? out_me_data_i[96] : 
                              (N2568)? out_me_data_i[128] : 
                              (N2570)? out_me_data_i[160] : 
                              (N2572)? out_me_data_i[192] : 
                              (N2574)? out_me_data_i[224] : 
                              (N2561)? out_me_data_i[256] : 
                              (N2563)? out_me_data_i[288] : 
                              (N2565)? out_me_data_i[320] : 
                              (N2567)? out_me_data_i[352] : 
                              (N2569)? out_me_data_i[384] : 
                              (N2571)? out_me_data_i[416] : 
                              (N2573)? out_me_data_i[448] : 
                              (N2575)? out_me_data_i[480] : 1'b0;
  assign { N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[3:0];
  assign { N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[7:4];
  assign { N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[11:8];
  assign { N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[15:12];
  assign { N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[19:16];
  assign { N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[23:20];
  assign { N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[27:24];
  assign { N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[31:28];
  assign { N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[35:32];
  assign { N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[39:36];
  assign { N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[43:40];
  assign { N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[47:44];
  assign { N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[51:48];
  assign { N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[55:52];
  assign { N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[59:56];
  assign { N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << fwd_sel[63:60];
  assign N2237 = N2 & N3;
  assign N2 = ~fwd_dpath_sel_r_52;
  assign N3 = ~fwd_dpath_sel_r_53;
  assign N924 = N4 & N5;
  assign N4 = ~bk_dpath_sel_r_8;
  assign N5 = ~bk_dpath_sel_r_9;
  assign N1986 = N6 & N7 & N8;
  assign N6 = ~fwd_dpath_sel_r_46;
  assign N7 = ~fwd_dpath_sel_r_44;
  assign N8 = ~fwd_dpath_sel_r_45;
  assign N1987 = fwd_dpath_sel_r_44 & N9;
  assign N9 = ~fwd_dpath_sel_r_45;
  assign N1988 = N10 & fwd_dpath_sel_r_45;
  assign N10 = ~fwd_dpath_sel_r_44;
  assign N1989 = fwd_dpath_sel_r_44 & fwd_dpath_sel_r_45;
  assign N1861 = N11 & N12 & N13;
  assign N11 = ~fwd_dpath_sel_r_42;
  assign N12 = ~fwd_dpath_sel_r_40;
  assign N13 = ~fwd_dpath_sel_r_41;
  assign N1862 = fwd_dpath_sel_r_42 & N14;
  assign N14 = ~fwd_dpath_sel_r_40;
  assign N1863 = N15 & fwd_dpath_sel_r_40 & N16;
  assign N15 = ~fwd_dpath_sel_r_42;
  assign N16 = ~fwd_dpath_sel_r_41;
  assign N1865 = N17 & fwd_dpath_sel_r_41;
  assign N17 = ~fwd_dpath_sel_r_40;
  assign N1866 = fwd_dpath_sel_r_40 & fwd_dpath_sel_r_41;
  assign N1864 = fwd_dpath_sel_r_42 & fwd_dpath_sel_r_40;
  assign N1736 = N18 & N19 & N20;
  assign N18 = ~fwd_dpath_sel_r_38;
  assign N19 = ~fwd_dpath_sel_r_36;
  assign N20 = ~fwd_dpath_sel_r_37;
  assign N1737 = fwd_dpath_sel_r_38 & N21 & N22;
  assign N21 = ~fwd_dpath_sel_r_36;
  assign N22 = ~fwd_dpath_sel_r_37;
  assign N1738 = N23 & fwd_dpath_sel_r_36 & N24;
  assign N23 = ~fwd_dpath_sel_r_38;
  assign N24 = ~fwd_dpath_sel_r_37;
  assign N1740 = N25 & N26 & fwd_dpath_sel_r_37;
  assign N25 = ~fwd_dpath_sel_r_38;
  assign N26 = ~fwd_dpath_sel_r_36;
  assign N1742 = fwd_dpath_sel_r_36 & fwd_dpath_sel_r_37;
  assign N1739 = fwd_dpath_sel_r_38 & fwd_dpath_sel_r_36;
  assign N1741 = fwd_dpath_sel_r_38 & fwd_dpath_sel_r_37;
  assign N1419 = N27 & N28 & N29;
  assign N27 = ~bk_dpath_sel_r_26;
  assign N28 = ~bk_dpath_sel_r_24;
  assign N29 = ~bk_dpath_sel_r_25;
  assign N1420 = bk_dpath_sel_r_26 & N30 & N31;
  assign N30 = ~bk_dpath_sel_r_24;
  assign N31 = ~bk_dpath_sel_r_25;
  assign N1421 = N32 & bk_dpath_sel_r_24 & N33;
  assign N32 = ~bk_dpath_sel_r_26;
  assign N33 = ~bk_dpath_sel_r_25;
  assign N1423 = N34 & N35 & bk_dpath_sel_r_25;
  assign N34 = ~bk_dpath_sel_r_26;
  assign N35 = ~bk_dpath_sel_r_24;
  assign N1425 = bk_dpath_sel_r_24 & bk_dpath_sel_r_25;
  assign N1422 = bk_dpath_sel_r_26 & bk_dpath_sel_r_24;
  assign N1424 = bk_dpath_sel_r_26 & bk_dpath_sel_r_25;
  assign N1295 = N36 & N37 & N38;
  assign N36 = ~bk_dpath_sel_r_22;
  assign N37 = ~bk_dpath_sel_r_20;
  assign N38 = ~bk_dpath_sel_r_21;
  assign N1296 = bk_dpath_sel_r_22 & N39;
  assign N39 = ~bk_dpath_sel_r_20;
  assign N1297 = N40 & bk_dpath_sel_r_20 & N41;
  assign N40 = ~bk_dpath_sel_r_22;
  assign N41 = ~bk_dpath_sel_r_21;
  assign N1299 = N42 & bk_dpath_sel_r_21;
  assign N42 = ~bk_dpath_sel_r_20;
  assign N1300 = bk_dpath_sel_r_20 & bk_dpath_sel_r_21;
  assign N1298 = bk_dpath_sel_r_22 & bk_dpath_sel_r_20;
  assign N1172 = N43 & N44 & N45;
  assign N43 = ~bk_dpath_sel_r_18;
  assign N44 = ~bk_dpath_sel_r_16;
  assign N45 = ~bk_dpath_sel_r_17;
  assign N1173 = bk_dpath_sel_r_16 & N46;
  assign N46 = ~bk_dpath_sel_r_17;
  assign N1174 = N47 & bk_dpath_sel_r_17;
  assign N47 = ~bk_dpath_sel_r_16;
  assign N1175 = bk_dpath_sel_r_16 & bk_dpath_sel_r_17;
  assign N1474 = N48 & N49 & (N50 & N51);
  assign N48 = ~fwd_dpath_sel_r[31];
  assign N49 = ~fwd_dpath_sel_r[30];
  assign N50 = ~fwd_dpath_sel_r[28];
  assign N51 = ~fwd_dpath_sel_r[29];
  assign N1475 = N52 & fwd_dpath_sel_r[28] & N53;
  assign N52 = ~fwd_dpath_sel_r[30];
  assign N53 = ~fwd_dpath_sel_r[29];
  assign N1476 = N54 & N55 & fwd_dpath_sel_r[29];
  assign N54 = ~fwd_dpath_sel_r[30];
  assign N55 = ~fwd_dpath_sel_r[28];
  assign N1477 = N56 & fwd_dpath_sel_r[28] & fwd_dpath_sel_r[29];
  assign N56 = ~fwd_dpath_sel_r[30];
  assign N1478 = fwd_dpath_sel_r[30] & N57 & N58;
  assign N57 = ~fwd_dpath_sel_r[28];
  assign N58 = ~fwd_dpath_sel_r[29];
  assign N1479 = fwd_dpath_sel_r[30] & fwd_dpath_sel_r[28] & N59;
  assign N59 = ~fwd_dpath_sel_r[29];
  assign N1480 = fwd_dpath_sel_r[30] & N60 & fwd_dpath_sel_r[29];
  assign N60 = ~fwd_dpath_sel_r[28];
  assign N1481 = fwd_dpath_sel_r[30] & fwd_dpath_sel_r[28] & fwd_dpath_sel_r[29];
  assign N1349 = N61 & N62 & (N63 & N64);
  assign N61 = ~fwd_dpath_sel_r[27];
  assign N62 = ~fwd_dpath_sel_r[26];
  assign N63 = ~fwd_dpath_sel_r[24];
  assign N64 = ~fwd_dpath_sel_r[25];
  assign N1350 = fwd_dpath_sel_r[27] & N65;
  assign N65 = ~fwd_dpath_sel_r[24];
  assign N1351 = N66 & N67 & (fwd_dpath_sel_r[24] & N68);
  assign N66 = ~fwd_dpath_sel_r[27];
  assign N67 = ~fwd_dpath_sel_r[26];
  assign N68 = ~fwd_dpath_sel_r[25];
  assign N1353 = N69 & N70 & fwd_dpath_sel_r[25];
  assign N69 = ~fwd_dpath_sel_r[26];
  assign N70 = ~fwd_dpath_sel_r[24];
  assign N1354 = N71 & fwd_dpath_sel_r[24] & fwd_dpath_sel_r[25];
  assign N71 = ~fwd_dpath_sel_r[26];
  assign N1355 = fwd_dpath_sel_r[26] & N72 & N73;
  assign N72 = ~fwd_dpath_sel_r[24];
  assign N73 = ~fwd_dpath_sel_r[25];
  assign N1356 = fwd_dpath_sel_r[26] & fwd_dpath_sel_r[24] & N74;
  assign N74 = ~fwd_dpath_sel_r[25];
  assign N1357 = fwd_dpath_sel_r[26] & N75 & fwd_dpath_sel_r[25];
  assign N75 = ~fwd_dpath_sel_r[24];
  assign N1358 = fwd_dpath_sel_r[26] & fwd_dpath_sel_r[24] & fwd_dpath_sel_r[25];
  assign N1352 = fwd_dpath_sel_r[27] & fwd_dpath_sel_r[24];
  assign N1224 = N76 & N77 & (N78 & N79);
  assign N76 = ~fwd_dpath_sel_r[23];
  assign N77 = ~fwd_dpath_sel_r[22];
  assign N78 = ~fwd_dpath_sel_r[20];
  assign N79 = ~fwd_dpath_sel_r[21];
  assign N1225 = fwd_dpath_sel_r[23] & N80 & N81;
  assign N80 = ~fwd_dpath_sel_r[20];
  assign N81 = ~fwd_dpath_sel_r[21];
  assign N1226 = N82 & N83 & (fwd_dpath_sel_r[20] & N84);
  assign N82 = ~fwd_dpath_sel_r[23];
  assign N83 = ~fwd_dpath_sel_r[22];
  assign N84 = ~fwd_dpath_sel_r[21];
  assign N1228 = N85 & N86 & (N87 & fwd_dpath_sel_r[21]);
  assign N85 = ~fwd_dpath_sel_r[23];
  assign N86 = ~fwd_dpath_sel_r[22];
  assign N87 = ~fwd_dpath_sel_r[20];
  assign N1230 = N88 & fwd_dpath_sel_r[20] & fwd_dpath_sel_r[21];
  assign N88 = ~fwd_dpath_sel_r[22];
  assign N1231 = fwd_dpath_sel_r[22] & N89 & N90;
  assign N89 = ~fwd_dpath_sel_r[20];
  assign N90 = ~fwd_dpath_sel_r[21];
  assign N1232 = fwd_dpath_sel_r[22] & fwd_dpath_sel_r[20] & N91;
  assign N91 = ~fwd_dpath_sel_r[21];
  assign N1233 = fwd_dpath_sel_r[22] & N92 & fwd_dpath_sel_r[21];
  assign N92 = ~fwd_dpath_sel_r[20];
  assign N1234 = fwd_dpath_sel_r[22] & fwd_dpath_sel_r[20] & fwd_dpath_sel_r[21];
  assign N1227 = fwd_dpath_sel_r[23] & fwd_dpath_sel_r[20];
  assign N1229 = fwd_dpath_sel_r[23] & fwd_dpath_sel_r[21];
  assign N1100 = N93 & N94 & (N95 & N96);
  assign N93 = ~fwd_dpath_sel_r[19];
  assign N94 = ~fwd_dpath_sel_r[18];
  assign N95 = ~fwd_dpath_sel_r[16];
  assign N96 = ~fwd_dpath_sel_r[17];
  assign N1101 = fwd_dpath_sel_r[19] & N97 & N98;
  assign N97 = ~fwd_dpath_sel_r[16];
  assign N98 = ~fwd_dpath_sel_r[17];
  assign N1102 = N99 & N100 & (fwd_dpath_sel_r[16] & N101);
  assign N99 = ~fwd_dpath_sel_r[19];
  assign N100 = ~fwd_dpath_sel_r[18];
  assign N101 = ~fwd_dpath_sel_r[17];
  assign N1104 = N102 & N103 & (N104 & fwd_dpath_sel_r[17]);
  assign N102 = ~fwd_dpath_sel_r[19];
  assign N103 = ~fwd_dpath_sel_r[18];
  assign N104 = ~fwd_dpath_sel_r[16];
  assign N1106 = N105 & N106 & (fwd_dpath_sel_r[16] & fwd_dpath_sel_r[17]);
  assign N105 = ~fwd_dpath_sel_r[19];
  assign N106 = ~fwd_dpath_sel_r[18];
  assign N1108 = fwd_dpath_sel_r[18] & N107 & N108;
  assign N107 = ~fwd_dpath_sel_r[16];
  assign N108 = ~fwd_dpath_sel_r[17];
  assign N1109 = fwd_dpath_sel_r[18] & fwd_dpath_sel_r[16] & N109;
  assign N109 = ~fwd_dpath_sel_r[17];
  assign N1110 = fwd_dpath_sel_r[18] & N110 & fwd_dpath_sel_r[17];
  assign N110 = ~fwd_dpath_sel_r[16];
  assign N1111 = fwd_dpath_sel_r[18] & fwd_dpath_sel_r[16] & fwd_dpath_sel_r[17];
  assign N1103 = fwd_dpath_sel_r[19] & fwd_dpath_sel_r[16] & N111;
  assign N111 = ~fwd_dpath_sel_r[17];
  assign N1105 = fwd_dpath_sel_r[19] & N112 & fwd_dpath_sel_r[17];
  assign N112 = ~fwd_dpath_sel_r[16];
  assign N1107 = fwd_dpath_sel_r[19] & fwd_dpath_sel_r[16] & fwd_dpath_sel_r[17];
  assign N973 = N113 & N114 & (N115 & N116);
  assign N113 = ~fwd_dpath_sel_r[15];
  assign N114 = ~fwd_dpath_sel_r[14];
  assign N115 = ~fwd_dpath_sel_r[12];
  assign N116 = ~fwd_dpath_sel_r[13];
  assign N974 = fwd_dpath_sel_r[15] & N117 & (N118 & N119);
  assign N117 = ~fwd_dpath_sel_r[14];
  assign N118 = ~fwd_dpath_sel_r[12];
  assign N119 = ~fwd_dpath_sel_r[13];
  assign N975 = N120 & N121 & (fwd_dpath_sel_r[12] & N122);
  assign N120 = ~fwd_dpath_sel_r[15];
  assign N121 = ~fwd_dpath_sel_r[14];
  assign N122 = ~fwd_dpath_sel_r[13];
  assign N977 = N123 & N124 & (N125 & fwd_dpath_sel_r[13]);
  assign N123 = ~fwd_dpath_sel_r[15];
  assign N124 = ~fwd_dpath_sel_r[14];
  assign N125 = ~fwd_dpath_sel_r[12];
  assign N979 = N126 & N127 & (fwd_dpath_sel_r[12] & fwd_dpath_sel_r[13]);
  assign N126 = ~fwd_dpath_sel_r[15];
  assign N127 = ~fwd_dpath_sel_r[14];
  assign N981 = N128 & fwd_dpath_sel_r[14] & (N129 & N130);
  assign N128 = ~fwd_dpath_sel_r[15];
  assign N129 = ~fwd_dpath_sel_r[12];
  assign N130 = ~fwd_dpath_sel_r[13];
  assign N983 = fwd_dpath_sel_r[14] & fwd_dpath_sel_r[12] & N131;
  assign N131 = ~fwd_dpath_sel_r[13];
  assign N984 = fwd_dpath_sel_r[14] & N132 & fwd_dpath_sel_r[13];
  assign N132 = ~fwd_dpath_sel_r[12];
  assign N985 = fwd_dpath_sel_r[14] & fwd_dpath_sel_r[12] & fwd_dpath_sel_r[13];
  assign N976 = fwd_dpath_sel_r[15] & fwd_dpath_sel_r[12] & N133;
  assign N133 = ~fwd_dpath_sel_r[13];
  assign N978 = fwd_dpath_sel_r[15] & N134 & fwd_dpath_sel_r[13];
  assign N134 = ~fwd_dpath_sel_r[12];
  assign N980 = fwd_dpath_sel_r[15] & fwd_dpath_sel_r[12] & fwd_dpath_sel_r[13];
  assign N982 = fwd_dpath_sel_r[15] & fwd_dpath_sel_r[14];
  assign N850 = N135 & N136 & (N137 & N138);
  assign N135 = ~fwd_dpath_sel_r[11];
  assign N136 = ~fwd_dpath_sel_r[10];
  assign N137 = ~fwd_dpath_sel_r[8];
  assign N138 = ~fwd_dpath_sel_r[9];
  assign N851 = fwd_dpath_sel_r[11] & N139 & (N140 & N141);
  assign N139 = ~fwd_dpath_sel_r[10];
  assign N140 = ~fwd_dpath_sel_r[8];
  assign N141 = ~fwd_dpath_sel_r[9];
  assign N852 = N142 & N143 & (fwd_dpath_sel_r[8] & N144);
  assign N142 = ~fwd_dpath_sel_r[11];
  assign N143 = ~fwd_dpath_sel_r[10];
  assign N144 = ~fwd_dpath_sel_r[9];
  assign N854 = N145 & N146 & (N147 & fwd_dpath_sel_r[9]);
  assign N145 = ~fwd_dpath_sel_r[11];
  assign N146 = ~fwd_dpath_sel_r[10];
  assign N147 = ~fwd_dpath_sel_r[8];
  assign N856 = N148 & N149 & (fwd_dpath_sel_r[8] & fwd_dpath_sel_r[9]);
  assign N148 = ~fwd_dpath_sel_r[11];
  assign N149 = ~fwd_dpath_sel_r[10];
  assign N858 = N150 & fwd_dpath_sel_r[10] & (N151 & N152);
  assign N150 = ~fwd_dpath_sel_r[11];
  assign N151 = ~fwd_dpath_sel_r[8];
  assign N152 = ~fwd_dpath_sel_r[9];
  assign N860 = N153 & fwd_dpath_sel_r[10] & (fwd_dpath_sel_r[8] & N154);
  assign N153 = ~fwd_dpath_sel_r[11];
  assign N154 = ~fwd_dpath_sel_r[9];
  assign N862 = fwd_dpath_sel_r[10] & N155 & fwd_dpath_sel_r[9];
  assign N155 = ~fwd_dpath_sel_r[8];
  assign N863 = fwd_dpath_sel_r[10] & fwd_dpath_sel_r[8] & fwd_dpath_sel_r[9];
  assign N853 = fwd_dpath_sel_r[11] & N156 & (fwd_dpath_sel_r[8] & N157);
  assign N156 = ~fwd_dpath_sel_r[10];
  assign N157 = ~fwd_dpath_sel_r[9];
  assign N855 = fwd_dpath_sel_r[11] & N158 & fwd_dpath_sel_r[9];
  assign N158 = ~fwd_dpath_sel_r[8];
  assign N857 = fwd_dpath_sel_r[11] & fwd_dpath_sel_r[8] & fwd_dpath_sel_r[9];
  assign N859 = fwd_dpath_sel_r[11] & fwd_dpath_sel_r[10] & N159;
  assign N159 = ~fwd_dpath_sel_r[8];
  assign N861 = fwd_dpath_sel_r[11] & fwd_dpath_sel_r[10] & fwd_dpath_sel_r[8];
  assign N726 = N160 & N161 & (N162 & N163);
  assign N160 = ~fwd_dpath_sel_r[7];
  assign N161 = ~fwd_dpath_sel_r[6];
  assign N162 = ~fwd_dpath_sel_r[4];
  assign N163 = ~fwd_dpath_sel_r[5];
  assign N727 = fwd_dpath_sel_r[7] & N164 & (N165 & N166);
  assign N164 = ~fwd_dpath_sel_r[6];
  assign N165 = ~fwd_dpath_sel_r[4];
  assign N166 = ~fwd_dpath_sel_r[5];
  assign N728 = N167 & N168 & (fwd_dpath_sel_r[4] & N169);
  assign N167 = ~fwd_dpath_sel_r[7];
  assign N168 = ~fwd_dpath_sel_r[6];
  assign N169 = ~fwd_dpath_sel_r[5];
  assign N730 = N170 & N171 & (N172 & fwd_dpath_sel_r[5]);
  assign N170 = ~fwd_dpath_sel_r[7];
  assign N171 = ~fwd_dpath_sel_r[6];
  assign N172 = ~fwd_dpath_sel_r[4];
  assign N732 = N173 & N174 & (fwd_dpath_sel_r[4] & fwd_dpath_sel_r[5]);
  assign N173 = ~fwd_dpath_sel_r[7];
  assign N174 = ~fwd_dpath_sel_r[6];
  assign N734 = N175 & fwd_dpath_sel_r[6] & (N176 & N177);
  assign N175 = ~fwd_dpath_sel_r[7];
  assign N176 = ~fwd_dpath_sel_r[4];
  assign N177 = ~fwd_dpath_sel_r[5];
  assign N736 = N178 & fwd_dpath_sel_r[6] & (fwd_dpath_sel_r[4] & N179);
  assign N178 = ~fwd_dpath_sel_r[7];
  assign N179 = ~fwd_dpath_sel_r[5];
  assign N738 = N180 & fwd_dpath_sel_r[6] & (N181 & fwd_dpath_sel_r[5]);
  assign N180 = ~fwd_dpath_sel_r[7];
  assign N181 = ~fwd_dpath_sel_r[4];
  assign N740 = fwd_dpath_sel_r[6] & fwd_dpath_sel_r[4] & fwd_dpath_sel_r[5];
  assign N729 = fwd_dpath_sel_r[7] & N182 & (fwd_dpath_sel_r[4] & N183);
  assign N182 = ~fwd_dpath_sel_r[6];
  assign N183 = ~fwd_dpath_sel_r[5];
  assign N731 = fwd_dpath_sel_r[7] & N184 & (N185 & fwd_dpath_sel_r[5]);
  assign N184 = ~fwd_dpath_sel_r[6];
  assign N185 = ~fwd_dpath_sel_r[4];
  assign N733 = fwd_dpath_sel_r[7] & fwd_dpath_sel_r[4] & fwd_dpath_sel_r[5];
  assign N735 = fwd_dpath_sel_r[7] & fwd_dpath_sel_r[6] & (N186 & N187);
  assign N186 = ~fwd_dpath_sel_r[4];
  assign N187 = ~fwd_dpath_sel_r[5];
  assign N737 = fwd_dpath_sel_r[7] & fwd_dpath_sel_r[6] & fwd_dpath_sel_r[4];
  assign N739 = fwd_dpath_sel_r[7] & fwd_dpath_sel_r[6] & fwd_dpath_sel_r[5];
  assign N2421 = N188 & N189 & (N190 & N191);
  assign N188 = ~bk_dpath_sel_r[59];
  assign N189 = ~bk_dpath_sel_r[58];
  assign N190 = ~bk_dpath_sel_r[56];
  assign N191 = ~bk_dpath_sel_r[57];
  assign N2422 = bk_dpath_sel_r[59] & N192 & (N193 & N194);
  assign N192 = ~bk_dpath_sel_r[58];
  assign N193 = ~bk_dpath_sel_r[56];
  assign N194 = ~bk_dpath_sel_r[57];
  assign N2423 = N195 & N196 & (bk_dpath_sel_r[56] & N197);
  assign N195 = ~bk_dpath_sel_r[59];
  assign N196 = ~bk_dpath_sel_r[58];
  assign N197 = ~bk_dpath_sel_r[57];
  assign N2425 = N198 & N199 & (N200 & bk_dpath_sel_r[57]);
  assign N198 = ~bk_dpath_sel_r[59];
  assign N199 = ~bk_dpath_sel_r[58];
  assign N200 = ~bk_dpath_sel_r[56];
  assign N2427 = N201 & N202 & (bk_dpath_sel_r[56] & bk_dpath_sel_r[57]);
  assign N201 = ~bk_dpath_sel_r[59];
  assign N202 = ~bk_dpath_sel_r[58];
  assign N2429 = N203 & bk_dpath_sel_r[58] & (N204 & N205);
  assign N203 = ~bk_dpath_sel_r[59];
  assign N204 = ~bk_dpath_sel_r[56];
  assign N205 = ~bk_dpath_sel_r[57];
  assign N2431 = N206 & bk_dpath_sel_r[58] & (bk_dpath_sel_r[56] & N207);
  assign N206 = ~bk_dpath_sel_r[59];
  assign N207 = ~bk_dpath_sel_r[57];
  assign N2433 = N208 & bk_dpath_sel_r[58] & (N209 & bk_dpath_sel_r[57]);
  assign N208 = ~bk_dpath_sel_r[59];
  assign N209 = ~bk_dpath_sel_r[56];
  assign N2435 = bk_dpath_sel_r[58] & bk_dpath_sel_r[56] & bk_dpath_sel_r[57];
  assign N2424 = bk_dpath_sel_r[59] & N210 & (bk_dpath_sel_r[56] & N211);
  assign N210 = ~bk_dpath_sel_r[58];
  assign N211 = ~bk_dpath_sel_r[57];
  assign N2426 = bk_dpath_sel_r[59] & N212 & (N213 & bk_dpath_sel_r[57]);
  assign N212 = ~bk_dpath_sel_r[58];
  assign N213 = ~bk_dpath_sel_r[56];
  assign N2428 = bk_dpath_sel_r[59] & bk_dpath_sel_r[56] & bk_dpath_sel_r[57];
  assign N2430 = bk_dpath_sel_r[59] & bk_dpath_sel_r[58] & (N214 & N215);
  assign N214 = ~bk_dpath_sel_r[56];
  assign N215 = ~bk_dpath_sel_r[57];
  assign N2432 = bk_dpath_sel_r[59] & bk_dpath_sel_r[58] & bk_dpath_sel_r[56];
  assign N2434 = bk_dpath_sel_r[59] & bk_dpath_sel_r[58] & bk_dpath_sel_r[57];
  assign N2298 = N216 & N217 & (N218 & N219);
  assign N216 = ~bk_dpath_sel_r[55];
  assign N217 = ~bk_dpath_sel_r[54];
  assign N218 = ~bk_dpath_sel_r[52];
  assign N219 = ~bk_dpath_sel_r[53];
  assign N2299 = bk_dpath_sel_r[55] & N220 & (N221 & N222);
  assign N220 = ~bk_dpath_sel_r[54];
  assign N221 = ~bk_dpath_sel_r[52];
  assign N222 = ~bk_dpath_sel_r[53];
  assign N2300 = N223 & N224 & (bk_dpath_sel_r[52] & N225);
  assign N223 = ~bk_dpath_sel_r[55];
  assign N224 = ~bk_dpath_sel_r[54];
  assign N225 = ~bk_dpath_sel_r[53];
  assign N2302 = N226 & N227 & (N228 & bk_dpath_sel_r[53]);
  assign N226 = ~bk_dpath_sel_r[55];
  assign N227 = ~bk_dpath_sel_r[54];
  assign N228 = ~bk_dpath_sel_r[52];
  assign N2304 = N229 & N230 & (bk_dpath_sel_r[52] & bk_dpath_sel_r[53]);
  assign N229 = ~bk_dpath_sel_r[55];
  assign N230 = ~bk_dpath_sel_r[54];
  assign N2306 = N231 & bk_dpath_sel_r[54] & (N232 & N233);
  assign N231 = ~bk_dpath_sel_r[55];
  assign N232 = ~bk_dpath_sel_r[52];
  assign N233 = ~bk_dpath_sel_r[53];
  assign N2308 = N234 & bk_dpath_sel_r[54] & (bk_dpath_sel_r[52] & N235);
  assign N234 = ~bk_dpath_sel_r[55];
  assign N235 = ~bk_dpath_sel_r[53];
  assign N2310 = bk_dpath_sel_r[54] & N236 & bk_dpath_sel_r[53];
  assign N236 = ~bk_dpath_sel_r[52];
  assign N2311 = bk_dpath_sel_r[54] & bk_dpath_sel_r[52] & bk_dpath_sel_r[53];
  assign N2301 = bk_dpath_sel_r[55] & N237 & (bk_dpath_sel_r[52] & N238);
  assign N237 = ~bk_dpath_sel_r[54];
  assign N238 = ~bk_dpath_sel_r[53];
  assign N2303 = bk_dpath_sel_r[55] & N239 & bk_dpath_sel_r[53];
  assign N239 = ~bk_dpath_sel_r[52];
  assign N2305 = bk_dpath_sel_r[55] & bk_dpath_sel_r[52] & bk_dpath_sel_r[53];
  assign N2307 = bk_dpath_sel_r[55] & bk_dpath_sel_r[54] & N240;
  assign N240 = ~bk_dpath_sel_r[52];
  assign N2309 = bk_dpath_sel_r[55] & bk_dpath_sel_r[54] & bk_dpath_sel_r[52];
  assign N2176 = N241 & N242 & (N243 & N244);
  assign N241 = ~bk_dpath_sel_r[51];
  assign N242 = ~bk_dpath_sel_r[50];
  assign N243 = ~bk_dpath_sel_r[48];
  assign N244 = ~bk_dpath_sel_r[49];
  assign N2177 = bk_dpath_sel_r[51] & N245 & (N246 & N247);
  assign N245 = ~bk_dpath_sel_r[50];
  assign N246 = ~bk_dpath_sel_r[48];
  assign N247 = ~bk_dpath_sel_r[49];
  assign N2178 = N248 & N249 & (bk_dpath_sel_r[48] & N250);
  assign N248 = ~bk_dpath_sel_r[51];
  assign N249 = ~bk_dpath_sel_r[50];
  assign N250 = ~bk_dpath_sel_r[49];
  assign N2180 = N251 & N252 & (N253 & bk_dpath_sel_r[49]);
  assign N251 = ~bk_dpath_sel_r[51];
  assign N252 = ~bk_dpath_sel_r[50];
  assign N253 = ~bk_dpath_sel_r[48];
  assign N2182 = N254 & N255 & (bk_dpath_sel_r[48] & bk_dpath_sel_r[49]);
  assign N254 = ~bk_dpath_sel_r[51];
  assign N255 = ~bk_dpath_sel_r[50];
  assign N2184 = N256 & bk_dpath_sel_r[50] & (N257 & N258);
  assign N256 = ~bk_dpath_sel_r[51];
  assign N257 = ~bk_dpath_sel_r[48];
  assign N258 = ~bk_dpath_sel_r[49];
  assign N2186 = bk_dpath_sel_r[50] & bk_dpath_sel_r[48] & N259;
  assign N259 = ~bk_dpath_sel_r[49];
  assign N2187 = bk_dpath_sel_r[50] & N260 & bk_dpath_sel_r[49];
  assign N260 = ~bk_dpath_sel_r[48];
  assign N2188 = bk_dpath_sel_r[50] & bk_dpath_sel_r[48] & bk_dpath_sel_r[49];
  assign N2179 = bk_dpath_sel_r[51] & bk_dpath_sel_r[48] & N261;
  assign N261 = ~bk_dpath_sel_r[49];
  assign N2181 = bk_dpath_sel_r[51] & N262 & bk_dpath_sel_r[49];
  assign N262 = ~bk_dpath_sel_r[48];
  assign N2183 = bk_dpath_sel_r[51] & bk_dpath_sel_r[48] & bk_dpath_sel_r[49];
  assign N2185 = bk_dpath_sel_r[51] & bk_dpath_sel_r[50];
  assign N2050 = N263 & N264 & (N265 & N266);
  assign N263 = ~bk_dpath_sel_r[47];
  assign N264 = ~bk_dpath_sel_r[46];
  assign N265 = ~bk_dpath_sel_r[44];
  assign N266 = ~bk_dpath_sel_r[45];
  assign N2051 = bk_dpath_sel_r[47] & N267 & N268;
  assign N267 = ~bk_dpath_sel_r[44];
  assign N268 = ~bk_dpath_sel_r[45];
  assign N2052 = N269 & N270 & (bk_dpath_sel_r[44] & N271);
  assign N269 = ~bk_dpath_sel_r[47];
  assign N270 = ~bk_dpath_sel_r[46];
  assign N271 = ~bk_dpath_sel_r[45];
  assign N2054 = N272 & N273 & (N274 & bk_dpath_sel_r[45]);
  assign N272 = ~bk_dpath_sel_r[47];
  assign N273 = ~bk_dpath_sel_r[46];
  assign N274 = ~bk_dpath_sel_r[44];
  assign N2056 = N275 & N276 & (bk_dpath_sel_r[44] & bk_dpath_sel_r[45]);
  assign N275 = ~bk_dpath_sel_r[47];
  assign N276 = ~bk_dpath_sel_r[46];
  assign N2058 = bk_dpath_sel_r[46] & N277 & N278;
  assign N277 = ~bk_dpath_sel_r[44];
  assign N278 = ~bk_dpath_sel_r[45];
  assign N2059 = bk_dpath_sel_r[46] & bk_dpath_sel_r[44] & N279;
  assign N279 = ~bk_dpath_sel_r[45];
  assign N2060 = bk_dpath_sel_r[46] & N280 & bk_dpath_sel_r[45];
  assign N280 = ~bk_dpath_sel_r[44];
  assign N2061 = bk_dpath_sel_r[46] & bk_dpath_sel_r[44] & bk_dpath_sel_r[45];
  assign N2053 = bk_dpath_sel_r[47] & bk_dpath_sel_r[44] & N281;
  assign N281 = ~bk_dpath_sel_r[45];
  assign N2055 = bk_dpath_sel_r[47] & N282 & bk_dpath_sel_r[45];
  assign N282 = ~bk_dpath_sel_r[44];
  assign N2057 = bk_dpath_sel_r[47] & bk_dpath_sel_r[44] & bk_dpath_sel_r[45];
  assign N1927 = N283 & N284 & (N285 & N286);
  assign N283 = ~bk_dpath_sel_r[43];
  assign N284 = ~bk_dpath_sel_r[42];
  assign N285 = ~bk_dpath_sel_r[40];
  assign N286 = ~bk_dpath_sel_r[41];
  assign N1928 = bk_dpath_sel_r[43] & N287 & N288;
  assign N287 = ~bk_dpath_sel_r[40];
  assign N288 = ~bk_dpath_sel_r[41];
  assign N1929 = N289 & N290 & (bk_dpath_sel_r[40] & N291);
  assign N289 = ~bk_dpath_sel_r[43];
  assign N290 = ~bk_dpath_sel_r[42];
  assign N291 = ~bk_dpath_sel_r[41];
  assign N1931 = N292 & N293 & (N294 & bk_dpath_sel_r[41]);
  assign N292 = ~bk_dpath_sel_r[43];
  assign N293 = ~bk_dpath_sel_r[42];
  assign N294 = ~bk_dpath_sel_r[40];
  assign N1933 = N295 & bk_dpath_sel_r[40] & bk_dpath_sel_r[41];
  assign N295 = ~bk_dpath_sel_r[42];
  assign N1934 = bk_dpath_sel_r[42] & N296 & N297;
  assign N296 = ~bk_dpath_sel_r[40];
  assign N297 = ~bk_dpath_sel_r[41];
  assign N1935 = bk_dpath_sel_r[42] & bk_dpath_sel_r[40] & N298;
  assign N298 = ~bk_dpath_sel_r[41];
  assign N1936 = bk_dpath_sel_r[42] & N299 & bk_dpath_sel_r[41];
  assign N299 = ~bk_dpath_sel_r[40];
  assign N1937 = bk_dpath_sel_r[42] & bk_dpath_sel_r[40] & bk_dpath_sel_r[41];
  assign N1930 = bk_dpath_sel_r[43] & bk_dpath_sel_r[40];
  assign N1932 = bk_dpath_sel_r[43] & bk_dpath_sel_r[41];
  assign N1803 = N300 & N301 & (N302 & N303);
  assign N300 = ~bk_dpath_sel_r[39];
  assign N301 = ~bk_dpath_sel_r[38];
  assign N302 = ~bk_dpath_sel_r[36];
  assign N303 = ~bk_dpath_sel_r[37];
  assign N1804 = bk_dpath_sel_r[39] & N304;
  assign N304 = ~bk_dpath_sel_r[36];
  assign N1805 = N305 & N306 & (bk_dpath_sel_r[36] & N307);
  assign N305 = ~bk_dpath_sel_r[39];
  assign N306 = ~bk_dpath_sel_r[38];
  assign N307 = ~bk_dpath_sel_r[37];
  assign N1807 = N308 & N309 & bk_dpath_sel_r[37];
  assign N308 = ~bk_dpath_sel_r[38];
  assign N309 = ~bk_dpath_sel_r[36];
  assign N1808 = N310 & bk_dpath_sel_r[36] & bk_dpath_sel_r[37];
  assign N310 = ~bk_dpath_sel_r[38];
  assign N1809 = bk_dpath_sel_r[38] & N311 & N312;
  assign N311 = ~bk_dpath_sel_r[36];
  assign N312 = ~bk_dpath_sel_r[37];
  assign N1810 = bk_dpath_sel_r[38] & bk_dpath_sel_r[36] & N313;
  assign N313 = ~bk_dpath_sel_r[37];
  assign N1811 = bk_dpath_sel_r[38] & N314 & bk_dpath_sel_r[37];
  assign N314 = ~bk_dpath_sel_r[36];
  assign N1812 = bk_dpath_sel_r[38] & bk_dpath_sel_r[36] & bk_dpath_sel_r[37];
  assign N1806 = bk_dpath_sel_r[39] & bk_dpath_sel_r[36];
  assign N1680 = N315 & N316 & (N317 & N318);
  assign N315 = ~bk_dpath_sel_r[35];
  assign N316 = ~bk_dpath_sel_r[34];
  assign N317 = ~bk_dpath_sel_r[32];
  assign N318 = ~bk_dpath_sel_r[33];
  assign N1681 = N319 & bk_dpath_sel_r[32] & N320;
  assign N319 = ~bk_dpath_sel_r[34];
  assign N320 = ~bk_dpath_sel_r[33];
  assign N1682 = N321 & N322 & bk_dpath_sel_r[33];
  assign N321 = ~bk_dpath_sel_r[34];
  assign N322 = ~bk_dpath_sel_r[32];
  assign N1683 = N323 & bk_dpath_sel_r[32] & bk_dpath_sel_r[33];
  assign N323 = ~bk_dpath_sel_r[34];
  assign N1684 = bk_dpath_sel_r[34] & N324 & N325;
  assign N324 = ~bk_dpath_sel_r[32];
  assign N325 = ~bk_dpath_sel_r[33];
  assign N1685 = bk_dpath_sel_r[34] & bk_dpath_sel_r[32] & N326;
  assign N326 = ~bk_dpath_sel_r[33];
  assign N1686 = bk_dpath_sel_r[34] & N327 & bk_dpath_sel_r[33];
  assign N327 = ~bk_dpath_sel_r[32];
  assign N1687 = bk_dpath_sel_r[34] & bk_dpath_sel_r[32] & bk_dpath_sel_r[33];
  assign in_data_o[447] = (N328)? in_data_i[447] : 
                          (N329)? in_data_i[479] : 
                          (N330)? in_data_i_15__31_ : 1'b0;
  assign N328 = N2237;
  assign N329 = fwd_dpath_sel_r_52;
  assign N330 = fwd_dpath_sel_r_53;
  assign in_data_o[446] = (N328)? in_data_i[446] : 
                          (N329)? in_data_i[478] : 
                          (N330)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[445] = (N328)? in_data_i[445] : 
                          (N329)? in_data_i[477] : 
                          (N330)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[444] = (N328)? in_data_i[444] : 
                          (N329)? in_data_i[476] : 
                          (N330)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[443] = (N328)? in_data_i[443] : 
                          (N329)? in_data_i[475] : 
                          (N330)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[442] = (N328)? in_data_i[442] : 
                          (N329)? in_data_i[474] : 
                          (N330)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[441] = (N328)? in_data_i[441] : 
                          (N329)? in_data_i[473] : 
                          (N330)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[440] = (N328)? in_data_i[440] : 
                          (N329)? in_data_i[472] : 
                          (N330)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[439] = (N328)? in_data_i[439] : 
                          (N329)? in_data_i[471] : 
                          (N330)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[438] = (N328)? in_data_i[438] : 
                          (N329)? in_data_i[470] : 
                          (N330)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[437] = (N328)? in_data_i[437] : 
                          (N329)? in_data_i[469] : 
                          (N330)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[436] = (N328)? in_data_i[436] : 
                          (N329)? in_data_i[468] : 
                          (N330)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[435] = (N328)? in_data_i[435] : 
                          (N329)? in_data_i[467] : 
                          (N330)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[434] = (N328)? in_data_i[434] : 
                          (N329)? in_data_i[466] : 
                          (N330)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[433] = (N328)? in_data_i[433] : 
                          (N329)? in_data_i[465] : 
                          (N330)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[432] = (N328)? in_data_i[432] : 
                          (N329)? in_data_i[464] : 
                          (N330)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[431] = (N328)? in_data_i[431] : 
                          (N329)? in_data_i[463] : 
                          (N330)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[430] = (N328)? in_data_i[430] : 
                          (N329)? in_data_i[462] : 
                          (N330)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[429] = (N328)? in_data_i[429] : 
                          (N329)? in_data_i[461] : 
                          (N330)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[428] = (N328)? in_data_i[428] : 
                          (N329)? in_data_i[460] : 
                          (N330)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[427] = (N328)? in_data_i[427] : 
                          (N329)? in_data_i[459] : 
                          (N330)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[426] = (N328)? in_data_i[426] : 
                          (N329)? in_data_i[458] : 
                          (N330)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[425] = (N328)? in_data_i[425] : 
                          (N329)? in_data_i[457] : 
                          (N330)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[424] = (N328)? in_data_i[424] : 
                          (N329)? in_data_i[456] : 
                          (N330)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[423] = (N328)? in_data_i[423] : 
                          (N329)? in_data_i[455] : 
                          (N330)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[422] = (N328)? in_data_i[422] : 
                          (N329)? in_data_i[454] : 
                          (N330)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[421] = (N328)? in_data_i[421] : 
                          (N329)? in_data_i[453] : 
                          (N330)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[420] = (N328)? in_data_i[420] : 
                          (N329)? in_data_i[452] : 
                          (N330)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[419] = (N328)? in_data_i[419] : 
                          (N329)? in_data_i[451] : 
                          (N330)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[418] = (N328)? in_data_i[418] : 
                          (N329)? in_data_i[450] : 
                          (N330)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[417] = (N328)? in_data_i[417] : 
                          (N329)? in_data_i[449] : 
                          (N330)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[416] = (N328)? in_data_i[416] : 
                          (N329)? in_data_i[448] : 
                          (N330)? in_data_i_15__0_ : 1'b0;
  assign out_me_data_o[95] = (N331)? out_me_data_i_0__31_ : 
                             (N332)? out_me_data_i[63] : 
                             (N333)? out_me_data_i[95] : 1'b0;
  assign N331 = N924;
  assign N332 = bk_dpath_sel_r_8;
  assign N333 = bk_dpath_sel_r_9;
  assign out_me_data_o[94] = (N331)? out_me_data_i_0__30_ : 
                             (N332)? out_me_data_i[62] : 
                             (N333)? out_me_data_i[94] : 1'b0;
  assign out_me_data_o[93] = (N331)? out_me_data_i_0__29_ : 
                             (N332)? out_me_data_i[61] : 
                             (N333)? out_me_data_i[93] : 1'b0;
  assign out_me_data_o[92] = (N331)? out_me_data_i_0__28_ : 
                             (N332)? out_me_data_i[60] : 
                             (N333)? out_me_data_i[92] : 1'b0;
  assign out_me_data_o[91] = (N331)? out_me_data_i_0__27_ : 
                             (N332)? out_me_data_i[59] : 
                             (N333)? out_me_data_i[91] : 1'b0;
  assign out_me_data_o[90] = (N331)? out_me_data_i_0__26_ : 
                             (N332)? out_me_data_i[58] : 
                             (N333)? out_me_data_i[90] : 1'b0;
  assign out_me_data_o[89] = (N331)? out_me_data_i_0__25_ : 
                             (N332)? out_me_data_i[57] : 
                             (N333)? out_me_data_i[89] : 1'b0;
  assign out_me_data_o[88] = (N331)? out_me_data_i_0__24_ : 
                             (N332)? out_me_data_i[56] : 
                             (N333)? out_me_data_i[88] : 1'b0;
  assign out_me_data_o[87] = (N331)? out_me_data_i_0__23_ : 
                             (N332)? out_me_data_i[55] : 
                             (N333)? out_me_data_i[87] : 1'b0;
  assign out_me_data_o[86] = (N331)? out_me_data_i_0__22_ : 
                             (N332)? out_me_data_i[54] : 
                             (N333)? out_me_data_i[86] : 1'b0;
  assign out_me_data_o[85] = (N331)? out_me_data_i_0__21_ : 
                             (N332)? out_me_data_i[53] : 
                             (N333)? out_me_data_i[85] : 1'b0;
  assign out_me_data_o[84] = (N331)? out_me_data_i_0__20_ : 
                             (N332)? out_me_data_i[52] : 
                             (N333)? out_me_data_i[84] : 1'b0;
  assign out_me_data_o[83] = (N331)? out_me_data_i_0__19_ : 
                             (N332)? out_me_data_i[51] : 
                             (N333)? out_me_data_i[83] : 1'b0;
  assign out_me_data_o[82] = (N331)? out_me_data_i_0__18_ : 
                             (N332)? out_me_data_i[50] : 
                             (N333)? out_me_data_i[82] : 1'b0;
  assign out_me_data_o[81] = (N331)? out_me_data_i_0__17_ : 
                             (N332)? out_me_data_i[49] : 
                             (N333)? out_me_data_i[81] : 1'b0;
  assign out_me_data_o[80] = (N331)? out_me_data_i_0__16_ : 
                             (N332)? out_me_data_i[48] : 
                             (N333)? out_me_data_i[80] : 1'b0;
  assign out_me_data_o[79] = (N331)? out_me_data_i_0__15_ : 
                             (N332)? out_me_data_i[47] : 
                             (N333)? out_me_data_i[79] : 1'b0;
  assign out_me_data_o[78] = (N331)? out_me_data_i_0__14_ : 
                             (N332)? out_me_data_i[46] : 
                             (N333)? out_me_data_i[78] : 1'b0;
  assign out_me_data_o[77] = (N331)? out_me_data_i_0__13_ : 
                             (N332)? out_me_data_i[45] : 
                             (N333)? out_me_data_i[77] : 1'b0;
  assign out_me_data_o[76] = (N331)? out_me_data_i_0__12_ : 
                             (N332)? out_me_data_i[44] : 
                             (N333)? out_me_data_i[76] : 1'b0;
  assign out_me_data_o[75] = (N331)? out_me_data_i_0__11_ : 
                             (N332)? out_me_data_i[43] : 
                             (N333)? out_me_data_i[75] : 1'b0;
  assign out_me_data_o[74] = (N331)? out_me_data_i_0__10_ : 
                             (N332)? out_me_data_i[42] : 
                             (N333)? out_me_data_i[74] : 1'b0;
  assign out_me_data_o[73] = (N331)? out_me_data_i_0__9_ : 
                             (N332)? out_me_data_i[41] : 
                             (N333)? out_me_data_i[73] : 1'b0;
  assign out_me_data_o[72] = (N331)? out_me_data_i_0__8_ : 
                             (N332)? out_me_data_i[40] : 
                             (N333)? out_me_data_i[72] : 1'b0;
  assign out_me_data_o[71] = (N331)? out_me_data_i_0__7_ : 
                             (N332)? out_me_data_i[39] : 
                             (N333)? out_me_data_i[71] : 1'b0;
  assign out_me_data_o[70] = (N331)? out_me_data_i_0__6_ : 
                             (N332)? out_me_data_i[38] : 
                             (N333)? out_me_data_i[70] : 1'b0;
  assign out_me_data_o[69] = (N331)? out_me_data_i_0__5_ : 
                             (N332)? out_me_data_i[37] : 
                             (N333)? out_me_data_i[69] : 1'b0;
  assign out_me_data_o[68] = (N331)? out_me_data_i_0__4_ : 
                             (N332)? out_me_data_i[36] : 
                             (N333)? out_me_data_i[68] : 1'b0;
  assign out_me_data_o[67] = (N331)? out_me_data_i_0__3_ : 
                             (N332)? out_me_data_i[35] : 
                             (N333)? out_me_data_i[67] : 1'b0;
  assign out_me_data_o[66] = (N331)? out_me_data_i_0__2_ : 
                             (N332)? out_me_data_i[34] : 
                             (N333)? out_me_data_i[66] : 1'b0;
  assign out_me_data_o[65] = (N331)? out_me_data_i_0__1_ : 
                             (N332)? out_me_data_i[33] : 
                             (N333)? out_me_data_i[65] : 1'b0;
  assign out_me_data_o[64] = (N331)? out_me_data_i_0__0_ : 
                             (N332)? out_me_data_i[32] : 
                             (N333)? out_me_data_i[64] : 1'b0;
  assign in_data_o[383] = (N334)? in_data_i[383] : 
                          (N335)? in_data_i[415] : 
                          (N336)? in_data_i[447] : 
                          (N337)? in_data_i[479] : 
                          (N338)? in_data_i_15__31_ : 1'b0;
  assign N334 = N1986;
  assign N335 = N1987;
  assign N336 = N1988;
  assign N337 = N1989;
  assign N338 = fwd_dpath_sel_r_46;
  assign in_data_o[382] = (N334)? in_data_i[382] : 
                          (N335)? in_data_i[414] : 
                          (N336)? in_data_i[446] : 
                          (N337)? in_data_i[478] : 
                          (N338)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[381] = (N334)? in_data_i[381] : 
                          (N335)? in_data_i[413] : 
                          (N336)? in_data_i[445] : 
                          (N337)? in_data_i[477] : 
                          (N338)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[380] = (N334)? in_data_i[380] : 
                          (N335)? in_data_i[412] : 
                          (N336)? in_data_i[444] : 
                          (N337)? in_data_i[476] : 
                          (N338)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[379] = (N334)? in_data_i[379] : 
                          (N335)? in_data_i[411] : 
                          (N336)? in_data_i[443] : 
                          (N337)? in_data_i[475] : 
                          (N338)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[378] = (N334)? in_data_i[378] : 
                          (N335)? in_data_i[410] : 
                          (N336)? in_data_i[442] : 
                          (N337)? in_data_i[474] : 
                          (N338)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[377] = (N334)? in_data_i[377] : 
                          (N335)? in_data_i[409] : 
                          (N336)? in_data_i[441] : 
                          (N337)? in_data_i[473] : 
                          (N338)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[376] = (N334)? in_data_i[376] : 
                          (N335)? in_data_i[408] : 
                          (N336)? in_data_i[440] : 
                          (N337)? in_data_i[472] : 
                          (N338)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[375] = (N334)? in_data_i[375] : 
                          (N335)? in_data_i[407] : 
                          (N336)? in_data_i[439] : 
                          (N337)? in_data_i[471] : 
                          (N338)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[374] = (N334)? in_data_i[374] : 
                          (N335)? in_data_i[406] : 
                          (N336)? in_data_i[438] : 
                          (N337)? in_data_i[470] : 
                          (N338)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[373] = (N334)? in_data_i[373] : 
                          (N335)? in_data_i[405] : 
                          (N336)? in_data_i[437] : 
                          (N337)? in_data_i[469] : 
                          (N338)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[372] = (N334)? in_data_i[372] : 
                          (N335)? in_data_i[404] : 
                          (N336)? in_data_i[436] : 
                          (N337)? in_data_i[468] : 
                          (N338)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[371] = (N334)? in_data_i[371] : 
                          (N335)? in_data_i[403] : 
                          (N336)? in_data_i[435] : 
                          (N337)? in_data_i[467] : 
                          (N338)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[370] = (N334)? in_data_i[370] : 
                          (N335)? in_data_i[402] : 
                          (N336)? in_data_i[434] : 
                          (N337)? in_data_i[466] : 
                          (N338)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[369] = (N334)? in_data_i[369] : 
                          (N335)? in_data_i[401] : 
                          (N336)? in_data_i[433] : 
                          (N337)? in_data_i[465] : 
                          (N338)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[368] = (N334)? in_data_i[368] : 
                          (N335)? in_data_i[400] : 
                          (N336)? in_data_i[432] : 
                          (N337)? in_data_i[464] : 
                          (N338)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[367] = (N334)? in_data_i[367] : 
                          (N335)? in_data_i[399] : 
                          (N336)? in_data_i[431] : 
                          (N337)? in_data_i[463] : 
                          (N338)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[366] = (N334)? in_data_i[366] : 
                          (N335)? in_data_i[398] : 
                          (N336)? in_data_i[430] : 
                          (N337)? in_data_i[462] : 
                          (N338)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[365] = (N334)? in_data_i[365] : 
                          (N335)? in_data_i[397] : 
                          (N336)? in_data_i[429] : 
                          (N337)? in_data_i[461] : 
                          (N338)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[364] = (N334)? in_data_i[364] : 
                          (N335)? in_data_i[396] : 
                          (N336)? in_data_i[428] : 
                          (N337)? in_data_i[460] : 
                          (N338)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[363] = (N334)? in_data_i[363] : 
                          (N335)? in_data_i[395] : 
                          (N336)? in_data_i[427] : 
                          (N337)? in_data_i[459] : 
                          (N338)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[362] = (N334)? in_data_i[362] : 
                          (N335)? in_data_i[394] : 
                          (N336)? in_data_i[426] : 
                          (N337)? in_data_i[458] : 
                          (N338)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[361] = (N334)? in_data_i[361] : 
                          (N335)? in_data_i[393] : 
                          (N336)? in_data_i[425] : 
                          (N337)? in_data_i[457] : 
                          (N338)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[360] = (N334)? in_data_i[360] : 
                          (N335)? in_data_i[392] : 
                          (N336)? in_data_i[424] : 
                          (N337)? in_data_i[456] : 
                          (N338)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[359] = (N334)? in_data_i[359] : 
                          (N335)? in_data_i[391] : 
                          (N336)? in_data_i[423] : 
                          (N337)? in_data_i[455] : 
                          (N338)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[358] = (N334)? in_data_i[358] : 
                          (N335)? in_data_i[390] : 
                          (N336)? in_data_i[422] : 
                          (N337)? in_data_i[454] : 
                          (N338)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[357] = (N334)? in_data_i[357] : 
                          (N335)? in_data_i[389] : 
                          (N336)? in_data_i[421] : 
                          (N337)? in_data_i[453] : 
                          (N338)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[356] = (N334)? in_data_i[356] : 
                          (N335)? in_data_i[388] : 
                          (N336)? in_data_i[420] : 
                          (N337)? in_data_i[452] : 
                          (N338)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[355] = (N334)? in_data_i[355] : 
                          (N335)? in_data_i[387] : 
                          (N336)? in_data_i[419] : 
                          (N337)? in_data_i[451] : 
                          (N338)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[354] = (N334)? in_data_i[354] : 
                          (N335)? in_data_i[386] : 
                          (N336)? in_data_i[418] : 
                          (N337)? in_data_i[450] : 
                          (N338)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[353] = (N334)? in_data_i[353] : 
                          (N335)? in_data_i[385] : 
                          (N336)? in_data_i[417] : 
                          (N337)? in_data_i[449] : 
                          (N338)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[352] = (N334)? in_data_i[352] : 
                          (N335)? in_data_i[384] : 
                          (N336)? in_data_i[416] : 
                          (N337)? in_data_i[448] : 
                          (N338)? in_data_i_15__0_ : 1'b0;
  assign in_data_o[351] = (N339)? in_data_i[351] : 
                          (N340)? in_data_i[383] : 
                          (N341)? in_data_i[415] : 
                          (N342)? in_data_i[447] : 
                          (N343)? in_data_i[479] : 
                          (N344)? in_data_i_15__31_ : 1'b0;
  assign N339 = N1861;
  assign N340 = N1863;
  assign N341 = N1865;
  assign N342 = N1866;
  assign N343 = N1862;
  assign N344 = N1864;
  assign in_data_o[350] = (N339)? in_data_i[350] : 
                          (N340)? in_data_i[382] : 
                          (N341)? in_data_i[414] : 
                          (N342)? in_data_i[446] : 
                          (N343)? in_data_i[478] : 
                          (N344)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[349] = (N339)? in_data_i[349] : 
                          (N340)? in_data_i[381] : 
                          (N341)? in_data_i[413] : 
                          (N342)? in_data_i[445] : 
                          (N343)? in_data_i[477] : 
                          (N344)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[348] = (N339)? in_data_i[348] : 
                          (N340)? in_data_i[380] : 
                          (N341)? in_data_i[412] : 
                          (N342)? in_data_i[444] : 
                          (N343)? in_data_i[476] : 
                          (N344)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[347] = (N339)? in_data_i[347] : 
                          (N340)? in_data_i[379] : 
                          (N341)? in_data_i[411] : 
                          (N342)? in_data_i[443] : 
                          (N343)? in_data_i[475] : 
                          (N344)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[346] = (N339)? in_data_i[346] : 
                          (N340)? in_data_i[378] : 
                          (N341)? in_data_i[410] : 
                          (N342)? in_data_i[442] : 
                          (N343)? in_data_i[474] : 
                          (N344)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[345] = (N339)? in_data_i[345] : 
                          (N340)? in_data_i[377] : 
                          (N341)? in_data_i[409] : 
                          (N342)? in_data_i[441] : 
                          (N343)? in_data_i[473] : 
                          (N344)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[344] = (N339)? in_data_i[344] : 
                          (N340)? in_data_i[376] : 
                          (N341)? in_data_i[408] : 
                          (N342)? in_data_i[440] : 
                          (N343)? in_data_i[472] : 
                          (N344)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[343] = (N339)? in_data_i[343] : 
                          (N340)? in_data_i[375] : 
                          (N341)? in_data_i[407] : 
                          (N342)? in_data_i[439] : 
                          (N343)? in_data_i[471] : 
                          (N344)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[342] = (N339)? in_data_i[342] : 
                          (N340)? in_data_i[374] : 
                          (N341)? in_data_i[406] : 
                          (N342)? in_data_i[438] : 
                          (N343)? in_data_i[470] : 
                          (N344)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[341] = (N339)? in_data_i[341] : 
                          (N340)? in_data_i[373] : 
                          (N341)? in_data_i[405] : 
                          (N342)? in_data_i[437] : 
                          (N343)? in_data_i[469] : 
                          (N344)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[340] = (N339)? in_data_i[340] : 
                          (N340)? in_data_i[372] : 
                          (N341)? in_data_i[404] : 
                          (N342)? in_data_i[436] : 
                          (N343)? in_data_i[468] : 
                          (N344)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[339] = (N339)? in_data_i[339] : 
                          (N340)? in_data_i[371] : 
                          (N341)? in_data_i[403] : 
                          (N342)? in_data_i[435] : 
                          (N343)? in_data_i[467] : 
                          (N344)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[338] = (N339)? in_data_i[338] : 
                          (N340)? in_data_i[370] : 
                          (N341)? in_data_i[402] : 
                          (N342)? in_data_i[434] : 
                          (N343)? in_data_i[466] : 
                          (N344)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[337] = (N339)? in_data_i[337] : 
                          (N340)? in_data_i[369] : 
                          (N341)? in_data_i[401] : 
                          (N342)? in_data_i[433] : 
                          (N343)? in_data_i[465] : 
                          (N344)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[336] = (N339)? in_data_i[336] : 
                          (N340)? in_data_i[368] : 
                          (N341)? in_data_i[400] : 
                          (N342)? in_data_i[432] : 
                          (N343)? in_data_i[464] : 
                          (N344)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[335] = (N339)? in_data_i[335] : 
                          (N340)? in_data_i[367] : 
                          (N341)? in_data_i[399] : 
                          (N342)? in_data_i[431] : 
                          (N343)? in_data_i[463] : 
                          (N344)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[334] = (N339)? in_data_i[334] : 
                          (N340)? in_data_i[366] : 
                          (N341)? in_data_i[398] : 
                          (N342)? in_data_i[430] : 
                          (N343)? in_data_i[462] : 
                          (N344)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[333] = (N339)? in_data_i[333] : 
                          (N340)? in_data_i[365] : 
                          (N341)? in_data_i[397] : 
                          (N342)? in_data_i[429] : 
                          (N343)? in_data_i[461] : 
                          (N344)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[332] = (N339)? in_data_i[332] : 
                          (N340)? in_data_i[364] : 
                          (N341)? in_data_i[396] : 
                          (N342)? in_data_i[428] : 
                          (N343)? in_data_i[460] : 
                          (N344)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[331] = (N339)? in_data_i[331] : 
                          (N340)? in_data_i[363] : 
                          (N341)? in_data_i[395] : 
                          (N342)? in_data_i[427] : 
                          (N343)? in_data_i[459] : 
                          (N344)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[330] = (N339)? in_data_i[330] : 
                          (N340)? in_data_i[362] : 
                          (N341)? in_data_i[394] : 
                          (N342)? in_data_i[426] : 
                          (N343)? in_data_i[458] : 
                          (N344)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[329] = (N339)? in_data_i[329] : 
                          (N340)? in_data_i[361] : 
                          (N341)? in_data_i[393] : 
                          (N342)? in_data_i[425] : 
                          (N343)? in_data_i[457] : 
                          (N344)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[328] = (N339)? in_data_i[328] : 
                          (N340)? in_data_i[360] : 
                          (N341)? in_data_i[392] : 
                          (N342)? in_data_i[424] : 
                          (N343)? in_data_i[456] : 
                          (N344)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[327] = (N339)? in_data_i[327] : 
                          (N340)? in_data_i[359] : 
                          (N341)? in_data_i[391] : 
                          (N342)? in_data_i[423] : 
                          (N343)? in_data_i[455] : 
                          (N344)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[326] = (N339)? in_data_i[326] : 
                          (N340)? in_data_i[358] : 
                          (N341)? in_data_i[390] : 
                          (N342)? in_data_i[422] : 
                          (N343)? in_data_i[454] : 
                          (N344)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[325] = (N339)? in_data_i[325] : 
                          (N340)? in_data_i[357] : 
                          (N341)? in_data_i[389] : 
                          (N342)? in_data_i[421] : 
                          (N343)? in_data_i[453] : 
                          (N344)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[324] = (N339)? in_data_i[324] : 
                          (N340)? in_data_i[356] : 
                          (N341)? in_data_i[388] : 
                          (N342)? in_data_i[420] : 
                          (N343)? in_data_i[452] : 
                          (N344)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[323] = (N339)? in_data_i[323] : 
                          (N340)? in_data_i[355] : 
                          (N341)? in_data_i[387] : 
                          (N342)? in_data_i[419] : 
                          (N343)? in_data_i[451] : 
                          (N344)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[322] = (N339)? in_data_i[322] : 
                          (N340)? in_data_i[354] : 
                          (N341)? in_data_i[386] : 
                          (N342)? in_data_i[418] : 
                          (N343)? in_data_i[450] : 
                          (N344)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[321] = (N339)? in_data_i[321] : 
                          (N340)? in_data_i[353] : 
                          (N341)? in_data_i[385] : 
                          (N342)? in_data_i[417] : 
                          (N343)? in_data_i[449] : 
                          (N344)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[320] = (N339)? in_data_i[320] : 
                          (N340)? in_data_i[352] : 
                          (N341)? in_data_i[384] : 
                          (N342)? in_data_i[416] : 
                          (N343)? in_data_i[448] : 
                          (N344)? in_data_i_15__0_ : 1'b0;
  assign in_data_o[319] = (N345)? in_data_i[319] : 
                          (N346)? in_data_i[351] : 
                          (N347)? in_data_i[383] : 
                          (N348)? in_data_i[415] : 
                          (N349)? in_data_i[447] : 
                          (N350)? in_data_i[479] : 
                          (N351)? in_data_i_15__31_ : 1'b0;
  assign N345 = N1736;
  assign N346 = N1738;
  assign N347 = N1740;
  assign N348 = N1742;
  assign N349 = N1737;
  assign N350 = N1739;
  assign N351 = N1741;
  assign in_data_o[318] = (N345)? in_data_i[318] : 
                          (N346)? in_data_i[350] : 
                          (N347)? in_data_i[382] : 
                          (N348)? in_data_i[414] : 
                          (N349)? in_data_i[446] : 
                          (N350)? in_data_i[478] : 
                          (N351)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[317] = (N345)? in_data_i[317] : 
                          (N346)? in_data_i[349] : 
                          (N347)? in_data_i[381] : 
                          (N348)? in_data_i[413] : 
                          (N349)? in_data_i[445] : 
                          (N350)? in_data_i[477] : 
                          (N351)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[316] = (N345)? in_data_i[316] : 
                          (N346)? in_data_i[348] : 
                          (N347)? in_data_i[380] : 
                          (N348)? in_data_i[412] : 
                          (N349)? in_data_i[444] : 
                          (N350)? in_data_i[476] : 
                          (N351)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[315] = (N345)? in_data_i[315] : 
                          (N346)? in_data_i[347] : 
                          (N347)? in_data_i[379] : 
                          (N348)? in_data_i[411] : 
                          (N349)? in_data_i[443] : 
                          (N350)? in_data_i[475] : 
                          (N351)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[314] = (N345)? in_data_i[314] : 
                          (N346)? in_data_i[346] : 
                          (N347)? in_data_i[378] : 
                          (N348)? in_data_i[410] : 
                          (N349)? in_data_i[442] : 
                          (N350)? in_data_i[474] : 
                          (N351)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[313] = (N345)? in_data_i[313] : 
                          (N346)? in_data_i[345] : 
                          (N347)? in_data_i[377] : 
                          (N348)? in_data_i[409] : 
                          (N349)? in_data_i[441] : 
                          (N350)? in_data_i[473] : 
                          (N351)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[312] = (N345)? in_data_i[312] : 
                          (N346)? in_data_i[344] : 
                          (N347)? in_data_i[376] : 
                          (N348)? in_data_i[408] : 
                          (N349)? in_data_i[440] : 
                          (N350)? in_data_i[472] : 
                          (N351)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[311] = (N345)? in_data_i[311] : 
                          (N346)? in_data_i[343] : 
                          (N347)? in_data_i[375] : 
                          (N348)? in_data_i[407] : 
                          (N349)? in_data_i[439] : 
                          (N350)? in_data_i[471] : 
                          (N351)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[310] = (N345)? in_data_i[310] : 
                          (N346)? in_data_i[342] : 
                          (N347)? in_data_i[374] : 
                          (N348)? in_data_i[406] : 
                          (N349)? in_data_i[438] : 
                          (N350)? in_data_i[470] : 
                          (N351)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[309] = (N345)? in_data_i[309] : 
                          (N346)? in_data_i[341] : 
                          (N347)? in_data_i[373] : 
                          (N348)? in_data_i[405] : 
                          (N349)? in_data_i[437] : 
                          (N350)? in_data_i[469] : 
                          (N351)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[308] = (N345)? in_data_i[308] : 
                          (N346)? in_data_i[340] : 
                          (N347)? in_data_i[372] : 
                          (N348)? in_data_i[404] : 
                          (N349)? in_data_i[436] : 
                          (N350)? in_data_i[468] : 
                          (N351)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[307] = (N345)? in_data_i[307] : 
                          (N346)? in_data_i[339] : 
                          (N347)? in_data_i[371] : 
                          (N348)? in_data_i[403] : 
                          (N349)? in_data_i[435] : 
                          (N350)? in_data_i[467] : 
                          (N351)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[306] = (N345)? in_data_i[306] : 
                          (N346)? in_data_i[338] : 
                          (N347)? in_data_i[370] : 
                          (N348)? in_data_i[402] : 
                          (N349)? in_data_i[434] : 
                          (N350)? in_data_i[466] : 
                          (N351)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[305] = (N345)? in_data_i[305] : 
                          (N346)? in_data_i[337] : 
                          (N347)? in_data_i[369] : 
                          (N348)? in_data_i[401] : 
                          (N349)? in_data_i[433] : 
                          (N350)? in_data_i[465] : 
                          (N351)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[304] = (N345)? in_data_i[304] : 
                          (N346)? in_data_i[336] : 
                          (N347)? in_data_i[368] : 
                          (N348)? in_data_i[400] : 
                          (N349)? in_data_i[432] : 
                          (N350)? in_data_i[464] : 
                          (N351)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[303] = (N345)? in_data_i[303] : 
                          (N346)? in_data_i[335] : 
                          (N347)? in_data_i[367] : 
                          (N348)? in_data_i[399] : 
                          (N349)? in_data_i[431] : 
                          (N350)? in_data_i[463] : 
                          (N351)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[302] = (N345)? in_data_i[302] : 
                          (N346)? in_data_i[334] : 
                          (N347)? in_data_i[366] : 
                          (N348)? in_data_i[398] : 
                          (N349)? in_data_i[430] : 
                          (N350)? in_data_i[462] : 
                          (N351)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[301] = (N345)? in_data_i[301] : 
                          (N346)? in_data_i[333] : 
                          (N347)? in_data_i[365] : 
                          (N348)? in_data_i[397] : 
                          (N349)? in_data_i[429] : 
                          (N350)? in_data_i[461] : 
                          (N351)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[300] = (N345)? in_data_i[300] : 
                          (N346)? in_data_i[332] : 
                          (N347)? in_data_i[364] : 
                          (N348)? in_data_i[396] : 
                          (N349)? in_data_i[428] : 
                          (N350)? in_data_i[460] : 
                          (N351)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[299] = (N345)? in_data_i[299] : 
                          (N346)? in_data_i[331] : 
                          (N347)? in_data_i[363] : 
                          (N348)? in_data_i[395] : 
                          (N349)? in_data_i[427] : 
                          (N350)? in_data_i[459] : 
                          (N351)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[298] = (N345)? in_data_i[298] : 
                          (N346)? in_data_i[330] : 
                          (N347)? in_data_i[362] : 
                          (N348)? in_data_i[394] : 
                          (N349)? in_data_i[426] : 
                          (N350)? in_data_i[458] : 
                          (N351)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[297] = (N345)? in_data_i[297] : 
                          (N346)? in_data_i[329] : 
                          (N347)? in_data_i[361] : 
                          (N348)? in_data_i[393] : 
                          (N349)? in_data_i[425] : 
                          (N350)? in_data_i[457] : 
                          (N351)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[296] = (N345)? in_data_i[296] : 
                          (N346)? in_data_i[328] : 
                          (N347)? in_data_i[360] : 
                          (N348)? in_data_i[392] : 
                          (N349)? in_data_i[424] : 
                          (N350)? in_data_i[456] : 
                          (N351)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[295] = (N345)? in_data_i[295] : 
                          (N346)? in_data_i[327] : 
                          (N347)? in_data_i[359] : 
                          (N348)? in_data_i[391] : 
                          (N349)? in_data_i[423] : 
                          (N350)? in_data_i[455] : 
                          (N351)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[294] = (N345)? in_data_i[294] : 
                          (N346)? in_data_i[326] : 
                          (N347)? in_data_i[358] : 
                          (N348)? in_data_i[390] : 
                          (N349)? in_data_i[422] : 
                          (N350)? in_data_i[454] : 
                          (N351)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[293] = (N345)? in_data_i[293] : 
                          (N346)? in_data_i[325] : 
                          (N347)? in_data_i[357] : 
                          (N348)? in_data_i[389] : 
                          (N349)? in_data_i[421] : 
                          (N350)? in_data_i[453] : 
                          (N351)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[292] = (N345)? in_data_i[292] : 
                          (N346)? in_data_i[324] : 
                          (N347)? in_data_i[356] : 
                          (N348)? in_data_i[388] : 
                          (N349)? in_data_i[420] : 
                          (N350)? in_data_i[452] : 
                          (N351)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[291] = (N345)? in_data_i[291] : 
                          (N346)? in_data_i[323] : 
                          (N347)? in_data_i[355] : 
                          (N348)? in_data_i[387] : 
                          (N349)? in_data_i[419] : 
                          (N350)? in_data_i[451] : 
                          (N351)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[290] = (N345)? in_data_i[290] : 
                          (N346)? in_data_i[322] : 
                          (N347)? in_data_i[354] : 
                          (N348)? in_data_i[386] : 
                          (N349)? in_data_i[418] : 
                          (N350)? in_data_i[450] : 
                          (N351)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[289] = (N345)? in_data_i[289] : 
                          (N346)? in_data_i[321] : 
                          (N347)? in_data_i[353] : 
                          (N348)? in_data_i[385] : 
                          (N349)? in_data_i[417] : 
                          (N350)? in_data_i[449] : 
                          (N351)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[288] = (N345)? in_data_i[288] : 
                          (N346)? in_data_i[320] : 
                          (N347)? in_data_i[352] : 
                          (N348)? in_data_i[384] : 
                          (N349)? in_data_i[416] : 
                          (N350)? in_data_i[448] : 
                          (N351)? in_data_i_15__0_ : 1'b0;
  assign out_me_data_o[223] = (N352)? out_me_data_i_0__31_ : 
                              (N353)? out_me_data_i[63] : 
                              (N354)? out_me_data_i[95] : 
                              (N355)? out_me_data_i[127] : 
                              (N356)? out_me_data_i[159] : 
                              (N357)? out_me_data_i[191] : 
                              (N358)? out_me_data_i[223] : 1'b0;
  assign N352 = N1419;
  assign N353 = N1421;
  assign N354 = N1423;
  assign N355 = N1425;
  assign N356 = N1420;
  assign N357 = N1422;
  assign N358 = N1424;
  assign out_me_data_o[222] = (N352)? out_me_data_i_0__30_ : 
                              (N353)? out_me_data_i[62] : 
                              (N354)? out_me_data_i[94] : 
                              (N355)? out_me_data_i[126] : 
                              (N356)? out_me_data_i[158] : 
                              (N357)? out_me_data_i[190] : 
                              (N358)? out_me_data_i[222] : 1'b0;
  assign out_me_data_o[221] = (N352)? out_me_data_i_0__29_ : 
                              (N353)? out_me_data_i[61] : 
                              (N354)? out_me_data_i[93] : 
                              (N355)? out_me_data_i[125] : 
                              (N356)? out_me_data_i[157] : 
                              (N357)? out_me_data_i[189] : 
                              (N358)? out_me_data_i[221] : 1'b0;
  assign out_me_data_o[220] = (N352)? out_me_data_i_0__28_ : 
                              (N353)? out_me_data_i[60] : 
                              (N354)? out_me_data_i[92] : 
                              (N355)? out_me_data_i[124] : 
                              (N356)? out_me_data_i[156] : 
                              (N357)? out_me_data_i[188] : 
                              (N358)? out_me_data_i[220] : 1'b0;
  assign out_me_data_o[219] = (N352)? out_me_data_i_0__27_ : 
                              (N353)? out_me_data_i[59] : 
                              (N354)? out_me_data_i[91] : 
                              (N355)? out_me_data_i[123] : 
                              (N356)? out_me_data_i[155] : 
                              (N357)? out_me_data_i[187] : 
                              (N358)? out_me_data_i[219] : 1'b0;
  assign out_me_data_o[218] = (N352)? out_me_data_i_0__26_ : 
                              (N353)? out_me_data_i[58] : 
                              (N354)? out_me_data_i[90] : 
                              (N355)? out_me_data_i[122] : 
                              (N356)? out_me_data_i[154] : 
                              (N357)? out_me_data_i[186] : 
                              (N358)? out_me_data_i[218] : 1'b0;
  assign out_me_data_o[217] = (N352)? out_me_data_i_0__25_ : 
                              (N353)? out_me_data_i[57] : 
                              (N354)? out_me_data_i[89] : 
                              (N355)? out_me_data_i[121] : 
                              (N356)? out_me_data_i[153] : 
                              (N357)? out_me_data_i[185] : 
                              (N358)? out_me_data_i[217] : 1'b0;
  assign out_me_data_o[216] = (N352)? out_me_data_i_0__24_ : 
                              (N353)? out_me_data_i[56] : 
                              (N354)? out_me_data_i[88] : 
                              (N355)? out_me_data_i[120] : 
                              (N356)? out_me_data_i[152] : 
                              (N357)? out_me_data_i[184] : 
                              (N358)? out_me_data_i[216] : 1'b0;
  assign out_me_data_o[215] = (N352)? out_me_data_i_0__23_ : 
                              (N353)? out_me_data_i[55] : 
                              (N354)? out_me_data_i[87] : 
                              (N355)? out_me_data_i[119] : 
                              (N356)? out_me_data_i[151] : 
                              (N357)? out_me_data_i[183] : 
                              (N358)? out_me_data_i[215] : 1'b0;
  assign out_me_data_o[214] = (N352)? out_me_data_i_0__22_ : 
                              (N353)? out_me_data_i[54] : 
                              (N354)? out_me_data_i[86] : 
                              (N355)? out_me_data_i[118] : 
                              (N356)? out_me_data_i[150] : 
                              (N357)? out_me_data_i[182] : 
                              (N358)? out_me_data_i[214] : 1'b0;
  assign out_me_data_o[213] = (N352)? out_me_data_i_0__21_ : 
                              (N353)? out_me_data_i[53] : 
                              (N354)? out_me_data_i[85] : 
                              (N355)? out_me_data_i[117] : 
                              (N356)? out_me_data_i[149] : 
                              (N357)? out_me_data_i[181] : 
                              (N358)? out_me_data_i[213] : 1'b0;
  assign out_me_data_o[212] = (N352)? out_me_data_i_0__20_ : 
                              (N353)? out_me_data_i[52] : 
                              (N354)? out_me_data_i[84] : 
                              (N355)? out_me_data_i[116] : 
                              (N356)? out_me_data_i[148] : 
                              (N357)? out_me_data_i[180] : 
                              (N358)? out_me_data_i[212] : 1'b0;
  assign out_me_data_o[211] = (N352)? out_me_data_i_0__19_ : 
                              (N353)? out_me_data_i[51] : 
                              (N354)? out_me_data_i[83] : 
                              (N355)? out_me_data_i[115] : 
                              (N356)? out_me_data_i[147] : 
                              (N357)? out_me_data_i[179] : 
                              (N358)? out_me_data_i[211] : 1'b0;
  assign out_me_data_o[210] = (N352)? out_me_data_i_0__18_ : 
                              (N353)? out_me_data_i[50] : 
                              (N354)? out_me_data_i[82] : 
                              (N355)? out_me_data_i[114] : 
                              (N356)? out_me_data_i[146] : 
                              (N357)? out_me_data_i[178] : 
                              (N358)? out_me_data_i[210] : 1'b0;
  assign out_me_data_o[209] = (N352)? out_me_data_i_0__17_ : 
                              (N353)? out_me_data_i[49] : 
                              (N354)? out_me_data_i[81] : 
                              (N355)? out_me_data_i[113] : 
                              (N356)? out_me_data_i[145] : 
                              (N357)? out_me_data_i[177] : 
                              (N358)? out_me_data_i[209] : 1'b0;
  assign out_me_data_o[208] = (N352)? out_me_data_i_0__16_ : 
                              (N353)? out_me_data_i[48] : 
                              (N354)? out_me_data_i[80] : 
                              (N355)? out_me_data_i[112] : 
                              (N356)? out_me_data_i[144] : 
                              (N357)? out_me_data_i[176] : 
                              (N358)? out_me_data_i[208] : 1'b0;
  assign out_me_data_o[207] = (N352)? out_me_data_i_0__15_ : 
                              (N353)? out_me_data_i[47] : 
                              (N354)? out_me_data_i[79] : 
                              (N355)? out_me_data_i[111] : 
                              (N356)? out_me_data_i[143] : 
                              (N357)? out_me_data_i[175] : 
                              (N358)? out_me_data_i[207] : 1'b0;
  assign out_me_data_o[206] = (N352)? out_me_data_i_0__14_ : 
                              (N353)? out_me_data_i[46] : 
                              (N354)? out_me_data_i[78] : 
                              (N355)? out_me_data_i[110] : 
                              (N356)? out_me_data_i[142] : 
                              (N357)? out_me_data_i[174] : 
                              (N358)? out_me_data_i[206] : 1'b0;
  assign out_me_data_o[205] = (N352)? out_me_data_i_0__13_ : 
                              (N353)? out_me_data_i[45] : 
                              (N354)? out_me_data_i[77] : 
                              (N355)? out_me_data_i[109] : 
                              (N356)? out_me_data_i[141] : 
                              (N357)? out_me_data_i[173] : 
                              (N358)? out_me_data_i[205] : 1'b0;
  assign out_me_data_o[204] = (N352)? out_me_data_i_0__12_ : 
                              (N353)? out_me_data_i[44] : 
                              (N354)? out_me_data_i[76] : 
                              (N355)? out_me_data_i[108] : 
                              (N356)? out_me_data_i[140] : 
                              (N357)? out_me_data_i[172] : 
                              (N358)? out_me_data_i[204] : 1'b0;
  assign out_me_data_o[203] = (N352)? out_me_data_i_0__11_ : 
                              (N353)? out_me_data_i[43] : 
                              (N354)? out_me_data_i[75] : 
                              (N355)? out_me_data_i[107] : 
                              (N356)? out_me_data_i[139] : 
                              (N357)? out_me_data_i[171] : 
                              (N358)? out_me_data_i[203] : 1'b0;
  assign out_me_data_o[202] = (N352)? out_me_data_i_0__10_ : 
                              (N353)? out_me_data_i[42] : 
                              (N354)? out_me_data_i[74] : 
                              (N355)? out_me_data_i[106] : 
                              (N356)? out_me_data_i[138] : 
                              (N357)? out_me_data_i[170] : 
                              (N358)? out_me_data_i[202] : 1'b0;
  assign out_me_data_o[201] = (N352)? out_me_data_i_0__9_ : 
                              (N353)? out_me_data_i[41] : 
                              (N354)? out_me_data_i[73] : 
                              (N355)? out_me_data_i[105] : 
                              (N356)? out_me_data_i[137] : 
                              (N357)? out_me_data_i[169] : 
                              (N358)? out_me_data_i[201] : 1'b0;
  assign out_me_data_o[200] = (N352)? out_me_data_i_0__8_ : 
                              (N353)? out_me_data_i[40] : 
                              (N354)? out_me_data_i[72] : 
                              (N355)? out_me_data_i[104] : 
                              (N356)? out_me_data_i[136] : 
                              (N357)? out_me_data_i[168] : 
                              (N358)? out_me_data_i[200] : 1'b0;
  assign out_me_data_o[199] = (N352)? out_me_data_i_0__7_ : 
                              (N353)? out_me_data_i[39] : 
                              (N354)? out_me_data_i[71] : 
                              (N355)? out_me_data_i[103] : 
                              (N356)? out_me_data_i[135] : 
                              (N357)? out_me_data_i[167] : 
                              (N358)? out_me_data_i[199] : 1'b0;
  assign out_me_data_o[198] = (N352)? out_me_data_i_0__6_ : 
                              (N353)? out_me_data_i[38] : 
                              (N354)? out_me_data_i[70] : 
                              (N355)? out_me_data_i[102] : 
                              (N356)? out_me_data_i[134] : 
                              (N357)? out_me_data_i[166] : 
                              (N358)? out_me_data_i[198] : 1'b0;
  assign out_me_data_o[197] = (N352)? out_me_data_i_0__5_ : 
                              (N353)? out_me_data_i[37] : 
                              (N354)? out_me_data_i[69] : 
                              (N355)? out_me_data_i[101] : 
                              (N356)? out_me_data_i[133] : 
                              (N357)? out_me_data_i[165] : 
                              (N358)? out_me_data_i[197] : 1'b0;
  assign out_me_data_o[196] = (N352)? out_me_data_i_0__4_ : 
                              (N353)? out_me_data_i[36] : 
                              (N354)? out_me_data_i[68] : 
                              (N355)? out_me_data_i[100] : 
                              (N356)? out_me_data_i[132] : 
                              (N357)? out_me_data_i[164] : 
                              (N358)? out_me_data_i[196] : 1'b0;
  assign out_me_data_o[195] = (N352)? out_me_data_i_0__3_ : 
                              (N353)? out_me_data_i[35] : 
                              (N354)? out_me_data_i[67] : 
                              (N355)? out_me_data_i[99] : 
                              (N356)? out_me_data_i[131] : 
                              (N357)? out_me_data_i[163] : 
                              (N358)? out_me_data_i[195] : 1'b0;
  assign out_me_data_o[194] = (N352)? out_me_data_i_0__2_ : 
                              (N353)? out_me_data_i[34] : 
                              (N354)? out_me_data_i[66] : 
                              (N355)? out_me_data_i[98] : 
                              (N356)? out_me_data_i[130] : 
                              (N357)? out_me_data_i[162] : 
                              (N358)? out_me_data_i[194] : 1'b0;
  assign out_me_data_o[193] = (N352)? out_me_data_i_0__1_ : 
                              (N353)? out_me_data_i[33] : 
                              (N354)? out_me_data_i[65] : 
                              (N355)? out_me_data_i[97] : 
                              (N356)? out_me_data_i[129] : 
                              (N357)? out_me_data_i[161] : 
                              (N358)? out_me_data_i[193] : 1'b0;
  assign out_me_data_o[192] = (N352)? out_me_data_i_0__0_ : 
                              (N353)? out_me_data_i[32] : 
                              (N354)? out_me_data_i[64] : 
                              (N355)? out_me_data_i[96] : 
                              (N356)? out_me_data_i[128] : 
                              (N357)? out_me_data_i[160] : 
                              (N358)? out_me_data_i[192] : 1'b0;
  assign out_me_data_o[191] = (N359)? out_me_data_i_0__31_ : 
                              (N360)? out_me_data_i[63] : 
                              (N361)? out_me_data_i[95] : 
                              (N362)? out_me_data_i[127] : 
                              (N363)? out_me_data_i[159] : 
                              (N364)? out_me_data_i[191] : 1'b0;
  assign N359 = N1295;
  assign N360 = N1297;
  assign N361 = N1299;
  assign N362 = N1300;
  assign N363 = N1296;
  assign N364 = N1298;
  assign out_me_data_o[190] = (N359)? out_me_data_i_0__30_ : 
                              (N360)? out_me_data_i[62] : 
                              (N361)? out_me_data_i[94] : 
                              (N362)? out_me_data_i[126] : 
                              (N363)? out_me_data_i[158] : 
                              (N364)? out_me_data_i[190] : 1'b0;
  assign out_me_data_o[189] = (N359)? out_me_data_i_0__29_ : 
                              (N360)? out_me_data_i[61] : 
                              (N361)? out_me_data_i[93] : 
                              (N362)? out_me_data_i[125] : 
                              (N363)? out_me_data_i[157] : 
                              (N364)? out_me_data_i[189] : 1'b0;
  assign out_me_data_o[188] = (N359)? out_me_data_i_0__28_ : 
                              (N360)? out_me_data_i[60] : 
                              (N361)? out_me_data_i[92] : 
                              (N362)? out_me_data_i[124] : 
                              (N363)? out_me_data_i[156] : 
                              (N364)? out_me_data_i[188] : 1'b0;
  assign out_me_data_o[187] = (N359)? out_me_data_i_0__27_ : 
                              (N360)? out_me_data_i[59] : 
                              (N361)? out_me_data_i[91] : 
                              (N362)? out_me_data_i[123] : 
                              (N363)? out_me_data_i[155] : 
                              (N364)? out_me_data_i[187] : 1'b0;
  assign out_me_data_o[186] = (N359)? out_me_data_i_0__26_ : 
                              (N360)? out_me_data_i[58] : 
                              (N361)? out_me_data_i[90] : 
                              (N362)? out_me_data_i[122] : 
                              (N363)? out_me_data_i[154] : 
                              (N364)? out_me_data_i[186] : 1'b0;
  assign out_me_data_o[185] = (N359)? out_me_data_i_0__25_ : 
                              (N360)? out_me_data_i[57] : 
                              (N361)? out_me_data_i[89] : 
                              (N362)? out_me_data_i[121] : 
                              (N363)? out_me_data_i[153] : 
                              (N364)? out_me_data_i[185] : 1'b0;
  assign out_me_data_o[184] = (N359)? out_me_data_i_0__24_ : 
                              (N360)? out_me_data_i[56] : 
                              (N361)? out_me_data_i[88] : 
                              (N362)? out_me_data_i[120] : 
                              (N363)? out_me_data_i[152] : 
                              (N364)? out_me_data_i[184] : 1'b0;
  assign out_me_data_o[183] = (N359)? out_me_data_i_0__23_ : 
                              (N360)? out_me_data_i[55] : 
                              (N361)? out_me_data_i[87] : 
                              (N362)? out_me_data_i[119] : 
                              (N363)? out_me_data_i[151] : 
                              (N364)? out_me_data_i[183] : 1'b0;
  assign out_me_data_o[182] = (N359)? out_me_data_i_0__22_ : 
                              (N360)? out_me_data_i[54] : 
                              (N361)? out_me_data_i[86] : 
                              (N362)? out_me_data_i[118] : 
                              (N363)? out_me_data_i[150] : 
                              (N364)? out_me_data_i[182] : 1'b0;
  assign out_me_data_o[181] = (N359)? out_me_data_i_0__21_ : 
                              (N360)? out_me_data_i[53] : 
                              (N361)? out_me_data_i[85] : 
                              (N362)? out_me_data_i[117] : 
                              (N363)? out_me_data_i[149] : 
                              (N364)? out_me_data_i[181] : 1'b0;
  assign out_me_data_o[180] = (N359)? out_me_data_i_0__20_ : 
                              (N360)? out_me_data_i[52] : 
                              (N361)? out_me_data_i[84] : 
                              (N362)? out_me_data_i[116] : 
                              (N363)? out_me_data_i[148] : 
                              (N364)? out_me_data_i[180] : 1'b0;
  assign out_me_data_o[179] = (N359)? out_me_data_i_0__19_ : 
                              (N360)? out_me_data_i[51] : 
                              (N361)? out_me_data_i[83] : 
                              (N362)? out_me_data_i[115] : 
                              (N363)? out_me_data_i[147] : 
                              (N364)? out_me_data_i[179] : 1'b0;
  assign out_me_data_o[178] = (N359)? out_me_data_i_0__18_ : 
                              (N360)? out_me_data_i[50] : 
                              (N361)? out_me_data_i[82] : 
                              (N362)? out_me_data_i[114] : 
                              (N363)? out_me_data_i[146] : 
                              (N364)? out_me_data_i[178] : 1'b0;
  assign out_me_data_o[177] = (N359)? out_me_data_i_0__17_ : 
                              (N360)? out_me_data_i[49] : 
                              (N361)? out_me_data_i[81] : 
                              (N362)? out_me_data_i[113] : 
                              (N363)? out_me_data_i[145] : 
                              (N364)? out_me_data_i[177] : 1'b0;
  assign out_me_data_o[176] = (N359)? out_me_data_i_0__16_ : 
                              (N360)? out_me_data_i[48] : 
                              (N361)? out_me_data_i[80] : 
                              (N362)? out_me_data_i[112] : 
                              (N363)? out_me_data_i[144] : 
                              (N364)? out_me_data_i[176] : 1'b0;
  assign out_me_data_o[175] = (N359)? out_me_data_i_0__15_ : 
                              (N360)? out_me_data_i[47] : 
                              (N361)? out_me_data_i[79] : 
                              (N362)? out_me_data_i[111] : 
                              (N363)? out_me_data_i[143] : 
                              (N364)? out_me_data_i[175] : 1'b0;
  assign out_me_data_o[174] = (N359)? out_me_data_i_0__14_ : 
                              (N360)? out_me_data_i[46] : 
                              (N361)? out_me_data_i[78] : 
                              (N362)? out_me_data_i[110] : 
                              (N363)? out_me_data_i[142] : 
                              (N364)? out_me_data_i[174] : 1'b0;
  assign out_me_data_o[173] = (N359)? out_me_data_i_0__13_ : 
                              (N360)? out_me_data_i[45] : 
                              (N361)? out_me_data_i[77] : 
                              (N362)? out_me_data_i[109] : 
                              (N363)? out_me_data_i[141] : 
                              (N364)? out_me_data_i[173] : 1'b0;
  assign out_me_data_o[172] = (N359)? out_me_data_i_0__12_ : 
                              (N360)? out_me_data_i[44] : 
                              (N361)? out_me_data_i[76] : 
                              (N362)? out_me_data_i[108] : 
                              (N363)? out_me_data_i[140] : 
                              (N364)? out_me_data_i[172] : 1'b0;
  assign out_me_data_o[171] = (N359)? out_me_data_i_0__11_ : 
                              (N360)? out_me_data_i[43] : 
                              (N361)? out_me_data_i[75] : 
                              (N362)? out_me_data_i[107] : 
                              (N363)? out_me_data_i[139] : 
                              (N364)? out_me_data_i[171] : 1'b0;
  assign out_me_data_o[170] = (N359)? out_me_data_i_0__10_ : 
                              (N360)? out_me_data_i[42] : 
                              (N361)? out_me_data_i[74] : 
                              (N362)? out_me_data_i[106] : 
                              (N363)? out_me_data_i[138] : 
                              (N364)? out_me_data_i[170] : 1'b0;
  assign out_me_data_o[169] = (N359)? out_me_data_i_0__9_ : 
                              (N360)? out_me_data_i[41] : 
                              (N361)? out_me_data_i[73] : 
                              (N362)? out_me_data_i[105] : 
                              (N363)? out_me_data_i[137] : 
                              (N364)? out_me_data_i[169] : 1'b0;
  assign out_me_data_o[168] = (N359)? out_me_data_i_0__8_ : 
                              (N360)? out_me_data_i[40] : 
                              (N361)? out_me_data_i[72] : 
                              (N362)? out_me_data_i[104] : 
                              (N363)? out_me_data_i[136] : 
                              (N364)? out_me_data_i[168] : 1'b0;
  assign out_me_data_o[167] = (N359)? out_me_data_i_0__7_ : 
                              (N360)? out_me_data_i[39] : 
                              (N361)? out_me_data_i[71] : 
                              (N362)? out_me_data_i[103] : 
                              (N363)? out_me_data_i[135] : 
                              (N364)? out_me_data_i[167] : 1'b0;
  assign out_me_data_o[166] = (N359)? out_me_data_i_0__6_ : 
                              (N360)? out_me_data_i[38] : 
                              (N361)? out_me_data_i[70] : 
                              (N362)? out_me_data_i[102] : 
                              (N363)? out_me_data_i[134] : 
                              (N364)? out_me_data_i[166] : 1'b0;
  assign out_me_data_o[165] = (N359)? out_me_data_i_0__5_ : 
                              (N360)? out_me_data_i[37] : 
                              (N361)? out_me_data_i[69] : 
                              (N362)? out_me_data_i[101] : 
                              (N363)? out_me_data_i[133] : 
                              (N364)? out_me_data_i[165] : 1'b0;
  assign out_me_data_o[164] = (N359)? out_me_data_i_0__4_ : 
                              (N360)? out_me_data_i[36] : 
                              (N361)? out_me_data_i[68] : 
                              (N362)? out_me_data_i[100] : 
                              (N363)? out_me_data_i[132] : 
                              (N364)? out_me_data_i[164] : 1'b0;
  assign out_me_data_o[163] = (N359)? out_me_data_i_0__3_ : 
                              (N360)? out_me_data_i[35] : 
                              (N361)? out_me_data_i[67] : 
                              (N362)? out_me_data_i[99] : 
                              (N363)? out_me_data_i[131] : 
                              (N364)? out_me_data_i[163] : 1'b0;
  assign out_me_data_o[162] = (N359)? out_me_data_i_0__2_ : 
                              (N360)? out_me_data_i[34] : 
                              (N361)? out_me_data_i[66] : 
                              (N362)? out_me_data_i[98] : 
                              (N363)? out_me_data_i[130] : 
                              (N364)? out_me_data_i[162] : 1'b0;
  assign out_me_data_o[161] = (N359)? out_me_data_i_0__1_ : 
                              (N360)? out_me_data_i[33] : 
                              (N361)? out_me_data_i[65] : 
                              (N362)? out_me_data_i[97] : 
                              (N363)? out_me_data_i[129] : 
                              (N364)? out_me_data_i[161] : 1'b0;
  assign out_me_data_o[160] = (N359)? out_me_data_i_0__0_ : 
                              (N360)? out_me_data_i[32] : 
                              (N361)? out_me_data_i[64] : 
                              (N362)? out_me_data_i[96] : 
                              (N363)? out_me_data_i[128] : 
                              (N364)? out_me_data_i[160] : 1'b0;
  assign out_me_data_o[159] = (N365)? out_me_data_i_0__31_ : 
                              (N366)? out_me_data_i[63] : 
                              (N367)? out_me_data_i[95] : 
                              (N368)? out_me_data_i[127] : 
                              (N369)? out_me_data_i[159] : 1'b0;
  assign N365 = N1172;
  assign N366 = N1173;
  assign N367 = N1174;
  assign N368 = N1175;
  assign N369 = bk_dpath_sel_r_18;
  assign out_me_data_o[158] = (N365)? out_me_data_i_0__30_ : 
                              (N366)? out_me_data_i[62] : 
                              (N367)? out_me_data_i[94] : 
                              (N368)? out_me_data_i[126] : 
                              (N369)? out_me_data_i[158] : 1'b0;
  assign out_me_data_o[157] = (N365)? out_me_data_i_0__29_ : 
                              (N366)? out_me_data_i[61] : 
                              (N367)? out_me_data_i[93] : 
                              (N368)? out_me_data_i[125] : 
                              (N369)? out_me_data_i[157] : 1'b0;
  assign out_me_data_o[156] = (N365)? out_me_data_i_0__28_ : 
                              (N366)? out_me_data_i[60] : 
                              (N367)? out_me_data_i[92] : 
                              (N368)? out_me_data_i[124] : 
                              (N369)? out_me_data_i[156] : 1'b0;
  assign out_me_data_o[155] = (N365)? out_me_data_i_0__27_ : 
                              (N366)? out_me_data_i[59] : 
                              (N367)? out_me_data_i[91] : 
                              (N368)? out_me_data_i[123] : 
                              (N369)? out_me_data_i[155] : 1'b0;
  assign out_me_data_o[154] = (N365)? out_me_data_i_0__26_ : 
                              (N366)? out_me_data_i[58] : 
                              (N367)? out_me_data_i[90] : 
                              (N368)? out_me_data_i[122] : 
                              (N369)? out_me_data_i[154] : 1'b0;
  assign out_me_data_o[153] = (N365)? out_me_data_i_0__25_ : 
                              (N366)? out_me_data_i[57] : 
                              (N367)? out_me_data_i[89] : 
                              (N368)? out_me_data_i[121] : 
                              (N369)? out_me_data_i[153] : 1'b0;
  assign out_me_data_o[152] = (N365)? out_me_data_i_0__24_ : 
                              (N366)? out_me_data_i[56] : 
                              (N367)? out_me_data_i[88] : 
                              (N368)? out_me_data_i[120] : 
                              (N369)? out_me_data_i[152] : 1'b0;
  assign out_me_data_o[151] = (N365)? out_me_data_i_0__23_ : 
                              (N366)? out_me_data_i[55] : 
                              (N367)? out_me_data_i[87] : 
                              (N368)? out_me_data_i[119] : 
                              (N369)? out_me_data_i[151] : 1'b0;
  assign out_me_data_o[150] = (N365)? out_me_data_i_0__22_ : 
                              (N366)? out_me_data_i[54] : 
                              (N367)? out_me_data_i[86] : 
                              (N368)? out_me_data_i[118] : 
                              (N369)? out_me_data_i[150] : 1'b0;
  assign out_me_data_o[149] = (N365)? out_me_data_i_0__21_ : 
                              (N366)? out_me_data_i[53] : 
                              (N367)? out_me_data_i[85] : 
                              (N368)? out_me_data_i[117] : 
                              (N369)? out_me_data_i[149] : 1'b0;
  assign out_me_data_o[148] = (N365)? out_me_data_i_0__20_ : 
                              (N366)? out_me_data_i[52] : 
                              (N367)? out_me_data_i[84] : 
                              (N368)? out_me_data_i[116] : 
                              (N369)? out_me_data_i[148] : 1'b0;
  assign out_me_data_o[147] = (N365)? out_me_data_i_0__19_ : 
                              (N366)? out_me_data_i[51] : 
                              (N367)? out_me_data_i[83] : 
                              (N368)? out_me_data_i[115] : 
                              (N369)? out_me_data_i[147] : 1'b0;
  assign out_me_data_o[146] = (N365)? out_me_data_i_0__18_ : 
                              (N366)? out_me_data_i[50] : 
                              (N367)? out_me_data_i[82] : 
                              (N368)? out_me_data_i[114] : 
                              (N369)? out_me_data_i[146] : 1'b0;
  assign out_me_data_o[145] = (N365)? out_me_data_i_0__17_ : 
                              (N366)? out_me_data_i[49] : 
                              (N367)? out_me_data_i[81] : 
                              (N368)? out_me_data_i[113] : 
                              (N369)? out_me_data_i[145] : 1'b0;
  assign out_me_data_o[144] = (N365)? out_me_data_i_0__16_ : 
                              (N366)? out_me_data_i[48] : 
                              (N367)? out_me_data_i[80] : 
                              (N368)? out_me_data_i[112] : 
                              (N369)? out_me_data_i[144] : 1'b0;
  assign out_me_data_o[143] = (N365)? out_me_data_i_0__15_ : 
                              (N366)? out_me_data_i[47] : 
                              (N367)? out_me_data_i[79] : 
                              (N368)? out_me_data_i[111] : 
                              (N369)? out_me_data_i[143] : 1'b0;
  assign out_me_data_o[142] = (N365)? out_me_data_i_0__14_ : 
                              (N366)? out_me_data_i[46] : 
                              (N367)? out_me_data_i[78] : 
                              (N368)? out_me_data_i[110] : 
                              (N369)? out_me_data_i[142] : 1'b0;
  assign out_me_data_o[141] = (N365)? out_me_data_i_0__13_ : 
                              (N366)? out_me_data_i[45] : 
                              (N367)? out_me_data_i[77] : 
                              (N368)? out_me_data_i[109] : 
                              (N369)? out_me_data_i[141] : 1'b0;
  assign out_me_data_o[140] = (N365)? out_me_data_i_0__12_ : 
                              (N366)? out_me_data_i[44] : 
                              (N367)? out_me_data_i[76] : 
                              (N368)? out_me_data_i[108] : 
                              (N369)? out_me_data_i[140] : 1'b0;
  assign out_me_data_o[139] = (N365)? out_me_data_i_0__11_ : 
                              (N366)? out_me_data_i[43] : 
                              (N367)? out_me_data_i[75] : 
                              (N368)? out_me_data_i[107] : 
                              (N369)? out_me_data_i[139] : 1'b0;
  assign out_me_data_o[138] = (N365)? out_me_data_i_0__10_ : 
                              (N366)? out_me_data_i[42] : 
                              (N367)? out_me_data_i[74] : 
                              (N368)? out_me_data_i[106] : 
                              (N369)? out_me_data_i[138] : 1'b0;
  assign out_me_data_o[137] = (N365)? out_me_data_i_0__9_ : 
                              (N366)? out_me_data_i[41] : 
                              (N367)? out_me_data_i[73] : 
                              (N368)? out_me_data_i[105] : 
                              (N369)? out_me_data_i[137] : 1'b0;
  assign out_me_data_o[136] = (N365)? out_me_data_i_0__8_ : 
                              (N366)? out_me_data_i[40] : 
                              (N367)? out_me_data_i[72] : 
                              (N368)? out_me_data_i[104] : 
                              (N369)? out_me_data_i[136] : 1'b0;
  assign out_me_data_o[135] = (N365)? out_me_data_i_0__7_ : 
                              (N366)? out_me_data_i[39] : 
                              (N367)? out_me_data_i[71] : 
                              (N368)? out_me_data_i[103] : 
                              (N369)? out_me_data_i[135] : 1'b0;
  assign out_me_data_o[134] = (N365)? out_me_data_i_0__6_ : 
                              (N366)? out_me_data_i[38] : 
                              (N367)? out_me_data_i[70] : 
                              (N368)? out_me_data_i[102] : 
                              (N369)? out_me_data_i[134] : 1'b0;
  assign out_me_data_o[133] = (N365)? out_me_data_i_0__5_ : 
                              (N366)? out_me_data_i[37] : 
                              (N367)? out_me_data_i[69] : 
                              (N368)? out_me_data_i[101] : 
                              (N369)? out_me_data_i[133] : 1'b0;
  assign out_me_data_o[132] = (N365)? out_me_data_i_0__4_ : 
                              (N366)? out_me_data_i[36] : 
                              (N367)? out_me_data_i[68] : 
                              (N368)? out_me_data_i[100] : 
                              (N369)? out_me_data_i[132] : 1'b0;
  assign out_me_data_o[131] = (N365)? out_me_data_i_0__3_ : 
                              (N366)? out_me_data_i[35] : 
                              (N367)? out_me_data_i[67] : 
                              (N368)? out_me_data_i[99] : 
                              (N369)? out_me_data_i[131] : 1'b0;
  assign out_me_data_o[130] = (N365)? out_me_data_i_0__2_ : 
                              (N366)? out_me_data_i[34] : 
                              (N367)? out_me_data_i[66] : 
                              (N368)? out_me_data_i[98] : 
                              (N369)? out_me_data_i[130] : 1'b0;
  assign out_me_data_o[129] = (N365)? out_me_data_i_0__1_ : 
                              (N366)? out_me_data_i[33] : 
                              (N367)? out_me_data_i[65] : 
                              (N368)? out_me_data_i[97] : 
                              (N369)? out_me_data_i[129] : 1'b0;
  assign out_me_data_o[128] = (N365)? out_me_data_i_0__0_ : 
                              (N366)? out_me_data_i[32] : 
                              (N367)? out_me_data_i[64] : 
                              (N368)? out_me_data_i[96] : 
                              (N369)? out_me_data_i[128] : 1'b0;
  assign in_data_o[255] = (N370)? in_data_i[255] : 
                          (N371)? in_data_i[287] : 
                          (N372)? in_data_i[319] : 
                          (N373)? in_data_i[351] : 
                          (N374)? in_data_i[383] : 
                          (N375)? in_data_i[415] : 
                          (N376)? in_data_i[447] : 
                          (N377)? in_data_i[479] : 
                          (N378)? in_data_i_15__31_ : 1'b0;
  assign N370 = N1474;
  assign N371 = N1475;
  assign N372 = N1476;
  assign N373 = N1477;
  assign N374 = N1478;
  assign N375 = N1479;
  assign N376 = N1480;
  assign N377 = N1481;
  assign N378 = fwd_dpath_sel_r[31];
  assign in_data_o[254] = (N370)? in_data_i[254] : 
                          (N371)? in_data_i[286] : 
                          (N372)? in_data_i[318] : 
                          (N373)? in_data_i[350] : 
                          (N374)? in_data_i[382] : 
                          (N375)? in_data_i[414] : 
                          (N376)? in_data_i[446] : 
                          (N377)? in_data_i[478] : 
                          (N378)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[253] = (N370)? in_data_i[253] : 
                          (N371)? in_data_i[285] : 
                          (N372)? in_data_i[317] : 
                          (N373)? in_data_i[349] : 
                          (N374)? in_data_i[381] : 
                          (N375)? in_data_i[413] : 
                          (N376)? in_data_i[445] : 
                          (N377)? in_data_i[477] : 
                          (N378)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[252] = (N370)? in_data_i[252] : 
                          (N371)? in_data_i[284] : 
                          (N372)? in_data_i[316] : 
                          (N373)? in_data_i[348] : 
                          (N374)? in_data_i[380] : 
                          (N375)? in_data_i[412] : 
                          (N376)? in_data_i[444] : 
                          (N377)? in_data_i[476] : 
                          (N378)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[251] = (N370)? in_data_i[251] : 
                          (N371)? in_data_i[283] : 
                          (N372)? in_data_i[315] : 
                          (N373)? in_data_i[347] : 
                          (N374)? in_data_i[379] : 
                          (N375)? in_data_i[411] : 
                          (N376)? in_data_i[443] : 
                          (N377)? in_data_i[475] : 
                          (N378)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[250] = (N370)? in_data_i[250] : 
                          (N371)? in_data_i[282] : 
                          (N372)? in_data_i[314] : 
                          (N373)? in_data_i[346] : 
                          (N374)? in_data_i[378] : 
                          (N375)? in_data_i[410] : 
                          (N376)? in_data_i[442] : 
                          (N377)? in_data_i[474] : 
                          (N378)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[249] = (N370)? in_data_i[249] : 
                          (N371)? in_data_i[281] : 
                          (N372)? in_data_i[313] : 
                          (N373)? in_data_i[345] : 
                          (N374)? in_data_i[377] : 
                          (N375)? in_data_i[409] : 
                          (N376)? in_data_i[441] : 
                          (N377)? in_data_i[473] : 
                          (N378)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[248] = (N370)? in_data_i[248] : 
                          (N371)? in_data_i[280] : 
                          (N372)? in_data_i[312] : 
                          (N373)? in_data_i[344] : 
                          (N374)? in_data_i[376] : 
                          (N375)? in_data_i[408] : 
                          (N376)? in_data_i[440] : 
                          (N377)? in_data_i[472] : 
                          (N378)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[247] = (N370)? in_data_i[247] : 
                          (N371)? in_data_i[279] : 
                          (N372)? in_data_i[311] : 
                          (N373)? in_data_i[343] : 
                          (N374)? in_data_i[375] : 
                          (N375)? in_data_i[407] : 
                          (N376)? in_data_i[439] : 
                          (N377)? in_data_i[471] : 
                          (N378)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[246] = (N370)? in_data_i[246] : 
                          (N371)? in_data_i[278] : 
                          (N372)? in_data_i[310] : 
                          (N373)? in_data_i[342] : 
                          (N374)? in_data_i[374] : 
                          (N375)? in_data_i[406] : 
                          (N376)? in_data_i[438] : 
                          (N377)? in_data_i[470] : 
                          (N378)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[245] = (N370)? in_data_i[245] : 
                          (N371)? in_data_i[277] : 
                          (N372)? in_data_i[309] : 
                          (N373)? in_data_i[341] : 
                          (N374)? in_data_i[373] : 
                          (N375)? in_data_i[405] : 
                          (N376)? in_data_i[437] : 
                          (N377)? in_data_i[469] : 
                          (N378)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[244] = (N370)? in_data_i[244] : 
                          (N371)? in_data_i[276] : 
                          (N372)? in_data_i[308] : 
                          (N373)? in_data_i[340] : 
                          (N374)? in_data_i[372] : 
                          (N375)? in_data_i[404] : 
                          (N376)? in_data_i[436] : 
                          (N377)? in_data_i[468] : 
                          (N378)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[243] = (N370)? in_data_i[243] : 
                          (N371)? in_data_i[275] : 
                          (N372)? in_data_i[307] : 
                          (N373)? in_data_i[339] : 
                          (N374)? in_data_i[371] : 
                          (N375)? in_data_i[403] : 
                          (N376)? in_data_i[435] : 
                          (N377)? in_data_i[467] : 
                          (N378)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[242] = (N370)? in_data_i[242] : 
                          (N371)? in_data_i[274] : 
                          (N372)? in_data_i[306] : 
                          (N373)? in_data_i[338] : 
                          (N374)? in_data_i[370] : 
                          (N375)? in_data_i[402] : 
                          (N376)? in_data_i[434] : 
                          (N377)? in_data_i[466] : 
                          (N378)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[241] = (N370)? in_data_i[241] : 
                          (N371)? in_data_i[273] : 
                          (N372)? in_data_i[305] : 
                          (N373)? in_data_i[337] : 
                          (N374)? in_data_i[369] : 
                          (N375)? in_data_i[401] : 
                          (N376)? in_data_i[433] : 
                          (N377)? in_data_i[465] : 
                          (N378)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[240] = (N370)? in_data_i[240] : 
                          (N371)? in_data_i[272] : 
                          (N372)? in_data_i[304] : 
                          (N373)? in_data_i[336] : 
                          (N374)? in_data_i[368] : 
                          (N375)? in_data_i[400] : 
                          (N376)? in_data_i[432] : 
                          (N377)? in_data_i[464] : 
                          (N378)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[239] = (N370)? in_data_i[239] : 
                          (N371)? in_data_i[271] : 
                          (N372)? in_data_i[303] : 
                          (N373)? in_data_i[335] : 
                          (N374)? in_data_i[367] : 
                          (N375)? in_data_i[399] : 
                          (N376)? in_data_i[431] : 
                          (N377)? in_data_i[463] : 
                          (N378)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[238] = (N370)? in_data_i[238] : 
                          (N371)? in_data_i[270] : 
                          (N372)? in_data_i[302] : 
                          (N373)? in_data_i[334] : 
                          (N374)? in_data_i[366] : 
                          (N375)? in_data_i[398] : 
                          (N376)? in_data_i[430] : 
                          (N377)? in_data_i[462] : 
                          (N378)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[237] = (N370)? in_data_i[237] : 
                          (N371)? in_data_i[269] : 
                          (N372)? in_data_i[301] : 
                          (N373)? in_data_i[333] : 
                          (N374)? in_data_i[365] : 
                          (N375)? in_data_i[397] : 
                          (N376)? in_data_i[429] : 
                          (N377)? in_data_i[461] : 
                          (N378)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[236] = (N370)? in_data_i[236] : 
                          (N371)? in_data_i[268] : 
                          (N372)? in_data_i[300] : 
                          (N373)? in_data_i[332] : 
                          (N374)? in_data_i[364] : 
                          (N375)? in_data_i[396] : 
                          (N376)? in_data_i[428] : 
                          (N377)? in_data_i[460] : 
                          (N378)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[235] = (N370)? in_data_i[235] : 
                          (N371)? in_data_i[267] : 
                          (N372)? in_data_i[299] : 
                          (N373)? in_data_i[331] : 
                          (N374)? in_data_i[363] : 
                          (N375)? in_data_i[395] : 
                          (N376)? in_data_i[427] : 
                          (N377)? in_data_i[459] : 
                          (N378)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[234] = (N370)? in_data_i[234] : 
                          (N371)? in_data_i[266] : 
                          (N372)? in_data_i[298] : 
                          (N373)? in_data_i[330] : 
                          (N374)? in_data_i[362] : 
                          (N375)? in_data_i[394] : 
                          (N376)? in_data_i[426] : 
                          (N377)? in_data_i[458] : 
                          (N378)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[233] = (N370)? in_data_i[233] : 
                          (N371)? in_data_i[265] : 
                          (N372)? in_data_i[297] : 
                          (N373)? in_data_i[329] : 
                          (N374)? in_data_i[361] : 
                          (N375)? in_data_i[393] : 
                          (N376)? in_data_i[425] : 
                          (N377)? in_data_i[457] : 
                          (N378)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[232] = (N370)? in_data_i[232] : 
                          (N371)? in_data_i[264] : 
                          (N372)? in_data_i[296] : 
                          (N373)? in_data_i[328] : 
                          (N374)? in_data_i[360] : 
                          (N375)? in_data_i[392] : 
                          (N376)? in_data_i[424] : 
                          (N377)? in_data_i[456] : 
                          (N378)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[231] = (N370)? in_data_i[231] : 
                          (N371)? in_data_i[263] : 
                          (N372)? in_data_i[295] : 
                          (N373)? in_data_i[327] : 
                          (N374)? in_data_i[359] : 
                          (N375)? in_data_i[391] : 
                          (N376)? in_data_i[423] : 
                          (N377)? in_data_i[455] : 
                          (N378)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[230] = (N370)? in_data_i[230] : 
                          (N371)? in_data_i[262] : 
                          (N372)? in_data_i[294] : 
                          (N373)? in_data_i[326] : 
                          (N374)? in_data_i[358] : 
                          (N375)? in_data_i[390] : 
                          (N376)? in_data_i[422] : 
                          (N377)? in_data_i[454] : 
                          (N378)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[229] = (N370)? in_data_i[229] : 
                          (N371)? in_data_i[261] : 
                          (N372)? in_data_i[293] : 
                          (N373)? in_data_i[325] : 
                          (N374)? in_data_i[357] : 
                          (N375)? in_data_i[389] : 
                          (N376)? in_data_i[421] : 
                          (N377)? in_data_i[453] : 
                          (N378)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[228] = (N370)? in_data_i[228] : 
                          (N371)? in_data_i[260] : 
                          (N372)? in_data_i[292] : 
                          (N373)? in_data_i[324] : 
                          (N374)? in_data_i[356] : 
                          (N375)? in_data_i[388] : 
                          (N376)? in_data_i[420] : 
                          (N377)? in_data_i[452] : 
                          (N378)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[227] = (N370)? in_data_i[227] : 
                          (N371)? in_data_i[259] : 
                          (N372)? in_data_i[291] : 
                          (N373)? in_data_i[323] : 
                          (N374)? in_data_i[355] : 
                          (N375)? in_data_i[387] : 
                          (N376)? in_data_i[419] : 
                          (N377)? in_data_i[451] : 
                          (N378)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[226] = (N370)? in_data_i[226] : 
                          (N371)? in_data_i[258] : 
                          (N372)? in_data_i[290] : 
                          (N373)? in_data_i[322] : 
                          (N374)? in_data_i[354] : 
                          (N375)? in_data_i[386] : 
                          (N376)? in_data_i[418] : 
                          (N377)? in_data_i[450] : 
                          (N378)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[225] = (N370)? in_data_i[225] : 
                          (N371)? in_data_i[257] : 
                          (N372)? in_data_i[289] : 
                          (N373)? in_data_i[321] : 
                          (N374)? in_data_i[353] : 
                          (N375)? in_data_i[385] : 
                          (N376)? in_data_i[417] : 
                          (N377)? in_data_i[449] : 
                          (N378)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[224] = (N370)? in_data_i[224] : 
                          (N371)? in_data_i[256] : 
                          (N372)? in_data_i[288] : 
                          (N373)? in_data_i[320] : 
                          (N374)? in_data_i[352] : 
                          (N375)? in_data_i[384] : 
                          (N376)? in_data_i[416] : 
                          (N377)? in_data_i[448] : 
                          (N378)? in_data_i_15__0_ : 1'b0;
  assign in_data_o[223] = (N379)? in_data_i[223] : 
                          (N380)? in_data_i[255] : 
                          (N381)? in_data_i[287] : 
                          (N382)? in_data_i[319] : 
                          (N383)? in_data_i[351] : 
                          (N384)? in_data_i[383] : 
                          (N385)? in_data_i[415] : 
                          (N386)? in_data_i[447] : 
                          (N387)? in_data_i[479] : 
                          (N388)? in_data_i_15__31_ : 1'b0;
  assign N379 = N1349;
  assign N380 = N1351;
  assign N381 = N1353;
  assign N382 = N1354;
  assign N383 = N1355;
  assign N384 = N1356;
  assign N385 = N1357;
  assign N386 = N1358;
  assign N387 = N1350;
  assign N388 = N1352;
  assign in_data_o[222] = (N379)? in_data_i[222] : 
                          (N380)? in_data_i[254] : 
                          (N381)? in_data_i[286] : 
                          (N382)? in_data_i[318] : 
                          (N383)? in_data_i[350] : 
                          (N384)? in_data_i[382] : 
                          (N385)? in_data_i[414] : 
                          (N386)? in_data_i[446] : 
                          (N387)? in_data_i[478] : 
                          (N388)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[221] = (N379)? in_data_i[221] : 
                          (N380)? in_data_i[253] : 
                          (N381)? in_data_i[285] : 
                          (N382)? in_data_i[317] : 
                          (N383)? in_data_i[349] : 
                          (N384)? in_data_i[381] : 
                          (N385)? in_data_i[413] : 
                          (N386)? in_data_i[445] : 
                          (N387)? in_data_i[477] : 
                          (N388)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[220] = (N379)? in_data_i[220] : 
                          (N380)? in_data_i[252] : 
                          (N381)? in_data_i[284] : 
                          (N382)? in_data_i[316] : 
                          (N383)? in_data_i[348] : 
                          (N384)? in_data_i[380] : 
                          (N385)? in_data_i[412] : 
                          (N386)? in_data_i[444] : 
                          (N387)? in_data_i[476] : 
                          (N388)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[219] = (N379)? in_data_i[219] : 
                          (N380)? in_data_i[251] : 
                          (N381)? in_data_i[283] : 
                          (N382)? in_data_i[315] : 
                          (N383)? in_data_i[347] : 
                          (N384)? in_data_i[379] : 
                          (N385)? in_data_i[411] : 
                          (N386)? in_data_i[443] : 
                          (N387)? in_data_i[475] : 
                          (N388)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[218] = (N379)? in_data_i[218] : 
                          (N380)? in_data_i[250] : 
                          (N381)? in_data_i[282] : 
                          (N382)? in_data_i[314] : 
                          (N383)? in_data_i[346] : 
                          (N384)? in_data_i[378] : 
                          (N385)? in_data_i[410] : 
                          (N386)? in_data_i[442] : 
                          (N387)? in_data_i[474] : 
                          (N388)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[217] = (N379)? in_data_i[217] : 
                          (N380)? in_data_i[249] : 
                          (N381)? in_data_i[281] : 
                          (N382)? in_data_i[313] : 
                          (N383)? in_data_i[345] : 
                          (N384)? in_data_i[377] : 
                          (N385)? in_data_i[409] : 
                          (N386)? in_data_i[441] : 
                          (N387)? in_data_i[473] : 
                          (N388)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[216] = (N379)? in_data_i[216] : 
                          (N380)? in_data_i[248] : 
                          (N381)? in_data_i[280] : 
                          (N382)? in_data_i[312] : 
                          (N383)? in_data_i[344] : 
                          (N384)? in_data_i[376] : 
                          (N385)? in_data_i[408] : 
                          (N386)? in_data_i[440] : 
                          (N387)? in_data_i[472] : 
                          (N388)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[215] = (N379)? in_data_i[215] : 
                          (N380)? in_data_i[247] : 
                          (N381)? in_data_i[279] : 
                          (N382)? in_data_i[311] : 
                          (N383)? in_data_i[343] : 
                          (N384)? in_data_i[375] : 
                          (N385)? in_data_i[407] : 
                          (N386)? in_data_i[439] : 
                          (N387)? in_data_i[471] : 
                          (N388)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[214] = (N379)? in_data_i[214] : 
                          (N380)? in_data_i[246] : 
                          (N381)? in_data_i[278] : 
                          (N382)? in_data_i[310] : 
                          (N383)? in_data_i[342] : 
                          (N384)? in_data_i[374] : 
                          (N385)? in_data_i[406] : 
                          (N386)? in_data_i[438] : 
                          (N387)? in_data_i[470] : 
                          (N388)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[213] = (N379)? in_data_i[213] : 
                          (N380)? in_data_i[245] : 
                          (N381)? in_data_i[277] : 
                          (N382)? in_data_i[309] : 
                          (N383)? in_data_i[341] : 
                          (N384)? in_data_i[373] : 
                          (N385)? in_data_i[405] : 
                          (N386)? in_data_i[437] : 
                          (N387)? in_data_i[469] : 
                          (N388)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[212] = (N379)? in_data_i[212] : 
                          (N380)? in_data_i[244] : 
                          (N381)? in_data_i[276] : 
                          (N382)? in_data_i[308] : 
                          (N383)? in_data_i[340] : 
                          (N384)? in_data_i[372] : 
                          (N385)? in_data_i[404] : 
                          (N386)? in_data_i[436] : 
                          (N387)? in_data_i[468] : 
                          (N388)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[211] = (N379)? in_data_i[211] : 
                          (N380)? in_data_i[243] : 
                          (N381)? in_data_i[275] : 
                          (N382)? in_data_i[307] : 
                          (N383)? in_data_i[339] : 
                          (N384)? in_data_i[371] : 
                          (N385)? in_data_i[403] : 
                          (N386)? in_data_i[435] : 
                          (N387)? in_data_i[467] : 
                          (N388)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[210] = (N379)? in_data_i[210] : 
                          (N380)? in_data_i[242] : 
                          (N381)? in_data_i[274] : 
                          (N382)? in_data_i[306] : 
                          (N383)? in_data_i[338] : 
                          (N384)? in_data_i[370] : 
                          (N385)? in_data_i[402] : 
                          (N386)? in_data_i[434] : 
                          (N387)? in_data_i[466] : 
                          (N388)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[209] = (N379)? in_data_i[209] : 
                          (N380)? in_data_i[241] : 
                          (N381)? in_data_i[273] : 
                          (N382)? in_data_i[305] : 
                          (N383)? in_data_i[337] : 
                          (N384)? in_data_i[369] : 
                          (N385)? in_data_i[401] : 
                          (N386)? in_data_i[433] : 
                          (N387)? in_data_i[465] : 
                          (N388)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[208] = (N379)? in_data_i[208] : 
                          (N380)? in_data_i[240] : 
                          (N381)? in_data_i[272] : 
                          (N382)? in_data_i[304] : 
                          (N383)? in_data_i[336] : 
                          (N384)? in_data_i[368] : 
                          (N385)? in_data_i[400] : 
                          (N386)? in_data_i[432] : 
                          (N387)? in_data_i[464] : 
                          (N388)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[207] = (N379)? in_data_i[207] : 
                          (N380)? in_data_i[239] : 
                          (N381)? in_data_i[271] : 
                          (N382)? in_data_i[303] : 
                          (N383)? in_data_i[335] : 
                          (N384)? in_data_i[367] : 
                          (N385)? in_data_i[399] : 
                          (N386)? in_data_i[431] : 
                          (N387)? in_data_i[463] : 
                          (N388)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[206] = (N379)? in_data_i[206] : 
                          (N380)? in_data_i[238] : 
                          (N381)? in_data_i[270] : 
                          (N382)? in_data_i[302] : 
                          (N383)? in_data_i[334] : 
                          (N384)? in_data_i[366] : 
                          (N385)? in_data_i[398] : 
                          (N386)? in_data_i[430] : 
                          (N387)? in_data_i[462] : 
                          (N388)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[205] = (N379)? in_data_i[205] : 
                          (N380)? in_data_i[237] : 
                          (N381)? in_data_i[269] : 
                          (N382)? in_data_i[301] : 
                          (N383)? in_data_i[333] : 
                          (N384)? in_data_i[365] : 
                          (N385)? in_data_i[397] : 
                          (N386)? in_data_i[429] : 
                          (N387)? in_data_i[461] : 
                          (N388)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[204] = (N379)? in_data_i[204] : 
                          (N380)? in_data_i[236] : 
                          (N381)? in_data_i[268] : 
                          (N382)? in_data_i[300] : 
                          (N383)? in_data_i[332] : 
                          (N384)? in_data_i[364] : 
                          (N385)? in_data_i[396] : 
                          (N386)? in_data_i[428] : 
                          (N387)? in_data_i[460] : 
                          (N388)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[203] = (N379)? in_data_i[203] : 
                          (N380)? in_data_i[235] : 
                          (N381)? in_data_i[267] : 
                          (N382)? in_data_i[299] : 
                          (N383)? in_data_i[331] : 
                          (N384)? in_data_i[363] : 
                          (N385)? in_data_i[395] : 
                          (N386)? in_data_i[427] : 
                          (N387)? in_data_i[459] : 
                          (N388)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[202] = (N379)? in_data_i[202] : 
                          (N380)? in_data_i[234] : 
                          (N381)? in_data_i[266] : 
                          (N382)? in_data_i[298] : 
                          (N383)? in_data_i[330] : 
                          (N384)? in_data_i[362] : 
                          (N385)? in_data_i[394] : 
                          (N386)? in_data_i[426] : 
                          (N387)? in_data_i[458] : 
                          (N388)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[201] = (N379)? in_data_i[201] : 
                          (N380)? in_data_i[233] : 
                          (N381)? in_data_i[265] : 
                          (N382)? in_data_i[297] : 
                          (N383)? in_data_i[329] : 
                          (N384)? in_data_i[361] : 
                          (N385)? in_data_i[393] : 
                          (N386)? in_data_i[425] : 
                          (N387)? in_data_i[457] : 
                          (N388)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[200] = (N379)? in_data_i[200] : 
                          (N380)? in_data_i[232] : 
                          (N381)? in_data_i[264] : 
                          (N382)? in_data_i[296] : 
                          (N383)? in_data_i[328] : 
                          (N384)? in_data_i[360] : 
                          (N385)? in_data_i[392] : 
                          (N386)? in_data_i[424] : 
                          (N387)? in_data_i[456] : 
                          (N388)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[199] = (N379)? in_data_i[199] : 
                          (N380)? in_data_i[231] : 
                          (N381)? in_data_i[263] : 
                          (N382)? in_data_i[295] : 
                          (N383)? in_data_i[327] : 
                          (N384)? in_data_i[359] : 
                          (N385)? in_data_i[391] : 
                          (N386)? in_data_i[423] : 
                          (N387)? in_data_i[455] : 
                          (N388)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[198] = (N379)? in_data_i[198] : 
                          (N380)? in_data_i[230] : 
                          (N381)? in_data_i[262] : 
                          (N382)? in_data_i[294] : 
                          (N383)? in_data_i[326] : 
                          (N384)? in_data_i[358] : 
                          (N385)? in_data_i[390] : 
                          (N386)? in_data_i[422] : 
                          (N387)? in_data_i[454] : 
                          (N388)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[197] = (N379)? in_data_i[197] : 
                          (N380)? in_data_i[229] : 
                          (N381)? in_data_i[261] : 
                          (N382)? in_data_i[293] : 
                          (N383)? in_data_i[325] : 
                          (N384)? in_data_i[357] : 
                          (N385)? in_data_i[389] : 
                          (N386)? in_data_i[421] : 
                          (N387)? in_data_i[453] : 
                          (N388)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[196] = (N379)? in_data_i[196] : 
                          (N380)? in_data_i[228] : 
                          (N381)? in_data_i[260] : 
                          (N382)? in_data_i[292] : 
                          (N383)? in_data_i[324] : 
                          (N384)? in_data_i[356] : 
                          (N385)? in_data_i[388] : 
                          (N386)? in_data_i[420] : 
                          (N387)? in_data_i[452] : 
                          (N388)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[195] = (N379)? in_data_i[195] : 
                          (N380)? in_data_i[227] : 
                          (N381)? in_data_i[259] : 
                          (N382)? in_data_i[291] : 
                          (N383)? in_data_i[323] : 
                          (N384)? in_data_i[355] : 
                          (N385)? in_data_i[387] : 
                          (N386)? in_data_i[419] : 
                          (N387)? in_data_i[451] : 
                          (N388)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[194] = (N379)? in_data_i[194] : 
                          (N380)? in_data_i[226] : 
                          (N381)? in_data_i[258] : 
                          (N382)? in_data_i[290] : 
                          (N383)? in_data_i[322] : 
                          (N384)? in_data_i[354] : 
                          (N385)? in_data_i[386] : 
                          (N386)? in_data_i[418] : 
                          (N387)? in_data_i[450] : 
                          (N388)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[193] = (N379)? in_data_i[193] : 
                          (N380)? in_data_i[225] : 
                          (N381)? in_data_i[257] : 
                          (N382)? in_data_i[289] : 
                          (N383)? in_data_i[321] : 
                          (N384)? in_data_i[353] : 
                          (N385)? in_data_i[385] : 
                          (N386)? in_data_i[417] : 
                          (N387)? in_data_i[449] : 
                          (N388)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[192] = (N379)? in_data_i[192] : 
                          (N380)? in_data_i[224] : 
                          (N381)? in_data_i[256] : 
                          (N382)? in_data_i[288] : 
                          (N383)? in_data_i[320] : 
                          (N384)? in_data_i[352] : 
                          (N385)? in_data_i[384] : 
                          (N386)? in_data_i[416] : 
                          (N387)? in_data_i[448] : 
                          (N388)? in_data_i_15__0_ : 1'b0;
  assign in_data_o[191] = (N389)? in_data_i[191] : 
                          (N390)? in_data_i[223] : 
                          (N391)? in_data_i[255] : 
                          (N392)? in_data_i[287] : 
                          (N393)? in_data_i[319] : 
                          (N394)? in_data_i[351] : 
                          (N395)? in_data_i[383] : 
                          (N396)? in_data_i[415] : 
                          (N397)? in_data_i[447] : 
                          (N398)? in_data_i[479] : 
                          (N399)? in_data_i_15__31_ : 1'b0;
  assign N389 = N1224;
  assign N390 = N1226;
  assign N391 = N1228;
  assign N392 = N1230;
  assign N393 = N1231;
  assign N394 = N1232;
  assign N395 = N1233;
  assign N396 = N1234;
  assign N397 = N1225;
  assign N398 = N1227;
  assign N399 = N1229;
  assign in_data_o[190] = (N389)? in_data_i[190] : 
                          (N390)? in_data_i[222] : 
                          (N391)? in_data_i[254] : 
                          (N392)? in_data_i[286] : 
                          (N393)? in_data_i[318] : 
                          (N394)? in_data_i[350] : 
                          (N395)? in_data_i[382] : 
                          (N396)? in_data_i[414] : 
                          (N397)? in_data_i[446] : 
                          (N398)? in_data_i[478] : 
                          (N399)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[189] = (N389)? in_data_i[189] : 
                          (N390)? in_data_i[221] : 
                          (N391)? in_data_i[253] : 
                          (N392)? in_data_i[285] : 
                          (N393)? in_data_i[317] : 
                          (N394)? in_data_i[349] : 
                          (N395)? in_data_i[381] : 
                          (N396)? in_data_i[413] : 
                          (N397)? in_data_i[445] : 
                          (N398)? in_data_i[477] : 
                          (N399)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[188] = (N389)? in_data_i[188] : 
                          (N390)? in_data_i[220] : 
                          (N391)? in_data_i[252] : 
                          (N392)? in_data_i[284] : 
                          (N393)? in_data_i[316] : 
                          (N394)? in_data_i[348] : 
                          (N395)? in_data_i[380] : 
                          (N396)? in_data_i[412] : 
                          (N397)? in_data_i[444] : 
                          (N398)? in_data_i[476] : 
                          (N399)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[187] = (N389)? in_data_i[187] : 
                          (N390)? in_data_i[219] : 
                          (N391)? in_data_i[251] : 
                          (N392)? in_data_i[283] : 
                          (N393)? in_data_i[315] : 
                          (N394)? in_data_i[347] : 
                          (N395)? in_data_i[379] : 
                          (N396)? in_data_i[411] : 
                          (N397)? in_data_i[443] : 
                          (N398)? in_data_i[475] : 
                          (N399)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[186] = (N389)? in_data_i[186] : 
                          (N390)? in_data_i[218] : 
                          (N391)? in_data_i[250] : 
                          (N392)? in_data_i[282] : 
                          (N393)? in_data_i[314] : 
                          (N394)? in_data_i[346] : 
                          (N395)? in_data_i[378] : 
                          (N396)? in_data_i[410] : 
                          (N397)? in_data_i[442] : 
                          (N398)? in_data_i[474] : 
                          (N399)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[185] = (N389)? in_data_i[185] : 
                          (N390)? in_data_i[217] : 
                          (N391)? in_data_i[249] : 
                          (N392)? in_data_i[281] : 
                          (N393)? in_data_i[313] : 
                          (N394)? in_data_i[345] : 
                          (N395)? in_data_i[377] : 
                          (N396)? in_data_i[409] : 
                          (N397)? in_data_i[441] : 
                          (N398)? in_data_i[473] : 
                          (N399)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[184] = (N389)? in_data_i[184] : 
                          (N390)? in_data_i[216] : 
                          (N391)? in_data_i[248] : 
                          (N392)? in_data_i[280] : 
                          (N393)? in_data_i[312] : 
                          (N394)? in_data_i[344] : 
                          (N395)? in_data_i[376] : 
                          (N396)? in_data_i[408] : 
                          (N397)? in_data_i[440] : 
                          (N398)? in_data_i[472] : 
                          (N399)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[183] = (N389)? in_data_i[183] : 
                          (N390)? in_data_i[215] : 
                          (N391)? in_data_i[247] : 
                          (N392)? in_data_i[279] : 
                          (N393)? in_data_i[311] : 
                          (N394)? in_data_i[343] : 
                          (N395)? in_data_i[375] : 
                          (N396)? in_data_i[407] : 
                          (N397)? in_data_i[439] : 
                          (N398)? in_data_i[471] : 
                          (N399)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[182] = (N389)? in_data_i[182] : 
                          (N390)? in_data_i[214] : 
                          (N391)? in_data_i[246] : 
                          (N392)? in_data_i[278] : 
                          (N393)? in_data_i[310] : 
                          (N394)? in_data_i[342] : 
                          (N395)? in_data_i[374] : 
                          (N396)? in_data_i[406] : 
                          (N397)? in_data_i[438] : 
                          (N398)? in_data_i[470] : 
                          (N399)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[181] = (N389)? in_data_i[181] : 
                          (N390)? in_data_i[213] : 
                          (N391)? in_data_i[245] : 
                          (N392)? in_data_i[277] : 
                          (N393)? in_data_i[309] : 
                          (N394)? in_data_i[341] : 
                          (N395)? in_data_i[373] : 
                          (N396)? in_data_i[405] : 
                          (N397)? in_data_i[437] : 
                          (N398)? in_data_i[469] : 
                          (N399)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[180] = (N389)? in_data_i[180] : 
                          (N390)? in_data_i[212] : 
                          (N391)? in_data_i[244] : 
                          (N392)? in_data_i[276] : 
                          (N393)? in_data_i[308] : 
                          (N394)? in_data_i[340] : 
                          (N395)? in_data_i[372] : 
                          (N396)? in_data_i[404] : 
                          (N397)? in_data_i[436] : 
                          (N398)? in_data_i[468] : 
                          (N399)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[179] = (N389)? in_data_i[179] : 
                          (N390)? in_data_i[211] : 
                          (N391)? in_data_i[243] : 
                          (N392)? in_data_i[275] : 
                          (N393)? in_data_i[307] : 
                          (N394)? in_data_i[339] : 
                          (N395)? in_data_i[371] : 
                          (N396)? in_data_i[403] : 
                          (N397)? in_data_i[435] : 
                          (N398)? in_data_i[467] : 
                          (N399)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[178] = (N389)? in_data_i[178] : 
                          (N390)? in_data_i[210] : 
                          (N391)? in_data_i[242] : 
                          (N392)? in_data_i[274] : 
                          (N393)? in_data_i[306] : 
                          (N394)? in_data_i[338] : 
                          (N395)? in_data_i[370] : 
                          (N396)? in_data_i[402] : 
                          (N397)? in_data_i[434] : 
                          (N398)? in_data_i[466] : 
                          (N399)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[177] = (N389)? in_data_i[177] : 
                          (N390)? in_data_i[209] : 
                          (N391)? in_data_i[241] : 
                          (N392)? in_data_i[273] : 
                          (N393)? in_data_i[305] : 
                          (N394)? in_data_i[337] : 
                          (N395)? in_data_i[369] : 
                          (N396)? in_data_i[401] : 
                          (N397)? in_data_i[433] : 
                          (N398)? in_data_i[465] : 
                          (N399)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[176] = (N389)? in_data_i[176] : 
                          (N390)? in_data_i[208] : 
                          (N391)? in_data_i[240] : 
                          (N392)? in_data_i[272] : 
                          (N393)? in_data_i[304] : 
                          (N394)? in_data_i[336] : 
                          (N395)? in_data_i[368] : 
                          (N396)? in_data_i[400] : 
                          (N397)? in_data_i[432] : 
                          (N398)? in_data_i[464] : 
                          (N399)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[175] = (N389)? in_data_i[175] : 
                          (N390)? in_data_i[207] : 
                          (N391)? in_data_i[239] : 
                          (N392)? in_data_i[271] : 
                          (N393)? in_data_i[303] : 
                          (N394)? in_data_i[335] : 
                          (N395)? in_data_i[367] : 
                          (N396)? in_data_i[399] : 
                          (N397)? in_data_i[431] : 
                          (N398)? in_data_i[463] : 
                          (N399)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[174] = (N389)? in_data_i[174] : 
                          (N390)? in_data_i[206] : 
                          (N391)? in_data_i[238] : 
                          (N392)? in_data_i[270] : 
                          (N393)? in_data_i[302] : 
                          (N394)? in_data_i[334] : 
                          (N395)? in_data_i[366] : 
                          (N396)? in_data_i[398] : 
                          (N397)? in_data_i[430] : 
                          (N398)? in_data_i[462] : 
                          (N399)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[173] = (N389)? in_data_i[173] : 
                          (N390)? in_data_i[205] : 
                          (N391)? in_data_i[237] : 
                          (N392)? in_data_i[269] : 
                          (N393)? in_data_i[301] : 
                          (N394)? in_data_i[333] : 
                          (N395)? in_data_i[365] : 
                          (N396)? in_data_i[397] : 
                          (N397)? in_data_i[429] : 
                          (N398)? in_data_i[461] : 
                          (N399)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[172] = (N389)? in_data_i[172] : 
                          (N390)? in_data_i[204] : 
                          (N391)? in_data_i[236] : 
                          (N392)? in_data_i[268] : 
                          (N393)? in_data_i[300] : 
                          (N394)? in_data_i[332] : 
                          (N395)? in_data_i[364] : 
                          (N396)? in_data_i[396] : 
                          (N397)? in_data_i[428] : 
                          (N398)? in_data_i[460] : 
                          (N399)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[171] = (N389)? in_data_i[171] : 
                          (N390)? in_data_i[203] : 
                          (N391)? in_data_i[235] : 
                          (N392)? in_data_i[267] : 
                          (N393)? in_data_i[299] : 
                          (N394)? in_data_i[331] : 
                          (N395)? in_data_i[363] : 
                          (N396)? in_data_i[395] : 
                          (N397)? in_data_i[427] : 
                          (N398)? in_data_i[459] : 
                          (N399)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[170] = (N389)? in_data_i[170] : 
                          (N390)? in_data_i[202] : 
                          (N391)? in_data_i[234] : 
                          (N392)? in_data_i[266] : 
                          (N393)? in_data_i[298] : 
                          (N394)? in_data_i[330] : 
                          (N395)? in_data_i[362] : 
                          (N396)? in_data_i[394] : 
                          (N397)? in_data_i[426] : 
                          (N398)? in_data_i[458] : 
                          (N399)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[169] = (N389)? in_data_i[169] : 
                          (N390)? in_data_i[201] : 
                          (N391)? in_data_i[233] : 
                          (N392)? in_data_i[265] : 
                          (N393)? in_data_i[297] : 
                          (N394)? in_data_i[329] : 
                          (N395)? in_data_i[361] : 
                          (N396)? in_data_i[393] : 
                          (N397)? in_data_i[425] : 
                          (N398)? in_data_i[457] : 
                          (N399)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[168] = (N389)? in_data_i[168] : 
                          (N390)? in_data_i[200] : 
                          (N391)? in_data_i[232] : 
                          (N392)? in_data_i[264] : 
                          (N393)? in_data_i[296] : 
                          (N394)? in_data_i[328] : 
                          (N395)? in_data_i[360] : 
                          (N396)? in_data_i[392] : 
                          (N397)? in_data_i[424] : 
                          (N398)? in_data_i[456] : 
                          (N399)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[167] = (N389)? in_data_i[167] : 
                          (N390)? in_data_i[199] : 
                          (N391)? in_data_i[231] : 
                          (N392)? in_data_i[263] : 
                          (N393)? in_data_i[295] : 
                          (N394)? in_data_i[327] : 
                          (N395)? in_data_i[359] : 
                          (N396)? in_data_i[391] : 
                          (N397)? in_data_i[423] : 
                          (N398)? in_data_i[455] : 
                          (N399)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[166] = (N389)? in_data_i[166] : 
                          (N390)? in_data_i[198] : 
                          (N391)? in_data_i[230] : 
                          (N392)? in_data_i[262] : 
                          (N393)? in_data_i[294] : 
                          (N394)? in_data_i[326] : 
                          (N395)? in_data_i[358] : 
                          (N396)? in_data_i[390] : 
                          (N397)? in_data_i[422] : 
                          (N398)? in_data_i[454] : 
                          (N399)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[165] = (N389)? in_data_i[165] : 
                          (N390)? in_data_i[197] : 
                          (N391)? in_data_i[229] : 
                          (N392)? in_data_i[261] : 
                          (N393)? in_data_i[293] : 
                          (N394)? in_data_i[325] : 
                          (N395)? in_data_i[357] : 
                          (N396)? in_data_i[389] : 
                          (N397)? in_data_i[421] : 
                          (N398)? in_data_i[453] : 
                          (N399)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[164] = (N389)? in_data_i[164] : 
                          (N390)? in_data_i[196] : 
                          (N391)? in_data_i[228] : 
                          (N392)? in_data_i[260] : 
                          (N393)? in_data_i[292] : 
                          (N394)? in_data_i[324] : 
                          (N395)? in_data_i[356] : 
                          (N396)? in_data_i[388] : 
                          (N397)? in_data_i[420] : 
                          (N398)? in_data_i[452] : 
                          (N399)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[163] = (N389)? in_data_i[163] : 
                          (N390)? in_data_i[195] : 
                          (N391)? in_data_i[227] : 
                          (N392)? in_data_i[259] : 
                          (N393)? in_data_i[291] : 
                          (N394)? in_data_i[323] : 
                          (N395)? in_data_i[355] : 
                          (N396)? in_data_i[387] : 
                          (N397)? in_data_i[419] : 
                          (N398)? in_data_i[451] : 
                          (N399)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[162] = (N389)? in_data_i[162] : 
                          (N390)? in_data_i[194] : 
                          (N391)? in_data_i[226] : 
                          (N392)? in_data_i[258] : 
                          (N393)? in_data_i[290] : 
                          (N394)? in_data_i[322] : 
                          (N395)? in_data_i[354] : 
                          (N396)? in_data_i[386] : 
                          (N397)? in_data_i[418] : 
                          (N398)? in_data_i[450] : 
                          (N399)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[161] = (N389)? in_data_i[161] : 
                          (N390)? in_data_i[193] : 
                          (N391)? in_data_i[225] : 
                          (N392)? in_data_i[257] : 
                          (N393)? in_data_i[289] : 
                          (N394)? in_data_i[321] : 
                          (N395)? in_data_i[353] : 
                          (N396)? in_data_i[385] : 
                          (N397)? in_data_i[417] : 
                          (N398)? in_data_i[449] : 
                          (N399)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[160] = (N389)? in_data_i[160] : 
                          (N390)? in_data_i[192] : 
                          (N391)? in_data_i[224] : 
                          (N392)? in_data_i[256] : 
                          (N393)? in_data_i[288] : 
                          (N394)? in_data_i[320] : 
                          (N395)? in_data_i[352] : 
                          (N396)? in_data_i[384] : 
                          (N397)? in_data_i[416] : 
                          (N398)? in_data_i[448] : 
                          (N399)? in_data_i_15__0_ : 1'b0;
  assign in_data_o[159] = (N400)? in_data_i[159] : 
                          (N401)? in_data_i[191] : 
                          (N402)? in_data_i[223] : 
                          (N403)? in_data_i[255] : 
                          (N404)? in_data_i[287] : 
                          (N405)? in_data_i[319] : 
                          (N406)? in_data_i[351] : 
                          (N407)? in_data_i[383] : 
                          (N408)? in_data_i[415] : 
                          (N409)? in_data_i[447] : 
                          (N410)? in_data_i[479] : 
                          (N411)? in_data_i_15__31_ : 1'b0;
  assign N400 = N1100;
  assign N401 = N1102;
  assign N402 = N1104;
  assign N403 = N1106;
  assign N404 = N1108;
  assign N405 = N1109;
  assign N406 = N1110;
  assign N407 = N1111;
  assign N408 = N1101;
  assign N409 = N1103;
  assign N410 = N1105;
  assign N411 = N1107;
  assign in_data_o[158] = (N400)? in_data_i[158] : 
                          (N401)? in_data_i[190] : 
                          (N402)? in_data_i[222] : 
                          (N403)? in_data_i[254] : 
                          (N404)? in_data_i[286] : 
                          (N405)? in_data_i[318] : 
                          (N406)? in_data_i[350] : 
                          (N407)? in_data_i[382] : 
                          (N408)? in_data_i[414] : 
                          (N409)? in_data_i[446] : 
                          (N410)? in_data_i[478] : 
                          (N411)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[157] = (N400)? in_data_i[157] : 
                          (N401)? in_data_i[189] : 
                          (N402)? in_data_i[221] : 
                          (N403)? in_data_i[253] : 
                          (N404)? in_data_i[285] : 
                          (N405)? in_data_i[317] : 
                          (N406)? in_data_i[349] : 
                          (N407)? in_data_i[381] : 
                          (N408)? in_data_i[413] : 
                          (N409)? in_data_i[445] : 
                          (N410)? in_data_i[477] : 
                          (N411)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[156] = (N400)? in_data_i[156] : 
                          (N401)? in_data_i[188] : 
                          (N402)? in_data_i[220] : 
                          (N403)? in_data_i[252] : 
                          (N404)? in_data_i[284] : 
                          (N405)? in_data_i[316] : 
                          (N406)? in_data_i[348] : 
                          (N407)? in_data_i[380] : 
                          (N408)? in_data_i[412] : 
                          (N409)? in_data_i[444] : 
                          (N410)? in_data_i[476] : 
                          (N411)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[155] = (N400)? in_data_i[155] : 
                          (N401)? in_data_i[187] : 
                          (N402)? in_data_i[219] : 
                          (N403)? in_data_i[251] : 
                          (N404)? in_data_i[283] : 
                          (N405)? in_data_i[315] : 
                          (N406)? in_data_i[347] : 
                          (N407)? in_data_i[379] : 
                          (N408)? in_data_i[411] : 
                          (N409)? in_data_i[443] : 
                          (N410)? in_data_i[475] : 
                          (N411)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[154] = (N400)? in_data_i[154] : 
                          (N401)? in_data_i[186] : 
                          (N402)? in_data_i[218] : 
                          (N403)? in_data_i[250] : 
                          (N404)? in_data_i[282] : 
                          (N405)? in_data_i[314] : 
                          (N406)? in_data_i[346] : 
                          (N407)? in_data_i[378] : 
                          (N408)? in_data_i[410] : 
                          (N409)? in_data_i[442] : 
                          (N410)? in_data_i[474] : 
                          (N411)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[153] = (N400)? in_data_i[153] : 
                          (N401)? in_data_i[185] : 
                          (N402)? in_data_i[217] : 
                          (N403)? in_data_i[249] : 
                          (N404)? in_data_i[281] : 
                          (N405)? in_data_i[313] : 
                          (N406)? in_data_i[345] : 
                          (N407)? in_data_i[377] : 
                          (N408)? in_data_i[409] : 
                          (N409)? in_data_i[441] : 
                          (N410)? in_data_i[473] : 
                          (N411)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[152] = (N400)? in_data_i[152] : 
                          (N401)? in_data_i[184] : 
                          (N402)? in_data_i[216] : 
                          (N403)? in_data_i[248] : 
                          (N404)? in_data_i[280] : 
                          (N405)? in_data_i[312] : 
                          (N406)? in_data_i[344] : 
                          (N407)? in_data_i[376] : 
                          (N408)? in_data_i[408] : 
                          (N409)? in_data_i[440] : 
                          (N410)? in_data_i[472] : 
                          (N411)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[151] = (N400)? in_data_i[151] : 
                          (N401)? in_data_i[183] : 
                          (N402)? in_data_i[215] : 
                          (N403)? in_data_i[247] : 
                          (N404)? in_data_i[279] : 
                          (N405)? in_data_i[311] : 
                          (N406)? in_data_i[343] : 
                          (N407)? in_data_i[375] : 
                          (N408)? in_data_i[407] : 
                          (N409)? in_data_i[439] : 
                          (N410)? in_data_i[471] : 
                          (N411)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[150] = (N400)? in_data_i[150] : 
                          (N401)? in_data_i[182] : 
                          (N402)? in_data_i[214] : 
                          (N403)? in_data_i[246] : 
                          (N404)? in_data_i[278] : 
                          (N405)? in_data_i[310] : 
                          (N406)? in_data_i[342] : 
                          (N407)? in_data_i[374] : 
                          (N408)? in_data_i[406] : 
                          (N409)? in_data_i[438] : 
                          (N410)? in_data_i[470] : 
                          (N411)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[149] = (N400)? in_data_i[149] : 
                          (N401)? in_data_i[181] : 
                          (N402)? in_data_i[213] : 
                          (N403)? in_data_i[245] : 
                          (N404)? in_data_i[277] : 
                          (N405)? in_data_i[309] : 
                          (N406)? in_data_i[341] : 
                          (N407)? in_data_i[373] : 
                          (N408)? in_data_i[405] : 
                          (N409)? in_data_i[437] : 
                          (N410)? in_data_i[469] : 
                          (N411)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[148] = (N400)? in_data_i[148] : 
                          (N401)? in_data_i[180] : 
                          (N402)? in_data_i[212] : 
                          (N403)? in_data_i[244] : 
                          (N404)? in_data_i[276] : 
                          (N405)? in_data_i[308] : 
                          (N406)? in_data_i[340] : 
                          (N407)? in_data_i[372] : 
                          (N408)? in_data_i[404] : 
                          (N409)? in_data_i[436] : 
                          (N410)? in_data_i[468] : 
                          (N411)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[147] = (N400)? in_data_i[147] : 
                          (N401)? in_data_i[179] : 
                          (N402)? in_data_i[211] : 
                          (N403)? in_data_i[243] : 
                          (N404)? in_data_i[275] : 
                          (N405)? in_data_i[307] : 
                          (N406)? in_data_i[339] : 
                          (N407)? in_data_i[371] : 
                          (N408)? in_data_i[403] : 
                          (N409)? in_data_i[435] : 
                          (N410)? in_data_i[467] : 
                          (N411)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[146] = (N400)? in_data_i[146] : 
                          (N401)? in_data_i[178] : 
                          (N402)? in_data_i[210] : 
                          (N403)? in_data_i[242] : 
                          (N404)? in_data_i[274] : 
                          (N405)? in_data_i[306] : 
                          (N406)? in_data_i[338] : 
                          (N407)? in_data_i[370] : 
                          (N408)? in_data_i[402] : 
                          (N409)? in_data_i[434] : 
                          (N410)? in_data_i[466] : 
                          (N411)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[145] = (N400)? in_data_i[145] : 
                          (N401)? in_data_i[177] : 
                          (N402)? in_data_i[209] : 
                          (N403)? in_data_i[241] : 
                          (N404)? in_data_i[273] : 
                          (N405)? in_data_i[305] : 
                          (N406)? in_data_i[337] : 
                          (N407)? in_data_i[369] : 
                          (N408)? in_data_i[401] : 
                          (N409)? in_data_i[433] : 
                          (N410)? in_data_i[465] : 
                          (N411)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[144] = (N400)? in_data_i[144] : 
                          (N401)? in_data_i[176] : 
                          (N402)? in_data_i[208] : 
                          (N403)? in_data_i[240] : 
                          (N404)? in_data_i[272] : 
                          (N405)? in_data_i[304] : 
                          (N406)? in_data_i[336] : 
                          (N407)? in_data_i[368] : 
                          (N408)? in_data_i[400] : 
                          (N409)? in_data_i[432] : 
                          (N410)? in_data_i[464] : 
                          (N411)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[143] = (N400)? in_data_i[143] : 
                          (N401)? in_data_i[175] : 
                          (N402)? in_data_i[207] : 
                          (N403)? in_data_i[239] : 
                          (N404)? in_data_i[271] : 
                          (N405)? in_data_i[303] : 
                          (N406)? in_data_i[335] : 
                          (N407)? in_data_i[367] : 
                          (N408)? in_data_i[399] : 
                          (N409)? in_data_i[431] : 
                          (N410)? in_data_i[463] : 
                          (N411)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[142] = (N400)? in_data_i[142] : 
                          (N401)? in_data_i[174] : 
                          (N402)? in_data_i[206] : 
                          (N403)? in_data_i[238] : 
                          (N404)? in_data_i[270] : 
                          (N405)? in_data_i[302] : 
                          (N406)? in_data_i[334] : 
                          (N407)? in_data_i[366] : 
                          (N408)? in_data_i[398] : 
                          (N409)? in_data_i[430] : 
                          (N410)? in_data_i[462] : 
                          (N411)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[141] = (N400)? in_data_i[141] : 
                          (N401)? in_data_i[173] : 
                          (N402)? in_data_i[205] : 
                          (N403)? in_data_i[237] : 
                          (N404)? in_data_i[269] : 
                          (N405)? in_data_i[301] : 
                          (N406)? in_data_i[333] : 
                          (N407)? in_data_i[365] : 
                          (N408)? in_data_i[397] : 
                          (N409)? in_data_i[429] : 
                          (N410)? in_data_i[461] : 
                          (N411)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[140] = (N400)? in_data_i[140] : 
                          (N401)? in_data_i[172] : 
                          (N402)? in_data_i[204] : 
                          (N403)? in_data_i[236] : 
                          (N404)? in_data_i[268] : 
                          (N405)? in_data_i[300] : 
                          (N406)? in_data_i[332] : 
                          (N407)? in_data_i[364] : 
                          (N408)? in_data_i[396] : 
                          (N409)? in_data_i[428] : 
                          (N410)? in_data_i[460] : 
                          (N411)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[139] = (N400)? in_data_i[139] : 
                          (N401)? in_data_i[171] : 
                          (N402)? in_data_i[203] : 
                          (N403)? in_data_i[235] : 
                          (N404)? in_data_i[267] : 
                          (N405)? in_data_i[299] : 
                          (N406)? in_data_i[331] : 
                          (N407)? in_data_i[363] : 
                          (N408)? in_data_i[395] : 
                          (N409)? in_data_i[427] : 
                          (N410)? in_data_i[459] : 
                          (N411)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[138] = (N400)? in_data_i[138] : 
                          (N401)? in_data_i[170] : 
                          (N402)? in_data_i[202] : 
                          (N403)? in_data_i[234] : 
                          (N404)? in_data_i[266] : 
                          (N405)? in_data_i[298] : 
                          (N406)? in_data_i[330] : 
                          (N407)? in_data_i[362] : 
                          (N408)? in_data_i[394] : 
                          (N409)? in_data_i[426] : 
                          (N410)? in_data_i[458] : 
                          (N411)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[137] = (N400)? in_data_i[137] : 
                          (N401)? in_data_i[169] : 
                          (N402)? in_data_i[201] : 
                          (N403)? in_data_i[233] : 
                          (N404)? in_data_i[265] : 
                          (N405)? in_data_i[297] : 
                          (N406)? in_data_i[329] : 
                          (N407)? in_data_i[361] : 
                          (N408)? in_data_i[393] : 
                          (N409)? in_data_i[425] : 
                          (N410)? in_data_i[457] : 
                          (N411)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[136] = (N400)? in_data_i[136] : 
                          (N401)? in_data_i[168] : 
                          (N402)? in_data_i[200] : 
                          (N403)? in_data_i[232] : 
                          (N404)? in_data_i[264] : 
                          (N405)? in_data_i[296] : 
                          (N406)? in_data_i[328] : 
                          (N407)? in_data_i[360] : 
                          (N408)? in_data_i[392] : 
                          (N409)? in_data_i[424] : 
                          (N410)? in_data_i[456] : 
                          (N411)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[135] = (N400)? in_data_i[135] : 
                          (N401)? in_data_i[167] : 
                          (N402)? in_data_i[199] : 
                          (N403)? in_data_i[231] : 
                          (N404)? in_data_i[263] : 
                          (N405)? in_data_i[295] : 
                          (N406)? in_data_i[327] : 
                          (N407)? in_data_i[359] : 
                          (N408)? in_data_i[391] : 
                          (N409)? in_data_i[423] : 
                          (N410)? in_data_i[455] : 
                          (N411)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[134] = (N400)? in_data_i[134] : 
                          (N401)? in_data_i[166] : 
                          (N402)? in_data_i[198] : 
                          (N403)? in_data_i[230] : 
                          (N404)? in_data_i[262] : 
                          (N405)? in_data_i[294] : 
                          (N406)? in_data_i[326] : 
                          (N407)? in_data_i[358] : 
                          (N408)? in_data_i[390] : 
                          (N409)? in_data_i[422] : 
                          (N410)? in_data_i[454] : 
                          (N411)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[133] = (N400)? in_data_i[133] : 
                          (N401)? in_data_i[165] : 
                          (N402)? in_data_i[197] : 
                          (N403)? in_data_i[229] : 
                          (N404)? in_data_i[261] : 
                          (N405)? in_data_i[293] : 
                          (N406)? in_data_i[325] : 
                          (N407)? in_data_i[357] : 
                          (N408)? in_data_i[389] : 
                          (N409)? in_data_i[421] : 
                          (N410)? in_data_i[453] : 
                          (N411)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[132] = (N400)? in_data_i[132] : 
                          (N401)? in_data_i[164] : 
                          (N402)? in_data_i[196] : 
                          (N403)? in_data_i[228] : 
                          (N404)? in_data_i[260] : 
                          (N405)? in_data_i[292] : 
                          (N406)? in_data_i[324] : 
                          (N407)? in_data_i[356] : 
                          (N408)? in_data_i[388] : 
                          (N409)? in_data_i[420] : 
                          (N410)? in_data_i[452] : 
                          (N411)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[131] = (N400)? in_data_i[131] : 
                          (N401)? in_data_i[163] : 
                          (N402)? in_data_i[195] : 
                          (N403)? in_data_i[227] : 
                          (N404)? in_data_i[259] : 
                          (N405)? in_data_i[291] : 
                          (N406)? in_data_i[323] : 
                          (N407)? in_data_i[355] : 
                          (N408)? in_data_i[387] : 
                          (N409)? in_data_i[419] : 
                          (N410)? in_data_i[451] : 
                          (N411)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[130] = (N400)? in_data_i[130] : 
                          (N401)? in_data_i[162] : 
                          (N402)? in_data_i[194] : 
                          (N403)? in_data_i[226] : 
                          (N404)? in_data_i[258] : 
                          (N405)? in_data_i[290] : 
                          (N406)? in_data_i[322] : 
                          (N407)? in_data_i[354] : 
                          (N408)? in_data_i[386] : 
                          (N409)? in_data_i[418] : 
                          (N410)? in_data_i[450] : 
                          (N411)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[129] = (N400)? in_data_i[129] : 
                          (N401)? in_data_i[161] : 
                          (N402)? in_data_i[193] : 
                          (N403)? in_data_i[225] : 
                          (N404)? in_data_i[257] : 
                          (N405)? in_data_i[289] : 
                          (N406)? in_data_i[321] : 
                          (N407)? in_data_i[353] : 
                          (N408)? in_data_i[385] : 
                          (N409)? in_data_i[417] : 
                          (N410)? in_data_i[449] : 
                          (N411)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[128] = (N400)? in_data_i[128] : 
                          (N401)? in_data_i[160] : 
                          (N402)? in_data_i[192] : 
                          (N403)? in_data_i[224] : 
                          (N404)? in_data_i[256] : 
                          (N405)? in_data_i[288] : 
                          (N406)? in_data_i[320] : 
                          (N407)? in_data_i[352] : 
                          (N408)? in_data_i[384] : 
                          (N409)? in_data_i[416] : 
                          (N410)? in_data_i[448] : 
                          (N411)? in_data_i_15__0_ : 1'b0;
  assign in_data_o[127] = (N412)? in_data_i[127] : 
                          (N413)? in_data_i[159] : 
                          (N414)? in_data_i[191] : 
                          (N415)? in_data_i[223] : 
                          (N416)? in_data_i[255] : 
                          (N417)? in_data_i[287] : 
                          (N418)? in_data_i[319] : 
                          (N419)? in_data_i[351] : 
                          (N420)? in_data_i[383] : 
                          (N421)? in_data_i[415] : 
                          (N422)? in_data_i[447] : 
                          (N423)? in_data_i[479] : 
                          (N424)? in_data_i_15__31_ : 1'b0;
  assign N412 = N973;
  assign N413 = N975;
  assign N414 = N977;
  assign N415 = N979;
  assign N416 = N981;
  assign N417 = N983;
  assign N418 = N984;
  assign N419 = N985;
  assign N420 = N974;
  assign N421 = N976;
  assign N422 = N978;
  assign N423 = N980;
  assign N424 = N982;
  assign in_data_o[126] = (N412)? in_data_i[126] : 
                          (N413)? in_data_i[158] : 
                          (N414)? in_data_i[190] : 
                          (N415)? in_data_i[222] : 
                          (N416)? in_data_i[254] : 
                          (N417)? in_data_i[286] : 
                          (N418)? in_data_i[318] : 
                          (N419)? in_data_i[350] : 
                          (N420)? in_data_i[382] : 
                          (N421)? in_data_i[414] : 
                          (N422)? in_data_i[446] : 
                          (N423)? in_data_i[478] : 
                          (N424)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[125] = (N412)? in_data_i[125] : 
                          (N413)? in_data_i[157] : 
                          (N414)? in_data_i[189] : 
                          (N415)? in_data_i[221] : 
                          (N416)? in_data_i[253] : 
                          (N417)? in_data_i[285] : 
                          (N418)? in_data_i[317] : 
                          (N419)? in_data_i[349] : 
                          (N420)? in_data_i[381] : 
                          (N421)? in_data_i[413] : 
                          (N422)? in_data_i[445] : 
                          (N423)? in_data_i[477] : 
                          (N424)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[124] = (N412)? in_data_i[124] : 
                          (N413)? in_data_i[156] : 
                          (N414)? in_data_i[188] : 
                          (N415)? in_data_i[220] : 
                          (N416)? in_data_i[252] : 
                          (N417)? in_data_i[284] : 
                          (N418)? in_data_i[316] : 
                          (N419)? in_data_i[348] : 
                          (N420)? in_data_i[380] : 
                          (N421)? in_data_i[412] : 
                          (N422)? in_data_i[444] : 
                          (N423)? in_data_i[476] : 
                          (N424)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[123] = (N412)? in_data_i[123] : 
                          (N413)? in_data_i[155] : 
                          (N414)? in_data_i[187] : 
                          (N415)? in_data_i[219] : 
                          (N416)? in_data_i[251] : 
                          (N417)? in_data_i[283] : 
                          (N418)? in_data_i[315] : 
                          (N419)? in_data_i[347] : 
                          (N420)? in_data_i[379] : 
                          (N421)? in_data_i[411] : 
                          (N422)? in_data_i[443] : 
                          (N423)? in_data_i[475] : 
                          (N424)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[122] = (N412)? in_data_i[122] : 
                          (N413)? in_data_i[154] : 
                          (N414)? in_data_i[186] : 
                          (N415)? in_data_i[218] : 
                          (N416)? in_data_i[250] : 
                          (N417)? in_data_i[282] : 
                          (N418)? in_data_i[314] : 
                          (N419)? in_data_i[346] : 
                          (N420)? in_data_i[378] : 
                          (N421)? in_data_i[410] : 
                          (N422)? in_data_i[442] : 
                          (N423)? in_data_i[474] : 
                          (N424)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[121] = (N412)? in_data_i[121] : 
                          (N413)? in_data_i[153] : 
                          (N414)? in_data_i[185] : 
                          (N415)? in_data_i[217] : 
                          (N416)? in_data_i[249] : 
                          (N417)? in_data_i[281] : 
                          (N418)? in_data_i[313] : 
                          (N419)? in_data_i[345] : 
                          (N420)? in_data_i[377] : 
                          (N421)? in_data_i[409] : 
                          (N422)? in_data_i[441] : 
                          (N423)? in_data_i[473] : 
                          (N424)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[120] = (N412)? in_data_i[120] : 
                          (N413)? in_data_i[152] : 
                          (N414)? in_data_i[184] : 
                          (N415)? in_data_i[216] : 
                          (N416)? in_data_i[248] : 
                          (N417)? in_data_i[280] : 
                          (N418)? in_data_i[312] : 
                          (N419)? in_data_i[344] : 
                          (N420)? in_data_i[376] : 
                          (N421)? in_data_i[408] : 
                          (N422)? in_data_i[440] : 
                          (N423)? in_data_i[472] : 
                          (N424)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[119] = (N412)? in_data_i[119] : 
                          (N413)? in_data_i[151] : 
                          (N414)? in_data_i[183] : 
                          (N415)? in_data_i[215] : 
                          (N416)? in_data_i[247] : 
                          (N417)? in_data_i[279] : 
                          (N418)? in_data_i[311] : 
                          (N419)? in_data_i[343] : 
                          (N420)? in_data_i[375] : 
                          (N421)? in_data_i[407] : 
                          (N422)? in_data_i[439] : 
                          (N423)? in_data_i[471] : 
                          (N424)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[118] = (N412)? in_data_i[118] : 
                          (N413)? in_data_i[150] : 
                          (N414)? in_data_i[182] : 
                          (N415)? in_data_i[214] : 
                          (N416)? in_data_i[246] : 
                          (N417)? in_data_i[278] : 
                          (N418)? in_data_i[310] : 
                          (N419)? in_data_i[342] : 
                          (N420)? in_data_i[374] : 
                          (N421)? in_data_i[406] : 
                          (N422)? in_data_i[438] : 
                          (N423)? in_data_i[470] : 
                          (N424)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[117] = (N412)? in_data_i[117] : 
                          (N413)? in_data_i[149] : 
                          (N414)? in_data_i[181] : 
                          (N415)? in_data_i[213] : 
                          (N416)? in_data_i[245] : 
                          (N417)? in_data_i[277] : 
                          (N418)? in_data_i[309] : 
                          (N419)? in_data_i[341] : 
                          (N420)? in_data_i[373] : 
                          (N421)? in_data_i[405] : 
                          (N422)? in_data_i[437] : 
                          (N423)? in_data_i[469] : 
                          (N424)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[116] = (N412)? in_data_i[116] : 
                          (N413)? in_data_i[148] : 
                          (N414)? in_data_i[180] : 
                          (N415)? in_data_i[212] : 
                          (N416)? in_data_i[244] : 
                          (N417)? in_data_i[276] : 
                          (N418)? in_data_i[308] : 
                          (N419)? in_data_i[340] : 
                          (N420)? in_data_i[372] : 
                          (N421)? in_data_i[404] : 
                          (N422)? in_data_i[436] : 
                          (N423)? in_data_i[468] : 
                          (N424)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[115] = (N412)? in_data_i[115] : 
                          (N413)? in_data_i[147] : 
                          (N414)? in_data_i[179] : 
                          (N415)? in_data_i[211] : 
                          (N416)? in_data_i[243] : 
                          (N417)? in_data_i[275] : 
                          (N418)? in_data_i[307] : 
                          (N419)? in_data_i[339] : 
                          (N420)? in_data_i[371] : 
                          (N421)? in_data_i[403] : 
                          (N422)? in_data_i[435] : 
                          (N423)? in_data_i[467] : 
                          (N424)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[114] = (N412)? in_data_i[114] : 
                          (N413)? in_data_i[146] : 
                          (N414)? in_data_i[178] : 
                          (N415)? in_data_i[210] : 
                          (N416)? in_data_i[242] : 
                          (N417)? in_data_i[274] : 
                          (N418)? in_data_i[306] : 
                          (N419)? in_data_i[338] : 
                          (N420)? in_data_i[370] : 
                          (N421)? in_data_i[402] : 
                          (N422)? in_data_i[434] : 
                          (N423)? in_data_i[466] : 
                          (N424)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[113] = (N412)? in_data_i[113] : 
                          (N413)? in_data_i[145] : 
                          (N414)? in_data_i[177] : 
                          (N415)? in_data_i[209] : 
                          (N416)? in_data_i[241] : 
                          (N417)? in_data_i[273] : 
                          (N418)? in_data_i[305] : 
                          (N419)? in_data_i[337] : 
                          (N420)? in_data_i[369] : 
                          (N421)? in_data_i[401] : 
                          (N422)? in_data_i[433] : 
                          (N423)? in_data_i[465] : 
                          (N424)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[112] = (N412)? in_data_i[112] : 
                          (N413)? in_data_i[144] : 
                          (N414)? in_data_i[176] : 
                          (N415)? in_data_i[208] : 
                          (N416)? in_data_i[240] : 
                          (N417)? in_data_i[272] : 
                          (N418)? in_data_i[304] : 
                          (N419)? in_data_i[336] : 
                          (N420)? in_data_i[368] : 
                          (N421)? in_data_i[400] : 
                          (N422)? in_data_i[432] : 
                          (N423)? in_data_i[464] : 
                          (N424)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[111] = (N412)? in_data_i[111] : 
                          (N413)? in_data_i[143] : 
                          (N414)? in_data_i[175] : 
                          (N415)? in_data_i[207] : 
                          (N416)? in_data_i[239] : 
                          (N417)? in_data_i[271] : 
                          (N418)? in_data_i[303] : 
                          (N419)? in_data_i[335] : 
                          (N420)? in_data_i[367] : 
                          (N421)? in_data_i[399] : 
                          (N422)? in_data_i[431] : 
                          (N423)? in_data_i[463] : 
                          (N424)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[110] = (N412)? in_data_i[110] : 
                          (N413)? in_data_i[142] : 
                          (N414)? in_data_i[174] : 
                          (N415)? in_data_i[206] : 
                          (N416)? in_data_i[238] : 
                          (N417)? in_data_i[270] : 
                          (N418)? in_data_i[302] : 
                          (N419)? in_data_i[334] : 
                          (N420)? in_data_i[366] : 
                          (N421)? in_data_i[398] : 
                          (N422)? in_data_i[430] : 
                          (N423)? in_data_i[462] : 
                          (N424)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[109] = (N412)? in_data_i[109] : 
                          (N413)? in_data_i[141] : 
                          (N414)? in_data_i[173] : 
                          (N415)? in_data_i[205] : 
                          (N416)? in_data_i[237] : 
                          (N417)? in_data_i[269] : 
                          (N418)? in_data_i[301] : 
                          (N419)? in_data_i[333] : 
                          (N420)? in_data_i[365] : 
                          (N421)? in_data_i[397] : 
                          (N422)? in_data_i[429] : 
                          (N423)? in_data_i[461] : 
                          (N424)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[108] = (N412)? in_data_i[108] : 
                          (N413)? in_data_i[140] : 
                          (N414)? in_data_i[172] : 
                          (N415)? in_data_i[204] : 
                          (N416)? in_data_i[236] : 
                          (N417)? in_data_i[268] : 
                          (N418)? in_data_i[300] : 
                          (N419)? in_data_i[332] : 
                          (N420)? in_data_i[364] : 
                          (N421)? in_data_i[396] : 
                          (N422)? in_data_i[428] : 
                          (N423)? in_data_i[460] : 
                          (N424)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[107] = (N412)? in_data_i[107] : 
                          (N413)? in_data_i[139] : 
                          (N414)? in_data_i[171] : 
                          (N415)? in_data_i[203] : 
                          (N416)? in_data_i[235] : 
                          (N417)? in_data_i[267] : 
                          (N418)? in_data_i[299] : 
                          (N419)? in_data_i[331] : 
                          (N420)? in_data_i[363] : 
                          (N421)? in_data_i[395] : 
                          (N422)? in_data_i[427] : 
                          (N423)? in_data_i[459] : 
                          (N424)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[106] = (N412)? in_data_i[106] : 
                          (N413)? in_data_i[138] : 
                          (N414)? in_data_i[170] : 
                          (N415)? in_data_i[202] : 
                          (N416)? in_data_i[234] : 
                          (N417)? in_data_i[266] : 
                          (N418)? in_data_i[298] : 
                          (N419)? in_data_i[330] : 
                          (N420)? in_data_i[362] : 
                          (N421)? in_data_i[394] : 
                          (N422)? in_data_i[426] : 
                          (N423)? in_data_i[458] : 
                          (N424)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[105] = (N412)? in_data_i[105] : 
                          (N413)? in_data_i[137] : 
                          (N414)? in_data_i[169] : 
                          (N415)? in_data_i[201] : 
                          (N416)? in_data_i[233] : 
                          (N417)? in_data_i[265] : 
                          (N418)? in_data_i[297] : 
                          (N419)? in_data_i[329] : 
                          (N420)? in_data_i[361] : 
                          (N421)? in_data_i[393] : 
                          (N422)? in_data_i[425] : 
                          (N423)? in_data_i[457] : 
                          (N424)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[104] = (N412)? in_data_i[104] : 
                          (N413)? in_data_i[136] : 
                          (N414)? in_data_i[168] : 
                          (N415)? in_data_i[200] : 
                          (N416)? in_data_i[232] : 
                          (N417)? in_data_i[264] : 
                          (N418)? in_data_i[296] : 
                          (N419)? in_data_i[328] : 
                          (N420)? in_data_i[360] : 
                          (N421)? in_data_i[392] : 
                          (N422)? in_data_i[424] : 
                          (N423)? in_data_i[456] : 
                          (N424)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[103] = (N412)? in_data_i[103] : 
                          (N413)? in_data_i[135] : 
                          (N414)? in_data_i[167] : 
                          (N415)? in_data_i[199] : 
                          (N416)? in_data_i[231] : 
                          (N417)? in_data_i[263] : 
                          (N418)? in_data_i[295] : 
                          (N419)? in_data_i[327] : 
                          (N420)? in_data_i[359] : 
                          (N421)? in_data_i[391] : 
                          (N422)? in_data_i[423] : 
                          (N423)? in_data_i[455] : 
                          (N424)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[102] = (N412)? in_data_i[102] : 
                          (N413)? in_data_i[134] : 
                          (N414)? in_data_i[166] : 
                          (N415)? in_data_i[198] : 
                          (N416)? in_data_i[230] : 
                          (N417)? in_data_i[262] : 
                          (N418)? in_data_i[294] : 
                          (N419)? in_data_i[326] : 
                          (N420)? in_data_i[358] : 
                          (N421)? in_data_i[390] : 
                          (N422)? in_data_i[422] : 
                          (N423)? in_data_i[454] : 
                          (N424)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[101] = (N412)? in_data_i[101] : 
                          (N413)? in_data_i[133] : 
                          (N414)? in_data_i[165] : 
                          (N415)? in_data_i[197] : 
                          (N416)? in_data_i[229] : 
                          (N417)? in_data_i[261] : 
                          (N418)? in_data_i[293] : 
                          (N419)? in_data_i[325] : 
                          (N420)? in_data_i[357] : 
                          (N421)? in_data_i[389] : 
                          (N422)? in_data_i[421] : 
                          (N423)? in_data_i[453] : 
                          (N424)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[100] = (N412)? in_data_i[100] : 
                          (N413)? in_data_i[132] : 
                          (N414)? in_data_i[164] : 
                          (N415)? in_data_i[196] : 
                          (N416)? in_data_i[228] : 
                          (N417)? in_data_i[260] : 
                          (N418)? in_data_i[292] : 
                          (N419)? in_data_i[324] : 
                          (N420)? in_data_i[356] : 
                          (N421)? in_data_i[388] : 
                          (N422)? in_data_i[420] : 
                          (N423)? in_data_i[452] : 
                          (N424)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[99] = (N412)? in_data_i[99] : 
                         (N413)? in_data_i[131] : 
                         (N414)? in_data_i[163] : 
                         (N415)? in_data_i[195] : 
                         (N416)? in_data_i[227] : 
                         (N417)? in_data_i[259] : 
                         (N418)? in_data_i[291] : 
                         (N419)? in_data_i[323] : 
                         (N420)? in_data_i[355] : 
                         (N421)? in_data_i[387] : 
                         (N422)? in_data_i[419] : 
                         (N423)? in_data_i[451] : 
                         (N424)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[98] = (N412)? in_data_i[98] : 
                         (N413)? in_data_i[130] : 
                         (N414)? in_data_i[162] : 
                         (N415)? in_data_i[194] : 
                         (N416)? in_data_i[226] : 
                         (N417)? in_data_i[258] : 
                         (N418)? in_data_i[290] : 
                         (N419)? in_data_i[322] : 
                         (N420)? in_data_i[354] : 
                         (N421)? in_data_i[386] : 
                         (N422)? in_data_i[418] : 
                         (N423)? in_data_i[450] : 
                         (N424)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[97] = (N412)? in_data_i[97] : 
                         (N413)? in_data_i[129] : 
                         (N414)? in_data_i[161] : 
                         (N415)? in_data_i[193] : 
                         (N416)? in_data_i[225] : 
                         (N417)? in_data_i[257] : 
                         (N418)? in_data_i[289] : 
                         (N419)? in_data_i[321] : 
                         (N420)? in_data_i[353] : 
                         (N421)? in_data_i[385] : 
                         (N422)? in_data_i[417] : 
                         (N423)? in_data_i[449] : 
                         (N424)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[96] = (N412)? in_data_i[96] : 
                         (N413)? in_data_i[128] : 
                         (N414)? in_data_i[160] : 
                         (N415)? in_data_i[192] : 
                         (N416)? in_data_i[224] : 
                         (N417)? in_data_i[256] : 
                         (N418)? in_data_i[288] : 
                         (N419)? in_data_i[320] : 
                         (N420)? in_data_i[352] : 
                         (N421)? in_data_i[384] : 
                         (N422)? in_data_i[416] : 
                         (N423)? in_data_i[448] : 
                         (N424)? in_data_i_15__0_ : 1'b0;
  assign in_data_o[95] = (N425)? in_data_i[95] : 
                         (N426)? in_data_i[127] : 
                         (N427)? in_data_i[159] : 
                         (N428)? in_data_i[191] : 
                         (N429)? in_data_i[223] : 
                         (N430)? in_data_i[255] : 
                         (N431)? in_data_i[287] : 
                         (N432)? in_data_i[319] : 
                         (N433)? in_data_i[351] : 
                         (N434)? in_data_i[383] : 
                         (N435)? in_data_i[415] : 
                         (N436)? in_data_i[447] : 
                         (N437)? in_data_i[479] : 
                         (N438)? in_data_i_15__31_ : 1'b0;
  assign N425 = N850;
  assign N426 = N852;
  assign N427 = N854;
  assign N428 = N856;
  assign N429 = N858;
  assign N430 = N860;
  assign N431 = N862;
  assign N432 = N863;
  assign N433 = N851;
  assign N434 = N853;
  assign N435 = N855;
  assign N436 = N857;
  assign N437 = N859;
  assign N438 = N861;
  assign in_data_o[94] = (N425)? in_data_i[94] : 
                         (N426)? in_data_i[126] : 
                         (N427)? in_data_i[158] : 
                         (N428)? in_data_i[190] : 
                         (N429)? in_data_i[222] : 
                         (N430)? in_data_i[254] : 
                         (N431)? in_data_i[286] : 
                         (N432)? in_data_i[318] : 
                         (N433)? in_data_i[350] : 
                         (N434)? in_data_i[382] : 
                         (N435)? in_data_i[414] : 
                         (N436)? in_data_i[446] : 
                         (N437)? in_data_i[478] : 
                         (N438)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[93] = (N425)? in_data_i[93] : 
                         (N426)? in_data_i[125] : 
                         (N427)? in_data_i[157] : 
                         (N428)? in_data_i[189] : 
                         (N429)? in_data_i[221] : 
                         (N430)? in_data_i[253] : 
                         (N431)? in_data_i[285] : 
                         (N432)? in_data_i[317] : 
                         (N433)? in_data_i[349] : 
                         (N434)? in_data_i[381] : 
                         (N435)? in_data_i[413] : 
                         (N436)? in_data_i[445] : 
                         (N437)? in_data_i[477] : 
                         (N438)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[92] = (N425)? in_data_i[92] : 
                         (N426)? in_data_i[124] : 
                         (N427)? in_data_i[156] : 
                         (N428)? in_data_i[188] : 
                         (N429)? in_data_i[220] : 
                         (N430)? in_data_i[252] : 
                         (N431)? in_data_i[284] : 
                         (N432)? in_data_i[316] : 
                         (N433)? in_data_i[348] : 
                         (N434)? in_data_i[380] : 
                         (N435)? in_data_i[412] : 
                         (N436)? in_data_i[444] : 
                         (N437)? in_data_i[476] : 
                         (N438)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[91] = (N425)? in_data_i[91] : 
                         (N426)? in_data_i[123] : 
                         (N427)? in_data_i[155] : 
                         (N428)? in_data_i[187] : 
                         (N429)? in_data_i[219] : 
                         (N430)? in_data_i[251] : 
                         (N431)? in_data_i[283] : 
                         (N432)? in_data_i[315] : 
                         (N433)? in_data_i[347] : 
                         (N434)? in_data_i[379] : 
                         (N435)? in_data_i[411] : 
                         (N436)? in_data_i[443] : 
                         (N437)? in_data_i[475] : 
                         (N438)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[90] = (N425)? in_data_i[90] : 
                         (N426)? in_data_i[122] : 
                         (N427)? in_data_i[154] : 
                         (N428)? in_data_i[186] : 
                         (N429)? in_data_i[218] : 
                         (N430)? in_data_i[250] : 
                         (N431)? in_data_i[282] : 
                         (N432)? in_data_i[314] : 
                         (N433)? in_data_i[346] : 
                         (N434)? in_data_i[378] : 
                         (N435)? in_data_i[410] : 
                         (N436)? in_data_i[442] : 
                         (N437)? in_data_i[474] : 
                         (N438)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[89] = (N425)? in_data_i[89] : 
                         (N426)? in_data_i[121] : 
                         (N427)? in_data_i[153] : 
                         (N428)? in_data_i[185] : 
                         (N429)? in_data_i[217] : 
                         (N430)? in_data_i[249] : 
                         (N431)? in_data_i[281] : 
                         (N432)? in_data_i[313] : 
                         (N433)? in_data_i[345] : 
                         (N434)? in_data_i[377] : 
                         (N435)? in_data_i[409] : 
                         (N436)? in_data_i[441] : 
                         (N437)? in_data_i[473] : 
                         (N438)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[88] = (N425)? in_data_i[88] : 
                         (N426)? in_data_i[120] : 
                         (N427)? in_data_i[152] : 
                         (N428)? in_data_i[184] : 
                         (N429)? in_data_i[216] : 
                         (N430)? in_data_i[248] : 
                         (N431)? in_data_i[280] : 
                         (N432)? in_data_i[312] : 
                         (N433)? in_data_i[344] : 
                         (N434)? in_data_i[376] : 
                         (N435)? in_data_i[408] : 
                         (N436)? in_data_i[440] : 
                         (N437)? in_data_i[472] : 
                         (N438)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[87] = (N425)? in_data_i[87] : 
                         (N426)? in_data_i[119] : 
                         (N427)? in_data_i[151] : 
                         (N428)? in_data_i[183] : 
                         (N429)? in_data_i[215] : 
                         (N430)? in_data_i[247] : 
                         (N431)? in_data_i[279] : 
                         (N432)? in_data_i[311] : 
                         (N433)? in_data_i[343] : 
                         (N434)? in_data_i[375] : 
                         (N435)? in_data_i[407] : 
                         (N436)? in_data_i[439] : 
                         (N437)? in_data_i[471] : 
                         (N438)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[86] = (N425)? in_data_i[86] : 
                         (N426)? in_data_i[118] : 
                         (N427)? in_data_i[150] : 
                         (N428)? in_data_i[182] : 
                         (N429)? in_data_i[214] : 
                         (N430)? in_data_i[246] : 
                         (N431)? in_data_i[278] : 
                         (N432)? in_data_i[310] : 
                         (N433)? in_data_i[342] : 
                         (N434)? in_data_i[374] : 
                         (N435)? in_data_i[406] : 
                         (N436)? in_data_i[438] : 
                         (N437)? in_data_i[470] : 
                         (N438)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[85] = (N425)? in_data_i[85] : 
                         (N426)? in_data_i[117] : 
                         (N427)? in_data_i[149] : 
                         (N428)? in_data_i[181] : 
                         (N429)? in_data_i[213] : 
                         (N430)? in_data_i[245] : 
                         (N431)? in_data_i[277] : 
                         (N432)? in_data_i[309] : 
                         (N433)? in_data_i[341] : 
                         (N434)? in_data_i[373] : 
                         (N435)? in_data_i[405] : 
                         (N436)? in_data_i[437] : 
                         (N437)? in_data_i[469] : 
                         (N438)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[84] = (N425)? in_data_i[84] : 
                         (N426)? in_data_i[116] : 
                         (N427)? in_data_i[148] : 
                         (N428)? in_data_i[180] : 
                         (N429)? in_data_i[212] : 
                         (N430)? in_data_i[244] : 
                         (N431)? in_data_i[276] : 
                         (N432)? in_data_i[308] : 
                         (N433)? in_data_i[340] : 
                         (N434)? in_data_i[372] : 
                         (N435)? in_data_i[404] : 
                         (N436)? in_data_i[436] : 
                         (N437)? in_data_i[468] : 
                         (N438)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[83] = (N425)? in_data_i[83] : 
                         (N426)? in_data_i[115] : 
                         (N427)? in_data_i[147] : 
                         (N428)? in_data_i[179] : 
                         (N429)? in_data_i[211] : 
                         (N430)? in_data_i[243] : 
                         (N431)? in_data_i[275] : 
                         (N432)? in_data_i[307] : 
                         (N433)? in_data_i[339] : 
                         (N434)? in_data_i[371] : 
                         (N435)? in_data_i[403] : 
                         (N436)? in_data_i[435] : 
                         (N437)? in_data_i[467] : 
                         (N438)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[82] = (N425)? in_data_i[82] : 
                         (N426)? in_data_i[114] : 
                         (N427)? in_data_i[146] : 
                         (N428)? in_data_i[178] : 
                         (N429)? in_data_i[210] : 
                         (N430)? in_data_i[242] : 
                         (N431)? in_data_i[274] : 
                         (N432)? in_data_i[306] : 
                         (N433)? in_data_i[338] : 
                         (N434)? in_data_i[370] : 
                         (N435)? in_data_i[402] : 
                         (N436)? in_data_i[434] : 
                         (N437)? in_data_i[466] : 
                         (N438)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[81] = (N425)? in_data_i[81] : 
                         (N426)? in_data_i[113] : 
                         (N427)? in_data_i[145] : 
                         (N428)? in_data_i[177] : 
                         (N429)? in_data_i[209] : 
                         (N430)? in_data_i[241] : 
                         (N431)? in_data_i[273] : 
                         (N432)? in_data_i[305] : 
                         (N433)? in_data_i[337] : 
                         (N434)? in_data_i[369] : 
                         (N435)? in_data_i[401] : 
                         (N436)? in_data_i[433] : 
                         (N437)? in_data_i[465] : 
                         (N438)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[80] = (N425)? in_data_i[80] : 
                         (N426)? in_data_i[112] : 
                         (N427)? in_data_i[144] : 
                         (N428)? in_data_i[176] : 
                         (N429)? in_data_i[208] : 
                         (N430)? in_data_i[240] : 
                         (N431)? in_data_i[272] : 
                         (N432)? in_data_i[304] : 
                         (N433)? in_data_i[336] : 
                         (N434)? in_data_i[368] : 
                         (N435)? in_data_i[400] : 
                         (N436)? in_data_i[432] : 
                         (N437)? in_data_i[464] : 
                         (N438)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[79] = (N425)? in_data_i[79] : 
                         (N426)? in_data_i[111] : 
                         (N427)? in_data_i[143] : 
                         (N428)? in_data_i[175] : 
                         (N429)? in_data_i[207] : 
                         (N430)? in_data_i[239] : 
                         (N431)? in_data_i[271] : 
                         (N432)? in_data_i[303] : 
                         (N433)? in_data_i[335] : 
                         (N434)? in_data_i[367] : 
                         (N435)? in_data_i[399] : 
                         (N436)? in_data_i[431] : 
                         (N437)? in_data_i[463] : 
                         (N438)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[78] = (N425)? in_data_i[78] : 
                         (N426)? in_data_i[110] : 
                         (N427)? in_data_i[142] : 
                         (N428)? in_data_i[174] : 
                         (N429)? in_data_i[206] : 
                         (N430)? in_data_i[238] : 
                         (N431)? in_data_i[270] : 
                         (N432)? in_data_i[302] : 
                         (N433)? in_data_i[334] : 
                         (N434)? in_data_i[366] : 
                         (N435)? in_data_i[398] : 
                         (N436)? in_data_i[430] : 
                         (N437)? in_data_i[462] : 
                         (N438)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[77] = (N425)? in_data_i[77] : 
                         (N426)? in_data_i[109] : 
                         (N427)? in_data_i[141] : 
                         (N428)? in_data_i[173] : 
                         (N429)? in_data_i[205] : 
                         (N430)? in_data_i[237] : 
                         (N431)? in_data_i[269] : 
                         (N432)? in_data_i[301] : 
                         (N433)? in_data_i[333] : 
                         (N434)? in_data_i[365] : 
                         (N435)? in_data_i[397] : 
                         (N436)? in_data_i[429] : 
                         (N437)? in_data_i[461] : 
                         (N438)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[76] = (N425)? in_data_i[76] : 
                         (N426)? in_data_i[108] : 
                         (N427)? in_data_i[140] : 
                         (N428)? in_data_i[172] : 
                         (N429)? in_data_i[204] : 
                         (N430)? in_data_i[236] : 
                         (N431)? in_data_i[268] : 
                         (N432)? in_data_i[300] : 
                         (N433)? in_data_i[332] : 
                         (N434)? in_data_i[364] : 
                         (N435)? in_data_i[396] : 
                         (N436)? in_data_i[428] : 
                         (N437)? in_data_i[460] : 
                         (N438)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[75] = (N425)? in_data_i[75] : 
                         (N426)? in_data_i[107] : 
                         (N427)? in_data_i[139] : 
                         (N428)? in_data_i[171] : 
                         (N429)? in_data_i[203] : 
                         (N430)? in_data_i[235] : 
                         (N431)? in_data_i[267] : 
                         (N432)? in_data_i[299] : 
                         (N433)? in_data_i[331] : 
                         (N434)? in_data_i[363] : 
                         (N435)? in_data_i[395] : 
                         (N436)? in_data_i[427] : 
                         (N437)? in_data_i[459] : 
                         (N438)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[74] = (N425)? in_data_i[74] : 
                         (N426)? in_data_i[106] : 
                         (N427)? in_data_i[138] : 
                         (N428)? in_data_i[170] : 
                         (N429)? in_data_i[202] : 
                         (N430)? in_data_i[234] : 
                         (N431)? in_data_i[266] : 
                         (N432)? in_data_i[298] : 
                         (N433)? in_data_i[330] : 
                         (N434)? in_data_i[362] : 
                         (N435)? in_data_i[394] : 
                         (N436)? in_data_i[426] : 
                         (N437)? in_data_i[458] : 
                         (N438)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[73] = (N425)? in_data_i[73] : 
                         (N426)? in_data_i[105] : 
                         (N427)? in_data_i[137] : 
                         (N428)? in_data_i[169] : 
                         (N429)? in_data_i[201] : 
                         (N430)? in_data_i[233] : 
                         (N431)? in_data_i[265] : 
                         (N432)? in_data_i[297] : 
                         (N433)? in_data_i[329] : 
                         (N434)? in_data_i[361] : 
                         (N435)? in_data_i[393] : 
                         (N436)? in_data_i[425] : 
                         (N437)? in_data_i[457] : 
                         (N438)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[72] = (N425)? in_data_i[72] : 
                         (N426)? in_data_i[104] : 
                         (N427)? in_data_i[136] : 
                         (N428)? in_data_i[168] : 
                         (N429)? in_data_i[200] : 
                         (N430)? in_data_i[232] : 
                         (N431)? in_data_i[264] : 
                         (N432)? in_data_i[296] : 
                         (N433)? in_data_i[328] : 
                         (N434)? in_data_i[360] : 
                         (N435)? in_data_i[392] : 
                         (N436)? in_data_i[424] : 
                         (N437)? in_data_i[456] : 
                         (N438)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[71] = (N425)? in_data_i[71] : 
                         (N426)? in_data_i[103] : 
                         (N427)? in_data_i[135] : 
                         (N428)? in_data_i[167] : 
                         (N429)? in_data_i[199] : 
                         (N430)? in_data_i[231] : 
                         (N431)? in_data_i[263] : 
                         (N432)? in_data_i[295] : 
                         (N433)? in_data_i[327] : 
                         (N434)? in_data_i[359] : 
                         (N435)? in_data_i[391] : 
                         (N436)? in_data_i[423] : 
                         (N437)? in_data_i[455] : 
                         (N438)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[70] = (N425)? in_data_i[70] : 
                         (N426)? in_data_i[102] : 
                         (N427)? in_data_i[134] : 
                         (N428)? in_data_i[166] : 
                         (N429)? in_data_i[198] : 
                         (N430)? in_data_i[230] : 
                         (N431)? in_data_i[262] : 
                         (N432)? in_data_i[294] : 
                         (N433)? in_data_i[326] : 
                         (N434)? in_data_i[358] : 
                         (N435)? in_data_i[390] : 
                         (N436)? in_data_i[422] : 
                         (N437)? in_data_i[454] : 
                         (N438)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[69] = (N425)? in_data_i[69] : 
                         (N426)? in_data_i[101] : 
                         (N427)? in_data_i[133] : 
                         (N428)? in_data_i[165] : 
                         (N429)? in_data_i[197] : 
                         (N430)? in_data_i[229] : 
                         (N431)? in_data_i[261] : 
                         (N432)? in_data_i[293] : 
                         (N433)? in_data_i[325] : 
                         (N434)? in_data_i[357] : 
                         (N435)? in_data_i[389] : 
                         (N436)? in_data_i[421] : 
                         (N437)? in_data_i[453] : 
                         (N438)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[68] = (N425)? in_data_i[68] : 
                         (N426)? in_data_i[100] : 
                         (N427)? in_data_i[132] : 
                         (N428)? in_data_i[164] : 
                         (N429)? in_data_i[196] : 
                         (N430)? in_data_i[228] : 
                         (N431)? in_data_i[260] : 
                         (N432)? in_data_i[292] : 
                         (N433)? in_data_i[324] : 
                         (N434)? in_data_i[356] : 
                         (N435)? in_data_i[388] : 
                         (N436)? in_data_i[420] : 
                         (N437)? in_data_i[452] : 
                         (N438)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[67] = (N425)? in_data_i[67] : 
                         (N426)? in_data_i[99] : 
                         (N427)? in_data_i[131] : 
                         (N428)? in_data_i[163] : 
                         (N429)? in_data_i[195] : 
                         (N430)? in_data_i[227] : 
                         (N431)? in_data_i[259] : 
                         (N432)? in_data_i[291] : 
                         (N433)? in_data_i[323] : 
                         (N434)? in_data_i[355] : 
                         (N435)? in_data_i[387] : 
                         (N436)? in_data_i[419] : 
                         (N437)? in_data_i[451] : 
                         (N438)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[66] = (N425)? in_data_i[66] : 
                         (N426)? in_data_i[98] : 
                         (N427)? in_data_i[130] : 
                         (N428)? in_data_i[162] : 
                         (N429)? in_data_i[194] : 
                         (N430)? in_data_i[226] : 
                         (N431)? in_data_i[258] : 
                         (N432)? in_data_i[290] : 
                         (N433)? in_data_i[322] : 
                         (N434)? in_data_i[354] : 
                         (N435)? in_data_i[386] : 
                         (N436)? in_data_i[418] : 
                         (N437)? in_data_i[450] : 
                         (N438)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[65] = (N425)? in_data_i[65] : 
                         (N426)? in_data_i[97] : 
                         (N427)? in_data_i[129] : 
                         (N428)? in_data_i[161] : 
                         (N429)? in_data_i[193] : 
                         (N430)? in_data_i[225] : 
                         (N431)? in_data_i[257] : 
                         (N432)? in_data_i[289] : 
                         (N433)? in_data_i[321] : 
                         (N434)? in_data_i[353] : 
                         (N435)? in_data_i[385] : 
                         (N436)? in_data_i[417] : 
                         (N437)? in_data_i[449] : 
                         (N438)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[64] = (N425)? in_data_i[64] : 
                         (N426)? in_data_i[96] : 
                         (N427)? in_data_i[128] : 
                         (N428)? in_data_i[160] : 
                         (N429)? in_data_i[192] : 
                         (N430)? in_data_i[224] : 
                         (N431)? in_data_i[256] : 
                         (N432)? in_data_i[288] : 
                         (N433)? in_data_i[320] : 
                         (N434)? in_data_i[352] : 
                         (N435)? in_data_i[384] : 
                         (N436)? in_data_i[416] : 
                         (N437)? in_data_i[448] : 
                         (N438)? in_data_i_15__0_ : 1'b0;
  assign in_data_o[63] = (N439)? in_data_i[63] : 
                         (N440)? in_data_i[95] : 
                         (N441)? in_data_i[127] : 
                         (N442)? in_data_i[159] : 
                         (N443)? in_data_i[191] : 
                         (N444)? in_data_i[223] : 
                         (N445)? in_data_i[255] : 
                         (N446)? in_data_i[287] : 
                         (N447)? in_data_i[319] : 
                         (N448)? in_data_i[351] : 
                         (N449)? in_data_i[383] : 
                         (N450)? in_data_i[415] : 
                         (N451)? in_data_i[447] : 
                         (N452)? in_data_i[479] : 
                         (N453)? in_data_i_15__31_ : 1'b0;
  assign N439 = N726;
  assign N440 = N728;
  assign N441 = N730;
  assign N442 = N732;
  assign N443 = N734;
  assign N444 = N736;
  assign N445 = N738;
  assign N446 = N740;
  assign N447 = N727;
  assign N448 = N729;
  assign N449 = N731;
  assign N450 = N733;
  assign N451 = N735;
  assign N452 = N737;
  assign N453 = N739;
  assign in_data_o[62] = (N439)? in_data_i[62] : 
                         (N440)? in_data_i[94] : 
                         (N441)? in_data_i[126] : 
                         (N442)? in_data_i[158] : 
                         (N443)? in_data_i[190] : 
                         (N444)? in_data_i[222] : 
                         (N445)? in_data_i[254] : 
                         (N446)? in_data_i[286] : 
                         (N447)? in_data_i[318] : 
                         (N448)? in_data_i[350] : 
                         (N449)? in_data_i[382] : 
                         (N450)? in_data_i[414] : 
                         (N451)? in_data_i[446] : 
                         (N452)? in_data_i[478] : 
                         (N453)? in_data_i_15__30_ : 1'b0;
  assign in_data_o[61] = (N439)? in_data_i[61] : 
                         (N440)? in_data_i[93] : 
                         (N441)? in_data_i[125] : 
                         (N442)? in_data_i[157] : 
                         (N443)? in_data_i[189] : 
                         (N444)? in_data_i[221] : 
                         (N445)? in_data_i[253] : 
                         (N446)? in_data_i[285] : 
                         (N447)? in_data_i[317] : 
                         (N448)? in_data_i[349] : 
                         (N449)? in_data_i[381] : 
                         (N450)? in_data_i[413] : 
                         (N451)? in_data_i[445] : 
                         (N452)? in_data_i[477] : 
                         (N453)? in_data_i_15__29_ : 1'b0;
  assign in_data_o[60] = (N439)? in_data_i[60] : 
                         (N440)? in_data_i[92] : 
                         (N441)? in_data_i[124] : 
                         (N442)? in_data_i[156] : 
                         (N443)? in_data_i[188] : 
                         (N444)? in_data_i[220] : 
                         (N445)? in_data_i[252] : 
                         (N446)? in_data_i[284] : 
                         (N447)? in_data_i[316] : 
                         (N448)? in_data_i[348] : 
                         (N449)? in_data_i[380] : 
                         (N450)? in_data_i[412] : 
                         (N451)? in_data_i[444] : 
                         (N452)? in_data_i[476] : 
                         (N453)? in_data_i_15__28_ : 1'b0;
  assign in_data_o[59] = (N439)? in_data_i[59] : 
                         (N440)? in_data_i[91] : 
                         (N441)? in_data_i[123] : 
                         (N442)? in_data_i[155] : 
                         (N443)? in_data_i[187] : 
                         (N444)? in_data_i[219] : 
                         (N445)? in_data_i[251] : 
                         (N446)? in_data_i[283] : 
                         (N447)? in_data_i[315] : 
                         (N448)? in_data_i[347] : 
                         (N449)? in_data_i[379] : 
                         (N450)? in_data_i[411] : 
                         (N451)? in_data_i[443] : 
                         (N452)? in_data_i[475] : 
                         (N453)? in_data_i_15__27_ : 1'b0;
  assign in_data_o[58] = (N439)? in_data_i[58] : 
                         (N440)? in_data_i[90] : 
                         (N441)? in_data_i[122] : 
                         (N442)? in_data_i[154] : 
                         (N443)? in_data_i[186] : 
                         (N444)? in_data_i[218] : 
                         (N445)? in_data_i[250] : 
                         (N446)? in_data_i[282] : 
                         (N447)? in_data_i[314] : 
                         (N448)? in_data_i[346] : 
                         (N449)? in_data_i[378] : 
                         (N450)? in_data_i[410] : 
                         (N451)? in_data_i[442] : 
                         (N452)? in_data_i[474] : 
                         (N453)? in_data_i_15__26_ : 1'b0;
  assign in_data_o[57] = (N439)? in_data_i[57] : 
                         (N440)? in_data_i[89] : 
                         (N441)? in_data_i[121] : 
                         (N442)? in_data_i[153] : 
                         (N443)? in_data_i[185] : 
                         (N444)? in_data_i[217] : 
                         (N445)? in_data_i[249] : 
                         (N446)? in_data_i[281] : 
                         (N447)? in_data_i[313] : 
                         (N448)? in_data_i[345] : 
                         (N449)? in_data_i[377] : 
                         (N450)? in_data_i[409] : 
                         (N451)? in_data_i[441] : 
                         (N452)? in_data_i[473] : 
                         (N453)? in_data_i_15__25_ : 1'b0;
  assign in_data_o[56] = (N439)? in_data_i[56] : 
                         (N440)? in_data_i[88] : 
                         (N441)? in_data_i[120] : 
                         (N442)? in_data_i[152] : 
                         (N443)? in_data_i[184] : 
                         (N444)? in_data_i[216] : 
                         (N445)? in_data_i[248] : 
                         (N446)? in_data_i[280] : 
                         (N447)? in_data_i[312] : 
                         (N448)? in_data_i[344] : 
                         (N449)? in_data_i[376] : 
                         (N450)? in_data_i[408] : 
                         (N451)? in_data_i[440] : 
                         (N452)? in_data_i[472] : 
                         (N453)? in_data_i_15__24_ : 1'b0;
  assign in_data_o[55] = (N439)? in_data_i[55] : 
                         (N440)? in_data_i[87] : 
                         (N441)? in_data_i[119] : 
                         (N442)? in_data_i[151] : 
                         (N443)? in_data_i[183] : 
                         (N444)? in_data_i[215] : 
                         (N445)? in_data_i[247] : 
                         (N446)? in_data_i[279] : 
                         (N447)? in_data_i[311] : 
                         (N448)? in_data_i[343] : 
                         (N449)? in_data_i[375] : 
                         (N450)? in_data_i[407] : 
                         (N451)? in_data_i[439] : 
                         (N452)? in_data_i[471] : 
                         (N453)? in_data_i_15__23_ : 1'b0;
  assign in_data_o[54] = (N439)? in_data_i[54] : 
                         (N440)? in_data_i[86] : 
                         (N441)? in_data_i[118] : 
                         (N442)? in_data_i[150] : 
                         (N443)? in_data_i[182] : 
                         (N444)? in_data_i[214] : 
                         (N445)? in_data_i[246] : 
                         (N446)? in_data_i[278] : 
                         (N447)? in_data_i[310] : 
                         (N448)? in_data_i[342] : 
                         (N449)? in_data_i[374] : 
                         (N450)? in_data_i[406] : 
                         (N451)? in_data_i[438] : 
                         (N452)? in_data_i[470] : 
                         (N453)? in_data_i_15__22_ : 1'b0;
  assign in_data_o[53] = (N439)? in_data_i[53] : 
                         (N440)? in_data_i[85] : 
                         (N441)? in_data_i[117] : 
                         (N442)? in_data_i[149] : 
                         (N443)? in_data_i[181] : 
                         (N444)? in_data_i[213] : 
                         (N445)? in_data_i[245] : 
                         (N446)? in_data_i[277] : 
                         (N447)? in_data_i[309] : 
                         (N448)? in_data_i[341] : 
                         (N449)? in_data_i[373] : 
                         (N450)? in_data_i[405] : 
                         (N451)? in_data_i[437] : 
                         (N452)? in_data_i[469] : 
                         (N453)? in_data_i_15__21_ : 1'b0;
  assign in_data_o[52] = (N439)? in_data_i[52] : 
                         (N440)? in_data_i[84] : 
                         (N441)? in_data_i[116] : 
                         (N442)? in_data_i[148] : 
                         (N443)? in_data_i[180] : 
                         (N444)? in_data_i[212] : 
                         (N445)? in_data_i[244] : 
                         (N446)? in_data_i[276] : 
                         (N447)? in_data_i[308] : 
                         (N448)? in_data_i[340] : 
                         (N449)? in_data_i[372] : 
                         (N450)? in_data_i[404] : 
                         (N451)? in_data_i[436] : 
                         (N452)? in_data_i[468] : 
                         (N453)? in_data_i_15__20_ : 1'b0;
  assign in_data_o[51] = (N439)? in_data_i[51] : 
                         (N440)? in_data_i[83] : 
                         (N441)? in_data_i[115] : 
                         (N442)? in_data_i[147] : 
                         (N443)? in_data_i[179] : 
                         (N444)? in_data_i[211] : 
                         (N445)? in_data_i[243] : 
                         (N446)? in_data_i[275] : 
                         (N447)? in_data_i[307] : 
                         (N448)? in_data_i[339] : 
                         (N449)? in_data_i[371] : 
                         (N450)? in_data_i[403] : 
                         (N451)? in_data_i[435] : 
                         (N452)? in_data_i[467] : 
                         (N453)? in_data_i_15__19_ : 1'b0;
  assign in_data_o[50] = (N439)? in_data_i[50] : 
                         (N440)? in_data_i[82] : 
                         (N441)? in_data_i[114] : 
                         (N442)? in_data_i[146] : 
                         (N443)? in_data_i[178] : 
                         (N444)? in_data_i[210] : 
                         (N445)? in_data_i[242] : 
                         (N446)? in_data_i[274] : 
                         (N447)? in_data_i[306] : 
                         (N448)? in_data_i[338] : 
                         (N449)? in_data_i[370] : 
                         (N450)? in_data_i[402] : 
                         (N451)? in_data_i[434] : 
                         (N452)? in_data_i[466] : 
                         (N453)? in_data_i_15__18_ : 1'b0;
  assign in_data_o[49] = (N439)? in_data_i[49] : 
                         (N440)? in_data_i[81] : 
                         (N441)? in_data_i[113] : 
                         (N442)? in_data_i[145] : 
                         (N443)? in_data_i[177] : 
                         (N444)? in_data_i[209] : 
                         (N445)? in_data_i[241] : 
                         (N446)? in_data_i[273] : 
                         (N447)? in_data_i[305] : 
                         (N448)? in_data_i[337] : 
                         (N449)? in_data_i[369] : 
                         (N450)? in_data_i[401] : 
                         (N451)? in_data_i[433] : 
                         (N452)? in_data_i[465] : 
                         (N453)? in_data_i_15__17_ : 1'b0;
  assign in_data_o[48] = (N439)? in_data_i[48] : 
                         (N440)? in_data_i[80] : 
                         (N441)? in_data_i[112] : 
                         (N442)? in_data_i[144] : 
                         (N443)? in_data_i[176] : 
                         (N444)? in_data_i[208] : 
                         (N445)? in_data_i[240] : 
                         (N446)? in_data_i[272] : 
                         (N447)? in_data_i[304] : 
                         (N448)? in_data_i[336] : 
                         (N449)? in_data_i[368] : 
                         (N450)? in_data_i[400] : 
                         (N451)? in_data_i[432] : 
                         (N452)? in_data_i[464] : 
                         (N453)? in_data_i_15__16_ : 1'b0;
  assign in_data_o[47] = (N439)? in_data_i[47] : 
                         (N440)? in_data_i[79] : 
                         (N441)? in_data_i[111] : 
                         (N442)? in_data_i[143] : 
                         (N443)? in_data_i[175] : 
                         (N444)? in_data_i[207] : 
                         (N445)? in_data_i[239] : 
                         (N446)? in_data_i[271] : 
                         (N447)? in_data_i[303] : 
                         (N448)? in_data_i[335] : 
                         (N449)? in_data_i[367] : 
                         (N450)? in_data_i[399] : 
                         (N451)? in_data_i[431] : 
                         (N452)? in_data_i[463] : 
                         (N453)? in_data_i_15__15_ : 1'b0;
  assign in_data_o[46] = (N439)? in_data_i[46] : 
                         (N440)? in_data_i[78] : 
                         (N441)? in_data_i[110] : 
                         (N442)? in_data_i[142] : 
                         (N443)? in_data_i[174] : 
                         (N444)? in_data_i[206] : 
                         (N445)? in_data_i[238] : 
                         (N446)? in_data_i[270] : 
                         (N447)? in_data_i[302] : 
                         (N448)? in_data_i[334] : 
                         (N449)? in_data_i[366] : 
                         (N450)? in_data_i[398] : 
                         (N451)? in_data_i[430] : 
                         (N452)? in_data_i[462] : 
                         (N453)? in_data_i_15__14_ : 1'b0;
  assign in_data_o[45] = (N439)? in_data_i[45] : 
                         (N440)? in_data_i[77] : 
                         (N441)? in_data_i[109] : 
                         (N442)? in_data_i[141] : 
                         (N443)? in_data_i[173] : 
                         (N444)? in_data_i[205] : 
                         (N445)? in_data_i[237] : 
                         (N446)? in_data_i[269] : 
                         (N447)? in_data_i[301] : 
                         (N448)? in_data_i[333] : 
                         (N449)? in_data_i[365] : 
                         (N450)? in_data_i[397] : 
                         (N451)? in_data_i[429] : 
                         (N452)? in_data_i[461] : 
                         (N453)? in_data_i_15__13_ : 1'b0;
  assign in_data_o[44] = (N439)? in_data_i[44] : 
                         (N440)? in_data_i[76] : 
                         (N441)? in_data_i[108] : 
                         (N442)? in_data_i[140] : 
                         (N443)? in_data_i[172] : 
                         (N444)? in_data_i[204] : 
                         (N445)? in_data_i[236] : 
                         (N446)? in_data_i[268] : 
                         (N447)? in_data_i[300] : 
                         (N448)? in_data_i[332] : 
                         (N449)? in_data_i[364] : 
                         (N450)? in_data_i[396] : 
                         (N451)? in_data_i[428] : 
                         (N452)? in_data_i[460] : 
                         (N453)? in_data_i_15__12_ : 1'b0;
  assign in_data_o[43] = (N439)? in_data_i[43] : 
                         (N440)? in_data_i[75] : 
                         (N441)? in_data_i[107] : 
                         (N442)? in_data_i[139] : 
                         (N443)? in_data_i[171] : 
                         (N444)? in_data_i[203] : 
                         (N445)? in_data_i[235] : 
                         (N446)? in_data_i[267] : 
                         (N447)? in_data_i[299] : 
                         (N448)? in_data_i[331] : 
                         (N449)? in_data_i[363] : 
                         (N450)? in_data_i[395] : 
                         (N451)? in_data_i[427] : 
                         (N452)? in_data_i[459] : 
                         (N453)? in_data_i_15__11_ : 1'b0;
  assign in_data_o[42] = (N439)? in_data_i[42] : 
                         (N440)? in_data_i[74] : 
                         (N441)? in_data_i[106] : 
                         (N442)? in_data_i[138] : 
                         (N443)? in_data_i[170] : 
                         (N444)? in_data_i[202] : 
                         (N445)? in_data_i[234] : 
                         (N446)? in_data_i[266] : 
                         (N447)? in_data_i[298] : 
                         (N448)? in_data_i[330] : 
                         (N449)? in_data_i[362] : 
                         (N450)? in_data_i[394] : 
                         (N451)? in_data_i[426] : 
                         (N452)? in_data_i[458] : 
                         (N453)? in_data_i_15__10_ : 1'b0;
  assign in_data_o[41] = (N439)? in_data_i[41] : 
                         (N440)? in_data_i[73] : 
                         (N441)? in_data_i[105] : 
                         (N442)? in_data_i[137] : 
                         (N443)? in_data_i[169] : 
                         (N444)? in_data_i[201] : 
                         (N445)? in_data_i[233] : 
                         (N446)? in_data_i[265] : 
                         (N447)? in_data_i[297] : 
                         (N448)? in_data_i[329] : 
                         (N449)? in_data_i[361] : 
                         (N450)? in_data_i[393] : 
                         (N451)? in_data_i[425] : 
                         (N452)? in_data_i[457] : 
                         (N453)? in_data_i_15__9_ : 1'b0;
  assign in_data_o[40] = (N439)? in_data_i[40] : 
                         (N440)? in_data_i[72] : 
                         (N441)? in_data_i[104] : 
                         (N442)? in_data_i[136] : 
                         (N443)? in_data_i[168] : 
                         (N444)? in_data_i[200] : 
                         (N445)? in_data_i[232] : 
                         (N446)? in_data_i[264] : 
                         (N447)? in_data_i[296] : 
                         (N448)? in_data_i[328] : 
                         (N449)? in_data_i[360] : 
                         (N450)? in_data_i[392] : 
                         (N451)? in_data_i[424] : 
                         (N452)? in_data_i[456] : 
                         (N453)? in_data_i_15__8_ : 1'b0;
  assign in_data_o[39] = (N439)? in_data_i[39] : 
                         (N440)? in_data_i[71] : 
                         (N441)? in_data_i[103] : 
                         (N442)? in_data_i[135] : 
                         (N443)? in_data_i[167] : 
                         (N444)? in_data_i[199] : 
                         (N445)? in_data_i[231] : 
                         (N446)? in_data_i[263] : 
                         (N447)? in_data_i[295] : 
                         (N448)? in_data_i[327] : 
                         (N449)? in_data_i[359] : 
                         (N450)? in_data_i[391] : 
                         (N451)? in_data_i[423] : 
                         (N452)? in_data_i[455] : 
                         (N453)? in_data_i_15__7_ : 1'b0;
  assign in_data_o[38] = (N439)? in_data_i[38] : 
                         (N440)? in_data_i[70] : 
                         (N441)? in_data_i[102] : 
                         (N442)? in_data_i[134] : 
                         (N443)? in_data_i[166] : 
                         (N444)? in_data_i[198] : 
                         (N445)? in_data_i[230] : 
                         (N446)? in_data_i[262] : 
                         (N447)? in_data_i[294] : 
                         (N448)? in_data_i[326] : 
                         (N449)? in_data_i[358] : 
                         (N450)? in_data_i[390] : 
                         (N451)? in_data_i[422] : 
                         (N452)? in_data_i[454] : 
                         (N453)? in_data_i_15__6_ : 1'b0;
  assign in_data_o[37] = (N439)? in_data_i[37] : 
                         (N440)? in_data_i[69] : 
                         (N441)? in_data_i[101] : 
                         (N442)? in_data_i[133] : 
                         (N443)? in_data_i[165] : 
                         (N444)? in_data_i[197] : 
                         (N445)? in_data_i[229] : 
                         (N446)? in_data_i[261] : 
                         (N447)? in_data_i[293] : 
                         (N448)? in_data_i[325] : 
                         (N449)? in_data_i[357] : 
                         (N450)? in_data_i[389] : 
                         (N451)? in_data_i[421] : 
                         (N452)? in_data_i[453] : 
                         (N453)? in_data_i_15__5_ : 1'b0;
  assign in_data_o[36] = (N439)? in_data_i[36] : 
                         (N440)? in_data_i[68] : 
                         (N441)? in_data_i[100] : 
                         (N442)? in_data_i[132] : 
                         (N443)? in_data_i[164] : 
                         (N444)? in_data_i[196] : 
                         (N445)? in_data_i[228] : 
                         (N446)? in_data_i[260] : 
                         (N447)? in_data_i[292] : 
                         (N448)? in_data_i[324] : 
                         (N449)? in_data_i[356] : 
                         (N450)? in_data_i[388] : 
                         (N451)? in_data_i[420] : 
                         (N452)? in_data_i[452] : 
                         (N453)? in_data_i_15__4_ : 1'b0;
  assign in_data_o[35] = (N439)? in_data_i[35] : 
                         (N440)? in_data_i[67] : 
                         (N441)? in_data_i[99] : 
                         (N442)? in_data_i[131] : 
                         (N443)? in_data_i[163] : 
                         (N444)? in_data_i[195] : 
                         (N445)? in_data_i[227] : 
                         (N446)? in_data_i[259] : 
                         (N447)? in_data_i[291] : 
                         (N448)? in_data_i[323] : 
                         (N449)? in_data_i[355] : 
                         (N450)? in_data_i[387] : 
                         (N451)? in_data_i[419] : 
                         (N452)? in_data_i[451] : 
                         (N453)? in_data_i_15__3_ : 1'b0;
  assign in_data_o[34] = (N439)? in_data_i[34] : 
                         (N440)? in_data_i[66] : 
                         (N441)? in_data_i[98] : 
                         (N442)? in_data_i[130] : 
                         (N443)? in_data_i[162] : 
                         (N444)? in_data_i[194] : 
                         (N445)? in_data_i[226] : 
                         (N446)? in_data_i[258] : 
                         (N447)? in_data_i[290] : 
                         (N448)? in_data_i[322] : 
                         (N449)? in_data_i[354] : 
                         (N450)? in_data_i[386] : 
                         (N451)? in_data_i[418] : 
                         (N452)? in_data_i[450] : 
                         (N453)? in_data_i_15__2_ : 1'b0;
  assign in_data_o[33] = (N439)? in_data_i[33] : 
                         (N440)? in_data_i[65] : 
                         (N441)? in_data_i[97] : 
                         (N442)? in_data_i[129] : 
                         (N443)? in_data_i[161] : 
                         (N444)? in_data_i[193] : 
                         (N445)? in_data_i[225] : 
                         (N446)? in_data_i[257] : 
                         (N447)? in_data_i[289] : 
                         (N448)? in_data_i[321] : 
                         (N449)? in_data_i[353] : 
                         (N450)? in_data_i[385] : 
                         (N451)? in_data_i[417] : 
                         (N452)? in_data_i[449] : 
                         (N453)? in_data_i_15__1_ : 1'b0;
  assign in_data_o[32] = (N439)? in_data_i[32] : 
                         (N440)? in_data_i[64] : 
                         (N441)? in_data_i[96] : 
                         (N442)? in_data_i[128] : 
                         (N443)? in_data_i[160] : 
                         (N444)? in_data_i[192] : 
                         (N445)? in_data_i[224] : 
                         (N446)? in_data_i[256] : 
                         (N447)? in_data_i[288] : 
                         (N448)? in_data_i[320] : 
                         (N449)? in_data_i[352] : 
                         (N450)? in_data_i[384] : 
                         (N451)? in_data_i[416] : 
                         (N452)? in_data_i[448] : 
                         (N453)? in_data_i_15__0_ : 1'b0;
  assign out_me_data_o[479] = (N454)? out_me_data_i_0__31_ : 
                              (N455)? out_me_data_i[63] : 
                              (N456)? out_me_data_i[95] : 
                              (N457)? out_me_data_i[127] : 
                              (N458)? out_me_data_i[159] : 
                              (N459)? out_me_data_i[191] : 
                              (N460)? out_me_data_i[223] : 
                              (N461)? out_me_data_i[255] : 
                              (N462)? out_me_data_i[287] : 
                              (N463)? out_me_data_i[319] : 
                              (N464)? out_me_data_i[351] : 
                              (N465)? out_me_data_i[383] : 
                              (N466)? out_me_data_i[415] : 
                              (N467)? out_me_data_i[447] : 
                              (N468)? out_me_data_i[479] : 1'b0;
  assign N454 = N2421;
  assign N455 = N2423;
  assign N456 = N2425;
  assign N457 = N2427;
  assign N458 = N2429;
  assign N459 = N2431;
  assign N460 = N2433;
  assign N461 = N2435;
  assign N462 = N2422;
  assign N463 = N2424;
  assign N464 = N2426;
  assign N465 = N2428;
  assign N466 = N2430;
  assign N467 = N2432;
  assign N468 = N2434;
  assign out_me_data_o[478] = (N454)? out_me_data_i_0__30_ : 
                              (N455)? out_me_data_i[62] : 
                              (N456)? out_me_data_i[94] : 
                              (N457)? out_me_data_i[126] : 
                              (N458)? out_me_data_i[158] : 
                              (N459)? out_me_data_i[190] : 
                              (N460)? out_me_data_i[222] : 
                              (N461)? out_me_data_i[254] : 
                              (N462)? out_me_data_i[286] : 
                              (N463)? out_me_data_i[318] : 
                              (N464)? out_me_data_i[350] : 
                              (N465)? out_me_data_i[382] : 
                              (N466)? out_me_data_i[414] : 
                              (N467)? out_me_data_i[446] : 
                              (N468)? out_me_data_i[478] : 1'b0;
  assign out_me_data_o[477] = (N454)? out_me_data_i_0__29_ : 
                              (N455)? out_me_data_i[61] : 
                              (N456)? out_me_data_i[93] : 
                              (N457)? out_me_data_i[125] : 
                              (N458)? out_me_data_i[157] : 
                              (N459)? out_me_data_i[189] : 
                              (N460)? out_me_data_i[221] : 
                              (N461)? out_me_data_i[253] : 
                              (N462)? out_me_data_i[285] : 
                              (N463)? out_me_data_i[317] : 
                              (N464)? out_me_data_i[349] : 
                              (N465)? out_me_data_i[381] : 
                              (N466)? out_me_data_i[413] : 
                              (N467)? out_me_data_i[445] : 
                              (N468)? out_me_data_i[477] : 1'b0;
  assign out_me_data_o[476] = (N454)? out_me_data_i_0__28_ : 
                              (N455)? out_me_data_i[60] : 
                              (N456)? out_me_data_i[92] : 
                              (N457)? out_me_data_i[124] : 
                              (N458)? out_me_data_i[156] : 
                              (N459)? out_me_data_i[188] : 
                              (N460)? out_me_data_i[220] : 
                              (N461)? out_me_data_i[252] : 
                              (N462)? out_me_data_i[284] : 
                              (N463)? out_me_data_i[316] : 
                              (N464)? out_me_data_i[348] : 
                              (N465)? out_me_data_i[380] : 
                              (N466)? out_me_data_i[412] : 
                              (N467)? out_me_data_i[444] : 
                              (N468)? out_me_data_i[476] : 1'b0;
  assign out_me_data_o[475] = (N454)? out_me_data_i_0__27_ : 
                              (N455)? out_me_data_i[59] : 
                              (N456)? out_me_data_i[91] : 
                              (N457)? out_me_data_i[123] : 
                              (N458)? out_me_data_i[155] : 
                              (N459)? out_me_data_i[187] : 
                              (N460)? out_me_data_i[219] : 
                              (N461)? out_me_data_i[251] : 
                              (N462)? out_me_data_i[283] : 
                              (N463)? out_me_data_i[315] : 
                              (N464)? out_me_data_i[347] : 
                              (N465)? out_me_data_i[379] : 
                              (N466)? out_me_data_i[411] : 
                              (N467)? out_me_data_i[443] : 
                              (N468)? out_me_data_i[475] : 1'b0;
  assign out_me_data_o[474] = (N454)? out_me_data_i_0__26_ : 
                              (N455)? out_me_data_i[58] : 
                              (N456)? out_me_data_i[90] : 
                              (N457)? out_me_data_i[122] : 
                              (N458)? out_me_data_i[154] : 
                              (N459)? out_me_data_i[186] : 
                              (N460)? out_me_data_i[218] : 
                              (N461)? out_me_data_i[250] : 
                              (N462)? out_me_data_i[282] : 
                              (N463)? out_me_data_i[314] : 
                              (N464)? out_me_data_i[346] : 
                              (N465)? out_me_data_i[378] : 
                              (N466)? out_me_data_i[410] : 
                              (N467)? out_me_data_i[442] : 
                              (N468)? out_me_data_i[474] : 1'b0;
  assign out_me_data_o[473] = (N454)? out_me_data_i_0__25_ : 
                              (N455)? out_me_data_i[57] : 
                              (N456)? out_me_data_i[89] : 
                              (N457)? out_me_data_i[121] : 
                              (N458)? out_me_data_i[153] : 
                              (N459)? out_me_data_i[185] : 
                              (N460)? out_me_data_i[217] : 
                              (N461)? out_me_data_i[249] : 
                              (N462)? out_me_data_i[281] : 
                              (N463)? out_me_data_i[313] : 
                              (N464)? out_me_data_i[345] : 
                              (N465)? out_me_data_i[377] : 
                              (N466)? out_me_data_i[409] : 
                              (N467)? out_me_data_i[441] : 
                              (N468)? out_me_data_i[473] : 1'b0;
  assign out_me_data_o[472] = (N454)? out_me_data_i_0__24_ : 
                              (N455)? out_me_data_i[56] : 
                              (N456)? out_me_data_i[88] : 
                              (N457)? out_me_data_i[120] : 
                              (N458)? out_me_data_i[152] : 
                              (N459)? out_me_data_i[184] : 
                              (N460)? out_me_data_i[216] : 
                              (N461)? out_me_data_i[248] : 
                              (N462)? out_me_data_i[280] : 
                              (N463)? out_me_data_i[312] : 
                              (N464)? out_me_data_i[344] : 
                              (N465)? out_me_data_i[376] : 
                              (N466)? out_me_data_i[408] : 
                              (N467)? out_me_data_i[440] : 
                              (N468)? out_me_data_i[472] : 1'b0;
  assign out_me_data_o[471] = (N454)? out_me_data_i_0__23_ : 
                              (N455)? out_me_data_i[55] : 
                              (N456)? out_me_data_i[87] : 
                              (N457)? out_me_data_i[119] : 
                              (N458)? out_me_data_i[151] : 
                              (N459)? out_me_data_i[183] : 
                              (N460)? out_me_data_i[215] : 
                              (N461)? out_me_data_i[247] : 
                              (N462)? out_me_data_i[279] : 
                              (N463)? out_me_data_i[311] : 
                              (N464)? out_me_data_i[343] : 
                              (N465)? out_me_data_i[375] : 
                              (N466)? out_me_data_i[407] : 
                              (N467)? out_me_data_i[439] : 
                              (N468)? out_me_data_i[471] : 1'b0;
  assign out_me_data_o[470] = (N454)? out_me_data_i_0__22_ : 
                              (N455)? out_me_data_i[54] : 
                              (N456)? out_me_data_i[86] : 
                              (N457)? out_me_data_i[118] : 
                              (N458)? out_me_data_i[150] : 
                              (N459)? out_me_data_i[182] : 
                              (N460)? out_me_data_i[214] : 
                              (N461)? out_me_data_i[246] : 
                              (N462)? out_me_data_i[278] : 
                              (N463)? out_me_data_i[310] : 
                              (N464)? out_me_data_i[342] : 
                              (N465)? out_me_data_i[374] : 
                              (N466)? out_me_data_i[406] : 
                              (N467)? out_me_data_i[438] : 
                              (N468)? out_me_data_i[470] : 1'b0;
  assign out_me_data_o[469] = (N454)? out_me_data_i_0__21_ : 
                              (N455)? out_me_data_i[53] : 
                              (N456)? out_me_data_i[85] : 
                              (N457)? out_me_data_i[117] : 
                              (N458)? out_me_data_i[149] : 
                              (N459)? out_me_data_i[181] : 
                              (N460)? out_me_data_i[213] : 
                              (N461)? out_me_data_i[245] : 
                              (N462)? out_me_data_i[277] : 
                              (N463)? out_me_data_i[309] : 
                              (N464)? out_me_data_i[341] : 
                              (N465)? out_me_data_i[373] : 
                              (N466)? out_me_data_i[405] : 
                              (N467)? out_me_data_i[437] : 
                              (N468)? out_me_data_i[469] : 1'b0;
  assign out_me_data_o[468] = (N454)? out_me_data_i_0__20_ : 
                              (N455)? out_me_data_i[52] : 
                              (N456)? out_me_data_i[84] : 
                              (N457)? out_me_data_i[116] : 
                              (N458)? out_me_data_i[148] : 
                              (N459)? out_me_data_i[180] : 
                              (N460)? out_me_data_i[212] : 
                              (N461)? out_me_data_i[244] : 
                              (N462)? out_me_data_i[276] : 
                              (N463)? out_me_data_i[308] : 
                              (N464)? out_me_data_i[340] : 
                              (N465)? out_me_data_i[372] : 
                              (N466)? out_me_data_i[404] : 
                              (N467)? out_me_data_i[436] : 
                              (N468)? out_me_data_i[468] : 1'b0;
  assign out_me_data_o[467] = (N454)? out_me_data_i_0__19_ : 
                              (N455)? out_me_data_i[51] : 
                              (N456)? out_me_data_i[83] : 
                              (N457)? out_me_data_i[115] : 
                              (N458)? out_me_data_i[147] : 
                              (N459)? out_me_data_i[179] : 
                              (N460)? out_me_data_i[211] : 
                              (N461)? out_me_data_i[243] : 
                              (N462)? out_me_data_i[275] : 
                              (N463)? out_me_data_i[307] : 
                              (N464)? out_me_data_i[339] : 
                              (N465)? out_me_data_i[371] : 
                              (N466)? out_me_data_i[403] : 
                              (N467)? out_me_data_i[435] : 
                              (N468)? out_me_data_i[467] : 1'b0;
  assign out_me_data_o[466] = (N454)? out_me_data_i_0__18_ : 
                              (N455)? out_me_data_i[50] : 
                              (N456)? out_me_data_i[82] : 
                              (N457)? out_me_data_i[114] : 
                              (N458)? out_me_data_i[146] : 
                              (N459)? out_me_data_i[178] : 
                              (N460)? out_me_data_i[210] : 
                              (N461)? out_me_data_i[242] : 
                              (N462)? out_me_data_i[274] : 
                              (N463)? out_me_data_i[306] : 
                              (N464)? out_me_data_i[338] : 
                              (N465)? out_me_data_i[370] : 
                              (N466)? out_me_data_i[402] : 
                              (N467)? out_me_data_i[434] : 
                              (N468)? out_me_data_i[466] : 1'b0;
  assign out_me_data_o[465] = (N454)? out_me_data_i_0__17_ : 
                              (N455)? out_me_data_i[49] : 
                              (N456)? out_me_data_i[81] : 
                              (N457)? out_me_data_i[113] : 
                              (N458)? out_me_data_i[145] : 
                              (N459)? out_me_data_i[177] : 
                              (N460)? out_me_data_i[209] : 
                              (N461)? out_me_data_i[241] : 
                              (N462)? out_me_data_i[273] : 
                              (N463)? out_me_data_i[305] : 
                              (N464)? out_me_data_i[337] : 
                              (N465)? out_me_data_i[369] : 
                              (N466)? out_me_data_i[401] : 
                              (N467)? out_me_data_i[433] : 
                              (N468)? out_me_data_i[465] : 1'b0;
  assign out_me_data_o[464] = (N454)? out_me_data_i_0__16_ : 
                              (N455)? out_me_data_i[48] : 
                              (N456)? out_me_data_i[80] : 
                              (N457)? out_me_data_i[112] : 
                              (N458)? out_me_data_i[144] : 
                              (N459)? out_me_data_i[176] : 
                              (N460)? out_me_data_i[208] : 
                              (N461)? out_me_data_i[240] : 
                              (N462)? out_me_data_i[272] : 
                              (N463)? out_me_data_i[304] : 
                              (N464)? out_me_data_i[336] : 
                              (N465)? out_me_data_i[368] : 
                              (N466)? out_me_data_i[400] : 
                              (N467)? out_me_data_i[432] : 
                              (N468)? out_me_data_i[464] : 1'b0;
  assign out_me_data_o[463] = (N454)? out_me_data_i_0__15_ : 
                              (N455)? out_me_data_i[47] : 
                              (N456)? out_me_data_i[79] : 
                              (N457)? out_me_data_i[111] : 
                              (N458)? out_me_data_i[143] : 
                              (N459)? out_me_data_i[175] : 
                              (N460)? out_me_data_i[207] : 
                              (N461)? out_me_data_i[239] : 
                              (N462)? out_me_data_i[271] : 
                              (N463)? out_me_data_i[303] : 
                              (N464)? out_me_data_i[335] : 
                              (N465)? out_me_data_i[367] : 
                              (N466)? out_me_data_i[399] : 
                              (N467)? out_me_data_i[431] : 
                              (N468)? out_me_data_i[463] : 1'b0;
  assign out_me_data_o[462] = (N454)? out_me_data_i_0__14_ : 
                              (N455)? out_me_data_i[46] : 
                              (N456)? out_me_data_i[78] : 
                              (N457)? out_me_data_i[110] : 
                              (N458)? out_me_data_i[142] : 
                              (N459)? out_me_data_i[174] : 
                              (N460)? out_me_data_i[206] : 
                              (N461)? out_me_data_i[238] : 
                              (N462)? out_me_data_i[270] : 
                              (N463)? out_me_data_i[302] : 
                              (N464)? out_me_data_i[334] : 
                              (N465)? out_me_data_i[366] : 
                              (N466)? out_me_data_i[398] : 
                              (N467)? out_me_data_i[430] : 
                              (N468)? out_me_data_i[462] : 1'b0;
  assign out_me_data_o[461] = (N454)? out_me_data_i_0__13_ : 
                              (N455)? out_me_data_i[45] : 
                              (N456)? out_me_data_i[77] : 
                              (N457)? out_me_data_i[109] : 
                              (N458)? out_me_data_i[141] : 
                              (N459)? out_me_data_i[173] : 
                              (N460)? out_me_data_i[205] : 
                              (N461)? out_me_data_i[237] : 
                              (N462)? out_me_data_i[269] : 
                              (N463)? out_me_data_i[301] : 
                              (N464)? out_me_data_i[333] : 
                              (N465)? out_me_data_i[365] : 
                              (N466)? out_me_data_i[397] : 
                              (N467)? out_me_data_i[429] : 
                              (N468)? out_me_data_i[461] : 1'b0;
  assign out_me_data_o[460] = (N454)? out_me_data_i_0__12_ : 
                              (N455)? out_me_data_i[44] : 
                              (N456)? out_me_data_i[76] : 
                              (N457)? out_me_data_i[108] : 
                              (N458)? out_me_data_i[140] : 
                              (N459)? out_me_data_i[172] : 
                              (N460)? out_me_data_i[204] : 
                              (N461)? out_me_data_i[236] : 
                              (N462)? out_me_data_i[268] : 
                              (N463)? out_me_data_i[300] : 
                              (N464)? out_me_data_i[332] : 
                              (N465)? out_me_data_i[364] : 
                              (N466)? out_me_data_i[396] : 
                              (N467)? out_me_data_i[428] : 
                              (N468)? out_me_data_i[460] : 1'b0;
  assign out_me_data_o[459] = (N454)? out_me_data_i_0__11_ : 
                              (N455)? out_me_data_i[43] : 
                              (N456)? out_me_data_i[75] : 
                              (N457)? out_me_data_i[107] : 
                              (N458)? out_me_data_i[139] : 
                              (N459)? out_me_data_i[171] : 
                              (N460)? out_me_data_i[203] : 
                              (N461)? out_me_data_i[235] : 
                              (N462)? out_me_data_i[267] : 
                              (N463)? out_me_data_i[299] : 
                              (N464)? out_me_data_i[331] : 
                              (N465)? out_me_data_i[363] : 
                              (N466)? out_me_data_i[395] : 
                              (N467)? out_me_data_i[427] : 
                              (N468)? out_me_data_i[459] : 1'b0;
  assign out_me_data_o[458] = (N454)? out_me_data_i_0__10_ : 
                              (N455)? out_me_data_i[42] : 
                              (N456)? out_me_data_i[74] : 
                              (N457)? out_me_data_i[106] : 
                              (N458)? out_me_data_i[138] : 
                              (N459)? out_me_data_i[170] : 
                              (N460)? out_me_data_i[202] : 
                              (N461)? out_me_data_i[234] : 
                              (N462)? out_me_data_i[266] : 
                              (N463)? out_me_data_i[298] : 
                              (N464)? out_me_data_i[330] : 
                              (N465)? out_me_data_i[362] : 
                              (N466)? out_me_data_i[394] : 
                              (N467)? out_me_data_i[426] : 
                              (N468)? out_me_data_i[458] : 1'b0;
  assign out_me_data_o[457] = (N454)? out_me_data_i_0__9_ : 
                              (N455)? out_me_data_i[41] : 
                              (N456)? out_me_data_i[73] : 
                              (N457)? out_me_data_i[105] : 
                              (N458)? out_me_data_i[137] : 
                              (N459)? out_me_data_i[169] : 
                              (N460)? out_me_data_i[201] : 
                              (N461)? out_me_data_i[233] : 
                              (N462)? out_me_data_i[265] : 
                              (N463)? out_me_data_i[297] : 
                              (N464)? out_me_data_i[329] : 
                              (N465)? out_me_data_i[361] : 
                              (N466)? out_me_data_i[393] : 
                              (N467)? out_me_data_i[425] : 
                              (N468)? out_me_data_i[457] : 1'b0;
  assign out_me_data_o[456] = (N454)? out_me_data_i_0__8_ : 
                              (N455)? out_me_data_i[40] : 
                              (N456)? out_me_data_i[72] : 
                              (N457)? out_me_data_i[104] : 
                              (N458)? out_me_data_i[136] : 
                              (N459)? out_me_data_i[168] : 
                              (N460)? out_me_data_i[200] : 
                              (N461)? out_me_data_i[232] : 
                              (N462)? out_me_data_i[264] : 
                              (N463)? out_me_data_i[296] : 
                              (N464)? out_me_data_i[328] : 
                              (N465)? out_me_data_i[360] : 
                              (N466)? out_me_data_i[392] : 
                              (N467)? out_me_data_i[424] : 
                              (N468)? out_me_data_i[456] : 1'b0;
  assign out_me_data_o[455] = (N454)? out_me_data_i_0__7_ : 
                              (N455)? out_me_data_i[39] : 
                              (N456)? out_me_data_i[71] : 
                              (N457)? out_me_data_i[103] : 
                              (N458)? out_me_data_i[135] : 
                              (N459)? out_me_data_i[167] : 
                              (N460)? out_me_data_i[199] : 
                              (N461)? out_me_data_i[231] : 
                              (N462)? out_me_data_i[263] : 
                              (N463)? out_me_data_i[295] : 
                              (N464)? out_me_data_i[327] : 
                              (N465)? out_me_data_i[359] : 
                              (N466)? out_me_data_i[391] : 
                              (N467)? out_me_data_i[423] : 
                              (N468)? out_me_data_i[455] : 1'b0;
  assign out_me_data_o[454] = (N454)? out_me_data_i_0__6_ : 
                              (N455)? out_me_data_i[38] : 
                              (N456)? out_me_data_i[70] : 
                              (N457)? out_me_data_i[102] : 
                              (N458)? out_me_data_i[134] : 
                              (N459)? out_me_data_i[166] : 
                              (N460)? out_me_data_i[198] : 
                              (N461)? out_me_data_i[230] : 
                              (N462)? out_me_data_i[262] : 
                              (N463)? out_me_data_i[294] : 
                              (N464)? out_me_data_i[326] : 
                              (N465)? out_me_data_i[358] : 
                              (N466)? out_me_data_i[390] : 
                              (N467)? out_me_data_i[422] : 
                              (N468)? out_me_data_i[454] : 1'b0;
  assign out_me_data_o[453] = (N454)? out_me_data_i_0__5_ : 
                              (N455)? out_me_data_i[37] : 
                              (N456)? out_me_data_i[69] : 
                              (N457)? out_me_data_i[101] : 
                              (N458)? out_me_data_i[133] : 
                              (N459)? out_me_data_i[165] : 
                              (N460)? out_me_data_i[197] : 
                              (N461)? out_me_data_i[229] : 
                              (N462)? out_me_data_i[261] : 
                              (N463)? out_me_data_i[293] : 
                              (N464)? out_me_data_i[325] : 
                              (N465)? out_me_data_i[357] : 
                              (N466)? out_me_data_i[389] : 
                              (N467)? out_me_data_i[421] : 
                              (N468)? out_me_data_i[453] : 1'b0;
  assign out_me_data_o[452] = (N454)? out_me_data_i_0__4_ : 
                              (N455)? out_me_data_i[36] : 
                              (N456)? out_me_data_i[68] : 
                              (N457)? out_me_data_i[100] : 
                              (N458)? out_me_data_i[132] : 
                              (N459)? out_me_data_i[164] : 
                              (N460)? out_me_data_i[196] : 
                              (N461)? out_me_data_i[228] : 
                              (N462)? out_me_data_i[260] : 
                              (N463)? out_me_data_i[292] : 
                              (N464)? out_me_data_i[324] : 
                              (N465)? out_me_data_i[356] : 
                              (N466)? out_me_data_i[388] : 
                              (N467)? out_me_data_i[420] : 
                              (N468)? out_me_data_i[452] : 1'b0;
  assign out_me_data_o[451] = (N454)? out_me_data_i_0__3_ : 
                              (N455)? out_me_data_i[35] : 
                              (N456)? out_me_data_i[67] : 
                              (N457)? out_me_data_i[99] : 
                              (N458)? out_me_data_i[131] : 
                              (N459)? out_me_data_i[163] : 
                              (N460)? out_me_data_i[195] : 
                              (N461)? out_me_data_i[227] : 
                              (N462)? out_me_data_i[259] : 
                              (N463)? out_me_data_i[291] : 
                              (N464)? out_me_data_i[323] : 
                              (N465)? out_me_data_i[355] : 
                              (N466)? out_me_data_i[387] : 
                              (N467)? out_me_data_i[419] : 
                              (N468)? out_me_data_i[451] : 1'b0;
  assign out_me_data_o[450] = (N454)? out_me_data_i_0__2_ : 
                              (N455)? out_me_data_i[34] : 
                              (N456)? out_me_data_i[66] : 
                              (N457)? out_me_data_i[98] : 
                              (N458)? out_me_data_i[130] : 
                              (N459)? out_me_data_i[162] : 
                              (N460)? out_me_data_i[194] : 
                              (N461)? out_me_data_i[226] : 
                              (N462)? out_me_data_i[258] : 
                              (N463)? out_me_data_i[290] : 
                              (N464)? out_me_data_i[322] : 
                              (N465)? out_me_data_i[354] : 
                              (N466)? out_me_data_i[386] : 
                              (N467)? out_me_data_i[418] : 
                              (N468)? out_me_data_i[450] : 1'b0;
  assign out_me_data_o[449] = (N454)? out_me_data_i_0__1_ : 
                              (N455)? out_me_data_i[33] : 
                              (N456)? out_me_data_i[65] : 
                              (N457)? out_me_data_i[97] : 
                              (N458)? out_me_data_i[129] : 
                              (N459)? out_me_data_i[161] : 
                              (N460)? out_me_data_i[193] : 
                              (N461)? out_me_data_i[225] : 
                              (N462)? out_me_data_i[257] : 
                              (N463)? out_me_data_i[289] : 
                              (N464)? out_me_data_i[321] : 
                              (N465)? out_me_data_i[353] : 
                              (N466)? out_me_data_i[385] : 
                              (N467)? out_me_data_i[417] : 
                              (N468)? out_me_data_i[449] : 1'b0;
  assign out_me_data_o[448] = (N454)? out_me_data_i_0__0_ : 
                              (N455)? out_me_data_i[32] : 
                              (N456)? out_me_data_i[64] : 
                              (N457)? out_me_data_i[96] : 
                              (N458)? out_me_data_i[128] : 
                              (N459)? out_me_data_i[160] : 
                              (N460)? out_me_data_i[192] : 
                              (N461)? out_me_data_i[224] : 
                              (N462)? out_me_data_i[256] : 
                              (N463)? out_me_data_i[288] : 
                              (N464)? out_me_data_i[320] : 
                              (N465)? out_me_data_i[352] : 
                              (N466)? out_me_data_i[384] : 
                              (N467)? out_me_data_i[416] : 
                              (N468)? out_me_data_i[448] : 1'b0;
  assign out_me_data_o[447] = (N469)? out_me_data_i_0__31_ : 
                              (N470)? out_me_data_i[63] : 
                              (N471)? out_me_data_i[95] : 
                              (N472)? out_me_data_i[127] : 
                              (N473)? out_me_data_i[159] : 
                              (N474)? out_me_data_i[191] : 
                              (N475)? out_me_data_i[223] : 
                              (N476)? out_me_data_i[255] : 
                              (N477)? out_me_data_i[287] : 
                              (N478)? out_me_data_i[319] : 
                              (N479)? out_me_data_i[351] : 
                              (N480)? out_me_data_i[383] : 
                              (N481)? out_me_data_i[415] : 
                              (N482)? out_me_data_i[447] : 1'b0;
  assign N469 = N2298;
  assign N470 = N2300;
  assign N471 = N2302;
  assign N472 = N2304;
  assign N473 = N2306;
  assign N474 = N2308;
  assign N475 = N2310;
  assign N476 = N2311;
  assign N477 = N2299;
  assign N478 = N2301;
  assign N479 = N2303;
  assign N480 = N2305;
  assign N481 = N2307;
  assign N482 = N2309;
  assign out_me_data_o[446] = (N469)? out_me_data_i_0__30_ : 
                              (N470)? out_me_data_i[62] : 
                              (N471)? out_me_data_i[94] : 
                              (N472)? out_me_data_i[126] : 
                              (N473)? out_me_data_i[158] : 
                              (N474)? out_me_data_i[190] : 
                              (N475)? out_me_data_i[222] : 
                              (N476)? out_me_data_i[254] : 
                              (N477)? out_me_data_i[286] : 
                              (N478)? out_me_data_i[318] : 
                              (N479)? out_me_data_i[350] : 
                              (N480)? out_me_data_i[382] : 
                              (N481)? out_me_data_i[414] : 
                              (N482)? out_me_data_i[446] : 1'b0;
  assign out_me_data_o[445] = (N469)? out_me_data_i_0__29_ : 
                              (N470)? out_me_data_i[61] : 
                              (N471)? out_me_data_i[93] : 
                              (N472)? out_me_data_i[125] : 
                              (N473)? out_me_data_i[157] : 
                              (N474)? out_me_data_i[189] : 
                              (N475)? out_me_data_i[221] : 
                              (N476)? out_me_data_i[253] : 
                              (N477)? out_me_data_i[285] : 
                              (N478)? out_me_data_i[317] : 
                              (N479)? out_me_data_i[349] : 
                              (N480)? out_me_data_i[381] : 
                              (N481)? out_me_data_i[413] : 
                              (N482)? out_me_data_i[445] : 1'b0;
  assign out_me_data_o[444] = (N469)? out_me_data_i_0__28_ : 
                              (N470)? out_me_data_i[60] : 
                              (N471)? out_me_data_i[92] : 
                              (N472)? out_me_data_i[124] : 
                              (N473)? out_me_data_i[156] : 
                              (N474)? out_me_data_i[188] : 
                              (N475)? out_me_data_i[220] : 
                              (N476)? out_me_data_i[252] : 
                              (N477)? out_me_data_i[284] : 
                              (N478)? out_me_data_i[316] : 
                              (N479)? out_me_data_i[348] : 
                              (N480)? out_me_data_i[380] : 
                              (N481)? out_me_data_i[412] : 
                              (N482)? out_me_data_i[444] : 1'b0;
  assign out_me_data_o[443] = (N469)? out_me_data_i_0__27_ : 
                              (N470)? out_me_data_i[59] : 
                              (N471)? out_me_data_i[91] : 
                              (N472)? out_me_data_i[123] : 
                              (N473)? out_me_data_i[155] : 
                              (N474)? out_me_data_i[187] : 
                              (N475)? out_me_data_i[219] : 
                              (N476)? out_me_data_i[251] : 
                              (N477)? out_me_data_i[283] : 
                              (N478)? out_me_data_i[315] : 
                              (N479)? out_me_data_i[347] : 
                              (N480)? out_me_data_i[379] : 
                              (N481)? out_me_data_i[411] : 
                              (N482)? out_me_data_i[443] : 1'b0;
  assign out_me_data_o[442] = (N469)? out_me_data_i_0__26_ : 
                              (N470)? out_me_data_i[58] : 
                              (N471)? out_me_data_i[90] : 
                              (N472)? out_me_data_i[122] : 
                              (N473)? out_me_data_i[154] : 
                              (N474)? out_me_data_i[186] : 
                              (N475)? out_me_data_i[218] : 
                              (N476)? out_me_data_i[250] : 
                              (N477)? out_me_data_i[282] : 
                              (N478)? out_me_data_i[314] : 
                              (N479)? out_me_data_i[346] : 
                              (N480)? out_me_data_i[378] : 
                              (N481)? out_me_data_i[410] : 
                              (N482)? out_me_data_i[442] : 1'b0;
  assign out_me_data_o[441] = (N469)? out_me_data_i_0__25_ : 
                              (N470)? out_me_data_i[57] : 
                              (N471)? out_me_data_i[89] : 
                              (N472)? out_me_data_i[121] : 
                              (N473)? out_me_data_i[153] : 
                              (N474)? out_me_data_i[185] : 
                              (N475)? out_me_data_i[217] : 
                              (N476)? out_me_data_i[249] : 
                              (N477)? out_me_data_i[281] : 
                              (N478)? out_me_data_i[313] : 
                              (N479)? out_me_data_i[345] : 
                              (N480)? out_me_data_i[377] : 
                              (N481)? out_me_data_i[409] : 
                              (N482)? out_me_data_i[441] : 1'b0;
  assign out_me_data_o[440] = (N469)? out_me_data_i_0__24_ : 
                              (N470)? out_me_data_i[56] : 
                              (N471)? out_me_data_i[88] : 
                              (N472)? out_me_data_i[120] : 
                              (N473)? out_me_data_i[152] : 
                              (N474)? out_me_data_i[184] : 
                              (N475)? out_me_data_i[216] : 
                              (N476)? out_me_data_i[248] : 
                              (N477)? out_me_data_i[280] : 
                              (N478)? out_me_data_i[312] : 
                              (N479)? out_me_data_i[344] : 
                              (N480)? out_me_data_i[376] : 
                              (N481)? out_me_data_i[408] : 
                              (N482)? out_me_data_i[440] : 1'b0;
  assign out_me_data_o[439] = (N469)? out_me_data_i_0__23_ : 
                              (N470)? out_me_data_i[55] : 
                              (N471)? out_me_data_i[87] : 
                              (N472)? out_me_data_i[119] : 
                              (N473)? out_me_data_i[151] : 
                              (N474)? out_me_data_i[183] : 
                              (N475)? out_me_data_i[215] : 
                              (N476)? out_me_data_i[247] : 
                              (N477)? out_me_data_i[279] : 
                              (N478)? out_me_data_i[311] : 
                              (N479)? out_me_data_i[343] : 
                              (N480)? out_me_data_i[375] : 
                              (N481)? out_me_data_i[407] : 
                              (N482)? out_me_data_i[439] : 1'b0;
  assign out_me_data_o[438] = (N469)? out_me_data_i_0__22_ : 
                              (N470)? out_me_data_i[54] : 
                              (N471)? out_me_data_i[86] : 
                              (N472)? out_me_data_i[118] : 
                              (N473)? out_me_data_i[150] : 
                              (N474)? out_me_data_i[182] : 
                              (N475)? out_me_data_i[214] : 
                              (N476)? out_me_data_i[246] : 
                              (N477)? out_me_data_i[278] : 
                              (N478)? out_me_data_i[310] : 
                              (N479)? out_me_data_i[342] : 
                              (N480)? out_me_data_i[374] : 
                              (N481)? out_me_data_i[406] : 
                              (N482)? out_me_data_i[438] : 1'b0;
  assign out_me_data_o[437] = (N469)? out_me_data_i_0__21_ : 
                              (N470)? out_me_data_i[53] : 
                              (N471)? out_me_data_i[85] : 
                              (N472)? out_me_data_i[117] : 
                              (N473)? out_me_data_i[149] : 
                              (N474)? out_me_data_i[181] : 
                              (N475)? out_me_data_i[213] : 
                              (N476)? out_me_data_i[245] : 
                              (N477)? out_me_data_i[277] : 
                              (N478)? out_me_data_i[309] : 
                              (N479)? out_me_data_i[341] : 
                              (N480)? out_me_data_i[373] : 
                              (N481)? out_me_data_i[405] : 
                              (N482)? out_me_data_i[437] : 1'b0;
  assign out_me_data_o[436] = (N469)? out_me_data_i_0__20_ : 
                              (N470)? out_me_data_i[52] : 
                              (N471)? out_me_data_i[84] : 
                              (N472)? out_me_data_i[116] : 
                              (N473)? out_me_data_i[148] : 
                              (N474)? out_me_data_i[180] : 
                              (N475)? out_me_data_i[212] : 
                              (N476)? out_me_data_i[244] : 
                              (N477)? out_me_data_i[276] : 
                              (N478)? out_me_data_i[308] : 
                              (N479)? out_me_data_i[340] : 
                              (N480)? out_me_data_i[372] : 
                              (N481)? out_me_data_i[404] : 
                              (N482)? out_me_data_i[436] : 1'b0;
  assign out_me_data_o[435] = (N469)? out_me_data_i_0__19_ : 
                              (N470)? out_me_data_i[51] : 
                              (N471)? out_me_data_i[83] : 
                              (N472)? out_me_data_i[115] : 
                              (N473)? out_me_data_i[147] : 
                              (N474)? out_me_data_i[179] : 
                              (N475)? out_me_data_i[211] : 
                              (N476)? out_me_data_i[243] : 
                              (N477)? out_me_data_i[275] : 
                              (N478)? out_me_data_i[307] : 
                              (N479)? out_me_data_i[339] : 
                              (N480)? out_me_data_i[371] : 
                              (N481)? out_me_data_i[403] : 
                              (N482)? out_me_data_i[435] : 1'b0;
  assign out_me_data_o[434] = (N469)? out_me_data_i_0__18_ : 
                              (N470)? out_me_data_i[50] : 
                              (N471)? out_me_data_i[82] : 
                              (N472)? out_me_data_i[114] : 
                              (N473)? out_me_data_i[146] : 
                              (N474)? out_me_data_i[178] : 
                              (N475)? out_me_data_i[210] : 
                              (N476)? out_me_data_i[242] : 
                              (N477)? out_me_data_i[274] : 
                              (N478)? out_me_data_i[306] : 
                              (N479)? out_me_data_i[338] : 
                              (N480)? out_me_data_i[370] : 
                              (N481)? out_me_data_i[402] : 
                              (N482)? out_me_data_i[434] : 1'b0;
  assign out_me_data_o[433] = (N469)? out_me_data_i_0__17_ : 
                              (N470)? out_me_data_i[49] : 
                              (N471)? out_me_data_i[81] : 
                              (N472)? out_me_data_i[113] : 
                              (N473)? out_me_data_i[145] : 
                              (N474)? out_me_data_i[177] : 
                              (N475)? out_me_data_i[209] : 
                              (N476)? out_me_data_i[241] : 
                              (N477)? out_me_data_i[273] : 
                              (N478)? out_me_data_i[305] : 
                              (N479)? out_me_data_i[337] : 
                              (N480)? out_me_data_i[369] : 
                              (N481)? out_me_data_i[401] : 
                              (N482)? out_me_data_i[433] : 1'b0;
  assign out_me_data_o[432] = (N469)? out_me_data_i_0__16_ : 
                              (N470)? out_me_data_i[48] : 
                              (N471)? out_me_data_i[80] : 
                              (N472)? out_me_data_i[112] : 
                              (N473)? out_me_data_i[144] : 
                              (N474)? out_me_data_i[176] : 
                              (N475)? out_me_data_i[208] : 
                              (N476)? out_me_data_i[240] : 
                              (N477)? out_me_data_i[272] : 
                              (N478)? out_me_data_i[304] : 
                              (N479)? out_me_data_i[336] : 
                              (N480)? out_me_data_i[368] : 
                              (N481)? out_me_data_i[400] : 
                              (N482)? out_me_data_i[432] : 1'b0;
  assign out_me_data_o[431] = (N469)? out_me_data_i_0__15_ : 
                              (N470)? out_me_data_i[47] : 
                              (N471)? out_me_data_i[79] : 
                              (N472)? out_me_data_i[111] : 
                              (N473)? out_me_data_i[143] : 
                              (N474)? out_me_data_i[175] : 
                              (N475)? out_me_data_i[207] : 
                              (N476)? out_me_data_i[239] : 
                              (N477)? out_me_data_i[271] : 
                              (N478)? out_me_data_i[303] : 
                              (N479)? out_me_data_i[335] : 
                              (N480)? out_me_data_i[367] : 
                              (N481)? out_me_data_i[399] : 
                              (N482)? out_me_data_i[431] : 1'b0;
  assign out_me_data_o[430] = (N469)? out_me_data_i_0__14_ : 
                              (N470)? out_me_data_i[46] : 
                              (N471)? out_me_data_i[78] : 
                              (N472)? out_me_data_i[110] : 
                              (N473)? out_me_data_i[142] : 
                              (N474)? out_me_data_i[174] : 
                              (N475)? out_me_data_i[206] : 
                              (N476)? out_me_data_i[238] : 
                              (N477)? out_me_data_i[270] : 
                              (N478)? out_me_data_i[302] : 
                              (N479)? out_me_data_i[334] : 
                              (N480)? out_me_data_i[366] : 
                              (N481)? out_me_data_i[398] : 
                              (N482)? out_me_data_i[430] : 1'b0;
  assign out_me_data_o[429] = (N469)? out_me_data_i_0__13_ : 
                              (N470)? out_me_data_i[45] : 
                              (N471)? out_me_data_i[77] : 
                              (N472)? out_me_data_i[109] : 
                              (N473)? out_me_data_i[141] : 
                              (N474)? out_me_data_i[173] : 
                              (N475)? out_me_data_i[205] : 
                              (N476)? out_me_data_i[237] : 
                              (N477)? out_me_data_i[269] : 
                              (N478)? out_me_data_i[301] : 
                              (N479)? out_me_data_i[333] : 
                              (N480)? out_me_data_i[365] : 
                              (N481)? out_me_data_i[397] : 
                              (N482)? out_me_data_i[429] : 1'b0;
  assign out_me_data_o[428] = (N469)? out_me_data_i_0__12_ : 
                              (N470)? out_me_data_i[44] : 
                              (N471)? out_me_data_i[76] : 
                              (N472)? out_me_data_i[108] : 
                              (N473)? out_me_data_i[140] : 
                              (N474)? out_me_data_i[172] : 
                              (N475)? out_me_data_i[204] : 
                              (N476)? out_me_data_i[236] : 
                              (N477)? out_me_data_i[268] : 
                              (N478)? out_me_data_i[300] : 
                              (N479)? out_me_data_i[332] : 
                              (N480)? out_me_data_i[364] : 
                              (N481)? out_me_data_i[396] : 
                              (N482)? out_me_data_i[428] : 1'b0;
  assign out_me_data_o[427] = (N469)? out_me_data_i_0__11_ : 
                              (N470)? out_me_data_i[43] : 
                              (N471)? out_me_data_i[75] : 
                              (N472)? out_me_data_i[107] : 
                              (N473)? out_me_data_i[139] : 
                              (N474)? out_me_data_i[171] : 
                              (N475)? out_me_data_i[203] : 
                              (N476)? out_me_data_i[235] : 
                              (N477)? out_me_data_i[267] : 
                              (N478)? out_me_data_i[299] : 
                              (N479)? out_me_data_i[331] : 
                              (N480)? out_me_data_i[363] : 
                              (N481)? out_me_data_i[395] : 
                              (N482)? out_me_data_i[427] : 1'b0;
  assign out_me_data_o[426] = (N469)? out_me_data_i_0__10_ : 
                              (N470)? out_me_data_i[42] : 
                              (N471)? out_me_data_i[74] : 
                              (N472)? out_me_data_i[106] : 
                              (N473)? out_me_data_i[138] : 
                              (N474)? out_me_data_i[170] : 
                              (N475)? out_me_data_i[202] : 
                              (N476)? out_me_data_i[234] : 
                              (N477)? out_me_data_i[266] : 
                              (N478)? out_me_data_i[298] : 
                              (N479)? out_me_data_i[330] : 
                              (N480)? out_me_data_i[362] : 
                              (N481)? out_me_data_i[394] : 
                              (N482)? out_me_data_i[426] : 1'b0;
  assign out_me_data_o[425] = (N469)? out_me_data_i_0__9_ : 
                              (N470)? out_me_data_i[41] : 
                              (N471)? out_me_data_i[73] : 
                              (N472)? out_me_data_i[105] : 
                              (N473)? out_me_data_i[137] : 
                              (N474)? out_me_data_i[169] : 
                              (N475)? out_me_data_i[201] : 
                              (N476)? out_me_data_i[233] : 
                              (N477)? out_me_data_i[265] : 
                              (N478)? out_me_data_i[297] : 
                              (N479)? out_me_data_i[329] : 
                              (N480)? out_me_data_i[361] : 
                              (N481)? out_me_data_i[393] : 
                              (N482)? out_me_data_i[425] : 1'b0;
  assign out_me_data_o[424] = (N469)? out_me_data_i_0__8_ : 
                              (N470)? out_me_data_i[40] : 
                              (N471)? out_me_data_i[72] : 
                              (N472)? out_me_data_i[104] : 
                              (N473)? out_me_data_i[136] : 
                              (N474)? out_me_data_i[168] : 
                              (N475)? out_me_data_i[200] : 
                              (N476)? out_me_data_i[232] : 
                              (N477)? out_me_data_i[264] : 
                              (N478)? out_me_data_i[296] : 
                              (N479)? out_me_data_i[328] : 
                              (N480)? out_me_data_i[360] : 
                              (N481)? out_me_data_i[392] : 
                              (N482)? out_me_data_i[424] : 1'b0;
  assign out_me_data_o[423] = (N469)? out_me_data_i_0__7_ : 
                              (N470)? out_me_data_i[39] : 
                              (N471)? out_me_data_i[71] : 
                              (N472)? out_me_data_i[103] : 
                              (N473)? out_me_data_i[135] : 
                              (N474)? out_me_data_i[167] : 
                              (N475)? out_me_data_i[199] : 
                              (N476)? out_me_data_i[231] : 
                              (N477)? out_me_data_i[263] : 
                              (N478)? out_me_data_i[295] : 
                              (N479)? out_me_data_i[327] : 
                              (N480)? out_me_data_i[359] : 
                              (N481)? out_me_data_i[391] : 
                              (N482)? out_me_data_i[423] : 1'b0;
  assign out_me_data_o[422] = (N469)? out_me_data_i_0__6_ : 
                              (N470)? out_me_data_i[38] : 
                              (N471)? out_me_data_i[70] : 
                              (N472)? out_me_data_i[102] : 
                              (N473)? out_me_data_i[134] : 
                              (N474)? out_me_data_i[166] : 
                              (N475)? out_me_data_i[198] : 
                              (N476)? out_me_data_i[230] : 
                              (N477)? out_me_data_i[262] : 
                              (N478)? out_me_data_i[294] : 
                              (N479)? out_me_data_i[326] : 
                              (N480)? out_me_data_i[358] : 
                              (N481)? out_me_data_i[390] : 
                              (N482)? out_me_data_i[422] : 1'b0;
  assign out_me_data_o[421] = (N469)? out_me_data_i_0__5_ : 
                              (N470)? out_me_data_i[37] : 
                              (N471)? out_me_data_i[69] : 
                              (N472)? out_me_data_i[101] : 
                              (N473)? out_me_data_i[133] : 
                              (N474)? out_me_data_i[165] : 
                              (N475)? out_me_data_i[197] : 
                              (N476)? out_me_data_i[229] : 
                              (N477)? out_me_data_i[261] : 
                              (N478)? out_me_data_i[293] : 
                              (N479)? out_me_data_i[325] : 
                              (N480)? out_me_data_i[357] : 
                              (N481)? out_me_data_i[389] : 
                              (N482)? out_me_data_i[421] : 1'b0;
  assign out_me_data_o[420] = (N469)? out_me_data_i_0__4_ : 
                              (N470)? out_me_data_i[36] : 
                              (N471)? out_me_data_i[68] : 
                              (N472)? out_me_data_i[100] : 
                              (N473)? out_me_data_i[132] : 
                              (N474)? out_me_data_i[164] : 
                              (N475)? out_me_data_i[196] : 
                              (N476)? out_me_data_i[228] : 
                              (N477)? out_me_data_i[260] : 
                              (N478)? out_me_data_i[292] : 
                              (N479)? out_me_data_i[324] : 
                              (N480)? out_me_data_i[356] : 
                              (N481)? out_me_data_i[388] : 
                              (N482)? out_me_data_i[420] : 1'b0;
  assign out_me_data_o[419] = (N469)? out_me_data_i_0__3_ : 
                              (N470)? out_me_data_i[35] : 
                              (N471)? out_me_data_i[67] : 
                              (N472)? out_me_data_i[99] : 
                              (N473)? out_me_data_i[131] : 
                              (N474)? out_me_data_i[163] : 
                              (N475)? out_me_data_i[195] : 
                              (N476)? out_me_data_i[227] : 
                              (N477)? out_me_data_i[259] : 
                              (N478)? out_me_data_i[291] : 
                              (N479)? out_me_data_i[323] : 
                              (N480)? out_me_data_i[355] : 
                              (N481)? out_me_data_i[387] : 
                              (N482)? out_me_data_i[419] : 1'b0;
  assign out_me_data_o[418] = (N469)? out_me_data_i_0__2_ : 
                              (N470)? out_me_data_i[34] : 
                              (N471)? out_me_data_i[66] : 
                              (N472)? out_me_data_i[98] : 
                              (N473)? out_me_data_i[130] : 
                              (N474)? out_me_data_i[162] : 
                              (N475)? out_me_data_i[194] : 
                              (N476)? out_me_data_i[226] : 
                              (N477)? out_me_data_i[258] : 
                              (N478)? out_me_data_i[290] : 
                              (N479)? out_me_data_i[322] : 
                              (N480)? out_me_data_i[354] : 
                              (N481)? out_me_data_i[386] : 
                              (N482)? out_me_data_i[418] : 1'b0;
  assign out_me_data_o[417] = (N469)? out_me_data_i_0__1_ : 
                              (N470)? out_me_data_i[33] : 
                              (N471)? out_me_data_i[65] : 
                              (N472)? out_me_data_i[97] : 
                              (N473)? out_me_data_i[129] : 
                              (N474)? out_me_data_i[161] : 
                              (N475)? out_me_data_i[193] : 
                              (N476)? out_me_data_i[225] : 
                              (N477)? out_me_data_i[257] : 
                              (N478)? out_me_data_i[289] : 
                              (N479)? out_me_data_i[321] : 
                              (N480)? out_me_data_i[353] : 
                              (N481)? out_me_data_i[385] : 
                              (N482)? out_me_data_i[417] : 1'b0;
  assign out_me_data_o[416] = (N469)? out_me_data_i_0__0_ : 
                              (N470)? out_me_data_i[32] : 
                              (N471)? out_me_data_i[64] : 
                              (N472)? out_me_data_i[96] : 
                              (N473)? out_me_data_i[128] : 
                              (N474)? out_me_data_i[160] : 
                              (N475)? out_me_data_i[192] : 
                              (N476)? out_me_data_i[224] : 
                              (N477)? out_me_data_i[256] : 
                              (N478)? out_me_data_i[288] : 
                              (N479)? out_me_data_i[320] : 
                              (N480)? out_me_data_i[352] : 
                              (N481)? out_me_data_i[384] : 
                              (N482)? out_me_data_i[416] : 1'b0;
  assign out_me_data_o[415] = (N483)? out_me_data_i_0__31_ : 
                              (N484)? out_me_data_i[63] : 
                              (N485)? out_me_data_i[95] : 
                              (N486)? out_me_data_i[127] : 
                              (N487)? out_me_data_i[159] : 
                              (N488)? out_me_data_i[191] : 
                              (N489)? out_me_data_i[223] : 
                              (N490)? out_me_data_i[255] : 
                              (N491)? out_me_data_i[287] : 
                              (N492)? out_me_data_i[319] : 
                              (N493)? out_me_data_i[351] : 
                              (N494)? out_me_data_i[383] : 
                              (N495)? out_me_data_i[415] : 1'b0;
  assign N483 = N2176;
  assign N484 = N2178;
  assign N485 = N2180;
  assign N486 = N2182;
  assign N487 = N2184;
  assign N488 = N2186;
  assign N489 = N2187;
  assign N490 = N2188;
  assign N491 = N2177;
  assign N492 = N2179;
  assign N493 = N2181;
  assign N494 = N2183;
  assign N495 = N2185;
  assign out_me_data_o[414] = (N483)? out_me_data_i_0__30_ : 
                              (N484)? out_me_data_i[62] : 
                              (N485)? out_me_data_i[94] : 
                              (N486)? out_me_data_i[126] : 
                              (N487)? out_me_data_i[158] : 
                              (N488)? out_me_data_i[190] : 
                              (N489)? out_me_data_i[222] : 
                              (N490)? out_me_data_i[254] : 
                              (N491)? out_me_data_i[286] : 
                              (N492)? out_me_data_i[318] : 
                              (N493)? out_me_data_i[350] : 
                              (N494)? out_me_data_i[382] : 
                              (N495)? out_me_data_i[414] : 1'b0;
  assign out_me_data_o[413] = (N483)? out_me_data_i_0__29_ : 
                              (N484)? out_me_data_i[61] : 
                              (N485)? out_me_data_i[93] : 
                              (N486)? out_me_data_i[125] : 
                              (N487)? out_me_data_i[157] : 
                              (N488)? out_me_data_i[189] : 
                              (N489)? out_me_data_i[221] : 
                              (N490)? out_me_data_i[253] : 
                              (N491)? out_me_data_i[285] : 
                              (N492)? out_me_data_i[317] : 
                              (N493)? out_me_data_i[349] : 
                              (N494)? out_me_data_i[381] : 
                              (N495)? out_me_data_i[413] : 1'b0;
  assign out_me_data_o[412] = (N483)? out_me_data_i_0__28_ : 
                              (N484)? out_me_data_i[60] : 
                              (N485)? out_me_data_i[92] : 
                              (N486)? out_me_data_i[124] : 
                              (N487)? out_me_data_i[156] : 
                              (N488)? out_me_data_i[188] : 
                              (N489)? out_me_data_i[220] : 
                              (N490)? out_me_data_i[252] : 
                              (N491)? out_me_data_i[284] : 
                              (N492)? out_me_data_i[316] : 
                              (N493)? out_me_data_i[348] : 
                              (N494)? out_me_data_i[380] : 
                              (N495)? out_me_data_i[412] : 1'b0;
  assign out_me_data_o[411] = (N483)? out_me_data_i_0__27_ : 
                              (N484)? out_me_data_i[59] : 
                              (N485)? out_me_data_i[91] : 
                              (N486)? out_me_data_i[123] : 
                              (N487)? out_me_data_i[155] : 
                              (N488)? out_me_data_i[187] : 
                              (N489)? out_me_data_i[219] : 
                              (N490)? out_me_data_i[251] : 
                              (N491)? out_me_data_i[283] : 
                              (N492)? out_me_data_i[315] : 
                              (N493)? out_me_data_i[347] : 
                              (N494)? out_me_data_i[379] : 
                              (N495)? out_me_data_i[411] : 1'b0;
  assign out_me_data_o[410] = (N483)? out_me_data_i_0__26_ : 
                              (N484)? out_me_data_i[58] : 
                              (N485)? out_me_data_i[90] : 
                              (N486)? out_me_data_i[122] : 
                              (N487)? out_me_data_i[154] : 
                              (N488)? out_me_data_i[186] : 
                              (N489)? out_me_data_i[218] : 
                              (N490)? out_me_data_i[250] : 
                              (N491)? out_me_data_i[282] : 
                              (N492)? out_me_data_i[314] : 
                              (N493)? out_me_data_i[346] : 
                              (N494)? out_me_data_i[378] : 
                              (N495)? out_me_data_i[410] : 1'b0;
  assign out_me_data_o[409] = (N483)? out_me_data_i_0__25_ : 
                              (N484)? out_me_data_i[57] : 
                              (N485)? out_me_data_i[89] : 
                              (N486)? out_me_data_i[121] : 
                              (N487)? out_me_data_i[153] : 
                              (N488)? out_me_data_i[185] : 
                              (N489)? out_me_data_i[217] : 
                              (N490)? out_me_data_i[249] : 
                              (N491)? out_me_data_i[281] : 
                              (N492)? out_me_data_i[313] : 
                              (N493)? out_me_data_i[345] : 
                              (N494)? out_me_data_i[377] : 
                              (N495)? out_me_data_i[409] : 1'b0;
  assign out_me_data_o[408] = (N483)? out_me_data_i_0__24_ : 
                              (N484)? out_me_data_i[56] : 
                              (N485)? out_me_data_i[88] : 
                              (N486)? out_me_data_i[120] : 
                              (N487)? out_me_data_i[152] : 
                              (N488)? out_me_data_i[184] : 
                              (N489)? out_me_data_i[216] : 
                              (N490)? out_me_data_i[248] : 
                              (N491)? out_me_data_i[280] : 
                              (N492)? out_me_data_i[312] : 
                              (N493)? out_me_data_i[344] : 
                              (N494)? out_me_data_i[376] : 
                              (N495)? out_me_data_i[408] : 1'b0;
  assign out_me_data_o[407] = (N483)? out_me_data_i_0__23_ : 
                              (N484)? out_me_data_i[55] : 
                              (N485)? out_me_data_i[87] : 
                              (N486)? out_me_data_i[119] : 
                              (N487)? out_me_data_i[151] : 
                              (N488)? out_me_data_i[183] : 
                              (N489)? out_me_data_i[215] : 
                              (N490)? out_me_data_i[247] : 
                              (N491)? out_me_data_i[279] : 
                              (N492)? out_me_data_i[311] : 
                              (N493)? out_me_data_i[343] : 
                              (N494)? out_me_data_i[375] : 
                              (N495)? out_me_data_i[407] : 1'b0;
  assign out_me_data_o[406] = (N483)? out_me_data_i_0__22_ : 
                              (N484)? out_me_data_i[54] : 
                              (N485)? out_me_data_i[86] : 
                              (N486)? out_me_data_i[118] : 
                              (N487)? out_me_data_i[150] : 
                              (N488)? out_me_data_i[182] : 
                              (N489)? out_me_data_i[214] : 
                              (N490)? out_me_data_i[246] : 
                              (N491)? out_me_data_i[278] : 
                              (N492)? out_me_data_i[310] : 
                              (N493)? out_me_data_i[342] : 
                              (N494)? out_me_data_i[374] : 
                              (N495)? out_me_data_i[406] : 1'b0;
  assign out_me_data_o[405] = (N483)? out_me_data_i_0__21_ : 
                              (N484)? out_me_data_i[53] : 
                              (N485)? out_me_data_i[85] : 
                              (N486)? out_me_data_i[117] : 
                              (N487)? out_me_data_i[149] : 
                              (N488)? out_me_data_i[181] : 
                              (N489)? out_me_data_i[213] : 
                              (N490)? out_me_data_i[245] : 
                              (N491)? out_me_data_i[277] : 
                              (N492)? out_me_data_i[309] : 
                              (N493)? out_me_data_i[341] : 
                              (N494)? out_me_data_i[373] : 
                              (N495)? out_me_data_i[405] : 1'b0;
  assign out_me_data_o[404] = (N483)? out_me_data_i_0__20_ : 
                              (N484)? out_me_data_i[52] : 
                              (N485)? out_me_data_i[84] : 
                              (N486)? out_me_data_i[116] : 
                              (N487)? out_me_data_i[148] : 
                              (N488)? out_me_data_i[180] : 
                              (N489)? out_me_data_i[212] : 
                              (N490)? out_me_data_i[244] : 
                              (N491)? out_me_data_i[276] : 
                              (N492)? out_me_data_i[308] : 
                              (N493)? out_me_data_i[340] : 
                              (N494)? out_me_data_i[372] : 
                              (N495)? out_me_data_i[404] : 1'b0;
  assign out_me_data_o[403] = (N483)? out_me_data_i_0__19_ : 
                              (N484)? out_me_data_i[51] : 
                              (N485)? out_me_data_i[83] : 
                              (N486)? out_me_data_i[115] : 
                              (N487)? out_me_data_i[147] : 
                              (N488)? out_me_data_i[179] : 
                              (N489)? out_me_data_i[211] : 
                              (N490)? out_me_data_i[243] : 
                              (N491)? out_me_data_i[275] : 
                              (N492)? out_me_data_i[307] : 
                              (N493)? out_me_data_i[339] : 
                              (N494)? out_me_data_i[371] : 
                              (N495)? out_me_data_i[403] : 1'b0;
  assign out_me_data_o[402] = (N483)? out_me_data_i_0__18_ : 
                              (N484)? out_me_data_i[50] : 
                              (N485)? out_me_data_i[82] : 
                              (N486)? out_me_data_i[114] : 
                              (N487)? out_me_data_i[146] : 
                              (N488)? out_me_data_i[178] : 
                              (N489)? out_me_data_i[210] : 
                              (N490)? out_me_data_i[242] : 
                              (N491)? out_me_data_i[274] : 
                              (N492)? out_me_data_i[306] : 
                              (N493)? out_me_data_i[338] : 
                              (N494)? out_me_data_i[370] : 
                              (N495)? out_me_data_i[402] : 1'b0;
  assign out_me_data_o[401] = (N483)? out_me_data_i_0__17_ : 
                              (N484)? out_me_data_i[49] : 
                              (N485)? out_me_data_i[81] : 
                              (N486)? out_me_data_i[113] : 
                              (N487)? out_me_data_i[145] : 
                              (N488)? out_me_data_i[177] : 
                              (N489)? out_me_data_i[209] : 
                              (N490)? out_me_data_i[241] : 
                              (N491)? out_me_data_i[273] : 
                              (N492)? out_me_data_i[305] : 
                              (N493)? out_me_data_i[337] : 
                              (N494)? out_me_data_i[369] : 
                              (N495)? out_me_data_i[401] : 1'b0;
  assign out_me_data_o[400] = (N483)? out_me_data_i_0__16_ : 
                              (N484)? out_me_data_i[48] : 
                              (N485)? out_me_data_i[80] : 
                              (N486)? out_me_data_i[112] : 
                              (N487)? out_me_data_i[144] : 
                              (N488)? out_me_data_i[176] : 
                              (N489)? out_me_data_i[208] : 
                              (N490)? out_me_data_i[240] : 
                              (N491)? out_me_data_i[272] : 
                              (N492)? out_me_data_i[304] : 
                              (N493)? out_me_data_i[336] : 
                              (N494)? out_me_data_i[368] : 
                              (N495)? out_me_data_i[400] : 1'b0;
  assign out_me_data_o[399] = (N483)? out_me_data_i_0__15_ : 
                              (N484)? out_me_data_i[47] : 
                              (N485)? out_me_data_i[79] : 
                              (N486)? out_me_data_i[111] : 
                              (N487)? out_me_data_i[143] : 
                              (N488)? out_me_data_i[175] : 
                              (N489)? out_me_data_i[207] : 
                              (N490)? out_me_data_i[239] : 
                              (N491)? out_me_data_i[271] : 
                              (N492)? out_me_data_i[303] : 
                              (N493)? out_me_data_i[335] : 
                              (N494)? out_me_data_i[367] : 
                              (N495)? out_me_data_i[399] : 1'b0;
  assign out_me_data_o[398] = (N483)? out_me_data_i_0__14_ : 
                              (N484)? out_me_data_i[46] : 
                              (N485)? out_me_data_i[78] : 
                              (N486)? out_me_data_i[110] : 
                              (N487)? out_me_data_i[142] : 
                              (N488)? out_me_data_i[174] : 
                              (N489)? out_me_data_i[206] : 
                              (N490)? out_me_data_i[238] : 
                              (N491)? out_me_data_i[270] : 
                              (N492)? out_me_data_i[302] : 
                              (N493)? out_me_data_i[334] : 
                              (N494)? out_me_data_i[366] : 
                              (N495)? out_me_data_i[398] : 1'b0;
  assign out_me_data_o[397] = (N483)? out_me_data_i_0__13_ : 
                              (N484)? out_me_data_i[45] : 
                              (N485)? out_me_data_i[77] : 
                              (N486)? out_me_data_i[109] : 
                              (N487)? out_me_data_i[141] : 
                              (N488)? out_me_data_i[173] : 
                              (N489)? out_me_data_i[205] : 
                              (N490)? out_me_data_i[237] : 
                              (N491)? out_me_data_i[269] : 
                              (N492)? out_me_data_i[301] : 
                              (N493)? out_me_data_i[333] : 
                              (N494)? out_me_data_i[365] : 
                              (N495)? out_me_data_i[397] : 1'b0;
  assign out_me_data_o[396] = (N483)? out_me_data_i_0__12_ : 
                              (N484)? out_me_data_i[44] : 
                              (N485)? out_me_data_i[76] : 
                              (N486)? out_me_data_i[108] : 
                              (N487)? out_me_data_i[140] : 
                              (N488)? out_me_data_i[172] : 
                              (N489)? out_me_data_i[204] : 
                              (N490)? out_me_data_i[236] : 
                              (N491)? out_me_data_i[268] : 
                              (N492)? out_me_data_i[300] : 
                              (N493)? out_me_data_i[332] : 
                              (N494)? out_me_data_i[364] : 
                              (N495)? out_me_data_i[396] : 1'b0;
  assign out_me_data_o[395] = (N483)? out_me_data_i_0__11_ : 
                              (N484)? out_me_data_i[43] : 
                              (N485)? out_me_data_i[75] : 
                              (N486)? out_me_data_i[107] : 
                              (N487)? out_me_data_i[139] : 
                              (N488)? out_me_data_i[171] : 
                              (N489)? out_me_data_i[203] : 
                              (N490)? out_me_data_i[235] : 
                              (N491)? out_me_data_i[267] : 
                              (N492)? out_me_data_i[299] : 
                              (N493)? out_me_data_i[331] : 
                              (N494)? out_me_data_i[363] : 
                              (N495)? out_me_data_i[395] : 1'b0;
  assign out_me_data_o[394] = (N483)? out_me_data_i_0__10_ : 
                              (N484)? out_me_data_i[42] : 
                              (N485)? out_me_data_i[74] : 
                              (N486)? out_me_data_i[106] : 
                              (N487)? out_me_data_i[138] : 
                              (N488)? out_me_data_i[170] : 
                              (N489)? out_me_data_i[202] : 
                              (N490)? out_me_data_i[234] : 
                              (N491)? out_me_data_i[266] : 
                              (N492)? out_me_data_i[298] : 
                              (N493)? out_me_data_i[330] : 
                              (N494)? out_me_data_i[362] : 
                              (N495)? out_me_data_i[394] : 1'b0;
  assign out_me_data_o[393] = (N483)? out_me_data_i_0__9_ : 
                              (N484)? out_me_data_i[41] : 
                              (N485)? out_me_data_i[73] : 
                              (N486)? out_me_data_i[105] : 
                              (N487)? out_me_data_i[137] : 
                              (N488)? out_me_data_i[169] : 
                              (N489)? out_me_data_i[201] : 
                              (N490)? out_me_data_i[233] : 
                              (N491)? out_me_data_i[265] : 
                              (N492)? out_me_data_i[297] : 
                              (N493)? out_me_data_i[329] : 
                              (N494)? out_me_data_i[361] : 
                              (N495)? out_me_data_i[393] : 1'b0;
  assign out_me_data_o[392] = (N483)? out_me_data_i_0__8_ : 
                              (N484)? out_me_data_i[40] : 
                              (N485)? out_me_data_i[72] : 
                              (N486)? out_me_data_i[104] : 
                              (N487)? out_me_data_i[136] : 
                              (N488)? out_me_data_i[168] : 
                              (N489)? out_me_data_i[200] : 
                              (N490)? out_me_data_i[232] : 
                              (N491)? out_me_data_i[264] : 
                              (N492)? out_me_data_i[296] : 
                              (N493)? out_me_data_i[328] : 
                              (N494)? out_me_data_i[360] : 
                              (N495)? out_me_data_i[392] : 1'b0;
  assign out_me_data_o[391] = (N483)? out_me_data_i_0__7_ : 
                              (N484)? out_me_data_i[39] : 
                              (N485)? out_me_data_i[71] : 
                              (N486)? out_me_data_i[103] : 
                              (N487)? out_me_data_i[135] : 
                              (N488)? out_me_data_i[167] : 
                              (N489)? out_me_data_i[199] : 
                              (N490)? out_me_data_i[231] : 
                              (N491)? out_me_data_i[263] : 
                              (N492)? out_me_data_i[295] : 
                              (N493)? out_me_data_i[327] : 
                              (N494)? out_me_data_i[359] : 
                              (N495)? out_me_data_i[391] : 1'b0;
  assign out_me_data_o[390] = (N483)? out_me_data_i_0__6_ : 
                              (N484)? out_me_data_i[38] : 
                              (N485)? out_me_data_i[70] : 
                              (N486)? out_me_data_i[102] : 
                              (N487)? out_me_data_i[134] : 
                              (N488)? out_me_data_i[166] : 
                              (N489)? out_me_data_i[198] : 
                              (N490)? out_me_data_i[230] : 
                              (N491)? out_me_data_i[262] : 
                              (N492)? out_me_data_i[294] : 
                              (N493)? out_me_data_i[326] : 
                              (N494)? out_me_data_i[358] : 
                              (N495)? out_me_data_i[390] : 1'b0;
  assign out_me_data_o[389] = (N483)? out_me_data_i_0__5_ : 
                              (N484)? out_me_data_i[37] : 
                              (N485)? out_me_data_i[69] : 
                              (N486)? out_me_data_i[101] : 
                              (N487)? out_me_data_i[133] : 
                              (N488)? out_me_data_i[165] : 
                              (N489)? out_me_data_i[197] : 
                              (N490)? out_me_data_i[229] : 
                              (N491)? out_me_data_i[261] : 
                              (N492)? out_me_data_i[293] : 
                              (N493)? out_me_data_i[325] : 
                              (N494)? out_me_data_i[357] : 
                              (N495)? out_me_data_i[389] : 1'b0;
  assign out_me_data_o[388] = (N483)? out_me_data_i_0__4_ : 
                              (N484)? out_me_data_i[36] : 
                              (N485)? out_me_data_i[68] : 
                              (N486)? out_me_data_i[100] : 
                              (N487)? out_me_data_i[132] : 
                              (N488)? out_me_data_i[164] : 
                              (N489)? out_me_data_i[196] : 
                              (N490)? out_me_data_i[228] : 
                              (N491)? out_me_data_i[260] : 
                              (N492)? out_me_data_i[292] : 
                              (N493)? out_me_data_i[324] : 
                              (N494)? out_me_data_i[356] : 
                              (N495)? out_me_data_i[388] : 1'b0;
  assign out_me_data_o[387] = (N483)? out_me_data_i_0__3_ : 
                              (N484)? out_me_data_i[35] : 
                              (N485)? out_me_data_i[67] : 
                              (N486)? out_me_data_i[99] : 
                              (N487)? out_me_data_i[131] : 
                              (N488)? out_me_data_i[163] : 
                              (N489)? out_me_data_i[195] : 
                              (N490)? out_me_data_i[227] : 
                              (N491)? out_me_data_i[259] : 
                              (N492)? out_me_data_i[291] : 
                              (N493)? out_me_data_i[323] : 
                              (N494)? out_me_data_i[355] : 
                              (N495)? out_me_data_i[387] : 1'b0;
  assign out_me_data_o[386] = (N483)? out_me_data_i_0__2_ : 
                              (N484)? out_me_data_i[34] : 
                              (N485)? out_me_data_i[66] : 
                              (N486)? out_me_data_i[98] : 
                              (N487)? out_me_data_i[130] : 
                              (N488)? out_me_data_i[162] : 
                              (N489)? out_me_data_i[194] : 
                              (N490)? out_me_data_i[226] : 
                              (N491)? out_me_data_i[258] : 
                              (N492)? out_me_data_i[290] : 
                              (N493)? out_me_data_i[322] : 
                              (N494)? out_me_data_i[354] : 
                              (N495)? out_me_data_i[386] : 1'b0;
  assign out_me_data_o[385] = (N483)? out_me_data_i_0__1_ : 
                              (N484)? out_me_data_i[33] : 
                              (N485)? out_me_data_i[65] : 
                              (N486)? out_me_data_i[97] : 
                              (N487)? out_me_data_i[129] : 
                              (N488)? out_me_data_i[161] : 
                              (N489)? out_me_data_i[193] : 
                              (N490)? out_me_data_i[225] : 
                              (N491)? out_me_data_i[257] : 
                              (N492)? out_me_data_i[289] : 
                              (N493)? out_me_data_i[321] : 
                              (N494)? out_me_data_i[353] : 
                              (N495)? out_me_data_i[385] : 1'b0;
  assign out_me_data_o[384] = (N483)? out_me_data_i_0__0_ : 
                              (N484)? out_me_data_i[32] : 
                              (N485)? out_me_data_i[64] : 
                              (N486)? out_me_data_i[96] : 
                              (N487)? out_me_data_i[128] : 
                              (N488)? out_me_data_i[160] : 
                              (N489)? out_me_data_i[192] : 
                              (N490)? out_me_data_i[224] : 
                              (N491)? out_me_data_i[256] : 
                              (N492)? out_me_data_i[288] : 
                              (N493)? out_me_data_i[320] : 
                              (N494)? out_me_data_i[352] : 
                              (N495)? out_me_data_i[384] : 1'b0;
  assign out_me_data_o[383] = (N496)? out_me_data_i_0__31_ : 
                              (N497)? out_me_data_i[63] : 
                              (N498)? out_me_data_i[95] : 
                              (N499)? out_me_data_i[127] : 
                              (N500)? out_me_data_i[159] : 
                              (N501)? out_me_data_i[191] : 
                              (N502)? out_me_data_i[223] : 
                              (N503)? out_me_data_i[255] : 
                              (N504)? out_me_data_i[287] : 
                              (N505)? out_me_data_i[319] : 
                              (N506)? out_me_data_i[351] : 
                              (N507)? out_me_data_i[383] : 1'b0;
  assign N496 = N2050;
  assign N497 = N2052;
  assign N498 = N2054;
  assign N499 = N2056;
  assign N500 = N2058;
  assign N501 = N2059;
  assign N502 = N2060;
  assign N503 = N2061;
  assign N504 = N2051;
  assign N505 = N2053;
  assign N506 = N2055;
  assign N507 = N2057;
  assign out_me_data_o[382] = (N496)? out_me_data_i_0__30_ : 
                              (N497)? out_me_data_i[62] : 
                              (N498)? out_me_data_i[94] : 
                              (N499)? out_me_data_i[126] : 
                              (N500)? out_me_data_i[158] : 
                              (N501)? out_me_data_i[190] : 
                              (N502)? out_me_data_i[222] : 
                              (N503)? out_me_data_i[254] : 
                              (N504)? out_me_data_i[286] : 
                              (N505)? out_me_data_i[318] : 
                              (N506)? out_me_data_i[350] : 
                              (N507)? out_me_data_i[382] : 1'b0;
  assign out_me_data_o[381] = (N496)? out_me_data_i_0__29_ : 
                              (N497)? out_me_data_i[61] : 
                              (N498)? out_me_data_i[93] : 
                              (N499)? out_me_data_i[125] : 
                              (N500)? out_me_data_i[157] : 
                              (N501)? out_me_data_i[189] : 
                              (N502)? out_me_data_i[221] : 
                              (N503)? out_me_data_i[253] : 
                              (N504)? out_me_data_i[285] : 
                              (N505)? out_me_data_i[317] : 
                              (N506)? out_me_data_i[349] : 
                              (N507)? out_me_data_i[381] : 1'b0;
  assign out_me_data_o[380] = (N496)? out_me_data_i_0__28_ : 
                              (N497)? out_me_data_i[60] : 
                              (N498)? out_me_data_i[92] : 
                              (N499)? out_me_data_i[124] : 
                              (N500)? out_me_data_i[156] : 
                              (N501)? out_me_data_i[188] : 
                              (N502)? out_me_data_i[220] : 
                              (N503)? out_me_data_i[252] : 
                              (N504)? out_me_data_i[284] : 
                              (N505)? out_me_data_i[316] : 
                              (N506)? out_me_data_i[348] : 
                              (N507)? out_me_data_i[380] : 1'b0;
  assign out_me_data_o[379] = (N496)? out_me_data_i_0__27_ : 
                              (N497)? out_me_data_i[59] : 
                              (N498)? out_me_data_i[91] : 
                              (N499)? out_me_data_i[123] : 
                              (N500)? out_me_data_i[155] : 
                              (N501)? out_me_data_i[187] : 
                              (N502)? out_me_data_i[219] : 
                              (N503)? out_me_data_i[251] : 
                              (N504)? out_me_data_i[283] : 
                              (N505)? out_me_data_i[315] : 
                              (N506)? out_me_data_i[347] : 
                              (N507)? out_me_data_i[379] : 1'b0;
  assign out_me_data_o[378] = (N496)? out_me_data_i_0__26_ : 
                              (N497)? out_me_data_i[58] : 
                              (N498)? out_me_data_i[90] : 
                              (N499)? out_me_data_i[122] : 
                              (N500)? out_me_data_i[154] : 
                              (N501)? out_me_data_i[186] : 
                              (N502)? out_me_data_i[218] : 
                              (N503)? out_me_data_i[250] : 
                              (N504)? out_me_data_i[282] : 
                              (N505)? out_me_data_i[314] : 
                              (N506)? out_me_data_i[346] : 
                              (N507)? out_me_data_i[378] : 1'b0;
  assign out_me_data_o[377] = (N496)? out_me_data_i_0__25_ : 
                              (N497)? out_me_data_i[57] : 
                              (N498)? out_me_data_i[89] : 
                              (N499)? out_me_data_i[121] : 
                              (N500)? out_me_data_i[153] : 
                              (N501)? out_me_data_i[185] : 
                              (N502)? out_me_data_i[217] : 
                              (N503)? out_me_data_i[249] : 
                              (N504)? out_me_data_i[281] : 
                              (N505)? out_me_data_i[313] : 
                              (N506)? out_me_data_i[345] : 
                              (N507)? out_me_data_i[377] : 1'b0;
  assign out_me_data_o[376] = (N496)? out_me_data_i_0__24_ : 
                              (N497)? out_me_data_i[56] : 
                              (N498)? out_me_data_i[88] : 
                              (N499)? out_me_data_i[120] : 
                              (N500)? out_me_data_i[152] : 
                              (N501)? out_me_data_i[184] : 
                              (N502)? out_me_data_i[216] : 
                              (N503)? out_me_data_i[248] : 
                              (N504)? out_me_data_i[280] : 
                              (N505)? out_me_data_i[312] : 
                              (N506)? out_me_data_i[344] : 
                              (N507)? out_me_data_i[376] : 1'b0;
  assign out_me_data_o[375] = (N496)? out_me_data_i_0__23_ : 
                              (N497)? out_me_data_i[55] : 
                              (N498)? out_me_data_i[87] : 
                              (N499)? out_me_data_i[119] : 
                              (N500)? out_me_data_i[151] : 
                              (N501)? out_me_data_i[183] : 
                              (N502)? out_me_data_i[215] : 
                              (N503)? out_me_data_i[247] : 
                              (N504)? out_me_data_i[279] : 
                              (N505)? out_me_data_i[311] : 
                              (N506)? out_me_data_i[343] : 
                              (N507)? out_me_data_i[375] : 1'b0;
  assign out_me_data_o[374] = (N496)? out_me_data_i_0__22_ : 
                              (N497)? out_me_data_i[54] : 
                              (N498)? out_me_data_i[86] : 
                              (N499)? out_me_data_i[118] : 
                              (N500)? out_me_data_i[150] : 
                              (N501)? out_me_data_i[182] : 
                              (N502)? out_me_data_i[214] : 
                              (N503)? out_me_data_i[246] : 
                              (N504)? out_me_data_i[278] : 
                              (N505)? out_me_data_i[310] : 
                              (N506)? out_me_data_i[342] : 
                              (N507)? out_me_data_i[374] : 1'b0;
  assign out_me_data_o[373] = (N496)? out_me_data_i_0__21_ : 
                              (N497)? out_me_data_i[53] : 
                              (N498)? out_me_data_i[85] : 
                              (N499)? out_me_data_i[117] : 
                              (N500)? out_me_data_i[149] : 
                              (N501)? out_me_data_i[181] : 
                              (N502)? out_me_data_i[213] : 
                              (N503)? out_me_data_i[245] : 
                              (N504)? out_me_data_i[277] : 
                              (N505)? out_me_data_i[309] : 
                              (N506)? out_me_data_i[341] : 
                              (N507)? out_me_data_i[373] : 1'b0;
  assign out_me_data_o[372] = (N496)? out_me_data_i_0__20_ : 
                              (N497)? out_me_data_i[52] : 
                              (N498)? out_me_data_i[84] : 
                              (N499)? out_me_data_i[116] : 
                              (N500)? out_me_data_i[148] : 
                              (N501)? out_me_data_i[180] : 
                              (N502)? out_me_data_i[212] : 
                              (N503)? out_me_data_i[244] : 
                              (N504)? out_me_data_i[276] : 
                              (N505)? out_me_data_i[308] : 
                              (N506)? out_me_data_i[340] : 
                              (N507)? out_me_data_i[372] : 1'b0;
  assign out_me_data_o[371] = (N496)? out_me_data_i_0__19_ : 
                              (N497)? out_me_data_i[51] : 
                              (N498)? out_me_data_i[83] : 
                              (N499)? out_me_data_i[115] : 
                              (N500)? out_me_data_i[147] : 
                              (N501)? out_me_data_i[179] : 
                              (N502)? out_me_data_i[211] : 
                              (N503)? out_me_data_i[243] : 
                              (N504)? out_me_data_i[275] : 
                              (N505)? out_me_data_i[307] : 
                              (N506)? out_me_data_i[339] : 
                              (N507)? out_me_data_i[371] : 1'b0;
  assign out_me_data_o[370] = (N496)? out_me_data_i_0__18_ : 
                              (N497)? out_me_data_i[50] : 
                              (N498)? out_me_data_i[82] : 
                              (N499)? out_me_data_i[114] : 
                              (N500)? out_me_data_i[146] : 
                              (N501)? out_me_data_i[178] : 
                              (N502)? out_me_data_i[210] : 
                              (N503)? out_me_data_i[242] : 
                              (N504)? out_me_data_i[274] : 
                              (N505)? out_me_data_i[306] : 
                              (N506)? out_me_data_i[338] : 
                              (N507)? out_me_data_i[370] : 1'b0;
  assign out_me_data_o[369] = (N496)? out_me_data_i_0__17_ : 
                              (N497)? out_me_data_i[49] : 
                              (N498)? out_me_data_i[81] : 
                              (N499)? out_me_data_i[113] : 
                              (N500)? out_me_data_i[145] : 
                              (N501)? out_me_data_i[177] : 
                              (N502)? out_me_data_i[209] : 
                              (N503)? out_me_data_i[241] : 
                              (N504)? out_me_data_i[273] : 
                              (N505)? out_me_data_i[305] : 
                              (N506)? out_me_data_i[337] : 
                              (N507)? out_me_data_i[369] : 1'b0;
  assign out_me_data_o[368] = (N496)? out_me_data_i_0__16_ : 
                              (N497)? out_me_data_i[48] : 
                              (N498)? out_me_data_i[80] : 
                              (N499)? out_me_data_i[112] : 
                              (N500)? out_me_data_i[144] : 
                              (N501)? out_me_data_i[176] : 
                              (N502)? out_me_data_i[208] : 
                              (N503)? out_me_data_i[240] : 
                              (N504)? out_me_data_i[272] : 
                              (N505)? out_me_data_i[304] : 
                              (N506)? out_me_data_i[336] : 
                              (N507)? out_me_data_i[368] : 1'b0;
  assign out_me_data_o[367] = (N496)? out_me_data_i_0__15_ : 
                              (N497)? out_me_data_i[47] : 
                              (N498)? out_me_data_i[79] : 
                              (N499)? out_me_data_i[111] : 
                              (N500)? out_me_data_i[143] : 
                              (N501)? out_me_data_i[175] : 
                              (N502)? out_me_data_i[207] : 
                              (N503)? out_me_data_i[239] : 
                              (N504)? out_me_data_i[271] : 
                              (N505)? out_me_data_i[303] : 
                              (N506)? out_me_data_i[335] : 
                              (N507)? out_me_data_i[367] : 1'b0;
  assign out_me_data_o[366] = (N496)? out_me_data_i_0__14_ : 
                              (N497)? out_me_data_i[46] : 
                              (N498)? out_me_data_i[78] : 
                              (N499)? out_me_data_i[110] : 
                              (N500)? out_me_data_i[142] : 
                              (N501)? out_me_data_i[174] : 
                              (N502)? out_me_data_i[206] : 
                              (N503)? out_me_data_i[238] : 
                              (N504)? out_me_data_i[270] : 
                              (N505)? out_me_data_i[302] : 
                              (N506)? out_me_data_i[334] : 
                              (N507)? out_me_data_i[366] : 1'b0;
  assign out_me_data_o[365] = (N496)? out_me_data_i_0__13_ : 
                              (N497)? out_me_data_i[45] : 
                              (N498)? out_me_data_i[77] : 
                              (N499)? out_me_data_i[109] : 
                              (N500)? out_me_data_i[141] : 
                              (N501)? out_me_data_i[173] : 
                              (N502)? out_me_data_i[205] : 
                              (N503)? out_me_data_i[237] : 
                              (N504)? out_me_data_i[269] : 
                              (N505)? out_me_data_i[301] : 
                              (N506)? out_me_data_i[333] : 
                              (N507)? out_me_data_i[365] : 1'b0;
  assign out_me_data_o[364] = (N496)? out_me_data_i_0__12_ : 
                              (N497)? out_me_data_i[44] : 
                              (N498)? out_me_data_i[76] : 
                              (N499)? out_me_data_i[108] : 
                              (N500)? out_me_data_i[140] : 
                              (N501)? out_me_data_i[172] : 
                              (N502)? out_me_data_i[204] : 
                              (N503)? out_me_data_i[236] : 
                              (N504)? out_me_data_i[268] : 
                              (N505)? out_me_data_i[300] : 
                              (N506)? out_me_data_i[332] : 
                              (N507)? out_me_data_i[364] : 1'b0;
  assign out_me_data_o[363] = (N496)? out_me_data_i_0__11_ : 
                              (N497)? out_me_data_i[43] : 
                              (N498)? out_me_data_i[75] : 
                              (N499)? out_me_data_i[107] : 
                              (N500)? out_me_data_i[139] : 
                              (N501)? out_me_data_i[171] : 
                              (N502)? out_me_data_i[203] : 
                              (N503)? out_me_data_i[235] : 
                              (N504)? out_me_data_i[267] : 
                              (N505)? out_me_data_i[299] : 
                              (N506)? out_me_data_i[331] : 
                              (N507)? out_me_data_i[363] : 1'b0;
  assign out_me_data_o[362] = (N496)? out_me_data_i_0__10_ : 
                              (N497)? out_me_data_i[42] : 
                              (N498)? out_me_data_i[74] : 
                              (N499)? out_me_data_i[106] : 
                              (N500)? out_me_data_i[138] : 
                              (N501)? out_me_data_i[170] : 
                              (N502)? out_me_data_i[202] : 
                              (N503)? out_me_data_i[234] : 
                              (N504)? out_me_data_i[266] : 
                              (N505)? out_me_data_i[298] : 
                              (N506)? out_me_data_i[330] : 
                              (N507)? out_me_data_i[362] : 1'b0;
  assign out_me_data_o[361] = (N496)? out_me_data_i_0__9_ : 
                              (N497)? out_me_data_i[41] : 
                              (N498)? out_me_data_i[73] : 
                              (N499)? out_me_data_i[105] : 
                              (N500)? out_me_data_i[137] : 
                              (N501)? out_me_data_i[169] : 
                              (N502)? out_me_data_i[201] : 
                              (N503)? out_me_data_i[233] : 
                              (N504)? out_me_data_i[265] : 
                              (N505)? out_me_data_i[297] : 
                              (N506)? out_me_data_i[329] : 
                              (N507)? out_me_data_i[361] : 1'b0;
  assign out_me_data_o[360] = (N496)? out_me_data_i_0__8_ : 
                              (N497)? out_me_data_i[40] : 
                              (N498)? out_me_data_i[72] : 
                              (N499)? out_me_data_i[104] : 
                              (N500)? out_me_data_i[136] : 
                              (N501)? out_me_data_i[168] : 
                              (N502)? out_me_data_i[200] : 
                              (N503)? out_me_data_i[232] : 
                              (N504)? out_me_data_i[264] : 
                              (N505)? out_me_data_i[296] : 
                              (N506)? out_me_data_i[328] : 
                              (N507)? out_me_data_i[360] : 1'b0;
  assign out_me_data_o[359] = (N496)? out_me_data_i_0__7_ : 
                              (N497)? out_me_data_i[39] : 
                              (N498)? out_me_data_i[71] : 
                              (N499)? out_me_data_i[103] : 
                              (N500)? out_me_data_i[135] : 
                              (N501)? out_me_data_i[167] : 
                              (N502)? out_me_data_i[199] : 
                              (N503)? out_me_data_i[231] : 
                              (N504)? out_me_data_i[263] : 
                              (N505)? out_me_data_i[295] : 
                              (N506)? out_me_data_i[327] : 
                              (N507)? out_me_data_i[359] : 1'b0;
  assign out_me_data_o[358] = (N496)? out_me_data_i_0__6_ : 
                              (N497)? out_me_data_i[38] : 
                              (N498)? out_me_data_i[70] : 
                              (N499)? out_me_data_i[102] : 
                              (N500)? out_me_data_i[134] : 
                              (N501)? out_me_data_i[166] : 
                              (N502)? out_me_data_i[198] : 
                              (N503)? out_me_data_i[230] : 
                              (N504)? out_me_data_i[262] : 
                              (N505)? out_me_data_i[294] : 
                              (N506)? out_me_data_i[326] : 
                              (N507)? out_me_data_i[358] : 1'b0;
  assign out_me_data_o[357] = (N496)? out_me_data_i_0__5_ : 
                              (N497)? out_me_data_i[37] : 
                              (N498)? out_me_data_i[69] : 
                              (N499)? out_me_data_i[101] : 
                              (N500)? out_me_data_i[133] : 
                              (N501)? out_me_data_i[165] : 
                              (N502)? out_me_data_i[197] : 
                              (N503)? out_me_data_i[229] : 
                              (N504)? out_me_data_i[261] : 
                              (N505)? out_me_data_i[293] : 
                              (N506)? out_me_data_i[325] : 
                              (N507)? out_me_data_i[357] : 1'b0;
  assign out_me_data_o[356] = (N496)? out_me_data_i_0__4_ : 
                              (N497)? out_me_data_i[36] : 
                              (N498)? out_me_data_i[68] : 
                              (N499)? out_me_data_i[100] : 
                              (N500)? out_me_data_i[132] : 
                              (N501)? out_me_data_i[164] : 
                              (N502)? out_me_data_i[196] : 
                              (N503)? out_me_data_i[228] : 
                              (N504)? out_me_data_i[260] : 
                              (N505)? out_me_data_i[292] : 
                              (N506)? out_me_data_i[324] : 
                              (N507)? out_me_data_i[356] : 1'b0;
  assign out_me_data_o[355] = (N496)? out_me_data_i_0__3_ : 
                              (N497)? out_me_data_i[35] : 
                              (N498)? out_me_data_i[67] : 
                              (N499)? out_me_data_i[99] : 
                              (N500)? out_me_data_i[131] : 
                              (N501)? out_me_data_i[163] : 
                              (N502)? out_me_data_i[195] : 
                              (N503)? out_me_data_i[227] : 
                              (N504)? out_me_data_i[259] : 
                              (N505)? out_me_data_i[291] : 
                              (N506)? out_me_data_i[323] : 
                              (N507)? out_me_data_i[355] : 1'b0;
  assign out_me_data_o[354] = (N496)? out_me_data_i_0__2_ : 
                              (N497)? out_me_data_i[34] : 
                              (N498)? out_me_data_i[66] : 
                              (N499)? out_me_data_i[98] : 
                              (N500)? out_me_data_i[130] : 
                              (N501)? out_me_data_i[162] : 
                              (N502)? out_me_data_i[194] : 
                              (N503)? out_me_data_i[226] : 
                              (N504)? out_me_data_i[258] : 
                              (N505)? out_me_data_i[290] : 
                              (N506)? out_me_data_i[322] : 
                              (N507)? out_me_data_i[354] : 1'b0;
  assign out_me_data_o[353] = (N496)? out_me_data_i_0__1_ : 
                              (N497)? out_me_data_i[33] : 
                              (N498)? out_me_data_i[65] : 
                              (N499)? out_me_data_i[97] : 
                              (N500)? out_me_data_i[129] : 
                              (N501)? out_me_data_i[161] : 
                              (N502)? out_me_data_i[193] : 
                              (N503)? out_me_data_i[225] : 
                              (N504)? out_me_data_i[257] : 
                              (N505)? out_me_data_i[289] : 
                              (N506)? out_me_data_i[321] : 
                              (N507)? out_me_data_i[353] : 1'b0;
  assign out_me_data_o[352] = (N496)? out_me_data_i_0__0_ : 
                              (N497)? out_me_data_i[32] : 
                              (N498)? out_me_data_i[64] : 
                              (N499)? out_me_data_i[96] : 
                              (N500)? out_me_data_i[128] : 
                              (N501)? out_me_data_i[160] : 
                              (N502)? out_me_data_i[192] : 
                              (N503)? out_me_data_i[224] : 
                              (N504)? out_me_data_i[256] : 
                              (N505)? out_me_data_i[288] : 
                              (N506)? out_me_data_i[320] : 
                              (N507)? out_me_data_i[352] : 1'b0;
  assign out_me_data_o[351] = (N508)? out_me_data_i_0__31_ : 
                              (N509)? out_me_data_i[63] : 
                              (N510)? out_me_data_i[95] : 
                              (N511)? out_me_data_i[127] : 
                              (N512)? out_me_data_i[159] : 
                              (N513)? out_me_data_i[191] : 
                              (N514)? out_me_data_i[223] : 
                              (N515)? out_me_data_i[255] : 
                              (N516)? out_me_data_i[287] : 
                              (N517)? out_me_data_i[319] : 
                              (N518)? out_me_data_i[351] : 1'b0;
  assign N508 = N1927;
  assign N509 = N1929;
  assign N510 = N1931;
  assign N511 = N1933;
  assign N512 = N1934;
  assign N513 = N1935;
  assign N514 = N1936;
  assign N515 = N1937;
  assign N516 = N1928;
  assign N517 = N1930;
  assign N518 = N1932;
  assign out_me_data_o[350] = (N508)? out_me_data_i_0__30_ : 
                              (N509)? out_me_data_i[62] : 
                              (N510)? out_me_data_i[94] : 
                              (N511)? out_me_data_i[126] : 
                              (N512)? out_me_data_i[158] : 
                              (N513)? out_me_data_i[190] : 
                              (N514)? out_me_data_i[222] : 
                              (N515)? out_me_data_i[254] : 
                              (N516)? out_me_data_i[286] : 
                              (N517)? out_me_data_i[318] : 
                              (N518)? out_me_data_i[350] : 1'b0;
  assign out_me_data_o[349] = (N508)? out_me_data_i_0__29_ : 
                              (N509)? out_me_data_i[61] : 
                              (N510)? out_me_data_i[93] : 
                              (N511)? out_me_data_i[125] : 
                              (N512)? out_me_data_i[157] : 
                              (N513)? out_me_data_i[189] : 
                              (N514)? out_me_data_i[221] : 
                              (N515)? out_me_data_i[253] : 
                              (N516)? out_me_data_i[285] : 
                              (N517)? out_me_data_i[317] : 
                              (N518)? out_me_data_i[349] : 1'b0;
  assign out_me_data_o[348] = (N508)? out_me_data_i_0__28_ : 
                              (N509)? out_me_data_i[60] : 
                              (N510)? out_me_data_i[92] : 
                              (N511)? out_me_data_i[124] : 
                              (N512)? out_me_data_i[156] : 
                              (N513)? out_me_data_i[188] : 
                              (N514)? out_me_data_i[220] : 
                              (N515)? out_me_data_i[252] : 
                              (N516)? out_me_data_i[284] : 
                              (N517)? out_me_data_i[316] : 
                              (N518)? out_me_data_i[348] : 1'b0;
  assign out_me_data_o[347] = (N508)? out_me_data_i_0__27_ : 
                              (N509)? out_me_data_i[59] : 
                              (N510)? out_me_data_i[91] : 
                              (N511)? out_me_data_i[123] : 
                              (N512)? out_me_data_i[155] : 
                              (N513)? out_me_data_i[187] : 
                              (N514)? out_me_data_i[219] : 
                              (N515)? out_me_data_i[251] : 
                              (N516)? out_me_data_i[283] : 
                              (N517)? out_me_data_i[315] : 
                              (N518)? out_me_data_i[347] : 1'b0;
  assign out_me_data_o[346] = (N508)? out_me_data_i_0__26_ : 
                              (N509)? out_me_data_i[58] : 
                              (N510)? out_me_data_i[90] : 
                              (N511)? out_me_data_i[122] : 
                              (N512)? out_me_data_i[154] : 
                              (N513)? out_me_data_i[186] : 
                              (N514)? out_me_data_i[218] : 
                              (N515)? out_me_data_i[250] : 
                              (N516)? out_me_data_i[282] : 
                              (N517)? out_me_data_i[314] : 
                              (N518)? out_me_data_i[346] : 1'b0;
  assign out_me_data_o[345] = (N508)? out_me_data_i_0__25_ : 
                              (N509)? out_me_data_i[57] : 
                              (N510)? out_me_data_i[89] : 
                              (N511)? out_me_data_i[121] : 
                              (N512)? out_me_data_i[153] : 
                              (N513)? out_me_data_i[185] : 
                              (N514)? out_me_data_i[217] : 
                              (N515)? out_me_data_i[249] : 
                              (N516)? out_me_data_i[281] : 
                              (N517)? out_me_data_i[313] : 
                              (N518)? out_me_data_i[345] : 1'b0;
  assign out_me_data_o[344] = (N508)? out_me_data_i_0__24_ : 
                              (N509)? out_me_data_i[56] : 
                              (N510)? out_me_data_i[88] : 
                              (N511)? out_me_data_i[120] : 
                              (N512)? out_me_data_i[152] : 
                              (N513)? out_me_data_i[184] : 
                              (N514)? out_me_data_i[216] : 
                              (N515)? out_me_data_i[248] : 
                              (N516)? out_me_data_i[280] : 
                              (N517)? out_me_data_i[312] : 
                              (N518)? out_me_data_i[344] : 1'b0;
  assign out_me_data_o[343] = (N508)? out_me_data_i_0__23_ : 
                              (N509)? out_me_data_i[55] : 
                              (N510)? out_me_data_i[87] : 
                              (N511)? out_me_data_i[119] : 
                              (N512)? out_me_data_i[151] : 
                              (N513)? out_me_data_i[183] : 
                              (N514)? out_me_data_i[215] : 
                              (N515)? out_me_data_i[247] : 
                              (N516)? out_me_data_i[279] : 
                              (N517)? out_me_data_i[311] : 
                              (N518)? out_me_data_i[343] : 1'b0;
  assign out_me_data_o[342] = (N508)? out_me_data_i_0__22_ : 
                              (N509)? out_me_data_i[54] : 
                              (N510)? out_me_data_i[86] : 
                              (N511)? out_me_data_i[118] : 
                              (N512)? out_me_data_i[150] : 
                              (N513)? out_me_data_i[182] : 
                              (N514)? out_me_data_i[214] : 
                              (N515)? out_me_data_i[246] : 
                              (N516)? out_me_data_i[278] : 
                              (N517)? out_me_data_i[310] : 
                              (N518)? out_me_data_i[342] : 1'b0;
  assign out_me_data_o[341] = (N508)? out_me_data_i_0__21_ : 
                              (N509)? out_me_data_i[53] : 
                              (N510)? out_me_data_i[85] : 
                              (N511)? out_me_data_i[117] : 
                              (N512)? out_me_data_i[149] : 
                              (N513)? out_me_data_i[181] : 
                              (N514)? out_me_data_i[213] : 
                              (N515)? out_me_data_i[245] : 
                              (N516)? out_me_data_i[277] : 
                              (N517)? out_me_data_i[309] : 
                              (N518)? out_me_data_i[341] : 1'b0;
  assign out_me_data_o[340] = (N508)? out_me_data_i_0__20_ : 
                              (N509)? out_me_data_i[52] : 
                              (N510)? out_me_data_i[84] : 
                              (N511)? out_me_data_i[116] : 
                              (N512)? out_me_data_i[148] : 
                              (N513)? out_me_data_i[180] : 
                              (N514)? out_me_data_i[212] : 
                              (N515)? out_me_data_i[244] : 
                              (N516)? out_me_data_i[276] : 
                              (N517)? out_me_data_i[308] : 
                              (N518)? out_me_data_i[340] : 1'b0;
  assign out_me_data_o[339] = (N508)? out_me_data_i_0__19_ : 
                              (N509)? out_me_data_i[51] : 
                              (N510)? out_me_data_i[83] : 
                              (N511)? out_me_data_i[115] : 
                              (N512)? out_me_data_i[147] : 
                              (N513)? out_me_data_i[179] : 
                              (N514)? out_me_data_i[211] : 
                              (N515)? out_me_data_i[243] : 
                              (N516)? out_me_data_i[275] : 
                              (N517)? out_me_data_i[307] : 
                              (N518)? out_me_data_i[339] : 1'b0;
  assign out_me_data_o[338] = (N508)? out_me_data_i_0__18_ : 
                              (N509)? out_me_data_i[50] : 
                              (N510)? out_me_data_i[82] : 
                              (N511)? out_me_data_i[114] : 
                              (N512)? out_me_data_i[146] : 
                              (N513)? out_me_data_i[178] : 
                              (N514)? out_me_data_i[210] : 
                              (N515)? out_me_data_i[242] : 
                              (N516)? out_me_data_i[274] : 
                              (N517)? out_me_data_i[306] : 
                              (N518)? out_me_data_i[338] : 1'b0;
  assign out_me_data_o[337] = (N508)? out_me_data_i_0__17_ : 
                              (N509)? out_me_data_i[49] : 
                              (N510)? out_me_data_i[81] : 
                              (N511)? out_me_data_i[113] : 
                              (N512)? out_me_data_i[145] : 
                              (N513)? out_me_data_i[177] : 
                              (N514)? out_me_data_i[209] : 
                              (N515)? out_me_data_i[241] : 
                              (N516)? out_me_data_i[273] : 
                              (N517)? out_me_data_i[305] : 
                              (N518)? out_me_data_i[337] : 1'b0;
  assign out_me_data_o[336] = (N508)? out_me_data_i_0__16_ : 
                              (N509)? out_me_data_i[48] : 
                              (N510)? out_me_data_i[80] : 
                              (N511)? out_me_data_i[112] : 
                              (N512)? out_me_data_i[144] : 
                              (N513)? out_me_data_i[176] : 
                              (N514)? out_me_data_i[208] : 
                              (N515)? out_me_data_i[240] : 
                              (N516)? out_me_data_i[272] : 
                              (N517)? out_me_data_i[304] : 
                              (N518)? out_me_data_i[336] : 1'b0;
  assign out_me_data_o[335] = (N508)? out_me_data_i_0__15_ : 
                              (N509)? out_me_data_i[47] : 
                              (N510)? out_me_data_i[79] : 
                              (N511)? out_me_data_i[111] : 
                              (N512)? out_me_data_i[143] : 
                              (N513)? out_me_data_i[175] : 
                              (N514)? out_me_data_i[207] : 
                              (N515)? out_me_data_i[239] : 
                              (N516)? out_me_data_i[271] : 
                              (N517)? out_me_data_i[303] : 
                              (N518)? out_me_data_i[335] : 1'b0;
  assign out_me_data_o[334] = (N508)? out_me_data_i_0__14_ : 
                              (N509)? out_me_data_i[46] : 
                              (N510)? out_me_data_i[78] : 
                              (N511)? out_me_data_i[110] : 
                              (N512)? out_me_data_i[142] : 
                              (N513)? out_me_data_i[174] : 
                              (N514)? out_me_data_i[206] : 
                              (N515)? out_me_data_i[238] : 
                              (N516)? out_me_data_i[270] : 
                              (N517)? out_me_data_i[302] : 
                              (N518)? out_me_data_i[334] : 1'b0;
  assign out_me_data_o[333] = (N508)? out_me_data_i_0__13_ : 
                              (N509)? out_me_data_i[45] : 
                              (N510)? out_me_data_i[77] : 
                              (N511)? out_me_data_i[109] : 
                              (N512)? out_me_data_i[141] : 
                              (N513)? out_me_data_i[173] : 
                              (N514)? out_me_data_i[205] : 
                              (N515)? out_me_data_i[237] : 
                              (N516)? out_me_data_i[269] : 
                              (N517)? out_me_data_i[301] : 
                              (N518)? out_me_data_i[333] : 1'b0;
  assign out_me_data_o[332] = (N508)? out_me_data_i_0__12_ : 
                              (N509)? out_me_data_i[44] : 
                              (N510)? out_me_data_i[76] : 
                              (N511)? out_me_data_i[108] : 
                              (N512)? out_me_data_i[140] : 
                              (N513)? out_me_data_i[172] : 
                              (N514)? out_me_data_i[204] : 
                              (N515)? out_me_data_i[236] : 
                              (N516)? out_me_data_i[268] : 
                              (N517)? out_me_data_i[300] : 
                              (N518)? out_me_data_i[332] : 1'b0;
  assign out_me_data_o[331] = (N508)? out_me_data_i_0__11_ : 
                              (N509)? out_me_data_i[43] : 
                              (N510)? out_me_data_i[75] : 
                              (N511)? out_me_data_i[107] : 
                              (N512)? out_me_data_i[139] : 
                              (N513)? out_me_data_i[171] : 
                              (N514)? out_me_data_i[203] : 
                              (N515)? out_me_data_i[235] : 
                              (N516)? out_me_data_i[267] : 
                              (N517)? out_me_data_i[299] : 
                              (N518)? out_me_data_i[331] : 1'b0;
  assign out_me_data_o[330] = (N508)? out_me_data_i_0__10_ : 
                              (N509)? out_me_data_i[42] : 
                              (N510)? out_me_data_i[74] : 
                              (N511)? out_me_data_i[106] : 
                              (N512)? out_me_data_i[138] : 
                              (N513)? out_me_data_i[170] : 
                              (N514)? out_me_data_i[202] : 
                              (N515)? out_me_data_i[234] : 
                              (N516)? out_me_data_i[266] : 
                              (N517)? out_me_data_i[298] : 
                              (N518)? out_me_data_i[330] : 1'b0;
  assign out_me_data_o[329] = (N508)? out_me_data_i_0__9_ : 
                              (N509)? out_me_data_i[41] : 
                              (N510)? out_me_data_i[73] : 
                              (N511)? out_me_data_i[105] : 
                              (N512)? out_me_data_i[137] : 
                              (N513)? out_me_data_i[169] : 
                              (N514)? out_me_data_i[201] : 
                              (N515)? out_me_data_i[233] : 
                              (N516)? out_me_data_i[265] : 
                              (N517)? out_me_data_i[297] : 
                              (N518)? out_me_data_i[329] : 1'b0;
  assign out_me_data_o[328] = (N508)? out_me_data_i_0__8_ : 
                              (N509)? out_me_data_i[40] : 
                              (N510)? out_me_data_i[72] : 
                              (N511)? out_me_data_i[104] : 
                              (N512)? out_me_data_i[136] : 
                              (N513)? out_me_data_i[168] : 
                              (N514)? out_me_data_i[200] : 
                              (N515)? out_me_data_i[232] : 
                              (N516)? out_me_data_i[264] : 
                              (N517)? out_me_data_i[296] : 
                              (N518)? out_me_data_i[328] : 1'b0;
  assign out_me_data_o[327] = (N508)? out_me_data_i_0__7_ : 
                              (N509)? out_me_data_i[39] : 
                              (N510)? out_me_data_i[71] : 
                              (N511)? out_me_data_i[103] : 
                              (N512)? out_me_data_i[135] : 
                              (N513)? out_me_data_i[167] : 
                              (N514)? out_me_data_i[199] : 
                              (N515)? out_me_data_i[231] : 
                              (N516)? out_me_data_i[263] : 
                              (N517)? out_me_data_i[295] : 
                              (N518)? out_me_data_i[327] : 1'b0;
  assign out_me_data_o[326] = (N508)? out_me_data_i_0__6_ : 
                              (N509)? out_me_data_i[38] : 
                              (N510)? out_me_data_i[70] : 
                              (N511)? out_me_data_i[102] : 
                              (N512)? out_me_data_i[134] : 
                              (N513)? out_me_data_i[166] : 
                              (N514)? out_me_data_i[198] : 
                              (N515)? out_me_data_i[230] : 
                              (N516)? out_me_data_i[262] : 
                              (N517)? out_me_data_i[294] : 
                              (N518)? out_me_data_i[326] : 1'b0;
  assign out_me_data_o[325] = (N508)? out_me_data_i_0__5_ : 
                              (N509)? out_me_data_i[37] : 
                              (N510)? out_me_data_i[69] : 
                              (N511)? out_me_data_i[101] : 
                              (N512)? out_me_data_i[133] : 
                              (N513)? out_me_data_i[165] : 
                              (N514)? out_me_data_i[197] : 
                              (N515)? out_me_data_i[229] : 
                              (N516)? out_me_data_i[261] : 
                              (N517)? out_me_data_i[293] : 
                              (N518)? out_me_data_i[325] : 1'b0;
  assign out_me_data_o[324] = (N508)? out_me_data_i_0__4_ : 
                              (N509)? out_me_data_i[36] : 
                              (N510)? out_me_data_i[68] : 
                              (N511)? out_me_data_i[100] : 
                              (N512)? out_me_data_i[132] : 
                              (N513)? out_me_data_i[164] : 
                              (N514)? out_me_data_i[196] : 
                              (N515)? out_me_data_i[228] : 
                              (N516)? out_me_data_i[260] : 
                              (N517)? out_me_data_i[292] : 
                              (N518)? out_me_data_i[324] : 1'b0;
  assign out_me_data_o[323] = (N508)? out_me_data_i_0__3_ : 
                              (N509)? out_me_data_i[35] : 
                              (N510)? out_me_data_i[67] : 
                              (N511)? out_me_data_i[99] : 
                              (N512)? out_me_data_i[131] : 
                              (N513)? out_me_data_i[163] : 
                              (N514)? out_me_data_i[195] : 
                              (N515)? out_me_data_i[227] : 
                              (N516)? out_me_data_i[259] : 
                              (N517)? out_me_data_i[291] : 
                              (N518)? out_me_data_i[323] : 1'b0;
  assign out_me_data_o[322] = (N508)? out_me_data_i_0__2_ : 
                              (N509)? out_me_data_i[34] : 
                              (N510)? out_me_data_i[66] : 
                              (N511)? out_me_data_i[98] : 
                              (N512)? out_me_data_i[130] : 
                              (N513)? out_me_data_i[162] : 
                              (N514)? out_me_data_i[194] : 
                              (N515)? out_me_data_i[226] : 
                              (N516)? out_me_data_i[258] : 
                              (N517)? out_me_data_i[290] : 
                              (N518)? out_me_data_i[322] : 1'b0;
  assign out_me_data_o[321] = (N508)? out_me_data_i_0__1_ : 
                              (N509)? out_me_data_i[33] : 
                              (N510)? out_me_data_i[65] : 
                              (N511)? out_me_data_i[97] : 
                              (N512)? out_me_data_i[129] : 
                              (N513)? out_me_data_i[161] : 
                              (N514)? out_me_data_i[193] : 
                              (N515)? out_me_data_i[225] : 
                              (N516)? out_me_data_i[257] : 
                              (N517)? out_me_data_i[289] : 
                              (N518)? out_me_data_i[321] : 1'b0;
  assign out_me_data_o[320] = (N508)? out_me_data_i_0__0_ : 
                              (N509)? out_me_data_i[32] : 
                              (N510)? out_me_data_i[64] : 
                              (N511)? out_me_data_i[96] : 
                              (N512)? out_me_data_i[128] : 
                              (N513)? out_me_data_i[160] : 
                              (N514)? out_me_data_i[192] : 
                              (N515)? out_me_data_i[224] : 
                              (N516)? out_me_data_i[256] : 
                              (N517)? out_me_data_i[288] : 
                              (N518)? out_me_data_i[320] : 1'b0;
  assign out_me_data_o[319] = (N519)? out_me_data_i_0__31_ : 
                              (N520)? out_me_data_i[63] : 
                              (N521)? out_me_data_i[95] : 
                              (N522)? out_me_data_i[127] : 
                              (N523)? out_me_data_i[159] : 
                              (N524)? out_me_data_i[191] : 
                              (N525)? out_me_data_i[223] : 
                              (N526)? out_me_data_i[255] : 
                              (N527)? out_me_data_i[287] : 
                              (N528)? out_me_data_i[319] : 1'b0;
  assign N519 = N1803;
  assign N520 = N1805;
  assign N521 = N1807;
  assign N522 = N1808;
  assign N523 = N1809;
  assign N524 = N1810;
  assign N525 = N1811;
  assign N526 = N1812;
  assign N527 = N1804;
  assign N528 = N1806;
  assign out_me_data_o[318] = (N519)? out_me_data_i_0__30_ : 
                              (N520)? out_me_data_i[62] : 
                              (N521)? out_me_data_i[94] : 
                              (N522)? out_me_data_i[126] : 
                              (N523)? out_me_data_i[158] : 
                              (N524)? out_me_data_i[190] : 
                              (N525)? out_me_data_i[222] : 
                              (N526)? out_me_data_i[254] : 
                              (N527)? out_me_data_i[286] : 
                              (N528)? out_me_data_i[318] : 1'b0;
  assign out_me_data_o[317] = (N519)? out_me_data_i_0__29_ : 
                              (N520)? out_me_data_i[61] : 
                              (N521)? out_me_data_i[93] : 
                              (N522)? out_me_data_i[125] : 
                              (N523)? out_me_data_i[157] : 
                              (N524)? out_me_data_i[189] : 
                              (N525)? out_me_data_i[221] : 
                              (N526)? out_me_data_i[253] : 
                              (N527)? out_me_data_i[285] : 
                              (N528)? out_me_data_i[317] : 1'b0;
  assign out_me_data_o[316] = (N519)? out_me_data_i_0__28_ : 
                              (N520)? out_me_data_i[60] : 
                              (N521)? out_me_data_i[92] : 
                              (N522)? out_me_data_i[124] : 
                              (N523)? out_me_data_i[156] : 
                              (N524)? out_me_data_i[188] : 
                              (N525)? out_me_data_i[220] : 
                              (N526)? out_me_data_i[252] : 
                              (N527)? out_me_data_i[284] : 
                              (N528)? out_me_data_i[316] : 1'b0;
  assign out_me_data_o[315] = (N519)? out_me_data_i_0__27_ : 
                              (N520)? out_me_data_i[59] : 
                              (N521)? out_me_data_i[91] : 
                              (N522)? out_me_data_i[123] : 
                              (N523)? out_me_data_i[155] : 
                              (N524)? out_me_data_i[187] : 
                              (N525)? out_me_data_i[219] : 
                              (N526)? out_me_data_i[251] : 
                              (N527)? out_me_data_i[283] : 
                              (N528)? out_me_data_i[315] : 1'b0;
  assign out_me_data_o[314] = (N519)? out_me_data_i_0__26_ : 
                              (N520)? out_me_data_i[58] : 
                              (N521)? out_me_data_i[90] : 
                              (N522)? out_me_data_i[122] : 
                              (N523)? out_me_data_i[154] : 
                              (N524)? out_me_data_i[186] : 
                              (N525)? out_me_data_i[218] : 
                              (N526)? out_me_data_i[250] : 
                              (N527)? out_me_data_i[282] : 
                              (N528)? out_me_data_i[314] : 1'b0;
  assign out_me_data_o[313] = (N519)? out_me_data_i_0__25_ : 
                              (N520)? out_me_data_i[57] : 
                              (N521)? out_me_data_i[89] : 
                              (N522)? out_me_data_i[121] : 
                              (N523)? out_me_data_i[153] : 
                              (N524)? out_me_data_i[185] : 
                              (N525)? out_me_data_i[217] : 
                              (N526)? out_me_data_i[249] : 
                              (N527)? out_me_data_i[281] : 
                              (N528)? out_me_data_i[313] : 1'b0;
  assign out_me_data_o[312] = (N519)? out_me_data_i_0__24_ : 
                              (N520)? out_me_data_i[56] : 
                              (N521)? out_me_data_i[88] : 
                              (N522)? out_me_data_i[120] : 
                              (N523)? out_me_data_i[152] : 
                              (N524)? out_me_data_i[184] : 
                              (N525)? out_me_data_i[216] : 
                              (N526)? out_me_data_i[248] : 
                              (N527)? out_me_data_i[280] : 
                              (N528)? out_me_data_i[312] : 1'b0;
  assign out_me_data_o[311] = (N519)? out_me_data_i_0__23_ : 
                              (N520)? out_me_data_i[55] : 
                              (N521)? out_me_data_i[87] : 
                              (N522)? out_me_data_i[119] : 
                              (N523)? out_me_data_i[151] : 
                              (N524)? out_me_data_i[183] : 
                              (N525)? out_me_data_i[215] : 
                              (N526)? out_me_data_i[247] : 
                              (N527)? out_me_data_i[279] : 
                              (N528)? out_me_data_i[311] : 1'b0;
  assign out_me_data_o[310] = (N519)? out_me_data_i_0__22_ : 
                              (N520)? out_me_data_i[54] : 
                              (N521)? out_me_data_i[86] : 
                              (N522)? out_me_data_i[118] : 
                              (N523)? out_me_data_i[150] : 
                              (N524)? out_me_data_i[182] : 
                              (N525)? out_me_data_i[214] : 
                              (N526)? out_me_data_i[246] : 
                              (N527)? out_me_data_i[278] : 
                              (N528)? out_me_data_i[310] : 1'b0;
  assign out_me_data_o[309] = (N519)? out_me_data_i_0__21_ : 
                              (N520)? out_me_data_i[53] : 
                              (N521)? out_me_data_i[85] : 
                              (N522)? out_me_data_i[117] : 
                              (N523)? out_me_data_i[149] : 
                              (N524)? out_me_data_i[181] : 
                              (N525)? out_me_data_i[213] : 
                              (N526)? out_me_data_i[245] : 
                              (N527)? out_me_data_i[277] : 
                              (N528)? out_me_data_i[309] : 1'b0;
  assign out_me_data_o[308] = (N519)? out_me_data_i_0__20_ : 
                              (N520)? out_me_data_i[52] : 
                              (N521)? out_me_data_i[84] : 
                              (N522)? out_me_data_i[116] : 
                              (N523)? out_me_data_i[148] : 
                              (N524)? out_me_data_i[180] : 
                              (N525)? out_me_data_i[212] : 
                              (N526)? out_me_data_i[244] : 
                              (N527)? out_me_data_i[276] : 
                              (N528)? out_me_data_i[308] : 1'b0;
  assign out_me_data_o[307] = (N519)? out_me_data_i_0__19_ : 
                              (N520)? out_me_data_i[51] : 
                              (N521)? out_me_data_i[83] : 
                              (N522)? out_me_data_i[115] : 
                              (N523)? out_me_data_i[147] : 
                              (N524)? out_me_data_i[179] : 
                              (N525)? out_me_data_i[211] : 
                              (N526)? out_me_data_i[243] : 
                              (N527)? out_me_data_i[275] : 
                              (N528)? out_me_data_i[307] : 1'b0;
  assign out_me_data_o[306] = (N519)? out_me_data_i_0__18_ : 
                              (N520)? out_me_data_i[50] : 
                              (N521)? out_me_data_i[82] : 
                              (N522)? out_me_data_i[114] : 
                              (N523)? out_me_data_i[146] : 
                              (N524)? out_me_data_i[178] : 
                              (N525)? out_me_data_i[210] : 
                              (N526)? out_me_data_i[242] : 
                              (N527)? out_me_data_i[274] : 
                              (N528)? out_me_data_i[306] : 1'b0;
  assign out_me_data_o[305] = (N519)? out_me_data_i_0__17_ : 
                              (N520)? out_me_data_i[49] : 
                              (N521)? out_me_data_i[81] : 
                              (N522)? out_me_data_i[113] : 
                              (N523)? out_me_data_i[145] : 
                              (N524)? out_me_data_i[177] : 
                              (N525)? out_me_data_i[209] : 
                              (N526)? out_me_data_i[241] : 
                              (N527)? out_me_data_i[273] : 
                              (N528)? out_me_data_i[305] : 1'b0;
  assign out_me_data_o[304] = (N519)? out_me_data_i_0__16_ : 
                              (N520)? out_me_data_i[48] : 
                              (N521)? out_me_data_i[80] : 
                              (N522)? out_me_data_i[112] : 
                              (N523)? out_me_data_i[144] : 
                              (N524)? out_me_data_i[176] : 
                              (N525)? out_me_data_i[208] : 
                              (N526)? out_me_data_i[240] : 
                              (N527)? out_me_data_i[272] : 
                              (N528)? out_me_data_i[304] : 1'b0;
  assign out_me_data_o[303] = (N519)? out_me_data_i_0__15_ : 
                              (N520)? out_me_data_i[47] : 
                              (N521)? out_me_data_i[79] : 
                              (N522)? out_me_data_i[111] : 
                              (N523)? out_me_data_i[143] : 
                              (N524)? out_me_data_i[175] : 
                              (N525)? out_me_data_i[207] : 
                              (N526)? out_me_data_i[239] : 
                              (N527)? out_me_data_i[271] : 
                              (N528)? out_me_data_i[303] : 1'b0;
  assign out_me_data_o[302] = (N519)? out_me_data_i_0__14_ : 
                              (N520)? out_me_data_i[46] : 
                              (N521)? out_me_data_i[78] : 
                              (N522)? out_me_data_i[110] : 
                              (N523)? out_me_data_i[142] : 
                              (N524)? out_me_data_i[174] : 
                              (N525)? out_me_data_i[206] : 
                              (N526)? out_me_data_i[238] : 
                              (N527)? out_me_data_i[270] : 
                              (N528)? out_me_data_i[302] : 1'b0;
  assign out_me_data_o[301] = (N519)? out_me_data_i_0__13_ : 
                              (N520)? out_me_data_i[45] : 
                              (N521)? out_me_data_i[77] : 
                              (N522)? out_me_data_i[109] : 
                              (N523)? out_me_data_i[141] : 
                              (N524)? out_me_data_i[173] : 
                              (N525)? out_me_data_i[205] : 
                              (N526)? out_me_data_i[237] : 
                              (N527)? out_me_data_i[269] : 
                              (N528)? out_me_data_i[301] : 1'b0;
  assign out_me_data_o[300] = (N519)? out_me_data_i_0__12_ : 
                              (N520)? out_me_data_i[44] : 
                              (N521)? out_me_data_i[76] : 
                              (N522)? out_me_data_i[108] : 
                              (N523)? out_me_data_i[140] : 
                              (N524)? out_me_data_i[172] : 
                              (N525)? out_me_data_i[204] : 
                              (N526)? out_me_data_i[236] : 
                              (N527)? out_me_data_i[268] : 
                              (N528)? out_me_data_i[300] : 1'b0;
  assign out_me_data_o[299] = (N519)? out_me_data_i_0__11_ : 
                              (N520)? out_me_data_i[43] : 
                              (N521)? out_me_data_i[75] : 
                              (N522)? out_me_data_i[107] : 
                              (N523)? out_me_data_i[139] : 
                              (N524)? out_me_data_i[171] : 
                              (N525)? out_me_data_i[203] : 
                              (N526)? out_me_data_i[235] : 
                              (N527)? out_me_data_i[267] : 
                              (N528)? out_me_data_i[299] : 1'b0;
  assign out_me_data_o[298] = (N519)? out_me_data_i_0__10_ : 
                              (N520)? out_me_data_i[42] : 
                              (N521)? out_me_data_i[74] : 
                              (N522)? out_me_data_i[106] : 
                              (N523)? out_me_data_i[138] : 
                              (N524)? out_me_data_i[170] : 
                              (N525)? out_me_data_i[202] : 
                              (N526)? out_me_data_i[234] : 
                              (N527)? out_me_data_i[266] : 
                              (N528)? out_me_data_i[298] : 1'b0;
  assign out_me_data_o[297] = (N519)? out_me_data_i_0__9_ : 
                              (N520)? out_me_data_i[41] : 
                              (N521)? out_me_data_i[73] : 
                              (N522)? out_me_data_i[105] : 
                              (N523)? out_me_data_i[137] : 
                              (N524)? out_me_data_i[169] : 
                              (N525)? out_me_data_i[201] : 
                              (N526)? out_me_data_i[233] : 
                              (N527)? out_me_data_i[265] : 
                              (N528)? out_me_data_i[297] : 1'b0;
  assign out_me_data_o[296] = (N519)? out_me_data_i_0__8_ : 
                              (N520)? out_me_data_i[40] : 
                              (N521)? out_me_data_i[72] : 
                              (N522)? out_me_data_i[104] : 
                              (N523)? out_me_data_i[136] : 
                              (N524)? out_me_data_i[168] : 
                              (N525)? out_me_data_i[200] : 
                              (N526)? out_me_data_i[232] : 
                              (N527)? out_me_data_i[264] : 
                              (N528)? out_me_data_i[296] : 1'b0;
  assign out_me_data_o[295] = (N519)? out_me_data_i_0__7_ : 
                              (N520)? out_me_data_i[39] : 
                              (N521)? out_me_data_i[71] : 
                              (N522)? out_me_data_i[103] : 
                              (N523)? out_me_data_i[135] : 
                              (N524)? out_me_data_i[167] : 
                              (N525)? out_me_data_i[199] : 
                              (N526)? out_me_data_i[231] : 
                              (N527)? out_me_data_i[263] : 
                              (N528)? out_me_data_i[295] : 1'b0;
  assign out_me_data_o[294] = (N519)? out_me_data_i_0__6_ : 
                              (N520)? out_me_data_i[38] : 
                              (N521)? out_me_data_i[70] : 
                              (N522)? out_me_data_i[102] : 
                              (N523)? out_me_data_i[134] : 
                              (N524)? out_me_data_i[166] : 
                              (N525)? out_me_data_i[198] : 
                              (N526)? out_me_data_i[230] : 
                              (N527)? out_me_data_i[262] : 
                              (N528)? out_me_data_i[294] : 1'b0;
  assign out_me_data_o[293] = (N519)? out_me_data_i_0__5_ : 
                              (N520)? out_me_data_i[37] : 
                              (N521)? out_me_data_i[69] : 
                              (N522)? out_me_data_i[101] : 
                              (N523)? out_me_data_i[133] : 
                              (N524)? out_me_data_i[165] : 
                              (N525)? out_me_data_i[197] : 
                              (N526)? out_me_data_i[229] : 
                              (N527)? out_me_data_i[261] : 
                              (N528)? out_me_data_i[293] : 1'b0;
  assign out_me_data_o[292] = (N519)? out_me_data_i_0__4_ : 
                              (N520)? out_me_data_i[36] : 
                              (N521)? out_me_data_i[68] : 
                              (N522)? out_me_data_i[100] : 
                              (N523)? out_me_data_i[132] : 
                              (N524)? out_me_data_i[164] : 
                              (N525)? out_me_data_i[196] : 
                              (N526)? out_me_data_i[228] : 
                              (N527)? out_me_data_i[260] : 
                              (N528)? out_me_data_i[292] : 1'b0;
  assign out_me_data_o[291] = (N519)? out_me_data_i_0__3_ : 
                              (N520)? out_me_data_i[35] : 
                              (N521)? out_me_data_i[67] : 
                              (N522)? out_me_data_i[99] : 
                              (N523)? out_me_data_i[131] : 
                              (N524)? out_me_data_i[163] : 
                              (N525)? out_me_data_i[195] : 
                              (N526)? out_me_data_i[227] : 
                              (N527)? out_me_data_i[259] : 
                              (N528)? out_me_data_i[291] : 1'b0;
  assign out_me_data_o[290] = (N519)? out_me_data_i_0__2_ : 
                              (N520)? out_me_data_i[34] : 
                              (N521)? out_me_data_i[66] : 
                              (N522)? out_me_data_i[98] : 
                              (N523)? out_me_data_i[130] : 
                              (N524)? out_me_data_i[162] : 
                              (N525)? out_me_data_i[194] : 
                              (N526)? out_me_data_i[226] : 
                              (N527)? out_me_data_i[258] : 
                              (N528)? out_me_data_i[290] : 1'b0;
  assign out_me_data_o[289] = (N519)? out_me_data_i_0__1_ : 
                              (N520)? out_me_data_i[33] : 
                              (N521)? out_me_data_i[65] : 
                              (N522)? out_me_data_i[97] : 
                              (N523)? out_me_data_i[129] : 
                              (N524)? out_me_data_i[161] : 
                              (N525)? out_me_data_i[193] : 
                              (N526)? out_me_data_i[225] : 
                              (N527)? out_me_data_i[257] : 
                              (N528)? out_me_data_i[289] : 1'b0;
  assign out_me_data_o[288] = (N519)? out_me_data_i_0__0_ : 
                              (N520)? out_me_data_i[32] : 
                              (N521)? out_me_data_i[64] : 
                              (N522)? out_me_data_i[96] : 
                              (N523)? out_me_data_i[128] : 
                              (N524)? out_me_data_i[160] : 
                              (N525)? out_me_data_i[192] : 
                              (N526)? out_me_data_i[224] : 
                              (N527)? out_me_data_i[256] : 
                              (N528)? out_me_data_i[288] : 1'b0;
  assign out_me_data_o[287] = (N529)? out_me_data_i_0__31_ : 
                              (N530)? out_me_data_i[63] : 
                              (N531)? out_me_data_i[95] : 
                              (N532)? out_me_data_i[127] : 
                              (N533)? out_me_data_i[159] : 
                              (N534)? out_me_data_i[191] : 
                              (N535)? out_me_data_i[223] : 
                              (N536)? out_me_data_i[255] : 
                              (N537)? out_me_data_i[287] : 1'b0;
  assign N529 = N1680;
  assign N530 = N1681;
  assign N531 = N1682;
  assign N532 = N1683;
  assign N533 = N1684;
  assign N534 = N1685;
  assign N535 = N1686;
  assign N536 = N1687;
  assign N537 = bk_dpath_sel_r[35];
  assign out_me_data_o[286] = (N529)? out_me_data_i_0__30_ : 
                              (N530)? out_me_data_i[62] : 
                              (N531)? out_me_data_i[94] : 
                              (N532)? out_me_data_i[126] : 
                              (N533)? out_me_data_i[158] : 
                              (N534)? out_me_data_i[190] : 
                              (N535)? out_me_data_i[222] : 
                              (N536)? out_me_data_i[254] : 
                              (N537)? out_me_data_i[286] : 1'b0;
  assign out_me_data_o[285] = (N529)? out_me_data_i_0__29_ : 
                              (N530)? out_me_data_i[61] : 
                              (N531)? out_me_data_i[93] : 
                              (N532)? out_me_data_i[125] : 
                              (N533)? out_me_data_i[157] : 
                              (N534)? out_me_data_i[189] : 
                              (N535)? out_me_data_i[221] : 
                              (N536)? out_me_data_i[253] : 
                              (N537)? out_me_data_i[285] : 1'b0;
  assign out_me_data_o[284] = (N529)? out_me_data_i_0__28_ : 
                              (N530)? out_me_data_i[60] : 
                              (N531)? out_me_data_i[92] : 
                              (N532)? out_me_data_i[124] : 
                              (N533)? out_me_data_i[156] : 
                              (N534)? out_me_data_i[188] : 
                              (N535)? out_me_data_i[220] : 
                              (N536)? out_me_data_i[252] : 
                              (N537)? out_me_data_i[284] : 1'b0;
  assign out_me_data_o[283] = (N529)? out_me_data_i_0__27_ : 
                              (N530)? out_me_data_i[59] : 
                              (N531)? out_me_data_i[91] : 
                              (N532)? out_me_data_i[123] : 
                              (N533)? out_me_data_i[155] : 
                              (N534)? out_me_data_i[187] : 
                              (N535)? out_me_data_i[219] : 
                              (N536)? out_me_data_i[251] : 
                              (N537)? out_me_data_i[283] : 1'b0;
  assign out_me_data_o[282] = (N529)? out_me_data_i_0__26_ : 
                              (N530)? out_me_data_i[58] : 
                              (N531)? out_me_data_i[90] : 
                              (N532)? out_me_data_i[122] : 
                              (N533)? out_me_data_i[154] : 
                              (N534)? out_me_data_i[186] : 
                              (N535)? out_me_data_i[218] : 
                              (N536)? out_me_data_i[250] : 
                              (N537)? out_me_data_i[282] : 1'b0;
  assign out_me_data_o[281] = (N529)? out_me_data_i_0__25_ : 
                              (N530)? out_me_data_i[57] : 
                              (N531)? out_me_data_i[89] : 
                              (N532)? out_me_data_i[121] : 
                              (N533)? out_me_data_i[153] : 
                              (N534)? out_me_data_i[185] : 
                              (N535)? out_me_data_i[217] : 
                              (N536)? out_me_data_i[249] : 
                              (N537)? out_me_data_i[281] : 1'b0;
  assign out_me_data_o[280] = (N529)? out_me_data_i_0__24_ : 
                              (N530)? out_me_data_i[56] : 
                              (N531)? out_me_data_i[88] : 
                              (N532)? out_me_data_i[120] : 
                              (N533)? out_me_data_i[152] : 
                              (N534)? out_me_data_i[184] : 
                              (N535)? out_me_data_i[216] : 
                              (N536)? out_me_data_i[248] : 
                              (N537)? out_me_data_i[280] : 1'b0;
  assign out_me_data_o[279] = (N529)? out_me_data_i_0__23_ : 
                              (N530)? out_me_data_i[55] : 
                              (N531)? out_me_data_i[87] : 
                              (N532)? out_me_data_i[119] : 
                              (N533)? out_me_data_i[151] : 
                              (N534)? out_me_data_i[183] : 
                              (N535)? out_me_data_i[215] : 
                              (N536)? out_me_data_i[247] : 
                              (N537)? out_me_data_i[279] : 1'b0;
  assign out_me_data_o[278] = (N529)? out_me_data_i_0__22_ : 
                              (N530)? out_me_data_i[54] : 
                              (N531)? out_me_data_i[86] : 
                              (N532)? out_me_data_i[118] : 
                              (N533)? out_me_data_i[150] : 
                              (N534)? out_me_data_i[182] : 
                              (N535)? out_me_data_i[214] : 
                              (N536)? out_me_data_i[246] : 
                              (N537)? out_me_data_i[278] : 1'b0;
  assign out_me_data_o[277] = (N529)? out_me_data_i_0__21_ : 
                              (N530)? out_me_data_i[53] : 
                              (N531)? out_me_data_i[85] : 
                              (N532)? out_me_data_i[117] : 
                              (N533)? out_me_data_i[149] : 
                              (N534)? out_me_data_i[181] : 
                              (N535)? out_me_data_i[213] : 
                              (N536)? out_me_data_i[245] : 
                              (N537)? out_me_data_i[277] : 1'b0;
  assign out_me_data_o[276] = (N529)? out_me_data_i_0__20_ : 
                              (N530)? out_me_data_i[52] : 
                              (N531)? out_me_data_i[84] : 
                              (N532)? out_me_data_i[116] : 
                              (N533)? out_me_data_i[148] : 
                              (N534)? out_me_data_i[180] : 
                              (N535)? out_me_data_i[212] : 
                              (N536)? out_me_data_i[244] : 
                              (N537)? out_me_data_i[276] : 1'b0;
  assign out_me_data_o[275] = (N529)? out_me_data_i_0__19_ : 
                              (N530)? out_me_data_i[51] : 
                              (N531)? out_me_data_i[83] : 
                              (N532)? out_me_data_i[115] : 
                              (N533)? out_me_data_i[147] : 
                              (N534)? out_me_data_i[179] : 
                              (N535)? out_me_data_i[211] : 
                              (N536)? out_me_data_i[243] : 
                              (N537)? out_me_data_i[275] : 1'b0;
  assign out_me_data_o[274] = (N529)? out_me_data_i_0__18_ : 
                              (N530)? out_me_data_i[50] : 
                              (N531)? out_me_data_i[82] : 
                              (N532)? out_me_data_i[114] : 
                              (N533)? out_me_data_i[146] : 
                              (N534)? out_me_data_i[178] : 
                              (N535)? out_me_data_i[210] : 
                              (N536)? out_me_data_i[242] : 
                              (N537)? out_me_data_i[274] : 1'b0;
  assign out_me_data_o[273] = (N529)? out_me_data_i_0__17_ : 
                              (N530)? out_me_data_i[49] : 
                              (N531)? out_me_data_i[81] : 
                              (N532)? out_me_data_i[113] : 
                              (N533)? out_me_data_i[145] : 
                              (N534)? out_me_data_i[177] : 
                              (N535)? out_me_data_i[209] : 
                              (N536)? out_me_data_i[241] : 
                              (N537)? out_me_data_i[273] : 1'b0;
  assign out_me_data_o[272] = (N529)? out_me_data_i_0__16_ : 
                              (N530)? out_me_data_i[48] : 
                              (N531)? out_me_data_i[80] : 
                              (N532)? out_me_data_i[112] : 
                              (N533)? out_me_data_i[144] : 
                              (N534)? out_me_data_i[176] : 
                              (N535)? out_me_data_i[208] : 
                              (N536)? out_me_data_i[240] : 
                              (N537)? out_me_data_i[272] : 1'b0;
  assign out_me_data_o[271] = (N529)? out_me_data_i_0__15_ : 
                              (N530)? out_me_data_i[47] : 
                              (N531)? out_me_data_i[79] : 
                              (N532)? out_me_data_i[111] : 
                              (N533)? out_me_data_i[143] : 
                              (N534)? out_me_data_i[175] : 
                              (N535)? out_me_data_i[207] : 
                              (N536)? out_me_data_i[239] : 
                              (N537)? out_me_data_i[271] : 1'b0;
  assign out_me_data_o[270] = (N529)? out_me_data_i_0__14_ : 
                              (N530)? out_me_data_i[46] : 
                              (N531)? out_me_data_i[78] : 
                              (N532)? out_me_data_i[110] : 
                              (N533)? out_me_data_i[142] : 
                              (N534)? out_me_data_i[174] : 
                              (N535)? out_me_data_i[206] : 
                              (N536)? out_me_data_i[238] : 
                              (N537)? out_me_data_i[270] : 1'b0;
  assign out_me_data_o[269] = (N529)? out_me_data_i_0__13_ : 
                              (N530)? out_me_data_i[45] : 
                              (N531)? out_me_data_i[77] : 
                              (N532)? out_me_data_i[109] : 
                              (N533)? out_me_data_i[141] : 
                              (N534)? out_me_data_i[173] : 
                              (N535)? out_me_data_i[205] : 
                              (N536)? out_me_data_i[237] : 
                              (N537)? out_me_data_i[269] : 1'b0;
  assign out_me_data_o[268] = (N529)? out_me_data_i_0__12_ : 
                              (N530)? out_me_data_i[44] : 
                              (N531)? out_me_data_i[76] : 
                              (N532)? out_me_data_i[108] : 
                              (N533)? out_me_data_i[140] : 
                              (N534)? out_me_data_i[172] : 
                              (N535)? out_me_data_i[204] : 
                              (N536)? out_me_data_i[236] : 
                              (N537)? out_me_data_i[268] : 1'b0;
  assign out_me_data_o[267] = (N529)? out_me_data_i_0__11_ : 
                              (N530)? out_me_data_i[43] : 
                              (N531)? out_me_data_i[75] : 
                              (N532)? out_me_data_i[107] : 
                              (N533)? out_me_data_i[139] : 
                              (N534)? out_me_data_i[171] : 
                              (N535)? out_me_data_i[203] : 
                              (N536)? out_me_data_i[235] : 
                              (N537)? out_me_data_i[267] : 1'b0;
  assign out_me_data_o[266] = (N529)? out_me_data_i_0__10_ : 
                              (N530)? out_me_data_i[42] : 
                              (N531)? out_me_data_i[74] : 
                              (N532)? out_me_data_i[106] : 
                              (N533)? out_me_data_i[138] : 
                              (N534)? out_me_data_i[170] : 
                              (N535)? out_me_data_i[202] : 
                              (N536)? out_me_data_i[234] : 
                              (N537)? out_me_data_i[266] : 1'b0;
  assign out_me_data_o[265] = (N529)? out_me_data_i_0__9_ : 
                              (N530)? out_me_data_i[41] : 
                              (N531)? out_me_data_i[73] : 
                              (N532)? out_me_data_i[105] : 
                              (N533)? out_me_data_i[137] : 
                              (N534)? out_me_data_i[169] : 
                              (N535)? out_me_data_i[201] : 
                              (N536)? out_me_data_i[233] : 
                              (N537)? out_me_data_i[265] : 1'b0;
  assign out_me_data_o[264] = (N529)? out_me_data_i_0__8_ : 
                              (N530)? out_me_data_i[40] : 
                              (N531)? out_me_data_i[72] : 
                              (N532)? out_me_data_i[104] : 
                              (N533)? out_me_data_i[136] : 
                              (N534)? out_me_data_i[168] : 
                              (N535)? out_me_data_i[200] : 
                              (N536)? out_me_data_i[232] : 
                              (N537)? out_me_data_i[264] : 1'b0;
  assign out_me_data_o[263] = (N529)? out_me_data_i_0__7_ : 
                              (N530)? out_me_data_i[39] : 
                              (N531)? out_me_data_i[71] : 
                              (N532)? out_me_data_i[103] : 
                              (N533)? out_me_data_i[135] : 
                              (N534)? out_me_data_i[167] : 
                              (N535)? out_me_data_i[199] : 
                              (N536)? out_me_data_i[231] : 
                              (N537)? out_me_data_i[263] : 1'b0;
  assign out_me_data_o[262] = (N529)? out_me_data_i_0__6_ : 
                              (N530)? out_me_data_i[38] : 
                              (N531)? out_me_data_i[70] : 
                              (N532)? out_me_data_i[102] : 
                              (N533)? out_me_data_i[134] : 
                              (N534)? out_me_data_i[166] : 
                              (N535)? out_me_data_i[198] : 
                              (N536)? out_me_data_i[230] : 
                              (N537)? out_me_data_i[262] : 1'b0;
  assign out_me_data_o[261] = (N529)? out_me_data_i_0__5_ : 
                              (N530)? out_me_data_i[37] : 
                              (N531)? out_me_data_i[69] : 
                              (N532)? out_me_data_i[101] : 
                              (N533)? out_me_data_i[133] : 
                              (N534)? out_me_data_i[165] : 
                              (N535)? out_me_data_i[197] : 
                              (N536)? out_me_data_i[229] : 
                              (N537)? out_me_data_i[261] : 1'b0;
  assign out_me_data_o[260] = (N529)? out_me_data_i_0__4_ : 
                              (N530)? out_me_data_i[36] : 
                              (N531)? out_me_data_i[68] : 
                              (N532)? out_me_data_i[100] : 
                              (N533)? out_me_data_i[132] : 
                              (N534)? out_me_data_i[164] : 
                              (N535)? out_me_data_i[196] : 
                              (N536)? out_me_data_i[228] : 
                              (N537)? out_me_data_i[260] : 1'b0;
  assign out_me_data_o[259] = (N529)? out_me_data_i_0__3_ : 
                              (N530)? out_me_data_i[35] : 
                              (N531)? out_me_data_i[67] : 
                              (N532)? out_me_data_i[99] : 
                              (N533)? out_me_data_i[131] : 
                              (N534)? out_me_data_i[163] : 
                              (N535)? out_me_data_i[195] : 
                              (N536)? out_me_data_i[227] : 
                              (N537)? out_me_data_i[259] : 1'b0;
  assign out_me_data_o[258] = (N529)? out_me_data_i_0__2_ : 
                              (N530)? out_me_data_i[34] : 
                              (N531)? out_me_data_i[66] : 
                              (N532)? out_me_data_i[98] : 
                              (N533)? out_me_data_i[130] : 
                              (N534)? out_me_data_i[162] : 
                              (N535)? out_me_data_i[194] : 
                              (N536)? out_me_data_i[226] : 
                              (N537)? out_me_data_i[258] : 1'b0;
  assign out_me_data_o[257] = (N529)? out_me_data_i_0__1_ : 
                              (N530)? out_me_data_i[33] : 
                              (N531)? out_me_data_i[65] : 
                              (N532)? out_me_data_i[97] : 
                              (N533)? out_me_data_i[129] : 
                              (N534)? out_me_data_i[161] : 
                              (N535)? out_me_data_i[193] : 
                              (N536)? out_me_data_i[225] : 
                              (N537)? out_me_data_i[257] : 1'b0;
  assign out_me_data_o[256] = (N529)? out_me_data_i_0__0_ : 
                              (N530)? out_me_data_i[32] : 
                              (N531)? out_me_data_i[64] : 
                              (N532)? out_me_data_i[96] : 
                              (N533)? out_me_data_i[128] : 
                              (N534)? out_me_data_i[160] : 
                              (N535)? out_me_data_i[192] : 
                              (N536)? out_me_data_i[224] : 
                              (N537)? out_me_data_i[256] : 1'b0;
  assign in_v_o[0] = N2604 | N2605;
  assign N2604 = N2602 | N2603;
  assign N2602 = N2600 | N2601;
  assign N2600 = N2598 | N2599;
  assign N2598 = N2596 | N2597;
  assign N2596 = N2594 | N2595;
  assign N2594 = N2592 | N2593;
  assign N2592 = N2590 | N2591;
  assign N2590 = N2588 | N2589;
  assign N2588 = N2586 | N2587;
  assign N2586 = N2584 | N2585;
  assign N2584 = N2582 | N2583;
  assign N2582 = N2580 | N2581;
  assign N2580 = N2578 | N2579;
  assign N2578 = N2576 | N2577;
  assign N2576 = in_v_i[15] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__15_ ;
  assign N2577 = in_v_i[14] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__14_ ;
  assign N2579 = in_v_i[13] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__13_ ;
  assign N2581 = in_v_i[12] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__12_ ;
  assign N2583 = in_v_i[11] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__11_ ;
  assign N2585 = in_v_i[10] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__10_ ;
  assign N2587 = in_v_i[9] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__9_ ;
  assign N2589 = in_v_i[8] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__8_ ;
  assign N2591 = in_v_i[7] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__7_ ;
  assign N2593 = in_v_i[6] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__6_ ;
  assign N2595 = in_v_i[5] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__5_ ;
  assign N2597 = in_v_i[4] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__4_ ;
  assign N2599 = in_v_i[3] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__3_ ;
  assign N2601 = in_v_i[2] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__2_ ;
  assign N2603 = in_v_i[1] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__1_ ;
  assign N2605 = in_v_i[0] & \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__0_ ;
  assign N554 = ~bk_sel_r[0];
  assign N555 = ~bk_sel_r[1];
  assign N556 = N554 & N555;
  assign N557 = N554 & bk_sel_r[1];
  assign N558 = bk_sel_r[0] & N555;
  assign N559 = bk_sel_r[0] & bk_sel_r[1];
  assign N560 = ~bk_sel_r[2];
  assign N561 = N556 & N560;
  assign N562 = N556 & bk_sel_r[2];
  assign N563 = N558 & N560;
  assign N564 = N558 & bk_sel_r[2];
  assign N565 = N557 & N560;
  assign N566 = N557 & bk_sel_r[2];
  assign N567 = N559 & N560;
  assign N568 = N559 & bk_sel_r[2];
  assign N569 = ~bk_sel_r[3];
  assign N570 = N561 & N569;
  assign N571 = N561 & bk_sel_r[3];
  assign N572 = N563 & N569;
  assign N573 = N563 & bk_sel_r[3];
  assign N574 = N565 & N569;
  assign N575 = N565 & bk_sel_r[3];
  assign N576 = N567 & N569;
  assign N577 = N567 & bk_sel_r[3];
  assign N578 = N562 & N569;
  assign N579 = N562 & bk_sel_r[3];
  assign N580 = N564 & N569;
  assign N581 = N564 & bk_sel_r[3];
  assign N582 = N566 & N569;
  assign N583 = N566 & bk_sel_r[3];
  assign N584 = N568 & N569;
  assign N585 = N568 & bk_sel_r[3];
  assign N586 = ~fwd_dpath_sel_r[0];
  assign N587 = ~fwd_dpath_sel_r[1];
  assign N588 = N586 & N587;
  assign N589 = N586 & fwd_dpath_sel_r[1];
  assign N590 = fwd_dpath_sel_r[0] & N587;
  assign N591 = fwd_dpath_sel_r[0] & fwd_dpath_sel_r[1];
  assign N592 = ~fwd_dpath_sel_r[2];
  assign N593 = N588 & N592;
  assign N594 = N588 & fwd_dpath_sel_r[2];
  assign N595 = N590 & N592;
  assign N596 = N590 & fwd_dpath_sel_r[2];
  assign N597 = N589 & N592;
  assign N598 = N589 & fwd_dpath_sel_r[2];
  assign N599 = N591 & N592;
  assign N600 = N591 & fwd_dpath_sel_r[2];
  assign N601 = ~fwd_dpath_sel_r[3];
  assign N602 = N593 & N601;
  assign N603 = N593 & fwd_dpath_sel_r[3];
  assign N604 = N595 & N601;
  assign N605 = N595 & fwd_dpath_sel_r[3];
  assign N606 = N597 & N601;
  assign N607 = N597 & fwd_dpath_sel_r[3];
  assign N608 = N599 & N601;
  assign N609 = N599 & fwd_dpath_sel_r[3];
  assign N610 = N594 & N601;
  assign N611 = N594 & fwd_dpath_sel_r[3];
  assign N612 = N596 & N601;
  assign N613 = N596 & fwd_dpath_sel_r[3];
  assign N614 = N598 & N601;
  assign N615 = N598 & fwd_dpath_sel_r[3];
  assign N616 = N600 & N601;
  assign N617 = N600 & fwd_dpath_sel_r[3];
  assign N618 = N554 & N555;
  assign N619 = N554 & bk_sel_r[1];
  assign N620 = bk_sel_r[0] & N555;
  assign N621 = bk_sel_r[0] & bk_sel_r[1];
  assign N622 = N618 & N560;
  assign N623 = N618 & bk_sel_r[2];
  assign N624 = N620 & N560;
  assign N625 = N620 & bk_sel_r[2];
  assign N626 = N619 & N560;
  assign N627 = N619 & bk_sel_r[2];
  assign N628 = N621 & N560;
  assign N629 = N621 & bk_sel_r[2];
  assign N630 = N622 & N569;
  assign N631 = N622 & bk_sel_r[3];
  assign N632 = N624 & N569;
  assign N633 = N624 & bk_sel_r[3];
  assign N634 = N626 & N569;
  assign N635 = N626 & bk_sel_r[3];
  assign N636 = N628 & N569;
  assign N637 = N628 & bk_sel_r[3];
  assign N638 = N623 & N569;
  assign N639 = N623 & bk_sel_r[3];
  assign N640 = N625 & N569;
  assign N641 = N625 & bk_sel_r[3];
  assign N642 = N627 & N569;
  assign N643 = N627 & bk_sel_r[3];
  assign N644 = N629 & N569;
  assign N645 = N629 & bk_sel_r[3];
  assign N646 = ~fwd_sel_r[0];
  assign N647 = ~fwd_sel_r[1];
  assign N648 = N646 & N647;
  assign N649 = N646 & fwd_sel_r[1];
  assign N650 = fwd_sel_r[0] & N647;
  assign N651 = fwd_sel_r[0] & fwd_sel_r[1];
  assign N652 = ~fwd_sel_r[2];
  assign N653 = N648 & N652;
  assign N654 = N648 & fwd_sel_r[2];
  assign N655 = N650 & N652;
  assign N656 = N650 & fwd_sel_r[2];
  assign N657 = N649 & N652;
  assign N658 = N649 & fwd_sel_r[2];
  assign N659 = N651 & N652;
  assign N660 = N651 & fwd_sel_r[2];
  assign N661 = ~fwd_sel_r[3];
  assign N662 = N653 & N661;
  assign N663 = N653 & fwd_sel_r[3];
  assign N664 = N655 & N661;
  assign N665 = N655 & fwd_sel_r[3];
  assign N666 = N657 & N661;
  assign N667 = N657 & fwd_sel_r[3];
  assign N668 = N659 & N661;
  assign N669 = N659 & fwd_sel_r[3];
  assign N670 = N654 & N661;
  assign N671 = N654 & fwd_sel_r[3];
  assign N672 = N656 & N661;
  assign N673 = N656 & fwd_sel_r[3];
  assign N674 = N658 & N661;
  assign N675 = N658 & fwd_sel_r[3];
  assign N676 = N660 & N661;
  assign N677 = N660 & fwd_sel_r[3];
  assign in_v_o[1] = N2634 | N2635;
  assign N2634 = N2632 | N2633;
  assign N2632 = N2630 | N2631;
  assign N2630 = N2628 | N2629;
  assign N2628 = N2626 | N2627;
  assign N2626 = N2624 | N2625;
  assign N2624 = N2622 | N2623;
  assign N2622 = N2620 | N2621;
  assign N2620 = N2618 | N2619;
  assign N2618 = N2616 | N2617;
  assign N2616 = N2614 | N2615;
  assign N2614 = N2612 | N2613;
  assign N2612 = N2610 | N2611;
  assign N2610 = N2608 | N2609;
  assign N2608 = N2606 | N2607;
  assign N2606 = in_v_i[15] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__15_ ;
  assign N2607 = in_v_i[14] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__14_ ;
  assign N2609 = in_v_i[13] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__13_ ;
  assign N2611 = in_v_i[12] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__12_ ;
  assign N2613 = in_v_i[11] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__11_ ;
  assign N2615 = in_v_i[10] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__10_ ;
  assign N2617 = in_v_i[9] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__9_ ;
  assign N2619 = in_v_i[8] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__8_ ;
  assign N2621 = in_v_i[7] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__7_ ;
  assign N2623 = in_v_i[6] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__6_ ;
  assign N2625 = in_v_i[5] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__5_ ;
  assign N2627 = in_v_i[4] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__4_ ;
  assign N2629 = in_v_i[3] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__3_ ;
  assign N2631 = in_v_i[2] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__2_ ;
  assign N2633 = in_v_i[1] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__1_ ;
  assign N2635 = in_v_i[0] & \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__0_ ;
  assign N694 = ~bk_sel_r[4];
  assign N695 = ~bk_sel_r[5];
  assign N696 = N694 & N695;
  assign N697 = N694 & bk_sel_r[5];
  assign N698 = bk_sel_r[4] & N695;
  assign N699 = bk_sel_r[4] & bk_sel_r[5];
  assign N700 = ~bk_sel_r[6];
  assign N701 = N696 & N700;
  assign N702 = N696 & bk_sel_r[6];
  assign N703 = N698 & N700;
  assign N704 = N698 & bk_sel_r[6];
  assign N705 = N697 & N700;
  assign N706 = N697 & bk_sel_r[6];
  assign N707 = N699 & N700;
  assign N708 = N699 & bk_sel_r[6];
  assign N709 = ~bk_sel_r[7];
  assign N710 = N701 & N709;
  assign N711 = N701 & bk_sel_r[7];
  assign N712 = N703 & N709;
  assign N713 = N703 & bk_sel_r[7];
  assign N714 = N705 & N709;
  assign N715 = N705 & bk_sel_r[7];
  assign N716 = N707 & N709;
  assign N717 = N707 & bk_sel_r[7];
  assign N718 = N702 & N709;
  assign N719 = N702 & bk_sel_r[7];
  assign N720 = N704 & N709;
  assign N721 = N704 & bk_sel_r[7];
  assign N722 = N706 & N709;
  assign N723 = N706 & bk_sel_r[7];
  assign N724 = N708 & N709;
  assign N725 = N708 & bk_sel_r[7];
  assign N741 = N694 & N695;
  assign N742 = N694 & bk_sel_r[5];
  assign N743 = bk_sel_r[4] & N695;
  assign N744 = bk_sel_r[4] & bk_sel_r[5];
  assign N745 = N741 & N700;
  assign N746 = N741 & bk_sel_r[6];
  assign N747 = N743 & N700;
  assign N748 = N743 & bk_sel_r[6];
  assign N749 = N742 & N700;
  assign N750 = N742 & bk_sel_r[6];
  assign N751 = N744 & N700;
  assign N752 = N744 & bk_sel_r[6];
  assign N753 = N745 & N709;
  assign N754 = N745 & bk_sel_r[7];
  assign N755 = N747 & N709;
  assign N756 = N747 & bk_sel_r[7];
  assign N757 = N749 & N709;
  assign N758 = N749 & bk_sel_r[7];
  assign N759 = N751 & N709;
  assign N760 = N751 & bk_sel_r[7];
  assign N761 = N746 & N709;
  assign N762 = N746 & bk_sel_r[7];
  assign N763 = N748 & N709;
  assign N764 = N748 & bk_sel_r[7];
  assign N765 = N750 & N709;
  assign N766 = N750 & bk_sel_r[7];
  assign N767 = N752 & N709;
  assign N768 = N752 & bk_sel_r[7];
  assign N769 = ~fwd_sel_r[4];
  assign N770 = ~fwd_sel_r[5];
  assign N771 = N769 & N770;
  assign N772 = N769 & fwd_sel_r[5];
  assign N773 = fwd_sel_r[4] & N770;
  assign N774 = fwd_sel_r[4] & fwd_sel_r[5];
  assign N775 = ~fwd_sel_r[6];
  assign N776 = N771 & N775;
  assign N777 = N771 & fwd_sel_r[6];
  assign N778 = N773 & N775;
  assign N779 = N773 & fwd_sel_r[6];
  assign N780 = N772 & N775;
  assign N781 = N772 & fwd_sel_r[6];
  assign N782 = N774 & N775;
  assign N783 = N774 & fwd_sel_r[6];
  assign N784 = ~fwd_sel_r[7];
  assign N785 = N776 & N784;
  assign N786 = N776 & fwd_sel_r[7];
  assign N787 = N778 & N784;
  assign N788 = N778 & fwd_sel_r[7];
  assign N789 = N780 & N784;
  assign N790 = N780 & fwd_sel_r[7];
  assign N791 = N782 & N784;
  assign N792 = N782 & fwd_sel_r[7];
  assign N793 = N777 & N784;
  assign N794 = N777 & fwd_sel_r[7];
  assign N795 = N779 & N784;
  assign N796 = N779 & fwd_sel_r[7];
  assign N797 = N781 & N784;
  assign N798 = N781 & fwd_sel_r[7];
  assign N799 = N783 & N784;
  assign N800 = N783 & fwd_sel_r[7];
  assign N801 = ~bk_dpath_sel_r_4;
  assign in_v_o[2] = N2664 | N2665;
  assign N2664 = N2662 | N2663;
  assign N2662 = N2660 | N2661;
  assign N2660 = N2658 | N2659;
  assign N2658 = N2656 | N2657;
  assign N2656 = N2654 | N2655;
  assign N2654 = N2652 | N2653;
  assign N2652 = N2650 | N2651;
  assign N2650 = N2648 | N2649;
  assign N2648 = N2646 | N2647;
  assign N2646 = N2644 | N2645;
  assign N2644 = N2642 | N2643;
  assign N2642 = N2640 | N2641;
  assign N2640 = N2638 | N2639;
  assign N2638 = N2636 | N2637;
  assign N2636 = in_v_i[15] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__15_ ;
  assign N2637 = in_v_i[14] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__14_ ;
  assign N2639 = in_v_i[13] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__13_ ;
  assign N2641 = in_v_i[12] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__12_ ;
  assign N2643 = in_v_i[11] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__11_ ;
  assign N2645 = in_v_i[10] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__10_ ;
  assign N2647 = in_v_i[9] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__9_ ;
  assign N2649 = in_v_i[8] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__8_ ;
  assign N2651 = in_v_i[7] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__7_ ;
  assign N2653 = in_v_i[6] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__6_ ;
  assign N2655 = in_v_i[5] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__5_ ;
  assign N2657 = in_v_i[4] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__4_ ;
  assign N2659 = in_v_i[3] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__3_ ;
  assign N2661 = in_v_i[2] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__2_ ;
  assign N2663 = in_v_i[1] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__1_ ;
  assign N2665 = in_v_i[0] & \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__0_ ;
  assign N818 = ~bk_sel_r[8];
  assign N819 = ~bk_sel_r[9];
  assign N820 = N818 & N819;
  assign N821 = N818 & bk_sel_r[9];
  assign N822 = bk_sel_r[8] & N819;
  assign N823 = bk_sel_r[8] & bk_sel_r[9];
  assign N824 = ~bk_sel_r[10];
  assign N825 = N820 & N824;
  assign N826 = N820 & bk_sel_r[10];
  assign N827 = N822 & N824;
  assign N828 = N822 & bk_sel_r[10];
  assign N829 = N821 & N824;
  assign N830 = N821 & bk_sel_r[10];
  assign N831 = N823 & N824;
  assign N832 = N823 & bk_sel_r[10];
  assign N833 = ~bk_sel_r[11];
  assign N834 = N825 & N833;
  assign N835 = N825 & bk_sel_r[11];
  assign N836 = N827 & N833;
  assign N837 = N827 & bk_sel_r[11];
  assign N838 = N829 & N833;
  assign N839 = N829 & bk_sel_r[11];
  assign N840 = N831 & N833;
  assign N841 = N831 & bk_sel_r[11];
  assign N842 = N826 & N833;
  assign N843 = N826 & bk_sel_r[11];
  assign N844 = N828 & N833;
  assign N845 = N828 & bk_sel_r[11];
  assign N846 = N830 & N833;
  assign N847 = N830 & bk_sel_r[11];
  assign N848 = N832 & N833;
  assign N849 = N832 & bk_sel_r[11];
  assign N864 = N818 & N819;
  assign N865 = N818 & bk_sel_r[9];
  assign N866 = bk_sel_r[8] & N819;
  assign N867 = bk_sel_r[8] & bk_sel_r[9];
  assign N868 = N864 & N824;
  assign N869 = N864 & bk_sel_r[10];
  assign N870 = N866 & N824;
  assign N871 = N866 & bk_sel_r[10];
  assign N872 = N865 & N824;
  assign N873 = N865 & bk_sel_r[10];
  assign N874 = N867 & N824;
  assign N875 = N867 & bk_sel_r[10];
  assign N876 = N868 & N833;
  assign N877 = N868 & bk_sel_r[11];
  assign N878 = N870 & N833;
  assign N879 = N870 & bk_sel_r[11];
  assign N880 = N872 & N833;
  assign N881 = N872 & bk_sel_r[11];
  assign N882 = N874 & N833;
  assign N883 = N874 & bk_sel_r[11];
  assign N884 = N869 & N833;
  assign N885 = N869 & bk_sel_r[11];
  assign N886 = N871 & N833;
  assign N887 = N871 & bk_sel_r[11];
  assign N888 = N873 & N833;
  assign N889 = N873 & bk_sel_r[11];
  assign N890 = N875 & N833;
  assign N891 = N875 & bk_sel_r[11];
  assign N892 = ~fwd_sel_r[8];
  assign N893 = ~fwd_sel_r[9];
  assign N894 = N892 & N893;
  assign N895 = N892 & fwd_sel_r[9];
  assign N896 = fwd_sel_r[8] & N893;
  assign N897 = fwd_sel_r[8] & fwd_sel_r[9];
  assign N898 = ~fwd_sel_r[10];
  assign N899 = N894 & N898;
  assign N900 = N894 & fwd_sel_r[10];
  assign N901 = N896 & N898;
  assign N902 = N896 & fwd_sel_r[10];
  assign N903 = N895 & N898;
  assign N904 = N895 & fwd_sel_r[10];
  assign N905 = N897 & N898;
  assign N906 = N897 & fwd_sel_r[10];
  assign N907 = ~fwd_sel_r[11];
  assign N908 = N899 & N907;
  assign N909 = N899 & fwd_sel_r[11];
  assign N910 = N901 & N907;
  assign N911 = N901 & fwd_sel_r[11];
  assign N912 = N903 & N907;
  assign N913 = N903 & fwd_sel_r[11];
  assign N914 = N905 & N907;
  assign N915 = N905 & fwd_sel_r[11];
  assign N916 = N900 & N907;
  assign N917 = N900 & fwd_sel_r[11];
  assign N918 = N902 & N907;
  assign N919 = N902 & fwd_sel_r[11];
  assign N920 = N904 & N907;
  assign N921 = N904 & fwd_sel_r[11];
  assign N922 = N906 & N907;
  assign N923 = N906 & fwd_sel_r[11];
  assign in_v_o[3] = N2694 | N2695;
  assign N2694 = N2692 | N2693;
  assign N2692 = N2690 | N2691;
  assign N2690 = N2688 | N2689;
  assign N2688 = N2686 | N2687;
  assign N2686 = N2684 | N2685;
  assign N2684 = N2682 | N2683;
  assign N2682 = N2680 | N2681;
  assign N2680 = N2678 | N2679;
  assign N2678 = N2676 | N2677;
  assign N2676 = N2674 | N2675;
  assign N2674 = N2672 | N2673;
  assign N2672 = N2670 | N2671;
  assign N2670 = N2668 | N2669;
  assign N2668 = N2666 | N2667;
  assign N2666 = in_v_i[15] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__15_ ;
  assign N2667 = in_v_i[14] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__14_ ;
  assign N2669 = in_v_i[13] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__13_ ;
  assign N2671 = in_v_i[12] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__12_ ;
  assign N2673 = in_v_i[11] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__11_ ;
  assign N2675 = in_v_i[10] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__10_ ;
  assign N2677 = in_v_i[9] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__9_ ;
  assign N2679 = in_v_i[8] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__8_ ;
  assign N2681 = in_v_i[7] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__7_ ;
  assign N2683 = in_v_i[6] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__6_ ;
  assign N2685 = in_v_i[5] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__5_ ;
  assign N2687 = in_v_i[4] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__4_ ;
  assign N2689 = in_v_i[3] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__3_ ;
  assign N2691 = in_v_i[2] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__2_ ;
  assign N2693 = in_v_i[1] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__1_ ;
  assign N2695 = in_v_i[0] & \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__0_ ;
  assign N941 = ~bk_sel_r[12];
  assign N942 = ~bk_sel_r[13];
  assign N943 = N941 & N942;
  assign N944 = N941 & bk_sel_r[13];
  assign N945 = bk_sel_r[12] & N942;
  assign N946 = bk_sel_r[12] & bk_sel_r[13];
  assign N947 = ~bk_sel_r[14];
  assign N948 = N943 & N947;
  assign N949 = N943 & bk_sel_r[14];
  assign N950 = N945 & N947;
  assign N951 = N945 & bk_sel_r[14];
  assign N952 = N944 & N947;
  assign N953 = N944 & bk_sel_r[14];
  assign N954 = N946 & N947;
  assign N955 = N946 & bk_sel_r[14];
  assign N956 = ~bk_sel_r[15];
  assign N957 = N948 & N956;
  assign N958 = N948 & bk_sel_r[15];
  assign N959 = N950 & N956;
  assign N960 = N950 & bk_sel_r[15];
  assign N961 = N952 & N956;
  assign N962 = N952 & bk_sel_r[15];
  assign N963 = N954 & N956;
  assign N964 = N954 & bk_sel_r[15];
  assign N965 = N949 & N956;
  assign N966 = N949 & bk_sel_r[15];
  assign N967 = N951 & N956;
  assign N968 = N951 & bk_sel_r[15];
  assign N969 = N953 & N956;
  assign N970 = N953 & bk_sel_r[15];
  assign N971 = N955 & N956;
  assign N972 = N955 & bk_sel_r[15];
  assign N986 = N941 & N942;
  assign N987 = N941 & bk_sel_r[13];
  assign N988 = bk_sel_r[12] & N942;
  assign N989 = bk_sel_r[12] & bk_sel_r[13];
  assign N990 = N986 & N947;
  assign N991 = N986 & bk_sel_r[14];
  assign N992 = N988 & N947;
  assign N993 = N988 & bk_sel_r[14];
  assign N994 = N987 & N947;
  assign N995 = N987 & bk_sel_r[14];
  assign N996 = N989 & N947;
  assign N997 = N989 & bk_sel_r[14];
  assign N998 = N990 & N956;
  assign N999 = N990 & bk_sel_r[15];
  assign N1000 = N992 & N956;
  assign N1001 = N992 & bk_sel_r[15];
  assign N1002 = N994 & N956;
  assign N1003 = N994 & bk_sel_r[15];
  assign N1004 = N996 & N956;
  assign N1005 = N996 & bk_sel_r[15];
  assign N1006 = N991 & N956;
  assign N1007 = N991 & bk_sel_r[15];
  assign N1008 = N993 & N956;
  assign N1009 = N993 & bk_sel_r[15];
  assign N1010 = N995 & N956;
  assign N1011 = N995 & bk_sel_r[15];
  assign N1012 = N997 & N956;
  assign N1013 = N997 & bk_sel_r[15];
  assign N1014 = ~fwd_sel_r[12];
  assign N1015 = ~fwd_sel_r[13];
  assign N1016 = N1014 & N1015;
  assign N1017 = N1014 & fwd_sel_r[13];
  assign N1018 = fwd_sel_r[12] & N1015;
  assign N1019 = fwd_sel_r[12] & fwd_sel_r[13];
  assign N1020 = ~fwd_sel_r[14];
  assign N1021 = N1016 & N1020;
  assign N1022 = N1016 & fwd_sel_r[14];
  assign N1023 = N1018 & N1020;
  assign N1024 = N1018 & fwd_sel_r[14];
  assign N1025 = N1017 & N1020;
  assign N1026 = N1017 & fwd_sel_r[14];
  assign N1027 = N1019 & N1020;
  assign N1028 = N1019 & fwd_sel_r[14];
  assign N1029 = ~fwd_sel_r[15];
  assign N1030 = N1021 & N1029;
  assign N1031 = N1021 & fwd_sel_r[15];
  assign N1032 = N1023 & N1029;
  assign N1033 = N1023 & fwd_sel_r[15];
  assign N1034 = N1025 & N1029;
  assign N1035 = N1025 & fwd_sel_r[15];
  assign N1036 = N1027 & N1029;
  assign N1037 = N1027 & fwd_sel_r[15];
  assign N1038 = N1022 & N1029;
  assign N1039 = N1022 & fwd_sel_r[15];
  assign N1040 = N1024 & N1029;
  assign N1041 = N1024 & fwd_sel_r[15];
  assign N1042 = N1026 & N1029;
  assign N1043 = N1026 & fwd_sel_r[15];
  assign N1044 = N1028 & N1029;
  assign N1045 = N1028 & fwd_sel_r[15];
  assign N1046 = ~bk_dpath_sel_r_12;
  assign N1047 = ~bk_dpath_sel_r_13;
  assign N1048 = N1046 & N1047;
  assign N1049 = N1046 & bk_dpath_sel_r_13;
  assign N1050 = bk_dpath_sel_r_12 & N1047;
  assign N1051 = bk_dpath_sel_r_12 & bk_dpath_sel_r_13;
  assign in_v_o[4] = N2724 | N2725;
  assign N2724 = N2722 | N2723;
  assign N2722 = N2720 | N2721;
  assign N2720 = N2718 | N2719;
  assign N2718 = N2716 | N2717;
  assign N2716 = N2714 | N2715;
  assign N2714 = N2712 | N2713;
  assign N2712 = N2710 | N2711;
  assign N2710 = N2708 | N2709;
  assign N2708 = N2706 | N2707;
  assign N2706 = N2704 | N2705;
  assign N2704 = N2702 | N2703;
  assign N2702 = N2700 | N2701;
  assign N2700 = N2698 | N2699;
  assign N2698 = N2696 | N2697;
  assign N2696 = in_v_i[15] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__15_ ;
  assign N2697 = in_v_i[14] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__14_ ;
  assign N2699 = in_v_i[13] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__13_ ;
  assign N2701 = in_v_i[12] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__12_ ;
  assign N2703 = in_v_i[11] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__11_ ;
  assign N2705 = in_v_i[10] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__10_ ;
  assign N2707 = in_v_i[9] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__9_ ;
  assign N2709 = in_v_i[8] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__8_ ;
  assign N2711 = in_v_i[7] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__7_ ;
  assign N2713 = in_v_i[6] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__6_ ;
  assign N2715 = in_v_i[5] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__5_ ;
  assign N2717 = in_v_i[4] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__4_ ;
  assign N2719 = in_v_i[3] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__3_ ;
  assign N2721 = in_v_i[2] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__2_ ;
  assign N2723 = in_v_i[1] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__1_ ;
  assign N2725 = in_v_i[0] & \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__0_ ;
  assign N1068 = ~bk_sel_r[16];
  assign N1069 = ~bk_sel_r[17];
  assign N1070 = N1068 & N1069;
  assign N1071 = N1068 & bk_sel_r[17];
  assign N1072 = bk_sel_r[16] & N1069;
  assign N1073 = bk_sel_r[16] & bk_sel_r[17];
  assign N1074 = ~bk_sel_r[18];
  assign N1075 = N1070 & N1074;
  assign N1076 = N1070 & bk_sel_r[18];
  assign N1077 = N1072 & N1074;
  assign N1078 = N1072 & bk_sel_r[18];
  assign N1079 = N1071 & N1074;
  assign N1080 = N1071 & bk_sel_r[18];
  assign N1081 = N1073 & N1074;
  assign N1082 = N1073 & bk_sel_r[18];
  assign N1083 = ~bk_sel_r[19];
  assign N1084 = N1075 & N1083;
  assign N1085 = N1075 & bk_sel_r[19];
  assign N1086 = N1077 & N1083;
  assign N1087 = N1077 & bk_sel_r[19];
  assign N1088 = N1079 & N1083;
  assign N1089 = N1079 & bk_sel_r[19];
  assign N1090 = N1081 & N1083;
  assign N1091 = N1081 & bk_sel_r[19];
  assign N1092 = N1076 & N1083;
  assign N1093 = N1076 & bk_sel_r[19];
  assign N1094 = N1078 & N1083;
  assign N1095 = N1078 & bk_sel_r[19];
  assign N1096 = N1080 & N1083;
  assign N1097 = N1080 & bk_sel_r[19];
  assign N1098 = N1082 & N1083;
  assign N1099 = N1082 & bk_sel_r[19];
  assign N1112 = N1068 & N1069;
  assign N1113 = N1068 & bk_sel_r[17];
  assign N1114 = bk_sel_r[16] & N1069;
  assign N1115 = bk_sel_r[16] & bk_sel_r[17];
  assign N1116 = N1112 & N1074;
  assign N1117 = N1112 & bk_sel_r[18];
  assign N1118 = N1114 & N1074;
  assign N1119 = N1114 & bk_sel_r[18];
  assign N1120 = N1113 & N1074;
  assign N1121 = N1113 & bk_sel_r[18];
  assign N1122 = N1115 & N1074;
  assign N1123 = N1115 & bk_sel_r[18];
  assign N1124 = N1116 & N1083;
  assign N1125 = N1116 & bk_sel_r[19];
  assign N1126 = N1118 & N1083;
  assign N1127 = N1118 & bk_sel_r[19];
  assign N1128 = N1120 & N1083;
  assign N1129 = N1120 & bk_sel_r[19];
  assign N1130 = N1122 & N1083;
  assign N1131 = N1122 & bk_sel_r[19];
  assign N1132 = N1117 & N1083;
  assign N1133 = N1117 & bk_sel_r[19];
  assign N1134 = N1119 & N1083;
  assign N1135 = N1119 & bk_sel_r[19];
  assign N1136 = N1121 & N1083;
  assign N1137 = N1121 & bk_sel_r[19];
  assign N1138 = N1123 & N1083;
  assign N1139 = N1123 & bk_sel_r[19];
  assign N1140 = ~fwd_sel_r[16];
  assign N1141 = ~fwd_sel_r[17];
  assign N1142 = N1140 & N1141;
  assign N1143 = N1140 & fwd_sel_r[17];
  assign N1144 = fwd_sel_r[16] & N1141;
  assign N1145 = fwd_sel_r[16] & fwd_sel_r[17];
  assign N1146 = ~fwd_sel_r[18];
  assign N1147 = N1142 & N1146;
  assign N1148 = N1142 & fwd_sel_r[18];
  assign N1149 = N1144 & N1146;
  assign N1150 = N1144 & fwd_sel_r[18];
  assign N1151 = N1143 & N1146;
  assign N1152 = N1143 & fwd_sel_r[18];
  assign N1153 = N1145 & N1146;
  assign N1154 = N1145 & fwd_sel_r[18];
  assign N1155 = ~fwd_sel_r[19];
  assign N1156 = N1147 & N1155;
  assign N1157 = N1147 & fwd_sel_r[19];
  assign N1158 = N1149 & N1155;
  assign N1159 = N1149 & fwd_sel_r[19];
  assign N1160 = N1151 & N1155;
  assign N1161 = N1151 & fwd_sel_r[19];
  assign N1162 = N1153 & N1155;
  assign N1163 = N1153 & fwd_sel_r[19];
  assign N1164 = N1148 & N1155;
  assign N1165 = N1148 & fwd_sel_r[19];
  assign N1166 = N1150 & N1155;
  assign N1167 = N1150 & fwd_sel_r[19];
  assign N1168 = N1152 & N1155;
  assign N1169 = N1152 & fwd_sel_r[19];
  assign N1170 = N1154 & N1155;
  assign N1171 = N1154 & fwd_sel_r[19];
  assign in_v_o[5] = N2754 | N2755;
  assign N2754 = N2752 | N2753;
  assign N2752 = N2750 | N2751;
  assign N2750 = N2748 | N2749;
  assign N2748 = N2746 | N2747;
  assign N2746 = N2744 | N2745;
  assign N2744 = N2742 | N2743;
  assign N2742 = N2740 | N2741;
  assign N2740 = N2738 | N2739;
  assign N2738 = N2736 | N2737;
  assign N2736 = N2734 | N2735;
  assign N2734 = N2732 | N2733;
  assign N2732 = N2730 | N2731;
  assign N2730 = N2728 | N2729;
  assign N2728 = N2726 | N2727;
  assign N2726 = in_v_i[15] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__15_ ;
  assign N2727 = in_v_i[14] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__14_ ;
  assign N2729 = in_v_i[13] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__13_ ;
  assign N2731 = in_v_i[12] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__12_ ;
  assign N2733 = in_v_i[11] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__11_ ;
  assign N2735 = in_v_i[10] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__10_ ;
  assign N2737 = in_v_i[9] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__9_ ;
  assign N2739 = in_v_i[8] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__8_ ;
  assign N2741 = in_v_i[7] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__7_ ;
  assign N2743 = in_v_i[6] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__6_ ;
  assign N2745 = in_v_i[5] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__5_ ;
  assign N2747 = in_v_i[4] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__4_ ;
  assign N2749 = in_v_i[3] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__3_ ;
  assign N2751 = in_v_i[2] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__2_ ;
  assign N2753 = in_v_i[1] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__1_ ;
  assign N2755 = in_v_i[0] & \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__0_ ;
  assign N1192 = ~bk_sel_r[20];
  assign N1193 = ~bk_sel_r[21];
  assign N1194 = N1192 & N1193;
  assign N1195 = N1192 & bk_sel_r[21];
  assign N1196 = bk_sel_r[20] & N1193;
  assign N1197 = bk_sel_r[20] & bk_sel_r[21];
  assign N1198 = ~bk_sel_r[22];
  assign N1199 = N1194 & N1198;
  assign N1200 = N1194 & bk_sel_r[22];
  assign N1201 = N1196 & N1198;
  assign N1202 = N1196 & bk_sel_r[22];
  assign N1203 = N1195 & N1198;
  assign N1204 = N1195 & bk_sel_r[22];
  assign N1205 = N1197 & N1198;
  assign N1206 = N1197 & bk_sel_r[22];
  assign N1207 = ~bk_sel_r[23];
  assign N1208 = N1199 & N1207;
  assign N1209 = N1199 & bk_sel_r[23];
  assign N1210 = N1201 & N1207;
  assign N1211 = N1201 & bk_sel_r[23];
  assign N1212 = N1203 & N1207;
  assign N1213 = N1203 & bk_sel_r[23];
  assign N1214 = N1205 & N1207;
  assign N1215 = N1205 & bk_sel_r[23];
  assign N1216 = N1200 & N1207;
  assign N1217 = N1200 & bk_sel_r[23];
  assign N1218 = N1202 & N1207;
  assign N1219 = N1202 & bk_sel_r[23];
  assign N1220 = N1204 & N1207;
  assign N1221 = N1204 & bk_sel_r[23];
  assign N1222 = N1206 & N1207;
  assign N1223 = N1206 & bk_sel_r[23];
  assign N1235 = N1192 & N1193;
  assign N1236 = N1192 & bk_sel_r[21];
  assign N1237 = bk_sel_r[20] & N1193;
  assign N1238 = bk_sel_r[20] & bk_sel_r[21];
  assign N1239 = N1235 & N1198;
  assign N1240 = N1235 & bk_sel_r[22];
  assign N1241 = N1237 & N1198;
  assign N1242 = N1237 & bk_sel_r[22];
  assign N1243 = N1236 & N1198;
  assign N1244 = N1236 & bk_sel_r[22];
  assign N1245 = N1238 & N1198;
  assign N1246 = N1238 & bk_sel_r[22];
  assign N1247 = N1239 & N1207;
  assign N1248 = N1239 & bk_sel_r[23];
  assign N1249 = N1241 & N1207;
  assign N1250 = N1241 & bk_sel_r[23];
  assign N1251 = N1243 & N1207;
  assign N1252 = N1243 & bk_sel_r[23];
  assign N1253 = N1245 & N1207;
  assign N1254 = N1245 & bk_sel_r[23];
  assign N1255 = N1240 & N1207;
  assign N1256 = N1240 & bk_sel_r[23];
  assign N1257 = N1242 & N1207;
  assign N1258 = N1242 & bk_sel_r[23];
  assign N1259 = N1244 & N1207;
  assign N1260 = N1244 & bk_sel_r[23];
  assign N1261 = N1246 & N1207;
  assign N1262 = N1246 & bk_sel_r[23];
  assign N1263 = ~fwd_sel_r[20];
  assign N1264 = ~fwd_sel_r[21];
  assign N1265 = N1263 & N1264;
  assign N1266 = N1263 & fwd_sel_r[21];
  assign N1267 = fwd_sel_r[20] & N1264;
  assign N1268 = fwd_sel_r[20] & fwd_sel_r[21];
  assign N1269 = ~fwd_sel_r[22];
  assign N1270 = N1265 & N1269;
  assign N1271 = N1265 & fwd_sel_r[22];
  assign N1272 = N1267 & N1269;
  assign N1273 = N1267 & fwd_sel_r[22];
  assign N1274 = N1266 & N1269;
  assign N1275 = N1266 & fwd_sel_r[22];
  assign N1276 = N1268 & N1269;
  assign N1277 = N1268 & fwd_sel_r[22];
  assign N1278 = ~fwd_sel_r[23];
  assign N1279 = N1270 & N1278;
  assign N1280 = N1270 & fwd_sel_r[23];
  assign N1281 = N1272 & N1278;
  assign N1282 = N1272 & fwd_sel_r[23];
  assign N1283 = N1274 & N1278;
  assign N1284 = N1274 & fwd_sel_r[23];
  assign N1285 = N1276 & N1278;
  assign N1286 = N1276 & fwd_sel_r[23];
  assign N1287 = N1271 & N1278;
  assign N1288 = N1271 & fwd_sel_r[23];
  assign N1289 = N1273 & N1278;
  assign N1290 = N1273 & fwd_sel_r[23];
  assign N1291 = N1275 & N1278;
  assign N1292 = N1275 & fwd_sel_r[23];
  assign N1293 = N1277 & N1278;
  assign N1294 = N1277 & fwd_sel_r[23];
  assign in_v_o[6] = N2784 | N2785;
  assign N2784 = N2782 | N2783;
  assign N2782 = N2780 | N2781;
  assign N2780 = N2778 | N2779;
  assign N2778 = N2776 | N2777;
  assign N2776 = N2774 | N2775;
  assign N2774 = N2772 | N2773;
  assign N2772 = N2770 | N2771;
  assign N2770 = N2768 | N2769;
  assign N2768 = N2766 | N2767;
  assign N2766 = N2764 | N2765;
  assign N2764 = N2762 | N2763;
  assign N2762 = N2760 | N2761;
  assign N2760 = N2758 | N2759;
  assign N2758 = N2756 | N2757;
  assign N2756 = in_v_i[15] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__15_ ;
  assign N2757 = in_v_i[14] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__14_ ;
  assign N2759 = in_v_i[13] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__13_ ;
  assign N2761 = in_v_i[12] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__12_ ;
  assign N2763 = in_v_i[11] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__11_ ;
  assign N2765 = in_v_i[10] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__10_ ;
  assign N2767 = in_v_i[9] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__9_ ;
  assign N2769 = in_v_i[8] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__8_ ;
  assign N2771 = in_v_i[7] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__7_ ;
  assign N2773 = in_v_i[6] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__6_ ;
  assign N2775 = in_v_i[5] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__5_ ;
  assign N2777 = in_v_i[4] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__4_ ;
  assign N2779 = in_v_i[3] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__3_ ;
  assign N2781 = in_v_i[2] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__2_ ;
  assign N2783 = in_v_i[1] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__1_ ;
  assign N2785 = in_v_i[0] & \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__0_ ;
  assign N1317 = ~bk_sel_r[24];
  assign N1318 = ~bk_sel_r[25];
  assign N1319 = N1317 & N1318;
  assign N1320 = N1317 & bk_sel_r[25];
  assign N1321 = bk_sel_r[24] & N1318;
  assign N1322 = bk_sel_r[24] & bk_sel_r[25];
  assign N1323 = ~bk_sel_r[26];
  assign N1324 = N1319 & N1323;
  assign N1325 = N1319 & bk_sel_r[26];
  assign N1326 = N1321 & N1323;
  assign N1327 = N1321 & bk_sel_r[26];
  assign N1328 = N1320 & N1323;
  assign N1329 = N1320 & bk_sel_r[26];
  assign N1330 = N1322 & N1323;
  assign N1331 = N1322 & bk_sel_r[26];
  assign N1332 = ~bk_sel_r[27];
  assign N1333 = N1324 & N1332;
  assign N1334 = N1324 & bk_sel_r[27];
  assign N1335 = N1326 & N1332;
  assign N1336 = N1326 & bk_sel_r[27];
  assign N1337 = N1328 & N1332;
  assign N1338 = N1328 & bk_sel_r[27];
  assign N1339 = N1330 & N1332;
  assign N1340 = N1330 & bk_sel_r[27];
  assign N1341 = N1325 & N1332;
  assign N1342 = N1325 & bk_sel_r[27];
  assign N1343 = N1327 & N1332;
  assign N1344 = N1327 & bk_sel_r[27];
  assign N1345 = N1329 & N1332;
  assign N1346 = N1329 & bk_sel_r[27];
  assign N1347 = N1331 & N1332;
  assign N1348 = N1331 & bk_sel_r[27];
  assign N1359 = N1317 & N1318;
  assign N1360 = N1317 & bk_sel_r[25];
  assign N1361 = bk_sel_r[24] & N1318;
  assign N1362 = bk_sel_r[24] & bk_sel_r[25];
  assign N1363 = N1359 & N1323;
  assign N1364 = N1359 & bk_sel_r[26];
  assign N1365 = N1361 & N1323;
  assign N1366 = N1361 & bk_sel_r[26];
  assign N1367 = N1360 & N1323;
  assign N1368 = N1360 & bk_sel_r[26];
  assign N1369 = N1362 & N1323;
  assign N1370 = N1362 & bk_sel_r[26];
  assign N1371 = N1363 & N1332;
  assign N1372 = N1363 & bk_sel_r[27];
  assign N1373 = N1365 & N1332;
  assign N1374 = N1365 & bk_sel_r[27];
  assign N1375 = N1367 & N1332;
  assign N1376 = N1367 & bk_sel_r[27];
  assign N1377 = N1369 & N1332;
  assign N1378 = N1369 & bk_sel_r[27];
  assign N1379 = N1364 & N1332;
  assign N1380 = N1364 & bk_sel_r[27];
  assign N1381 = N1366 & N1332;
  assign N1382 = N1366 & bk_sel_r[27];
  assign N1383 = N1368 & N1332;
  assign N1384 = N1368 & bk_sel_r[27];
  assign N1385 = N1370 & N1332;
  assign N1386 = N1370 & bk_sel_r[27];
  assign N1387 = ~fwd_sel_r[24];
  assign N1388 = ~fwd_sel_r[25];
  assign N1389 = N1387 & N1388;
  assign N1390 = N1387 & fwd_sel_r[25];
  assign N1391 = fwd_sel_r[24] & N1388;
  assign N1392 = fwd_sel_r[24] & fwd_sel_r[25];
  assign N1393 = ~fwd_sel_r[26];
  assign N1394 = N1389 & N1393;
  assign N1395 = N1389 & fwd_sel_r[26];
  assign N1396 = N1391 & N1393;
  assign N1397 = N1391 & fwd_sel_r[26];
  assign N1398 = N1390 & N1393;
  assign N1399 = N1390 & fwd_sel_r[26];
  assign N1400 = N1392 & N1393;
  assign N1401 = N1392 & fwd_sel_r[26];
  assign N1402 = ~fwd_sel_r[27];
  assign N1403 = N1394 & N1402;
  assign N1404 = N1394 & fwd_sel_r[27];
  assign N1405 = N1396 & N1402;
  assign N1406 = N1396 & fwd_sel_r[27];
  assign N1407 = N1398 & N1402;
  assign N1408 = N1398 & fwd_sel_r[27];
  assign N1409 = N1400 & N1402;
  assign N1410 = N1400 & fwd_sel_r[27];
  assign N1411 = N1395 & N1402;
  assign N1412 = N1395 & fwd_sel_r[27];
  assign N1413 = N1397 & N1402;
  assign N1414 = N1397 & fwd_sel_r[27];
  assign N1415 = N1399 & N1402;
  assign N1416 = N1399 & fwd_sel_r[27];
  assign N1417 = N1401 & N1402;
  assign N1418 = N1401 & fwd_sel_r[27];
  assign in_v_o[7] = N2814 | N2815;
  assign N2814 = N2812 | N2813;
  assign N2812 = N2810 | N2811;
  assign N2810 = N2808 | N2809;
  assign N2808 = N2806 | N2807;
  assign N2806 = N2804 | N2805;
  assign N2804 = N2802 | N2803;
  assign N2802 = N2800 | N2801;
  assign N2800 = N2798 | N2799;
  assign N2798 = N2796 | N2797;
  assign N2796 = N2794 | N2795;
  assign N2794 = N2792 | N2793;
  assign N2792 = N2790 | N2791;
  assign N2790 = N2788 | N2789;
  assign N2788 = N2786 | N2787;
  assign N2786 = in_v_i[15] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__15_ ;
  assign N2787 = in_v_i[14] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__14_ ;
  assign N2789 = in_v_i[13] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__13_ ;
  assign N2791 = in_v_i[12] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__12_ ;
  assign N2793 = in_v_i[11] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__11_ ;
  assign N2795 = in_v_i[10] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__10_ ;
  assign N2797 = in_v_i[9] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__9_ ;
  assign N2799 = in_v_i[8] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__8_ ;
  assign N2801 = in_v_i[7] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__7_ ;
  assign N2803 = in_v_i[6] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__6_ ;
  assign N2805 = in_v_i[5] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__5_ ;
  assign N2807 = in_v_i[4] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__4_ ;
  assign N2809 = in_v_i[3] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__3_ ;
  assign N2811 = in_v_i[2] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__2_ ;
  assign N2813 = in_v_i[1] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__1_ ;
  assign N2815 = in_v_i[0] & \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__0_ ;
  assign N1442 = ~bk_sel_r[28];
  assign N1443 = ~bk_sel_r[29];
  assign N1444 = N1442 & N1443;
  assign N1445 = N1442 & bk_sel_r[29];
  assign N1446 = bk_sel_r[28] & N1443;
  assign N1447 = bk_sel_r[28] & bk_sel_r[29];
  assign N1448 = ~bk_sel_r[30];
  assign N1449 = N1444 & N1448;
  assign N1450 = N1444 & bk_sel_r[30];
  assign N1451 = N1446 & N1448;
  assign N1452 = N1446 & bk_sel_r[30];
  assign N1453 = N1445 & N1448;
  assign N1454 = N1445 & bk_sel_r[30];
  assign N1455 = N1447 & N1448;
  assign N1456 = N1447 & bk_sel_r[30];
  assign N1457 = ~bk_sel_r[31];
  assign N1458 = N1449 & N1457;
  assign N1459 = N1449 & bk_sel_r[31];
  assign N1460 = N1451 & N1457;
  assign N1461 = N1451 & bk_sel_r[31];
  assign N1462 = N1453 & N1457;
  assign N1463 = N1453 & bk_sel_r[31];
  assign N1464 = N1455 & N1457;
  assign N1465 = N1455 & bk_sel_r[31];
  assign N1466 = N1450 & N1457;
  assign N1467 = N1450 & bk_sel_r[31];
  assign N1468 = N1452 & N1457;
  assign N1469 = N1452 & bk_sel_r[31];
  assign N1470 = N1454 & N1457;
  assign N1471 = N1454 & bk_sel_r[31];
  assign N1472 = N1456 & N1457;
  assign N1473 = N1456 & bk_sel_r[31];
  assign N1482 = N1442 & N1443;
  assign N1483 = N1442 & bk_sel_r[29];
  assign N1484 = bk_sel_r[28] & N1443;
  assign N1485 = bk_sel_r[28] & bk_sel_r[29];
  assign N1486 = N1482 & N1448;
  assign N1487 = N1482 & bk_sel_r[30];
  assign N1488 = N1484 & N1448;
  assign N1489 = N1484 & bk_sel_r[30];
  assign N1490 = N1483 & N1448;
  assign N1491 = N1483 & bk_sel_r[30];
  assign N1492 = N1485 & N1448;
  assign N1493 = N1485 & bk_sel_r[30];
  assign N1494 = N1486 & N1457;
  assign N1495 = N1486 & bk_sel_r[31];
  assign N1496 = N1488 & N1457;
  assign N1497 = N1488 & bk_sel_r[31];
  assign N1498 = N1490 & N1457;
  assign N1499 = N1490 & bk_sel_r[31];
  assign N1500 = N1492 & N1457;
  assign N1501 = N1492 & bk_sel_r[31];
  assign N1502 = N1487 & N1457;
  assign N1503 = N1487 & bk_sel_r[31];
  assign N1504 = N1489 & N1457;
  assign N1505 = N1489 & bk_sel_r[31];
  assign N1506 = N1491 & N1457;
  assign N1507 = N1491 & bk_sel_r[31];
  assign N1508 = N1493 & N1457;
  assign N1509 = N1493 & bk_sel_r[31];
  assign N1510 = ~fwd_sel_r[28];
  assign N1511 = ~fwd_sel_r[29];
  assign N1512 = N1510 & N1511;
  assign N1513 = N1510 & fwd_sel_r[29];
  assign N1514 = fwd_sel_r[28] & N1511;
  assign N1515 = fwd_sel_r[28] & fwd_sel_r[29];
  assign N1516 = ~fwd_sel_r[30];
  assign N1517 = N1512 & N1516;
  assign N1518 = N1512 & fwd_sel_r[30];
  assign N1519 = N1514 & N1516;
  assign N1520 = N1514 & fwd_sel_r[30];
  assign N1521 = N1513 & N1516;
  assign N1522 = N1513 & fwd_sel_r[30];
  assign N1523 = N1515 & N1516;
  assign N1524 = N1515 & fwd_sel_r[30];
  assign N1525 = ~fwd_sel_r[31];
  assign N1526 = N1517 & N1525;
  assign N1527 = N1517 & fwd_sel_r[31];
  assign N1528 = N1519 & N1525;
  assign N1529 = N1519 & fwd_sel_r[31];
  assign N1530 = N1521 & N1525;
  assign N1531 = N1521 & fwd_sel_r[31];
  assign N1532 = N1523 & N1525;
  assign N1533 = N1523 & fwd_sel_r[31];
  assign N1534 = N1518 & N1525;
  assign N1535 = N1518 & fwd_sel_r[31];
  assign N1536 = N1520 & N1525;
  assign N1537 = N1520 & fwd_sel_r[31];
  assign N1538 = N1522 & N1525;
  assign N1539 = N1522 & fwd_sel_r[31];
  assign N1540 = N1524 & N1525;
  assign N1541 = N1524 & fwd_sel_r[31];
  assign N1542 = ~bk_dpath_sel_r_28;
  assign N1543 = ~bk_dpath_sel_r_29;
  assign N1544 = N1542 & N1543;
  assign N1545 = N1542 & bk_dpath_sel_r_29;
  assign N1546 = bk_dpath_sel_r_28 & N1543;
  assign N1547 = bk_dpath_sel_r_28 & bk_dpath_sel_r_29;
  assign N1548 = ~bk_dpath_sel_r_30;
  assign N1549 = N1544 & N1548;
  assign N1550 = N1544 & bk_dpath_sel_r_30;
  assign N1551 = N1546 & N1548;
  assign N1552 = N1546 & bk_dpath_sel_r_30;
  assign N1553 = N1545 & N1548;
  assign N1554 = N1545 & bk_dpath_sel_r_30;
  assign N1555 = N1547 & N1548;
  assign N1556 = N1547 & bk_dpath_sel_r_30;
  assign in_v_o[8] = N2844 | N2845;
  assign N2844 = N2842 | N2843;
  assign N2842 = N2840 | N2841;
  assign N2840 = N2838 | N2839;
  assign N2838 = N2836 | N2837;
  assign N2836 = N2834 | N2835;
  assign N2834 = N2832 | N2833;
  assign N2832 = N2830 | N2831;
  assign N2830 = N2828 | N2829;
  assign N2828 = N2826 | N2827;
  assign N2826 = N2824 | N2825;
  assign N2824 = N2822 | N2823;
  assign N2822 = N2820 | N2821;
  assign N2820 = N2818 | N2819;
  assign N2818 = N2816 | N2817;
  assign N2816 = in_v_i[15] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__15_ ;
  assign N2817 = in_v_i[14] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__14_ ;
  assign N2819 = in_v_i[13] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__13_ ;
  assign N2821 = in_v_i[12] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__12_ ;
  assign N2823 = in_v_i[11] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__11_ ;
  assign N2825 = in_v_i[10] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__10_ ;
  assign N2827 = in_v_i[9] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__9_ ;
  assign N2829 = in_v_i[8] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__8_ ;
  assign N2831 = in_v_i[7] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__7_ ;
  assign N2833 = in_v_i[6] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__6_ ;
  assign N2835 = in_v_i[5] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__5_ ;
  assign N2837 = in_v_i[4] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__4_ ;
  assign N2839 = in_v_i[3] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__3_ ;
  assign N2841 = in_v_i[2] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__2_ ;
  assign N2843 = in_v_i[1] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__1_ ;
  assign N2845 = in_v_i[0] & \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__0_ ;
  assign N1573 = ~bk_sel_r[32];
  assign N1574 = ~bk_sel_r[33];
  assign N1575 = N1573 & N1574;
  assign N1576 = N1573 & bk_sel_r[33];
  assign N1577 = bk_sel_r[32] & N1574;
  assign N1578 = bk_sel_r[32] & bk_sel_r[33];
  assign N1579 = ~bk_sel_r[34];
  assign N1580 = N1575 & N1579;
  assign N1581 = N1575 & bk_sel_r[34];
  assign N1582 = N1577 & N1579;
  assign N1583 = N1577 & bk_sel_r[34];
  assign N1584 = N1576 & N1579;
  assign N1585 = N1576 & bk_sel_r[34];
  assign N1586 = N1578 & N1579;
  assign N1587 = N1578 & bk_sel_r[34];
  assign N1588 = ~bk_sel_r[35];
  assign N1589 = N1580 & N1588;
  assign N1590 = N1580 & bk_sel_r[35];
  assign N1591 = N1582 & N1588;
  assign N1592 = N1582 & bk_sel_r[35];
  assign N1593 = N1584 & N1588;
  assign N1594 = N1584 & bk_sel_r[35];
  assign N1595 = N1586 & N1588;
  assign N1596 = N1586 & bk_sel_r[35];
  assign N1597 = N1581 & N1588;
  assign N1598 = N1581 & bk_sel_r[35];
  assign N1599 = N1583 & N1588;
  assign N1600 = N1583 & bk_sel_r[35];
  assign N1601 = N1585 & N1588;
  assign N1602 = N1585 & bk_sel_r[35];
  assign N1603 = N1587 & N1588;
  assign N1604 = N1587 & bk_sel_r[35];
  assign N1605 = ~fwd_dpath_sel_r[32];
  assign N1606 = ~fwd_dpath_sel_r[33];
  assign N1607 = N1605 & N1606;
  assign N1608 = N1605 & fwd_dpath_sel_r[33];
  assign N1609 = fwd_dpath_sel_r[32] & N1606;
  assign N1610 = fwd_dpath_sel_r[32] & fwd_dpath_sel_r[33];
  assign N1611 = ~fwd_dpath_sel_r[34];
  assign N1612 = N1607 & N1611;
  assign N1613 = N1607 & fwd_dpath_sel_r[34];
  assign N1614 = N1609 & N1611;
  assign N1615 = N1609 & fwd_dpath_sel_r[34];
  assign N1616 = N1608 & N1611;
  assign N1617 = N1608 & fwd_dpath_sel_r[34];
  assign N1618 = N1610 & N1611;
  assign N1619 = N1610 & fwd_dpath_sel_r[34];
  assign N1620 = N1573 & N1574;
  assign N1621 = N1573 & bk_sel_r[33];
  assign N1622 = bk_sel_r[32] & N1574;
  assign N1623 = bk_sel_r[32] & bk_sel_r[33];
  assign N1624 = N1620 & N1579;
  assign N1625 = N1620 & bk_sel_r[34];
  assign N1626 = N1622 & N1579;
  assign N1627 = N1622 & bk_sel_r[34];
  assign N1628 = N1621 & N1579;
  assign N1629 = N1621 & bk_sel_r[34];
  assign N1630 = N1623 & N1579;
  assign N1631 = N1623 & bk_sel_r[34];
  assign N1632 = N1624 & N1588;
  assign N1633 = N1624 & bk_sel_r[35];
  assign N1634 = N1626 & N1588;
  assign N1635 = N1626 & bk_sel_r[35];
  assign N1636 = N1628 & N1588;
  assign N1637 = N1628 & bk_sel_r[35];
  assign N1638 = N1630 & N1588;
  assign N1639 = N1630 & bk_sel_r[35];
  assign N1640 = N1625 & N1588;
  assign N1641 = N1625 & bk_sel_r[35];
  assign N1642 = N1627 & N1588;
  assign N1643 = N1627 & bk_sel_r[35];
  assign N1644 = N1629 & N1588;
  assign N1645 = N1629 & bk_sel_r[35];
  assign N1646 = N1631 & N1588;
  assign N1647 = N1631 & bk_sel_r[35];
  assign N1648 = ~fwd_sel_r[32];
  assign N1649 = ~fwd_sel_r[33];
  assign N1650 = N1648 & N1649;
  assign N1651 = N1648 & fwd_sel_r[33];
  assign N1652 = fwd_sel_r[32] & N1649;
  assign N1653 = fwd_sel_r[32] & fwd_sel_r[33];
  assign N1654 = ~fwd_sel_r[34];
  assign N1655 = N1650 & N1654;
  assign N1656 = N1650 & fwd_sel_r[34];
  assign N1657 = N1652 & N1654;
  assign N1658 = N1652 & fwd_sel_r[34];
  assign N1659 = N1651 & N1654;
  assign N1660 = N1651 & fwd_sel_r[34];
  assign N1661 = N1653 & N1654;
  assign N1662 = N1653 & fwd_sel_r[34];
  assign N1663 = ~fwd_sel_r[35];
  assign N1664 = N1655 & N1663;
  assign N1665 = N1655 & fwd_sel_r[35];
  assign N1666 = N1657 & N1663;
  assign N1667 = N1657 & fwd_sel_r[35];
  assign N1668 = N1659 & N1663;
  assign N1669 = N1659 & fwd_sel_r[35];
  assign N1670 = N1661 & N1663;
  assign N1671 = N1661 & fwd_sel_r[35];
  assign N1672 = N1656 & N1663;
  assign N1673 = N1656 & fwd_sel_r[35];
  assign N1674 = N1658 & N1663;
  assign N1675 = N1658 & fwd_sel_r[35];
  assign N1676 = N1660 & N1663;
  assign N1677 = N1660 & fwd_sel_r[35];
  assign N1678 = N1662 & N1663;
  assign N1679 = N1662 & fwd_sel_r[35];
  assign in_v_o[9] = N2874 | N2875;
  assign N2874 = N2872 | N2873;
  assign N2872 = N2870 | N2871;
  assign N2870 = N2868 | N2869;
  assign N2868 = N2866 | N2867;
  assign N2866 = N2864 | N2865;
  assign N2864 = N2862 | N2863;
  assign N2862 = N2860 | N2861;
  assign N2860 = N2858 | N2859;
  assign N2858 = N2856 | N2857;
  assign N2856 = N2854 | N2855;
  assign N2854 = N2852 | N2853;
  assign N2852 = N2850 | N2851;
  assign N2850 = N2848 | N2849;
  assign N2848 = N2846 | N2847;
  assign N2846 = in_v_i[15] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__15_ ;
  assign N2847 = in_v_i[14] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__14_ ;
  assign N2849 = in_v_i[13] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__13_ ;
  assign N2851 = in_v_i[12] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__12_ ;
  assign N2853 = in_v_i[11] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__11_ ;
  assign N2855 = in_v_i[10] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__10_ ;
  assign N2857 = in_v_i[9] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__9_ ;
  assign N2859 = in_v_i[8] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__8_ ;
  assign N2861 = in_v_i[7] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__7_ ;
  assign N2863 = in_v_i[6] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__6_ ;
  assign N2865 = in_v_i[5] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__5_ ;
  assign N2867 = in_v_i[4] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__4_ ;
  assign N2869 = in_v_i[3] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__3_ ;
  assign N2871 = in_v_i[2] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__2_ ;
  assign N2873 = in_v_i[1] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__1_ ;
  assign N2875 = in_v_i[0] & \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__0_ ;
  assign N1704 = ~bk_sel_r[36];
  assign N1705 = ~bk_sel_r[37];
  assign N1706 = N1704 & N1705;
  assign N1707 = N1704 & bk_sel_r[37];
  assign N1708 = bk_sel_r[36] & N1705;
  assign N1709 = bk_sel_r[36] & bk_sel_r[37];
  assign N1710 = ~bk_sel_r[38];
  assign N1711 = N1706 & N1710;
  assign N1712 = N1706 & bk_sel_r[38];
  assign N1713 = N1708 & N1710;
  assign N1714 = N1708 & bk_sel_r[38];
  assign N1715 = N1707 & N1710;
  assign N1716 = N1707 & bk_sel_r[38];
  assign N1717 = N1709 & N1710;
  assign N1718 = N1709 & bk_sel_r[38];
  assign N1719 = ~bk_sel_r[39];
  assign N1720 = N1711 & N1719;
  assign N1721 = N1711 & bk_sel_r[39];
  assign N1722 = N1713 & N1719;
  assign N1723 = N1713 & bk_sel_r[39];
  assign N1724 = N1715 & N1719;
  assign N1725 = N1715 & bk_sel_r[39];
  assign N1726 = N1717 & N1719;
  assign N1727 = N1717 & bk_sel_r[39];
  assign N1728 = N1712 & N1719;
  assign N1729 = N1712 & bk_sel_r[39];
  assign N1730 = N1714 & N1719;
  assign N1731 = N1714 & bk_sel_r[39];
  assign N1732 = N1716 & N1719;
  assign N1733 = N1716 & bk_sel_r[39];
  assign N1734 = N1718 & N1719;
  assign N1735 = N1718 & bk_sel_r[39];
  assign N1743 = N1704 & N1705;
  assign N1744 = N1704 & bk_sel_r[37];
  assign N1745 = bk_sel_r[36] & N1705;
  assign N1746 = bk_sel_r[36] & bk_sel_r[37];
  assign N1747 = N1743 & N1710;
  assign N1748 = N1743 & bk_sel_r[38];
  assign N1749 = N1745 & N1710;
  assign N1750 = N1745 & bk_sel_r[38];
  assign N1751 = N1744 & N1710;
  assign N1752 = N1744 & bk_sel_r[38];
  assign N1753 = N1746 & N1710;
  assign N1754 = N1746 & bk_sel_r[38];
  assign N1755 = N1747 & N1719;
  assign N1756 = N1747 & bk_sel_r[39];
  assign N1757 = N1749 & N1719;
  assign N1758 = N1749 & bk_sel_r[39];
  assign N1759 = N1751 & N1719;
  assign N1760 = N1751 & bk_sel_r[39];
  assign N1761 = N1753 & N1719;
  assign N1762 = N1753 & bk_sel_r[39];
  assign N1763 = N1748 & N1719;
  assign N1764 = N1748 & bk_sel_r[39];
  assign N1765 = N1750 & N1719;
  assign N1766 = N1750 & bk_sel_r[39];
  assign N1767 = N1752 & N1719;
  assign N1768 = N1752 & bk_sel_r[39];
  assign N1769 = N1754 & N1719;
  assign N1770 = N1754 & bk_sel_r[39];
  assign N1771 = ~fwd_sel_r[36];
  assign N1772 = ~fwd_sel_r[37];
  assign N1773 = N1771 & N1772;
  assign N1774 = N1771 & fwd_sel_r[37];
  assign N1775 = fwd_sel_r[36] & N1772;
  assign N1776 = fwd_sel_r[36] & fwd_sel_r[37];
  assign N1777 = ~fwd_sel_r[38];
  assign N1778 = N1773 & N1777;
  assign N1779 = N1773 & fwd_sel_r[38];
  assign N1780 = N1775 & N1777;
  assign N1781 = N1775 & fwd_sel_r[38];
  assign N1782 = N1774 & N1777;
  assign N1783 = N1774 & fwd_sel_r[38];
  assign N1784 = N1776 & N1777;
  assign N1785 = N1776 & fwd_sel_r[38];
  assign N1786 = ~fwd_sel_r[39];
  assign N1787 = N1778 & N1786;
  assign N1788 = N1778 & fwd_sel_r[39];
  assign N1789 = N1780 & N1786;
  assign N1790 = N1780 & fwd_sel_r[39];
  assign N1791 = N1782 & N1786;
  assign N1792 = N1782 & fwd_sel_r[39];
  assign N1793 = N1784 & N1786;
  assign N1794 = N1784 & fwd_sel_r[39];
  assign N1795 = N1779 & N1786;
  assign N1796 = N1779 & fwd_sel_r[39];
  assign N1797 = N1781 & N1786;
  assign N1798 = N1781 & fwd_sel_r[39];
  assign N1799 = N1783 & N1786;
  assign N1800 = N1783 & fwd_sel_r[39];
  assign N1801 = N1785 & N1786;
  assign N1802 = N1785 & fwd_sel_r[39];
  assign in_v_o[10] = N2904 | N2905;
  assign N2904 = N2902 | N2903;
  assign N2902 = N2900 | N2901;
  assign N2900 = N2898 | N2899;
  assign N2898 = N2896 | N2897;
  assign N2896 = N2894 | N2895;
  assign N2894 = N2892 | N2893;
  assign N2892 = N2890 | N2891;
  assign N2890 = N2888 | N2889;
  assign N2888 = N2886 | N2887;
  assign N2886 = N2884 | N2885;
  assign N2884 = N2882 | N2883;
  assign N2882 = N2880 | N2881;
  assign N2880 = N2878 | N2879;
  assign N2878 = N2876 | N2877;
  assign N2876 = in_v_i[15] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__15_ ;
  assign N2877 = in_v_i[14] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__14_ ;
  assign N2879 = in_v_i[13] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__13_ ;
  assign N2881 = in_v_i[12] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__12_ ;
  assign N2883 = in_v_i[11] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__11_ ;
  assign N2885 = in_v_i[10] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__10_ ;
  assign N2887 = in_v_i[9] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__9_ ;
  assign N2889 = in_v_i[8] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__8_ ;
  assign N2891 = in_v_i[7] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__7_ ;
  assign N2893 = in_v_i[6] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__6_ ;
  assign N2895 = in_v_i[5] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__5_ ;
  assign N2897 = in_v_i[4] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__4_ ;
  assign N2899 = in_v_i[3] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__3_ ;
  assign N2901 = in_v_i[2] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__2_ ;
  assign N2903 = in_v_i[1] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__1_ ;
  assign N2905 = in_v_i[0] & \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__0_ ;
  assign N1829 = ~bk_sel_r[40];
  assign N1830 = ~bk_sel_r[41];
  assign N1831 = N1829 & N1830;
  assign N1832 = N1829 & bk_sel_r[41];
  assign N1833 = bk_sel_r[40] & N1830;
  assign N1834 = bk_sel_r[40] & bk_sel_r[41];
  assign N1835 = ~bk_sel_r[42];
  assign N1836 = N1831 & N1835;
  assign N1837 = N1831 & bk_sel_r[42];
  assign N1838 = N1833 & N1835;
  assign N1839 = N1833 & bk_sel_r[42];
  assign N1840 = N1832 & N1835;
  assign N1841 = N1832 & bk_sel_r[42];
  assign N1842 = N1834 & N1835;
  assign N1843 = N1834 & bk_sel_r[42];
  assign N1844 = ~bk_sel_r[43];
  assign N1845 = N1836 & N1844;
  assign N1846 = N1836 & bk_sel_r[43];
  assign N1847 = N1838 & N1844;
  assign N1848 = N1838 & bk_sel_r[43];
  assign N1849 = N1840 & N1844;
  assign N1850 = N1840 & bk_sel_r[43];
  assign N1851 = N1842 & N1844;
  assign N1852 = N1842 & bk_sel_r[43];
  assign N1853 = N1837 & N1844;
  assign N1854 = N1837 & bk_sel_r[43];
  assign N1855 = N1839 & N1844;
  assign N1856 = N1839 & bk_sel_r[43];
  assign N1857 = N1841 & N1844;
  assign N1858 = N1841 & bk_sel_r[43];
  assign N1859 = N1843 & N1844;
  assign N1860 = N1843 & bk_sel_r[43];
  assign N1867 = N1829 & N1830;
  assign N1868 = N1829 & bk_sel_r[41];
  assign N1869 = bk_sel_r[40] & N1830;
  assign N1870 = bk_sel_r[40] & bk_sel_r[41];
  assign N1871 = N1867 & N1835;
  assign N1872 = N1867 & bk_sel_r[42];
  assign N1873 = N1869 & N1835;
  assign N1874 = N1869 & bk_sel_r[42];
  assign N1875 = N1868 & N1835;
  assign N1876 = N1868 & bk_sel_r[42];
  assign N1877 = N1870 & N1835;
  assign N1878 = N1870 & bk_sel_r[42];
  assign N1879 = N1871 & N1844;
  assign N1880 = N1871 & bk_sel_r[43];
  assign N1881 = N1873 & N1844;
  assign N1882 = N1873 & bk_sel_r[43];
  assign N1883 = N1875 & N1844;
  assign N1884 = N1875 & bk_sel_r[43];
  assign N1885 = N1877 & N1844;
  assign N1886 = N1877 & bk_sel_r[43];
  assign N1887 = N1872 & N1844;
  assign N1888 = N1872 & bk_sel_r[43];
  assign N1889 = N1874 & N1844;
  assign N1890 = N1874 & bk_sel_r[43];
  assign N1891 = N1876 & N1844;
  assign N1892 = N1876 & bk_sel_r[43];
  assign N1893 = N1878 & N1844;
  assign N1894 = N1878 & bk_sel_r[43];
  assign N1895 = ~fwd_sel_r[40];
  assign N1896 = ~fwd_sel_r[41];
  assign N1897 = N1895 & N1896;
  assign N1898 = N1895 & fwd_sel_r[41];
  assign N1899 = fwd_sel_r[40] & N1896;
  assign N1900 = fwd_sel_r[40] & fwd_sel_r[41];
  assign N1901 = ~fwd_sel_r[42];
  assign N1902 = N1897 & N1901;
  assign N1903 = N1897 & fwd_sel_r[42];
  assign N1904 = N1899 & N1901;
  assign N1905 = N1899 & fwd_sel_r[42];
  assign N1906 = N1898 & N1901;
  assign N1907 = N1898 & fwd_sel_r[42];
  assign N1908 = N1900 & N1901;
  assign N1909 = N1900 & fwd_sel_r[42];
  assign N1910 = ~fwd_sel_r[43];
  assign N1911 = N1902 & N1910;
  assign N1912 = N1902 & fwd_sel_r[43];
  assign N1913 = N1904 & N1910;
  assign N1914 = N1904 & fwd_sel_r[43];
  assign N1915 = N1906 & N1910;
  assign N1916 = N1906 & fwd_sel_r[43];
  assign N1917 = N1908 & N1910;
  assign N1918 = N1908 & fwd_sel_r[43];
  assign N1919 = N1903 & N1910;
  assign N1920 = N1903 & fwd_sel_r[43];
  assign N1921 = N1905 & N1910;
  assign N1922 = N1905 & fwd_sel_r[43];
  assign N1923 = N1907 & N1910;
  assign N1924 = N1907 & fwd_sel_r[43];
  assign N1925 = N1909 & N1910;
  assign N1926 = N1909 & fwd_sel_r[43];
  assign in_v_o[11] = N2934 | N2935;
  assign N2934 = N2932 | N2933;
  assign N2932 = N2930 | N2931;
  assign N2930 = N2928 | N2929;
  assign N2928 = N2926 | N2927;
  assign N2926 = N2924 | N2925;
  assign N2924 = N2922 | N2923;
  assign N2922 = N2920 | N2921;
  assign N2920 = N2918 | N2919;
  assign N2918 = N2916 | N2917;
  assign N2916 = N2914 | N2915;
  assign N2914 = N2912 | N2913;
  assign N2912 = N2910 | N2911;
  assign N2910 = N2908 | N2909;
  assign N2908 = N2906 | N2907;
  assign N2906 = in_v_i[15] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__15_ ;
  assign N2907 = in_v_i[14] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__14_ ;
  assign N2909 = in_v_i[13] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__13_ ;
  assign N2911 = in_v_i[12] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__12_ ;
  assign N2913 = in_v_i[11] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__11_ ;
  assign N2915 = in_v_i[10] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__10_ ;
  assign N2917 = in_v_i[9] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__9_ ;
  assign N2919 = in_v_i[8] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__8_ ;
  assign N2921 = in_v_i[7] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__7_ ;
  assign N2923 = in_v_i[6] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__6_ ;
  assign N2925 = in_v_i[5] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__5_ ;
  assign N2927 = in_v_i[4] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__4_ ;
  assign N2929 = in_v_i[3] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__3_ ;
  assign N2931 = in_v_i[2] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__2_ ;
  assign N2933 = in_v_i[1] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__1_ ;
  assign N2935 = in_v_i[0] & \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__0_ ;
  assign N1954 = ~bk_sel_r[44];
  assign N1955 = ~bk_sel_r[45];
  assign N1956 = N1954 & N1955;
  assign N1957 = N1954 & bk_sel_r[45];
  assign N1958 = bk_sel_r[44] & N1955;
  assign N1959 = bk_sel_r[44] & bk_sel_r[45];
  assign N1960 = ~bk_sel_r[46];
  assign N1961 = N1956 & N1960;
  assign N1962 = N1956 & bk_sel_r[46];
  assign N1963 = N1958 & N1960;
  assign N1964 = N1958 & bk_sel_r[46];
  assign N1965 = N1957 & N1960;
  assign N1966 = N1957 & bk_sel_r[46];
  assign N1967 = N1959 & N1960;
  assign N1968 = N1959 & bk_sel_r[46];
  assign N1969 = ~bk_sel_r[47];
  assign N1970 = N1961 & N1969;
  assign N1971 = N1961 & bk_sel_r[47];
  assign N1972 = N1963 & N1969;
  assign N1973 = N1963 & bk_sel_r[47];
  assign N1974 = N1965 & N1969;
  assign N1975 = N1965 & bk_sel_r[47];
  assign N1976 = N1967 & N1969;
  assign N1977 = N1967 & bk_sel_r[47];
  assign N1978 = N1962 & N1969;
  assign N1979 = N1962 & bk_sel_r[47];
  assign N1980 = N1964 & N1969;
  assign N1981 = N1964 & bk_sel_r[47];
  assign N1982 = N1966 & N1969;
  assign N1983 = N1966 & bk_sel_r[47];
  assign N1984 = N1968 & N1969;
  assign N1985 = N1968 & bk_sel_r[47];
  assign N1990 = N1954 & N1955;
  assign N1991 = N1954 & bk_sel_r[45];
  assign N1992 = bk_sel_r[44] & N1955;
  assign N1993 = bk_sel_r[44] & bk_sel_r[45];
  assign N1994 = N1990 & N1960;
  assign N1995 = N1990 & bk_sel_r[46];
  assign N1996 = N1992 & N1960;
  assign N1997 = N1992 & bk_sel_r[46];
  assign N1998 = N1991 & N1960;
  assign N1999 = N1991 & bk_sel_r[46];
  assign N2000 = N1993 & N1960;
  assign N2001 = N1993 & bk_sel_r[46];
  assign N2002 = N1994 & N1969;
  assign N2003 = N1994 & bk_sel_r[47];
  assign N2004 = N1996 & N1969;
  assign N2005 = N1996 & bk_sel_r[47];
  assign N2006 = N1998 & N1969;
  assign N2007 = N1998 & bk_sel_r[47];
  assign N2008 = N2000 & N1969;
  assign N2009 = N2000 & bk_sel_r[47];
  assign N2010 = N1995 & N1969;
  assign N2011 = N1995 & bk_sel_r[47];
  assign N2012 = N1997 & N1969;
  assign N2013 = N1997 & bk_sel_r[47];
  assign N2014 = N1999 & N1969;
  assign N2015 = N1999 & bk_sel_r[47];
  assign N2016 = N2001 & N1969;
  assign N2017 = N2001 & bk_sel_r[47];
  assign N2018 = ~fwd_sel_r[44];
  assign N2019 = ~fwd_sel_r[45];
  assign N2020 = N2018 & N2019;
  assign N2021 = N2018 & fwd_sel_r[45];
  assign N2022 = fwd_sel_r[44] & N2019;
  assign N2023 = fwd_sel_r[44] & fwd_sel_r[45];
  assign N2024 = ~fwd_sel_r[46];
  assign N2025 = N2020 & N2024;
  assign N2026 = N2020 & fwd_sel_r[46];
  assign N2027 = N2022 & N2024;
  assign N2028 = N2022 & fwd_sel_r[46];
  assign N2029 = N2021 & N2024;
  assign N2030 = N2021 & fwd_sel_r[46];
  assign N2031 = N2023 & N2024;
  assign N2032 = N2023 & fwd_sel_r[46];
  assign N2033 = ~fwd_sel_r[47];
  assign N2034 = N2025 & N2033;
  assign N2035 = N2025 & fwd_sel_r[47];
  assign N2036 = N2027 & N2033;
  assign N2037 = N2027 & fwd_sel_r[47];
  assign N2038 = N2029 & N2033;
  assign N2039 = N2029 & fwd_sel_r[47];
  assign N2040 = N2031 & N2033;
  assign N2041 = N2031 & fwd_sel_r[47];
  assign N2042 = N2026 & N2033;
  assign N2043 = N2026 & fwd_sel_r[47];
  assign N2044 = N2028 & N2033;
  assign N2045 = N2028 & fwd_sel_r[47];
  assign N2046 = N2030 & N2033;
  assign N2047 = N2030 & fwd_sel_r[47];
  assign N2048 = N2032 & N2033;
  assign N2049 = N2032 & fwd_sel_r[47];
  assign in_v_o[12] = N2964 | N2965;
  assign N2964 = N2962 | N2963;
  assign N2962 = N2960 | N2961;
  assign N2960 = N2958 | N2959;
  assign N2958 = N2956 | N2957;
  assign N2956 = N2954 | N2955;
  assign N2954 = N2952 | N2953;
  assign N2952 = N2950 | N2951;
  assign N2950 = N2948 | N2949;
  assign N2948 = N2946 | N2947;
  assign N2946 = N2944 | N2945;
  assign N2944 = N2942 | N2943;
  assign N2942 = N2940 | N2941;
  assign N2940 = N2938 | N2939;
  assign N2938 = N2936 | N2937;
  assign N2936 = in_v_i[15] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__15_ ;
  assign N2937 = in_v_i[14] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__14_ ;
  assign N2939 = in_v_i[13] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__13_ ;
  assign N2941 = in_v_i[12] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__12_ ;
  assign N2943 = in_v_i[11] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__11_ ;
  assign N2945 = in_v_i[10] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__10_ ;
  assign N2947 = in_v_i[9] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__9_ ;
  assign N2949 = in_v_i[8] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__8_ ;
  assign N2951 = in_v_i[7] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__7_ ;
  assign N2953 = in_v_i[6] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__6_ ;
  assign N2955 = in_v_i[5] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__5_ ;
  assign N2957 = in_v_i[4] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__4_ ;
  assign N2959 = in_v_i[3] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__3_ ;
  assign N2961 = in_v_i[2] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__2_ ;
  assign N2963 = in_v_i[1] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__1_ ;
  assign N2965 = in_v_i[0] & \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__0_ ;
  assign N2078 = ~bk_sel_r[48];
  assign N2079 = ~bk_sel_r[49];
  assign N2080 = N2078 & N2079;
  assign N2081 = N2078 & bk_sel_r[49];
  assign N2082 = bk_sel_r[48] & N2079;
  assign N2083 = bk_sel_r[48] & bk_sel_r[49];
  assign N2084 = ~bk_sel_r[50];
  assign N2085 = N2080 & N2084;
  assign N2086 = N2080 & bk_sel_r[50];
  assign N2087 = N2082 & N2084;
  assign N2088 = N2082 & bk_sel_r[50];
  assign N2089 = N2081 & N2084;
  assign N2090 = N2081 & bk_sel_r[50];
  assign N2091 = N2083 & N2084;
  assign N2092 = N2083 & bk_sel_r[50];
  assign N2093 = ~bk_sel_r[51];
  assign N2094 = N2085 & N2093;
  assign N2095 = N2085 & bk_sel_r[51];
  assign N2096 = N2087 & N2093;
  assign N2097 = N2087 & bk_sel_r[51];
  assign N2098 = N2089 & N2093;
  assign N2099 = N2089 & bk_sel_r[51];
  assign N2100 = N2091 & N2093;
  assign N2101 = N2091 & bk_sel_r[51];
  assign N2102 = N2086 & N2093;
  assign N2103 = N2086 & bk_sel_r[51];
  assign N2104 = N2088 & N2093;
  assign N2105 = N2088 & bk_sel_r[51];
  assign N2106 = N2090 & N2093;
  assign N2107 = N2090 & bk_sel_r[51];
  assign N2108 = N2092 & N2093;
  assign N2109 = N2092 & bk_sel_r[51];
  assign N2110 = ~fwd_dpath_sel_r_48;
  assign N2111 = ~fwd_dpath_sel_r_49;
  assign N2112 = N2110 & N2111;
  assign N2113 = N2110 & fwd_dpath_sel_r_49;
  assign N2114 = fwd_dpath_sel_r_48 & N2111;
  assign N2115 = fwd_dpath_sel_r_48 & fwd_dpath_sel_r_49;
  assign N2116 = N2078 & N2079;
  assign N2117 = N2078 & bk_sel_r[49];
  assign N2118 = bk_sel_r[48] & N2079;
  assign N2119 = bk_sel_r[48] & bk_sel_r[49];
  assign N2120 = N2116 & N2084;
  assign N2121 = N2116 & bk_sel_r[50];
  assign N2122 = N2118 & N2084;
  assign N2123 = N2118 & bk_sel_r[50];
  assign N2124 = N2117 & N2084;
  assign N2125 = N2117 & bk_sel_r[50];
  assign N2126 = N2119 & N2084;
  assign N2127 = N2119 & bk_sel_r[50];
  assign N2128 = N2120 & N2093;
  assign N2129 = N2120 & bk_sel_r[51];
  assign N2130 = N2122 & N2093;
  assign N2131 = N2122 & bk_sel_r[51];
  assign N2132 = N2124 & N2093;
  assign N2133 = N2124 & bk_sel_r[51];
  assign N2134 = N2126 & N2093;
  assign N2135 = N2126 & bk_sel_r[51];
  assign N2136 = N2121 & N2093;
  assign N2137 = N2121 & bk_sel_r[51];
  assign N2138 = N2123 & N2093;
  assign N2139 = N2123 & bk_sel_r[51];
  assign N2140 = N2125 & N2093;
  assign N2141 = N2125 & bk_sel_r[51];
  assign N2142 = N2127 & N2093;
  assign N2143 = N2127 & bk_sel_r[51];
  assign N2144 = ~fwd_sel_r[48];
  assign N2145 = ~fwd_sel_r[49];
  assign N2146 = N2144 & N2145;
  assign N2147 = N2144 & fwd_sel_r[49];
  assign N2148 = fwd_sel_r[48] & N2145;
  assign N2149 = fwd_sel_r[48] & fwd_sel_r[49];
  assign N2150 = ~fwd_sel_r[50];
  assign N2151 = N2146 & N2150;
  assign N2152 = N2146 & fwd_sel_r[50];
  assign N2153 = N2148 & N2150;
  assign N2154 = N2148 & fwd_sel_r[50];
  assign N2155 = N2147 & N2150;
  assign N2156 = N2147 & fwd_sel_r[50];
  assign N2157 = N2149 & N2150;
  assign N2158 = N2149 & fwd_sel_r[50];
  assign N2159 = ~fwd_sel_r[51];
  assign N2160 = N2151 & N2159;
  assign N2161 = N2151 & fwd_sel_r[51];
  assign N2162 = N2153 & N2159;
  assign N2163 = N2153 & fwd_sel_r[51];
  assign N2164 = N2155 & N2159;
  assign N2165 = N2155 & fwd_sel_r[51];
  assign N2166 = N2157 & N2159;
  assign N2167 = N2157 & fwd_sel_r[51];
  assign N2168 = N2152 & N2159;
  assign N2169 = N2152 & fwd_sel_r[51];
  assign N2170 = N2154 & N2159;
  assign N2171 = N2154 & fwd_sel_r[51];
  assign N2172 = N2156 & N2159;
  assign N2173 = N2156 & fwd_sel_r[51];
  assign N2174 = N2158 & N2159;
  assign N2175 = N2158 & fwd_sel_r[51];
  assign in_v_o[13] = N2994 | N2995;
  assign N2994 = N2992 | N2993;
  assign N2992 = N2990 | N2991;
  assign N2990 = N2988 | N2989;
  assign N2988 = N2986 | N2987;
  assign N2986 = N2984 | N2985;
  assign N2984 = N2982 | N2983;
  assign N2982 = N2980 | N2981;
  assign N2980 = N2978 | N2979;
  assign N2978 = N2976 | N2977;
  assign N2976 = N2974 | N2975;
  assign N2974 = N2972 | N2973;
  assign N2972 = N2970 | N2971;
  assign N2970 = N2968 | N2969;
  assign N2968 = N2966 | N2967;
  assign N2966 = in_v_i[15] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__15_ ;
  assign N2967 = in_v_i[14] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__14_ ;
  assign N2969 = in_v_i[13] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__13_ ;
  assign N2971 = in_v_i[12] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__12_ ;
  assign N2973 = in_v_i[11] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__11_ ;
  assign N2975 = in_v_i[10] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__10_ ;
  assign N2977 = in_v_i[9] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__9_ ;
  assign N2979 = in_v_i[8] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__8_ ;
  assign N2981 = in_v_i[7] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__7_ ;
  assign N2983 = in_v_i[6] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__6_ ;
  assign N2985 = in_v_i[5] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__5_ ;
  assign N2987 = in_v_i[4] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__4_ ;
  assign N2989 = in_v_i[3] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__3_ ;
  assign N2991 = in_v_i[2] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__2_ ;
  assign N2993 = in_v_i[1] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__1_ ;
  assign N2995 = in_v_i[0] & \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__0_ ;
  assign N2205 = ~bk_sel_r[52];
  assign N2206 = ~bk_sel_r[53];
  assign N2207 = N2205 & N2206;
  assign N2208 = N2205 & bk_sel_r[53];
  assign N2209 = bk_sel_r[52] & N2206;
  assign N2210 = bk_sel_r[52] & bk_sel_r[53];
  assign N2211 = ~bk_sel_r[54];
  assign N2212 = N2207 & N2211;
  assign N2213 = N2207 & bk_sel_r[54];
  assign N2214 = N2209 & N2211;
  assign N2215 = N2209 & bk_sel_r[54];
  assign N2216 = N2208 & N2211;
  assign N2217 = N2208 & bk_sel_r[54];
  assign N2218 = N2210 & N2211;
  assign N2219 = N2210 & bk_sel_r[54];
  assign N2220 = ~bk_sel_r[55];
  assign N2221 = N2212 & N2220;
  assign N2222 = N2212 & bk_sel_r[55];
  assign N2223 = N2214 & N2220;
  assign N2224 = N2214 & bk_sel_r[55];
  assign N2225 = N2216 & N2220;
  assign N2226 = N2216 & bk_sel_r[55];
  assign N2227 = N2218 & N2220;
  assign N2228 = N2218 & bk_sel_r[55];
  assign N2229 = N2213 & N2220;
  assign N2230 = N2213 & bk_sel_r[55];
  assign N2231 = N2215 & N2220;
  assign N2232 = N2215 & bk_sel_r[55];
  assign N2233 = N2217 & N2220;
  assign N2234 = N2217 & bk_sel_r[55];
  assign N2235 = N2219 & N2220;
  assign N2236 = N2219 & bk_sel_r[55];
  assign N2238 = N2205 & N2206;
  assign N2239 = N2205 & bk_sel_r[53];
  assign N2240 = bk_sel_r[52] & N2206;
  assign N2241 = bk_sel_r[52] & bk_sel_r[53];
  assign N2242 = N2238 & N2211;
  assign N2243 = N2238 & bk_sel_r[54];
  assign N2244 = N2240 & N2211;
  assign N2245 = N2240 & bk_sel_r[54];
  assign N2246 = N2239 & N2211;
  assign N2247 = N2239 & bk_sel_r[54];
  assign N2248 = N2241 & N2211;
  assign N2249 = N2241 & bk_sel_r[54];
  assign N2250 = N2242 & N2220;
  assign N2251 = N2242 & bk_sel_r[55];
  assign N2252 = N2244 & N2220;
  assign N2253 = N2244 & bk_sel_r[55];
  assign N2254 = N2246 & N2220;
  assign N2255 = N2246 & bk_sel_r[55];
  assign N2256 = N2248 & N2220;
  assign N2257 = N2248 & bk_sel_r[55];
  assign N2258 = N2243 & N2220;
  assign N2259 = N2243 & bk_sel_r[55];
  assign N2260 = N2245 & N2220;
  assign N2261 = N2245 & bk_sel_r[55];
  assign N2262 = N2247 & N2220;
  assign N2263 = N2247 & bk_sel_r[55];
  assign N2264 = N2249 & N2220;
  assign N2265 = N2249 & bk_sel_r[55];
  assign N2266 = ~fwd_sel_r[52];
  assign N2267 = ~fwd_sel_r[53];
  assign N2268 = N2266 & N2267;
  assign N2269 = N2266 & fwd_sel_r[53];
  assign N2270 = fwd_sel_r[52] & N2267;
  assign N2271 = fwd_sel_r[52] & fwd_sel_r[53];
  assign N2272 = ~fwd_sel_r[54];
  assign N2273 = N2268 & N2272;
  assign N2274 = N2268 & fwd_sel_r[54];
  assign N2275 = N2270 & N2272;
  assign N2276 = N2270 & fwd_sel_r[54];
  assign N2277 = N2269 & N2272;
  assign N2278 = N2269 & fwd_sel_r[54];
  assign N2279 = N2271 & N2272;
  assign N2280 = N2271 & fwd_sel_r[54];
  assign N2281 = ~fwd_sel_r[55];
  assign N2282 = N2273 & N2281;
  assign N2283 = N2273 & fwd_sel_r[55];
  assign N2284 = N2275 & N2281;
  assign N2285 = N2275 & fwd_sel_r[55];
  assign N2286 = N2277 & N2281;
  assign N2287 = N2277 & fwd_sel_r[55];
  assign N2288 = N2279 & N2281;
  assign N2289 = N2279 & fwd_sel_r[55];
  assign N2290 = N2274 & N2281;
  assign N2291 = N2274 & fwd_sel_r[55];
  assign N2292 = N2276 & N2281;
  assign N2293 = N2276 & fwd_sel_r[55];
  assign N2294 = N2278 & N2281;
  assign N2295 = N2278 & fwd_sel_r[55];
  assign N2296 = N2280 & N2281;
  assign N2297 = N2280 & fwd_sel_r[55];
  assign in_v_o[14] = N3024 | N3025;
  assign N3024 = N3022 | N3023;
  assign N3022 = N3020 | N3021;
  assign N3020 = N3018 | N3019;
  assign N3018 = N3016 | N3017;
  assign N3016 = N3014 | N3015;
  assign N3014 = N3012 | N3013;
  assign N3012 = N3010 | N3011;
  assign N3010 = N3008 | N3009;
  assign N3008 = N3006 | N3007;
  assign N3006 = N3004 | N3005;
  assign N3004 = N3002 | N3003;
  assign N3002 = N3000 | N3001;
  assign N3000 = N2998 | N2999;
  assign N2998 = N2996 | N2997;
  assign N2996 = in_v_i[15] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__15_ ;
  assign N2997 = in_v_i[14] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__14_ ;
  assign N2999 = in_v_i[13] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__13_ ;
  assign N3001 = in_v_i[12] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__12_ ;
  assign N3003 = in_v_i[11] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__11_ ;
  assign N3005 = in_v_i[10] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__10_ ;
  assign N3007 = in_v_i[9] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__9_ ;
  assign N3009 = in_v_i[8] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__8_ ;
  assign N3011 = in_v_i[7] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__7_ ;
  assign N3013 = in_v_i[6] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__6_ ;
  assign N3015 = in_v_i[5] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__5_ ;
  assign N3017 = in_v_i[4] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__4_ ;
  assign N3019 = in_v_i[3] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__3_ ;
  assign N3021 = in_v_i[2] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__2_ ;
  assign N3023 = in_v_i[1] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__1_ ;
  assign N3025 = in_v_i[0] & \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__0_ ;
  assign N2328 = ~bk_sel_r[56];
  assign N2329 = ~bk_sel_r[57];
  assign N2330 = N2328 & N2329;
  assign N2331 = N2328 & bk_sel_r[57];
  assign N2332 = bk_sel_r[56] & N2329;
  assign N2333 = bk_sel_r[56] & bk_sel_r[57];
  assign N2334 = ~bk_sel_r[58];
  assign N2335 = N2330 & N2334;
  assign N2336 = N2330 & bk_sel_r[58];
  assign N2337 = N2332 & N2334;
  assign N2338 = N2332 & bk_sel_r[58];
  assign N2339 = N2331 & N2334;
  assign N2340 = N2331 & bk_sel_r[58];
  assign N2341 = N2333 & N2334;
  assign N2342 = N2333 & bk_sel_r[58];
  assign N2343 = ~bk_sel_r[59];
  assign N2344 = N2335 & N2343;
  assign N2345 = N2335 & bk_sel_r[59];
  assign N2346 = N2337 & N2343;
  assign N2347 = N2337 & bk_sel_r[59];
  assign N2348 = N2339 & N2343;
  assign N2349 = N2339 & bk_sel_r[59];
  assign N2350 = N2341 & N2343;
  assign N2351 = N2341 & bk_sel_r[59];
  assign N2352 = N2336 & N2343;
  assign N2353 = N2336 & bk_sel_r[59];
  assign N2354 = N2338 & N2343;
  assign N2355 = N2338 & bk_sel_r[59];
  assign N2356 = N2340 & N2343;
  assign N2357 = N2340 & bk_sel_r[59];
  assign N2358 = N2342 & N2343;
  assign N2359 = N2342 & bk_sel_r[59];
  assign N2360 = ~fwd_dpath_sel_r_56;
  assign N2361 = N2328 & N2329;
  assign N2362 = N2328 & bk_sel_r[57];
  assign N2363 = bk_sel_r[56] & N2329;
  assign N2364 = bk_sel_r[56] & bk_sel_r[57];
  assign N2365 = N2361 & N2334;
  assign N2366 = N2361 & bk_sel_r[58];
  assign N2367 = N2363 & N2334;
  assign N2368 = N2363 & bk_sel_r[58];
  assign N2369 = N2362 & N2334;
  assign N2370 = N2362 & bk_sel_r[58];
  assign N2371 = N2364 & N2334;
  assign N2372 = N2364 & bk_sel_r[58];
  assign N2373 = N2365 & N2343;
  assign N2374 = N2365 & bk_sel_r[59];
  assign N2375 = N2367 & N2343;
  assign N2376 = N2367 & bk_sel_r[59];
  assign N2377 = N2369 & N2343;
  assign N2378 = N2369 & bk_sel_r[59];
  assign N2379 = N2371 & N2343;
  assign N2380 = N2371 & bk_sel_r[59];
  assign N2381 = N2366 & N2343;
  assign N2382 = N2366 & bk_sel_r[59];
  assign N2383 = N2368 & N2343;
  assign N2384 = N2368 & bk_sel_r[59];
  assign N2385 = N2370 & N2343;
  assign N2386 = N2370 & bk_sel_r[59];
  assign N2387 = N2372 & N2343;
  assign N2388 = N2372 & bk_sel_r[59];
  assign N2389 = ~fwd_sel_r[56];
  assign N2390 = ~fwd_sel_r[57];
  assign N2391 = N2389 & N2390;
  assign N2392 = N2389 & fwd_sel_r[57];
  assign N2393 = fwd_sel_r[56] & N2390;
  assign N2394 = fwd_sel_r[56] & fwd_sel_r[57];
  assign N2395 = ~fwd_sel_r[58];
  assign N2396 = N2391 & N2395;
  assign N2397 = N2391 & fwd_sel_r[58];
  assign N2398 = N2393 & N2395;
  assign N2399 = N2393 & fwd_sel_r[58];
  assign N2400 = N2392 & N2395;
  assign N2401 = N2392 & fwd_sel_r[58];
  assign N2402 = N2394 & N2395;
  assign N2403 = N2394 & fwd_sel_r[58];
  assign N2404 = ~fwd_sel_r[59];
  assign N2405 = N2396 & N2404;
  assign N2406 = N2396 & fwd_sel_r[59];
  assign N2407 = N2398 & N2404;
  assign N2408 = N2398 & fwd_sel_r[59];
  assign N2409 = N2400 & N2404;
  assign N2410 = N2400 & fwd_sel_r[59];
  assign N2411 = N2402 & N2404;
  assign N2412 = N2402 & fwd_sel_r[59];
  assign N2413 = N2397 & N2404;
  assign N2414 = N2397 & fwd_sel_r[59];
  assign N2415 = N2399 & N2404;
  assign N2416 = N2399 & fwd_sel_r[59];
  assign N2417 = N2401 & N2404;
  assign N2418 = N2401 & fwd_sel_r[59];
  assign N2419 = N2403 & N2404;
  assign N2420 = N2403 & fwd_sel_r[59];
  assign in_v_o[15] = N3054 | N3055;
  assign N3054 = N3052 | N3053;
  assign N3052 = N3050 | N3051;
  assign N3050 = N3048 | N3049;
  assign N3048 = N3046 | N3047;
  assign N3046 = N3044 | N3045;
  assign N3044 = N3042 | N3043;
  assign N3042 = N3040 | N3041;
  assign N3040 = N3038 | N3039;
  assign N3038 = N3036 | N3037;
  assign N3036 = N3034 | N3035;
  assign N3034 = N3032 | N3033;
  assign N3032 = N3030 | N3031;
  assign N3030 = N3028 | N3029;
  assign N3028 = N3026 | N3027;
  assign N3026 = in_v_i[15] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__15_ ;
  assign N3027 = in_v_i[14] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__14_ ;
  assign N3029 = in_v_i[13] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__13_ ;
  assign N3031 = in_v_i[12] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__12_ ;
  assign N3033 = in_v_i[11] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__11_ ;
  assign N3035 = in_v_i[10] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__10_ ;
  assign N3037 = in_v_i[9] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__9_ ;
  assign N3039 = in_v_i[8] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__8_ ;
  assign N3041 = in_v_i[7] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__7_ ;
  assign N3043 = in_v_i[6] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__6_ ;
  assign N3045 = in_v_i[5] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__5_ ;
  assign N3047 = in_v_i[4] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__4_ ;
  assign N3049 = in_v_i[3] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__3_ ;
  assign N3051 = in_v_i[2] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__2_ ;
  assign N3053 = in_v_i[1] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__1_ ;
  assign N3055 = in_v_i[0] & \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__0_ ;
  assign N2452 = ~bk_sel_r[60];
  assign N2453 = ~bk_sel_r[61];
  assign N2454 = N2452 & N2453;
  assign N2455 = N2452 & bk_sel_r[61];
  assign N2456 = bk_sel_r[60] & N2453;
  assign N2457 = bk_sel_r[60] & bk_sel_r[61];
  assign N2458 = ~bk_sel_r[62];
  assign N2459 = N2454 & N2458;
  assign N2460 = N2454 & bk_sel_r[62];
  assign N2461 = N2456 & N2458;
  assign N2462 = N2456 & bk_sel_r[62];
  assign N2463 = N2455 & N2458;
  assign N2464 = N2455 & bk_sel_r[62];
  assign N2465 = N2457 & N2458;
  assign N2466 = N2457 & bk_sel_r[62];
  assign N2467 = ~bk_sel_r[63];
  assign N2468 = N2459 & N2467;
  assign N2469 = N2459 & bk_sel_r[63];
  assign N2470 = N2461 & N2467;
  assign N2471 = N2461 & bk_sel_r[63];
  assign N2472 = N2463 & N2467;
  assign N2473 = N2463 & bk_sel_r[63];
  assign N2474 = N2465 & N2467;
  assign N2475 = N2465 & bk_sel_r[63];
  assign N2476 = N2460 & N2467;
  assign N2477 = N2460 & bk_sel_r[63];
  assign N2478 = N2462 & N2467;
  assign N2479 = N2462 & bk_sel_r[63];
  assign N2480 = N2464 & N2467;
  assign N2481 = N2464 & bk_sel_r[63];
  assign N2482 = N2466 & N2467;
  assign N2483 = N2466 & bk_sel_r[63];
  assign N2484 = N2452 & N2453;
  assign N2485 = N2452 & bk_sel_r[61];
  assign N2486 = bk_sel_r[60] & N2453;
  assign N2487 = bk_sel_r[60] & bk_sel_r[61];
  assign N2488 = N2484 & N2458;
  assign N2489 = N2484 & bk_sel_r[62];
  assign N2490 = N2486 & N2458;
  assign N2491 = N2486 & bk_sel_r[62];
  assign N2492 = N2485 & N2458;
  assign N2493 = N2485 & bk_sel_r[62];
  assign N2494 = N2487 & N2458;
  assign N2495 = N2487 & bk_sel_r[62];
  assign N2496 = N2488 & N2467;
  assign N2497 = N2488 & bk_sel_r[63];
  assign N2498 = N2490 & N2467;
  assign N2499 = N2490 & bk_sel_r[63];
  assign N2500 = N2492 & N2467;
  assign N2501 = N2492 & bk_sel_r[63];
  assign N2502 = N2494 & N2467;
  assign N2503 = N2494 & bk_sel_r[63];
  assign N2504 = N2489 & N2467;
  assign N2505 = N2489 & bk_sel_r[63];
  assign N2506 = N2491 & N2467;
  assign N2507 = N2491 & bk_sel_r[63];
  assign N2508 = N2493 & N2467;
  assign N2509 = N2493 & bk_sel_r[63];
  assign N2510 = N2495 & N2467;
  assign N2511 = N2495 & bk_sel_r[63];
  assign N2512 = ~fwd_sel_r[60];
  assign N2513 = ~fwd_sel_r[61];
  assign N2514 = N2512 & N2513;
  assign N2515 = N2512 & fwd_sel_r[61];
  assign N2516 = fwd_sel_r[60] & N2513;
  assign N2517 = fwd_sel_r[60] & fwd_sel_r[61];
  assign N2518 = ~fwd_sel_r[62];
  assign N2519 = N2514 & N2518;
  assign N2520 = N2514 & fwd_sel_r[62];
  assign N2521 = N2516 & N2518;
  assign N2522 = N2516 & fwd_sel_r[62];
  assign N2523 = N2515 & N2518;
  assign N2524 = N2515 & fwd_sel_r[62];
  assign N2525 = N2517 & N2518;
  assign N2526 = N2517 & fwd_sel_r[62];
  assign N2527 = ~fwd_sel_r[63];
  assign N2528 = N2519 & N2527;
  assign N2529 = N2519 & fwd_sel_r[63];
  assign N2530 = N2521 & N2527;
  assign N2531 = N2521 & fwd_sel_r[63];
  assign N2532 = N2523 & N2527;
  assign N2533 = N2523 & fwd_sel_r[63];
  assign N2534 = N2525 & N2527;
  assign N2535 = N2525 & fwd_sel_r[63];
  assign N2536 = N2520 & N2527;
  assign N2537 = N2520 & fwd_sel_r[63];
  assign N2538 = N2522 & N2527;
  assign N2539 = N2522 & fwd_sel_r[63];
  assign N2540 = N2524 & N2527;
  assign N2541 = N2524 & fwd_sel_r[63];
  assign N2542 = N2526 & N2527;
  assign N2543 = N2526 & fwd_sel_r[63];
  assign N2544 = ~bk_dpath_sel_r[60];
  assign N2545 = ~bk_dpath_sel_r[61];
  assign N2546 = N2544 & N2545;
  assign N2547 = N2544 & bk_dpath_sel_r[61];
  assign N2548 = bk_dpath_sel_r[60] & N2545;
  assign N2549 = bk_dpath_sel_r[60] & bk_dpath_sel_r[61];
  assign N2550 = ~bk_dpath_sel_r[62];
  assign N2551 = N2546 & N2550;
  assign N2552 = N2546 & bk_dpath_sel_r[62];
  assign N2553 = N2548 & N2550;
  assign N2554 = N2548 & bk_dpath_sel_r[62];
  assign N2555 = N2547 & N2550;
  assign N2556 = N2547 & bk_dpath_sel_r[62];
  assign N2557 = N2549 & N2550;
  assign N2558 = N2549 & bk_dpath_sel_r[62];
  assign N2559 = ~bk_dpath_sel_r[63];
  assign N2560 = N2551 & N2559;
  assign N2561 = N2551 & bk_dpath_sel_r[63];
  assign N2562 = N2553 & N2559;
  assign N2563 = N2553 & bk_dpath_sel_r[63];
  assign N2564 = N2555 & N2559;
  assign N2565 = N2555 & bk_dpath_sel_r[63];
  assign N2566 = N2557 & N2559;
  assign N2567 = N2557 & bk_dpath_sel_r[63];
  assign N2568 = N2552 & N2559;
  assign N2569 = N2552 & bk_dpath_sel_r[63];
  assign N2570 = N2554 & N2559;
  assign N2571 = N2554 & bk_dpath_sel_r[63];
  assign N2572 = N2556 & N2559;
  assign N2573 = N2556 & bk_dpath_sel_r[63];
  assign N2574 = N2558 & N2559;
  assign N2575 = N2558 & bk_dpath_sel_r[63];

  always @(posedge clk_i) begin
    if(1'b1) begin
      fwd_sel_r_63_sv2v_reg <= fwd_sel[63];
      fwd_sel_r_62_sv2v_reg <= fwd_sel[62];
      fwd_sel_r_61_sv2v_reg <= fwd_sel[61];
      fwd_sel_r_60_sv2v_reg <= fwd_sel[60];
      fwd_sel_r_59_sv2v_reg <= fwd_sel[59];
      fwd_sel_r_58_sv2v_reg <= fwd_sel[58];
      fwd_sel_r_57_sv2v_reg <= fwd_sel[57];
      fwd_sel_r_56_sv2v_reg <= fwd_sel[56];
      fwd_sel_r_55_sv2v_reg <= fwd_sel[55];
      fwd_sel_r_54_sv2v_reg <= fwd_sel[54];
      fwd_sel_r_53_sv2v_reg <= fwd_sel[53];
      fwd_sel_r_52_sv2v_reg <= fwd_sel[52];
      fwd_sel_r_51_sv2v_reg <= fwd_sel[51];
      fwd_sel_r_50_sv2v_reg <= fwd_sel[50];
      fwd_sel_r_49_sv2v_reg <= fwd_sel[49];
      fwd_sel_r_48_sv2v_reg <= fwd_sel[48];
      fwd_sel_r_47_sv2v_reg <= fwd_sel[47];
      fwd_sel_r_46_sv2v_reg <= fwd_sel[46];
      fwd_sel_r_45_sv2v_reg <= fwd_sel[45];
      fwd_sel_r_44_sv2v_reg <= fwd_sel[44];
      fwd_sel_r_43_sv2v_reg <= fwd_sel[43];
      fwd_sel_r_42_sv2v_reg <= fwd_sel[42];
      fwd_sel_r_41_sv2v_reg <= fwd_sel[41];
      fwd_sel_r_40_sv2v_reg <= fwd_sel[40];
      fwd_sel_r_39_sv2v_reg <= fwd_sel[39];
      fwd_sel_r_38_sv2v_reg <= fwd_sel[38];
      fwd_sel_r_37_sv2v_reg <= fwd_sel[37];
      fwd_sel_r_36_sv2v_reg <= fwd_sel[36];
      fwd_sel_r_35_sv2v_reg <= fwd_sel[35];
      fwd_sel_r_34_sv2v_reg <= fwd_sel[34];
      fwd_sel_r_33_sv2v_reg <= fwd_sel[33];
      fwd_sel_r_32_sv2v_reg <= fwd_sel[32];
      fwd_sel_r_31_sv2v_reg <= fwd_sel[31];
      fwd_sel_r_30_sv2v_reg <= fwd_sel[30];
      fwd_sel_r_29_sv2v_reg <= fwd_sel[29];
      fwd_sel_r_28_sv2v_reg <= fwd_sel[28];
      fwd_sel_r_27_sv2v_reg <= fwd_sel[27];
      fwd_sel_r_26_sv2v_reg <= fwd_sel[26];
      fwd_sel_r_25_sv2v_reg <= fwd_sel[25];
      fwd_sel_r_24_sv2v_reg <= fwd_sel[24];
      fwd_sel_r_23_sv2v_reg <= fwd_sel[23];
      fwd_sel_r_22_sv2v_reg <= fwd_sel[22];
      fwd_sel_r_21_sv2v_reg <= fwd_sel[21];
      fwd_sel_r_20_sv2v_reg <= fwd_sel[20];
      fwd_sel_r_19_sv2v_reg <= fwd_sel[19];
      fwd_sel_r_18_sv2v_reg <= fwd_sel[18];
      fwd_sel_r_17_sv2v_reg <= fwd_sel[17];
      fwd_sel_r_16_sv2v_reg <= fwd_sel[16];
      fwd_sel_r_15_sv2v_reg <= fwd_sel[15];
      fwd_sel_r_14_sv2v_reg <= fwd_sel[14];
      fwd_sel_r_13_sv2v_reg <= fwd_sel[13];
      fwd_sel_r_12_sv2v_reg <= fwd_sel[12];
      fwd_sel_r_11_sv2v_reg <= fwd_sel[11];
      fwd_sel_r_10_sv2v_reg <= fwd_sel[10];
      fwd_sel_r_9_sv2v_reg <= fwd_sel[9];
      fwd_sel_r_8_sv2v_reg <= fwd_sel[8];
      fwd_sel_r_7_sv2v_reg <= fwd_sel[7];
      fwd_sel_r_6_sv2v_reg <= fwd_sel[6];
      fwd_sel_r_5_sv2v_reg <= fwd_sel[5];
      fwd_sel_r_4_sv2v_reg <= fwd_sel[4];
      fwd_sel_r_3_sv2v_reg <= fwd_sel[3];
      fwd_sel_r_2_sv2v_reg <= fwd_sel[2];
      fwd_sel_r_1_sv2v_reg <= fwd_sel[1];
      fwd_sel_r_0_sv2v_reg <= fwd_sel[0];
      fwd_dpath_sel_r_56_sv2v_reg <= fwd_dpath_sel[56];
      fwd_dpath_sel_r_53_sv2v_reg <= fwd_dpath_sel[53];
      fwd_dpath_sel_r_52_sv2v_reg <= fwd_dpath_sel[52];
      fwd_dpath_sel_r_49_sv2v_reg <= fwd_dpath_sel[49];
      fwd_dpath_sel_r_48_sv2v_reg <= fwd_dpath_sel[48];
      fwd_dpath_sel_r_46_sv2v_reg <= fwd_dpath_sel[46];
      fwd_dpath_sel_r_45_sv2v_reg <= fwd_dpath_sel[45];
      fwd_dpath_sel_r_44_sv2v_reg <= fwd_dpath_sel[44];
      fwd_dpath_sel_r_42_sv2v_reg <= fwd_dpath_sel[42];
      fwd_dpath_sel_r_41_sv2v_reg <= fwd_dpath_sel[41];
      fwd_dpath_sel_r_40_sv2v_reg <= fwd_dpath_sel[40];
      fwd_dpath_sel_r_38_sv2v_reg <= fwd_dpath_sel[38];
      fwd_dpath_sel_r_37_sv2v_reg <= fwd_dpath_sel[37];
      fwd_dpath_sel_r_36_sv2v_reg <= fwd_dpath_sel[36];
      fwd_dpath_sel_r_34_sv2v_reg <= fwd_dpath_sel[34];
      fwd_dpath_sel_r_33_sv2v_reg <= fwd_dpath_sel[33];
      fwd_dpath_sel_r_32_sv2v_reg <= fwd_dpath_sel[32];
      fwd_dpath_sel_r_31_sv2v_reg <= fwd_dpath_sel[31];
      fwd_dpath_sel_r_30_sv2v_reg <= fwd_dpath_sel[30];
      fwd_dpath_sel_r_29_sv2v_reg <= fwd_dpath_sel[29];
      fwd_dpath_sel_r_28_sv2v_reg <= fwd_dpath_sel[28];
      fwd_dpath_sel_r_27_sv2v_reg <= fwd_dpath_sel[27];
      fwd_dpath_sel_r_26_sv2v_reg <= fwd_dpath_sel[26];
      fwd_dpath_sel_r_25_sv2v_reg <= fwd_dpath_sel[25];
      fwd_dpath_sel_r_24_sv2v_reg <= fwd_dpath_sel[24];
      fwd_dpath_sel_r_23_sv2v_reg <= fwd_dpath_sel[23];
      fwd_dpath_sel_r_22_sv2v_reg <= fwd_dpath_sel[22];
      fwd_dpath_sel_r_21_sv2v_reg <= fwd_dpath_sel[21];
      fwd_dpath_sel_r_20_sv2v_reg <= fwd_dpath_sel[20];
      fwd_dpath_sel_r_19_sv2v_reg <= fwd_dpath_sel[19];
      fwd_dpath_sel_r_18_sv2v_reg <= fwd_dpath_sel[18];
      fwd_dpath_sel_r_17_sv2v_reg <= fwd_dpath_sel[17];
      fwd_dpath_sel_r_16_sv2v_reg <= fwd_dpath_sel[16];
      fwd_dpath_sel_r_15_sv2v_reg <= fwd_dpath_sel[15];
      fwd_dpath_sel_r_14_sv2v_reg <= fwd_dpath_sel[14];
      fwd_dpath_sel_r_13_sv2v_reg <= fwd_dpath_sel[13];
      fwd_dpath_sel_r_12_sv2v_reg <= fwd_dpath_sel[12];
      fwd_dpath_sel_r_11_sv2v_reg <= fwd_dpath_sel[11];
      fwd_dpath_sel_r_10_sv2v_reg <= fwd_dpath_sel[10];
      fwd_dpath_sel_r_9_sv2v_reg <= fwd_dpath_sel[9];
      fwd_dpath_sel_r_8_sv2v_reg <= fwd_dpath_sel[8];
      fwd_dpath_sel_r_7_sv2v_reg <= fwd_dpath_sel[7];
      fwd_dpath_sel_r_6_sv2v_reg <= fwd_dpath_sel[6];
      fwd_dpath_sel_r_5_sv2v_reg <= fwd_dpath_sel[5];
      fwd_dpath_sel_r_4_sv2v_reg <= fwd_dpath_sel[4];
      fwd_dpath_sel_r_3_sv2v_reg <= fwd_dpath_sel[3];
      fwd_dpath_sel_r_2_sv2v_reg <= fwd_dpath_sel[2];
      fwd_dpath_sel_r_1_sv2v_reg <= fwd_dpath_sel[1];
      fwd_dpath_sel_r_0_sv2v_reg <= fwd_dpath_sel[0];
      bk_sel_r_63_sv2v_reg <= bk_sel[63];
      bk_sel_r_62_sv2v_reg <= bk_sel[62];
      bk_sel_r_61_sv2v_reg <= bk_sel[61];
      bk_sel_r_60_sv2v_reg <= bk_sel[60];
      bk_sel_r_59_sv2v_reg <= bk_sel[59];
      bk_sel_r_58_sv2v_reg <= bk_sel[58];
      bk_sel_r_57_sv2v_reg <= bk_sel[57];
      bk_sel_r_56_sv2v_reg <= bk_sel[56];
      bk_sel_r_55_sv2v_reg <= bk_sel[55];
      bk_sel_r_54_sv2v_reg <= bk_sel[54];
      bk_sel_r_53_sv2v_reg <= bk_sel[53];
      bk_sel_r_52_sv2v_reg <= bk_sel[52];
      bk_sel_r_51_sv2v_reg <= bk_sel[51];
      bk_sel_r_50_sv2v_reg <= bk_sel[50];
      bk_sel_r_49_sv2v_reg <= bk_sel[49];
      bk_sel_r_48_sv2v_reg <= bk_sel[48];
      bk_sel_r_47_sv2v_reg <= bk_sel[47];
      bk_sel_r_46_sv2v_reg <= bk_sel[46];
      bk_sel_r_45_sv2v_reg <= bk_sel[45];
      bk_sel_r_44_sv2v_reg <= bk_sel[44];
      bk_sel_r_43_sv2v_reg <= bk_sel[43];
      bk_sel_r_42_sv2v_reg <= bk_sel[42];
      bk_sel_r_41_sv2v_reg <= bk_sel[41];
      bk_sel_r_40_sv2v_reg <= bk_sel[40];
      bk_sel_r_39_sv2v_reg <= bk_sel[39];
      bk_sel_r_38_sv2v_reg <= bk_sel[38];
      bk_sel_r_37_sv2v_reg <= bk_sel[37];
      bk_sel_r_36_sv2v_reg <= bk_sel[36];
      bk_sel_r_35_sv2v_reg <= bk_sel[35];
      bk_sel_r_34_sv2v_reg <= bk_sel[34];
      bk_sel_r_33_sv2v_reg <= bk_sel[33];
      bk_sel_r_32_sv2v_reg <= bk_sel[32];
      bk_sel_r_31_sv2v_reg <= bk_sel[31];
      bk_sel_r_30_sv2v_reg <= bk_sel[30];
      bk_sel_r_29_sv2v_reg <= bk_sel[29];
      bk_sel_r_28_sv2v_reg <= bk_sel[28];
      bk_sel_r_27_sv2v_reg <= bk_sel[27];
      bk_sel_r_26_sv2v_reg <= bk_sel[26];
      bk_sel_r_25_sv2v_reg <= bk_sel[25];
      bk_sel_r_24_sv2v_reg <= bk_sel[24];
      bk_sel_r_23_sv2v_reg <= bk_sel[23];
      bk_sel_r_22_sv2v_reg <= bk_sel[22];
      bk_sel_r_21_sv2v_reg <= bk_sel[21];
      bk_sel_r_20_sv2v_reg <= bk_sel[20];
      bk_sel_r_19_sv2v_reg <= bk_sel[19];
      bk_sel_r_18_sv2v_reg <= bk_sel[18];
      bk_sel_r_17_sv2v_reg <= bk_sel[17];
      bk_sel_r_16_sv2v_reg <= bk_sel[16];
      bk_sel_r_15_sv2v_reg <= bk_sel[15];
      bk_sel_r_14_sv2v_reg <= bk_sel[14];
      bk_sel_r_13_sv2v_reg <= bk_sel[13];
      bk_sel_r_12_sv2v_reg <= bk_sel[12];
      bk_sel_r_11_sv2v_reg <= bk_sel[11];
      bk_sel_r_10_sv2v_reg <= bk_sel[10];
      bk_sel_r_9_sv2v_reg <= bk_sel[9];
      bk_sel_r_8_sv2v_reg <= bk_sel[8];
      bk_sel_r_7_sv2v_reg <= bk_sel[7];
      bk_sel_r_6_sv2v_reg <= bk_sel[6];
      bk_sel_r_5_sv2v_reg <= bk_sel[5];
      bk_sel_r_4_sv2v_reg <= bk_sel[4];
      bk_sel_r_3_sv2v_reg <= bk_sel[3];
      bk_sel_r_2_sv2v_reg <= bk_sel[2];
      bk_sel_r_1_sv2v_reg <= bk_sel[1];
      bk_sel_r_0_sv2v_reg <= bk_sel[0];
      bk_dpath_sel_r_63_sv2v_reg <= bk_dpath_sel[63];
      bk_dpath_sel_r_62_sv2v_reg <= bk_dpath_sel[62];
      bk_dpath_sel_r_61_sv2v_reg <= bk_dpath_sel[61];
      bk_dpath_sel_r_60_sv2v_reg <= bk_dpath_sel[60];
      bk_dpath_sel_r_59_sv2v_reg <= bk_dpath_sel[59];
      bk_dpath_sel_r_58_sv2v_reg <= bk_dpath_sel[58];
      bk_dpath_sel_r_57_sv2v_reg <= bk_dpath_sel[57];
      bk_dpath_sel_r_56_sv2v_reg <= bk_dpath_sel[56];
      bk_dpath_sel_r_55_sv2v_reg <= bk_dpath_sel[55];
      bk_dpath_sel_r_54_sv2v_reg <= bk_dpath_sel[54];
      bk_dpath_sel_r_53_sv2v_reg <= bk_dpath_sel[53];
      bk_dpath_sel_r_52_sv2v_reg <= bk_dpath_sel[52];
      bk_dpath_sel_r_51_sv2v_reg <= bk_dpath_sel[51];
      bk_dpath_sel_r_50_sv2v_reg <= bk_dpath_sel[50];
      bk_dpath_sel_r_49_sv2v_reg <= bk_dpath_sel[49];
      bk_dpath_sel_r_48_sv2v_reg <= bk_dpath_sel[48];
      bk_dpath_sel_r_47_sv2v_reg <= bk_dpath_sel[47];
      bk_dpath_sel_r_46_sv2v_reg <= bk_dpath_sel[46];
      bk_dpath_sel_r_45_sv2v_reg <= bk_dpath_sel[45];
      bk_dpath_sel_r_44_sv2v_reg <= bk_dpath_sel[44];
      bk_dpath_sel_r_43_sv2v_reg <= bk_dpath_sel[43];
      bk_dpath_sel_r_42_sv2v_reg <= bk_dpath_sel[42];
      bk_dpath_sel_r_41_sv2v_reg <= bk_dpath_sel[41];
      bk_dpath_sel_r_40_sv2v_reg <= bk_dpath_sel[40];
      bk_dpath_sel_r_39_sv2v_reg <= bk_dpath_sel[39];
      bk_dpath_sel_r_38_sv2v_reg <= bk_dpath_sel[38];
      bk_dpath_sel_r_37_sv2v_reg <= bk_dpath_sel[37];
      bk_dpath_sel_r_36_sv2v_reg <= bk_dpath_sel[36];
      bk_dpath_sel_r_35_sv2v_reg <= bk_dpath_sel[35];
      bk_dpath_sel_r_34_sv2v_reg <= bk_dpath_sel[34];
      bk_dpath_sel_r_33_sv2v_reg <= bk_dpath_sel[33];
      bk_dpath_sel_r_32_sv2v_reg <= bk_dpath_sel[32];
      bk_dpath_sel_r_30_sv2v_reg <= bk_dpath_sel[30];
      bk_dpath_sel_r_29_sv2v_reg <= bk_dpath_sel[29];
      bk_dpath_sel_r_28_sv2v_reg <= bk_dpath_sel[28];
      bk_dpath_sel_r_26_sv2v_reg <= bk_dpath_sel[26];
      bk_dpath_sel_r_25_sv2v_reg <= bk_dpath_sel[25];
      bk_dpath_sel_r_24_sv2v_reg <= bk_dpath_sel[24];
      bk_dpath_sel_r_22_sv2v_reg <= bk_dpath_sel[22];
      bk_dpath_sel_r_21_sv2v_reg <= bk_dpath_sel[21];
      bk_dpath_sel_r_20_sv2v_reg <= bk_dpath_sel[20];
      bk_dpath_sel_r_18_sv2v_reg <= bk_dpath_sel[18];
      bk_dpath_sel_r_17_sv2v_reg <= bk_dpath_sel[17];
      bk_dpath_sel_r_16_sv2v_reg <= bk_dpath_sel[16];
      bk_dpath_sel_r_13_sv2v_reg <= bk_dpath_sel[13];
      bk_dpath_sel_r_12_sv2v_reg <= bk_dpath_sel[12];
      bk_dpath_sel_r_9_sv2v_reg <= bk_dpath_sel[9];
      bk_dpath_sel_r_8_sv2v_reg <= bk_dpath_sel[8];
      bk_dpath_sel_r_4_sv2v_reg <= bk_dpath_sel[4];
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__15__sv2v_reg  <= N553;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__14__sv2v_reg  <= N552;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__13__sv2v_reg  <= N551;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__12__sv2v_reg  <= N550;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__11__sv2v_reg  <= N549;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__10__sv2v_reg  <= N548;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__9__sv2v_reg  <= N547;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__8__sv2v_reg  <= N546;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__7__sv2v_reg  <= N545;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__6__sv2v_reg  <= N544;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__5__sv2v_reg  <= N543;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__4__sv2v_reg  <= N542;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__3__sv2v_reg  <= N541;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__2__sv2v_reg  <= N540;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__1__sv2v_reg  <= N539;
      \sbox_0_.fi1hot.fwd_sel_one_hot_r_0__0__sv2v_reg  <= N538;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__15__sv2v_reg  <= N693;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__14__sv2v_reg  <= N692;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__13__sv2v_reg  <= N691;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__12__sv2v_reg  <= N690;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__11__sv2v_reg  <= N689;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__10__sv2v_reg  <= N688;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__9__sv2v_reg  <= N687;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__8__sv2v_reg  <= N686;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__7__sv2v_reg  <= N685;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__6__sv2v_reg  <= N684;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__5__sv2v_reg  <= N683;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__4__sv2v_reg  <= N682;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__3__sv2v_reg  <= N681;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__2__sv2v_reg  <= N680;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__1__sv2v_reg  <= N679;
      \sbox_1_.fi1hot.fwd_sel_one_hot_r_1__0__sv2v_reg  <= N678;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__15__sv2v_reg  <= N817;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__14__sv2v_reg  <= N816;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__13__sv2v_reg  <= N815;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__12__sv2v_reg  <= N814;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__11__sv2v_reg  <= N813;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__10__sv2v_reg  <= N812;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__9__sv2v_reg  <= N811;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__8__sv2v_reg  <= N810;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__7__sv2v_reg  <= N809;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__6__sv2v_reg  <= N808;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__5__sv2v_reg  <= N807;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__4__sv2v_reg  <= N806;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__3__sv2v_reg  <= N805;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__2__sv2v_reg  <= N804;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__1__sv2v_reg  <= N803;
      \sbox_2_.fi1hot.fwd_sel_one_hot_r_2__0__sv2v_reg  <= N802;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__15__sv2v_reg  <= N940;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__14__sv2v_reg  <= N939;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__13__sv2v_reg  <= N938;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__12__sv2v_reg  <= N937;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__11__sv2v_reg  <= N936;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__10__sv2v_reg  <= N935;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__9__sv2v_reg  <= N934;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__8__sv2v_reg  <= N933;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__7__sv2v_reg  <= N932;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__6__sv2v_reg  <= N931;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__5__sv2v_reg  <= N930;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__4__sv2v_reg  <= N929;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__3__sv2v_reg  <= N928;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__2__sv2v_reg  <= N927;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__1__sv2v_reg  <= N926;
      \sbox_3_.fi1hot.fwd_sel_one_hot_r_3__0__sv2v_reg  <= N925;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__15__sv2v_reg  <= N1067;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__14__sv2v_reg  <= N1066;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__13__sv2v_reg  <= N1065;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__12__sv2v_reg  <= N1064;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__11__sv2v_reg  <= N1063;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__10__sv2v_reg  <= N1062;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__9__sv2v_reg  <= N1061;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__8__sv2v_reg  <= N1060;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__7__sv2v_reg  <= N1059;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__6__sv2v_reg  <= N1058;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__5__sv2v_reg  <= N1057;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__4__sv2v_reg  <= N1056;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__3__sv2v_reg  <= N1055;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__2__sv2v_reg  <= N1054;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__1__sv2v_reg  <= N1053;
      \sbox_4_.fi1hot.fwd_sel_one_hot_r_4__0__sv2v_reg  <= N1052;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__15__sv2v_reg  <= N1191;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__14__sv2v_reg  <= N1190;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__13__sv2v_reg  <= N1189;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__12__sv2v_reg  <= N1188;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__11__sv2v_reg  <= N1187;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__10__sv2v_reg  <= N1186;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__9__sv2v_reg  <= N1185;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__8__sv2v_reg  <= N1184;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__7__sv2v_reg  <= N1183;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__6__sv2v_reg  <= N1182;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__5__sv2v_reg  <= N1181;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__4__sv2v_reg  <= N1180;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__3__sv2v_reg  <= N1179;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__2__sv2v_reg  <= N1178;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__1__sv2v_reg  <= N1177;
      \sbox_5_.fi1hot.fwd_sel_one_hot_r_5__0__sv2v_reg  <= N1176;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__15__sv2v_reg  <= N1316;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__14__sv2v_reg  <= N1315;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__13__sv2v_reg  <= N1314;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__12__sv2v_reg  <= N1313;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__11__sv2v_reg  <= N1312;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__10__sv2v_reg  <= N1311;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__9__sv2v_reg  <= N1310;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__8__sv2v_reg  <= N1309;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__7__sv2v_reg  <= N1308;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__6__sv2v_reg  <= N1307;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__5__sv2v_reg  <= N1306;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__4__sv2v_reg  <= N1305;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__3__sv2v_reg  <= N1304;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__2__sv2v_reg  <= N1303;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__1__sv2v_reg  <= N1302;
      \sbox_6_.fi1hot.fwd_sel_one_hot_r_6__0__sv2v_reg  <= N1301;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__15__sv2v_reg  <= N1441;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__14__sv2v_reg  <= N1440;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__13__sv2v_reg  <= N1439;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__12__sv2v_reg  <= N1438;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__11__sv2v_reg  <= N1437;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__10__sv2v_reg  <= N1436;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__9__sv2v_reg  <= N1435;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__8__sv2v_reg  <= N1434;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__7__sv2v_reg  <= N1433;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__6__sv2v_reg  <= N1432;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__5__sv2v_reg  <= N1431;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__4__sv2v_reg  <= N1430;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__3__sv2v_reg  <= N1429;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__2__sv2v_reg  <= N1428;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__1__sv2v_reg  <= N1427;
      \sbox_7_.fi1hot.fwd_sel_one_hot_r_7__0__sv2v_reg  <= N1426;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__15__sv2v_reg  <= N1572;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__14__sv2v_reg  <= N1571;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__13__sv2v_reg  <= N1570;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__12__sv2v_reg  <= N1569;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__11__sv2v_reg  <= N1568;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__10__sv2v_reg  <= N1567;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__9__sv2v_reg  <= N1566;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__8__sv2v_reg  <= N1565;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__7__sv2v_reg  <= N1564;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__6__sv2v_reg  <= N1563;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__5__sv2v_reg  <= N1562;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__4__sv2v_reg  <= N1561;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__3__sv2v_reg  <= N1560;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__2__sv2v_reg  <= N1559;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__1__sv2v_reg  <= N1558;
      \sbox_8_.fi1hot.fwd_sel_one_hot_r_8__0__sv2v_reg  <= N1557;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__15__sv2v_reg  <= N1703;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__14__sv2v_reg  <= N1702;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__13__sv2v_reg  <= N1701;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__12__sv2v_reg  <= N1700;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__11__sv2v_reg  <= N1699;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__10__sv2v_reg  <= N1698;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__9__sv2v_reg  <= N1697;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__8__sv2v_reg  <= N1696;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__7__sv2v_reg  <= N1695;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__6__sv2v_reg  <= N1694;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__5__sv2v_reg  <= N1693;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__4__sv2v_reg  <= N1692;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__3__sv2v_reg  <= N1691;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__2__sv2v_reg  <= N1690;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__1__sv2v_reg  <= N1689;
      \sbox_9_.fi1hot.fwd_sel_one_hot_r_9__0__sv2v_reg  <= N1688;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__15__sv2v_reg  <= N1828;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__14__sv2v_reg  <= N1827;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__13__sv2v_reg  <= N1826;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__12__sv2v_reg  <= N1825;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__11__sv2v_reg  <= N1824;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__10__sv2v_reg  <= N1823;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__9__sv2v_reg  <= N1822;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__8__sv2v_reg  <= N1821;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__7__sv2v_reg  <= N1820;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__6__sv2v_reg  <= N1819;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__5__sv2v_reg  <= N1818;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__4__sv2v_reg  <= N1817;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__3__sv2v_reg  <= N1816;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__2__sv2v_reg  <= N1815;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__1__sv2v_reg  <= N1814;
      \sbox_10_.fi1hot.fwd_sel_one_hot_r_10__0__sv2v_reg  <= N1813;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__15__sv2v_reg  <= N1953;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__14__sv2v_reg  <= N1952;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__13__sv2v_reg  <= N1951;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__12__sv2v_reg  <= N1950;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__11__sv2v_reg  <= N1949;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__10__sv2v_reg  <= N1948;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__9__sv2v_reg  <= N1947;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__8__sv2v_reg  <= N1946;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__7__sv2v_reg  <= N1945;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__6__sv2v_reg  <= N1944;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__5__sv2v_reg  <= N1943;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__4__sv2v_reg  <= N1942;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__3__sv2v_reg  <= N1941;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__2__sv2v_reg  <= N1940;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__1__sv2v_reg  <= N1939;
      \sbox_11_.fi1hot.fwd_sel_one_hot_r_11__0__sv2v_reg  <= N1938;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__15__sv2v_reg  <= N2077;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__14__sv2v_reg  <= N2076;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__13__sv2v_reg  <= N2075;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__12__sv2v_reg  <= N2074;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__11__sv2v_reg  <= N2073;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__10__sv2v_reg  <= N2072;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__9__sv2v_reg  <= N2071;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__8__sv2v_reg  <= N2070;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__7__sv2v_reg  <= N2069;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__6__sv2v_reg  <= N2068;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__5__sv2v_reg  <= N2067;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__4__sv2v_reg  <= N2066;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__3__sv2v_reg  <= N2065;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__2__sv2v_reg  <= N2064;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__1__sv2v_reg  <= N2063;
      \sbox_12_.fi1hot.fwd_sel_one_hot_r_12__0__sv2v_reg  <= N2062;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__15__sv2v_reg  <= N2204;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__14__sv2v_reg  <= N2203;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__13__sv2v_reg  <= N2202;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__12__sv2v_reg  <= N2201;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__11__sv2v_reg  <= N2200;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__10__sv2v_reg  <= N2199;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__9__sv2v_reg  <= N2198;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__8__sv2v_reg  <= N2197;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__7__sv2v_reg  <= N2196;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__6__sv2v_reg  <= N2195;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__5__sv2v_reg  <= N2194;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__4__sv2v_reg  <= N2193;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__3__sv2v_reg  <= N2192;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__2__sv2v_reg  <= N2191;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__1__sv2v_reg  <= N2190;
      \sbox_13_.fi1hot.fwd_sel_one_hot_r_13__0__sv2v_reg  <= N2189;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__15__sv2v_reg  <= N2327;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__14__sv2v_reg  <= N2326;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__13__sv2v_reg  <= N2325;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__12__sv2v_reg  <= N2324;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__11__sv2v_reg  <= N2323;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__10__sv2v_reg  <= N2322;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__9__sv2v_reg  <= N2321;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__8__sv2v_reg  <= N2320;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__7__sv2v_reg  <= N2319;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__6__sv2v_reg  <= N2318;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__5__sv2v_reg  <= N2317;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__4__sv2v_reg  <= N2316;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__3__sv2v_reg  <= N2315;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__2__sv2v_reg  <= N2314;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__1__sv2v_reg  <= N2313;
      \sbox_14_.fi1hot.fwd_sel_one_hot_r_14__0__sv2v_reg  <= N2312;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__15__sv2v_reg  <= N2451;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__14__sv2v_reg  <= N2450;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__13__sv2v_reg  <= N2449;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__12__sv2v_reg  <= N2448;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__11__sv2v_reg  <= N2447;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__10__sv2v_reg  <= N2446;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__9__sv2v_reg  <= N2445;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__8__sv2v_reg  <= N2444;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__7__sv2v_reg  <= N2443;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__6__sv2v_reg  <= N2442;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__5__sv2v_reg  <= N2441;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__4__sv2v_reg  <= N2440;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__3__sv2v_reg  <= N2439;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__2__sv2v_reg  <= N2438;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__1__sv2v_reg  <= N2437;
      \sbox_15_.fi1hot.fwd_sel_one_hot_r_15__0__sv2v_reg  <= N2436;
    end 
  end


endmodule

