

module top
(
  clk_i,
  reset_i,
  dma_data_o,
  dma_data_v_o,
  dma_data_ready_i,
  app_rd_data_valid_i,
  app_rd_data_end_i,
  app_rd_data_i
);

  output [31:0] dma_data_o;
  input [31:0] app_rd_data_i;
  input clk_i;
  input reset_i;
  input dma_data_ready_i;
  input app_rd_data_valid_i;
  input app_rd_data_end_i;
  output dma_data_v_o;

  bsg_cache_to_dram_ctrl_rx
  wrapper
  (
    .dma_data_o(dma_data_o),
    .app_rd_data_i(app_rd_data_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .dma_data_ready_i(dma_data_ready_i),
    .app_rd_data_valid_i(app_rd_data_valid_i),
    .app_rd_data_end_i(app_rd_data_end_i),
    .dma_data_v_o(dma_data_v_o)
  );


endmodule



module bsg_serial_in_parallel_out_width_p32_els_p3_out_els_p2
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_cnt_i
);

  input [31:0] data_i;
  output [1:0] valid_o;
  output [63:0] data_o;
  input [1:0] yumi_cnt_i;
  input clk_i;
  input reset_i;
  input valid_i;
  output ready_o;
  wire [1:0] valid_o,num_els_r,num_els_n;
  wire [63:0] data_o;
  wire ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,data_n_3__31_,data_n_3__30_,data_n_3__29_,
  data_n_3__28_,data_n_3__27_,data_n_3__26_,data_n_3__25_,data_n_3__24_,data_n_3__23_,
  data_n_3__22_,data_n_3__21_,data_n_3__20_,data_n_3__19_,data_n_3__18_,
  data_n_3__17_,data_n_3__16_,data_n_3__15_,data_n_3__14_,data_n_3__13_,data_n_3__12_,
  data_n_3__11_,data_n_3__10_,data_n_3__9_,data_n_3__8_,data_n_3__7_,data_n_3__6_,
  data_n_3__5_,data_n_3__4_,data_n_3__3_,data_n_3__2_,data_n_3__1_,data_n_3__0_,
  data_n_2__31_,data_n_2__30_,data_n_2__29_,data_n_2__28_,data_n_2__27_,data_n_2__26_,
  data_n_2__25_,data_n_2__24_,data_n_2__23_,data_n_2__22_,data_n_2__21_,data_n_2__20_,
  data_n_2__19_,data_n_2__18_,data_n_2__17_,data_n_2__16_,data_n_2__15_,
  data_n_2__14_,data_n_2__13_,data_n_2__12_,data_n_2__11_,data_n_2__10_,data_n_2__9_,
  data_n_2__8_,data_n_2__7_,data_n_2__6_,data_n_2__5_,data_n_2__4_,data_n_2__3_,
  data_n_2__2_,data_n_2__1_,data_n_2__0_,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60;
  wire [2:0] valid_r,valid_nn;
  wire [95:0] data_r,data_nn;
  wire [3:2] valid_n;
  reg valid_r_2_sv2v_reg,valid_r_1_sv2v_reg,valid_r_0_sv2v_reg,num_els_r_1_sv2v_reg,
  num_els_r_0_sv2v_reg,data_r_95_sv2v_reg,data_r_94_sv2v_reg,data_r_93_sv2v_reg,
  data_r_92_sv2v_reg,data_r_91_sv2v_reg,data_r_90_sv2v_reg,data_r_89_sv2v_reg,
  data_r_88_sv2v_reg,data_r_87_sv2v_reg,data_r_86_sv2v_reg,data_r_85_sv2v_reg,
  data_r_84_sv2v_reg,data_r_83_sv2v_reg,data_r_82_sv2v_reg,data_r_81_sv2v_reg,
  data_r_80_sv2v_reg,data_r_79_sv2v_reg,data_r_78_sv2v_reg,data_r_77_sv2v_reg,data_r_76_sv2v_reg,
  data_r_75_sv2v_reg,data_r_74_sv2v_reg,data_r_73_sv2v_reg,data_r_72_sv2v_reg,
  data_r_71_sv2v_reg,data_r_70_sv2v_reg,data_r_69_sv2v_reg,data_r_68_sv2v_reg,
  data_r_67_sv2v_reg,data_r_66_sv2v_reg,data_r_65_sv2v_reg,data_r_64_sv2v_reg,
  data_r_63_sv2v_reg,data_r_62_sv2v_reg,data_r_61_sv2v_reg,data_r_60_sv2v_reg,
  data_r_59_sv2v_reg,data_r_58_sv2v_reg,data_r_57_sv2v_reg,data_r_56_sv2v_reg,data_r_55_sv2v_reg,
  data_r_54_sv2v_reg,data_r_53_sv2v_reg,data_r_52_sv2v_reg,data_r_51_sv2v_reg,
  data_r_50_sv2v_reg,data_r_49_sv2v_reg,data_r_48_sv2v_reg,data_r_47_sv2v_reg,
  data_r_46_sv2v_reg,data_r_45_sv2v_reg,data_r_44_sv2v_reg,data_r_43_sv2v_reg,
  data_r_42_sv2v_reg,data_r_41_sv2v_reg,data_r_40_sv2v_reg,data_r_39_sv2v_reg,
  data_r_38_sv2v_reg,data_r_37_sv2v_reg,data_r_36_sv2v_reg,data_r_35_sv2v_reg,data_r_34_sv2v_reg,
  data_r_33_sv2v_reg,data_r_32_sv2v_reg,data_r_31_sv2v_reg,data_r_30_sv2v_reg,
  data_r_29_sv2v_reg,data_r_28_sv2v_reg,data_r_27_sv2v_reg,data_r_26_sv2v_reg,
  data_r_25_sv2v_reg,data_r_24_sv2v_reg,data_r_23_sv2v_reg,data_r_22_sv2v_reg,
  data_r_21_sv2v_reg,data_r_20_sv2v_reg,data_r_19_sv2v_reg,data_r_18_sv2v_reg,data_r_17_sv2v_reg,
  data_r_16_sv2v_reg,data_r_15_sv2v_reg,data_r_14_sv2v_reg,data_r_13_sv2v_reg,
  data_r_12_sv2v_reg,data_r_11_sv2v_reg,data_r_10_sv2v_reg,data_r_9_sv2v_reg,
  data_r_8_sv2v_reg,data_r_7_sv2v_reg,data_r_6_sv2v_reg,data_r_5_sv2v_reg,
  data_r_4_sv2v_reg,data_r_3_sv2v_reg,data_r_2_sv2v_reg,data_r_1_sv2v_reg,data_r_0_sv2v_reg;
  assign valid_r[2] = valid_r_2_sv2v_reg;
  assign valid_r[1] = valid_r_1_sv2v_reg;
  assign valid_r[0] = valid_r_0_sv2v_reg;
  assign num_els_r[1] = num_els_r_1_sv2v_reg;
  assign num_els_r[0] = num_els_r_0_sv2v_reg;
  assign data_r[95] = data_r_95_sv2v_reg;
  assign data_r[94] = data_r_94_sv2v_reg;
  assign data_r[93] = data_r_93_sv2v_reg;
  assign data_r[92] = data_r_92_sv2v_reg;
  assign data_r[91] = data_r_91_sv2v_reg;
  assign data_r[90] = data_r_90_sv2v_reg;
  assign data_r[89] = data_r_89_sv2v_reg;
  assign data_r[88] = data_r_88_sv2v_reg;
  assign data_r[87] = data_r_87_sv2v_reg;
  assign data_r[86] = data_r_86_sv2v_reg;
  assign data_r[85] = data_r_85_sv2v_reg;
  assign data_r[84] = data_r_84_sv2v_reg;
  assign data_r[83] = data_r_83_sv2v_reg;
  assign data_r[82] = data_r_82_sv2v_reg;
  assign data_r[81] = data_r_81_sv2v_reg;
  assign data_r[80] = data_r_80_sv2v_reg;
  assign data_r[79] = data_r_79_sv2v_reg;
  assign data_r[78] = data_r_78_sv2v_reg;
  assign data_r[77] = data_r_77_sv2v_reg;
  assign data_r[76] = data_r_76_sv2v_reg;
  assign data_r[75] = data_r_75_sv2v_reg;
  assign data_r[74] = data_r_74_sv2v_reg;
  assign data_r[73] = data_r_73_sv2v_reg;
  assign data_r[72] = data_r_72_sv2v_reg;
  assign data_r[71] = data_r_71_sv2v_reg;
  assign data_r[70] = data_r_70_sv2v_reg;
  assign data_r[69] = data_r_69_sv2v_reg;
  assign data_r[68] = data_r_68_sv2v_reg;
  assign data_r[67] = data_r_67_sv2v_reg;
  assign data_r[66] = data_r_66_sv2v_reg;
  assign data_r[65] = data_r_65_sv2v_reg;
  assign data_r[64] = data_r_64_sv2v_reg;
  assign data_r[63] = data_r_63_sv2v_reg;
  assign data_r[62] = data_r_62_sv2v_reg;
  assign data_r[61] = data_r_61_sv2v_reg;
  assign data_r[60] = data_r_60_sv2v_reg;
  assign data_r[59] = data_r_59_sv2v_reg;
  assign data_r[58] = data_r_58_sv2v_reg;
  assign data_r[57] = data_r_57_sv2v_reg;
  assign data_r[56] = data_r_56_sv2v_reg;
  assign data_r[55] = data_r_55_sv2v_reg;
  assign data_r[54] = data_r_54_sv2v_reg;
  assign data_r[53] = data_r_53_sv2v_reg;
  assign data_r[52] = data_r_52_sv2v_reg;
  assign data_r[51] = data_r_51_sv2v_reg;
  assign data_r[50] = data_r_50_sv2v_reg;
  assign data_r[49] = data_r_49_sv2v_reg;
  assign data_r[48] = data_r_48_sv2v_reg;
  assign data_r[47] = data_r_47_sv2v_reg;
  assign data_r[46] = data_r_46_sv2v_reg;
  assign data_r[45] = data_r_45_sv2v_reg;
  assign data_r[44] = data_r_44_sv2v_reg;
  assign data_r[43] = data_r_43_sv2v_reg;
  assign data_r[42] = data_r_42_sv2v_reg;
  assign data_r[41] = data_r_41_sv2v_reg;
  assign data_r[40] = data_r_40_sv2v_reg;
  assign data_r[39] = data_r_39_sv2v_reg;
  assign data_r[38] = data_r_38_sv2v_reg;
  assign data_r[37] = data_r_37_sv2v_reg;
  assign data_r[36] = data_r_36_sv2v_reg;
  assign data_r[35] = data_r_35_sv2v_reg;
  assign data_r[34] = data_r_34_sv2v_reg;
  assign data_r[33] = data_r_33_sv2v_reg;
  assign data_r[32] = data_r_32_sv2v_reg;
  assign data_r[31] = data_r_31_sv2v_reg;
  assign data_r[30] = data_r_30_sv2v_reg;
  assign data_r[29] = data_r_29_sv2v_reg;
  assign data_r[28] = data_r_28_sv2v_reg;
  assign data_r[27] = data_r_27_sv2v_reg;
  assign data_r[26] = data_r_26_sv2v_reg;
  assign data_r[25] = data_r_25_sv2v_reg;
  assign data_r[24] = data_r_24_sv2v_reg;
  assign data_r[23] = data_r_23_sv2v_reg;
  assign data_r[22] = data_r_22_sv2v_reg;
  assign data_r[21] = data_r_21_sv2v_reg;
  assign data_r[20] = data_r_20_sv2v_reg;
  assign data_r[19] = data_r_19_sv2v_reg;
  assign data_r[18] = data_r_18_sv2v_reg;
  assign data_r[17] = data_r_17_sv2v_reg;
  assign data_r[16] = data_r_16_sv2v_reg;
  assign data_r[15] = data_r_15_sv2v_reg;
  assign data_r[14] = data_r_14_sv2v_reg;
  assign data_r[13] = data_r_13_sv2v_reg;
  assign data_r[12] = data_r_12_sv2v_reg;
  assign data_r[11] = data_r_11_sv2v_reg;
  assign data_r[10] = data_r_10_sv2v_reg;
  assign data_r[9] = data_r_9_sv2v_reg;
  assign data_r[8] = data_r_8_sv2v_reg;
  assign data_r[7] = data_r_7_sv2v_reg;
  assign data_r[6] = data_r_6_sv2v_reg;
  assign data_r[5] = data_r_5_sv2v_reg;
  assign data_r[4] = data_r_4_sv2v_reg;
  assign data_r[3] = data_r_3_sv2v_reg;
  assign data_r[2] = data_r_2_sv2v_reg;
  assign data_r[1] = data_r_1_sv2v_reg;
  assign data_r[0] = data_r_0_sv2v_reg;
  assign N60 = N52 | N55;
  assign { N28, N27 } = num_els_r + N26;
  assign num_els_n = { N28, N27 } - yumi_cnt_i;
  assign N32 = num_els_r[0] & num_els_r[1];
  assign N31 = N0 & num_els_r[1];
  assign N0 = ~num_els_r[0];
  assign N30 = num_els_r[0] & N1;
  assign N1 = ~num_els_r[1];
  assign N29 = N2 & N3;
  assign N2 = ~num_els_r[0];
  assign N3 = ~num_els_r[1];
  assign N40 = num_els_r[0] & num_els_r[1];
  assign N39 = N4 & num_els_r[1];
  assign N4 = ~num_els_r[0];
  assign N38 = num_els_r[0] & N5;
  assign N5 = ~num_els_r[1];
  assign N37 = N6 & N7;
  assign N6 = ~num_els_r[0];
  assign N7 = ~num_els_r[1];
  assign N52 = yumi_cnt_i[0] & yumi_cnt_i[1];
  assign N55 = N8 & yumi_cnt_i[1];
  assign N8 = ~yumi_cnt_i[0];
  assign N54 = yumi_cnt_i[0] & N9;
  assign N9 = ~yumi_cnt_i[1];
  assign N53 = N10 & N11;
  assign N10 = ~yumi_cnt_i[0];
  assign N11 = ~yumi_cnt_i[1];
  assign { data_o[0:0], data_o[1:1], data_o[2:2], data_o[3:3], data_o[4:4], data_o[5:5], data_o[6:6], data_o[7:7], data_o[8:8], data_o[9:9], data_o[10:10], data_o[11:11], data_o[12:12], data_o[13:13], data_o[14:14], data_o[15:15], data_o[16:16], data_o[17:17], data_o[18:18], data_o[19:19], data_o[20:20], data_o[21:21], data_o[22:22], data_o[23:23], data_o[24:24], data_o[25:25], data_o[26:26], data_o[27:27], data_o[28:28], data_o[29:29], data_o[30:30], data_o[31:31] } = (N12)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N33)? { data_r[0:0], data_r[1:1], data_r[2:2], data_r[3:3], data_r[4:4], data_r[5:5], data_r[6:6], data_r[7:7], data_r[8:8], data_r[9:9], data_r[10:10], data_r[11:11], data_r[12:12], data_r[13:13], data_r[14:14], data_r[15:15], data_r[16:16], data_r[17:17], data_r[18:18], data_r[19:19], data_r[20:20], data_r[21:21], data_r[22:22], data_r[23:23], data_r[24:24], data_r[25:25], data_r[26:26], data_r[27:27], data_r[28:28], data_r[29:29], data_r[30:30], data_r[31:31] } : 1'b0;
  assign N12 = N29;
  assign { data_o[32:32], data_o[33:33], data_o[34:34], data_o[35:35], data_o[36:36], data_o[37:37], data_o[38:38], data_o[39:39], data_o[40:40], data_o[41:41], data_o[42:42], data_o[43:43], data_o[44:44], data_o[45:45], data_o[46:46], data_o[47:47], data_o[48:48], data_o[49:49], data_o[50:50], data_o[51:51], data_o[52:52], data_o[53:53], data_o[54:54], data_o[55:55], data_o[56:56], data_o[57:57], data_o[58:58], data_o[59:59], data_o[60:60], data_o[61:61], data_o[62:62], data_o[63:63] } = (N13)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N34)? { data_r[32:32], data_r[33:33], data_r[34:34], data_r[35:35], data_r[36:36], data_r[37:37], data_r[38:38], data_r[39:39], data_r[40:40], data_r[41:41], data_r[42:42], data_r[43:43], data_r[44:44], data_r[45:45], data_r[46:46], data_r[47:47], data_r[48:48], data_r[49:49], data_r[50:50], data_r[51:51], data_r[52:52], data_r[53:53], data_r[54:54], data_r[55:55], data_r[56:56], data_r[57:57], data_r[58:58], data_r[59:59], data_r[60:60], data_r[61:61], data_r[62:62], data_r[63:63] } : 1'b0;
  assign N13 = N30;
  assign { data_n_2__0_, data_n_2__1_, data_n_2__2_, data_n_2__3_, data_n_2__4_, data_n_2__5_, data_n_2__6_, data_n_2__7_, data_n_2__8_, data_n_2__9_, data_n_2__10_, data_n_2__11_, data_n_2__12_, data_n_2__13_, data_n_2__14_, data_n_2__15_, data_n_2__16_, data_n_2__17_, data_n_2__18_, data_n_2__19_, data_n_2__20_, data_n_2__21_, data_n_2__22_, data_n_2__23_, data_n_2__24_, data_n_2__25_, data_n_2__26_, data_n_2__27_, data_n_2__28_, data_n_2__29_, data_n_2__30_, data_n_2__31_ } = (N14)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N35)? { data_r[64:64], data_r[65:65], data_r[66:66], data_r[67:67], data_r[68:68], data_r[69:69], data_r[70:70], data_r[71:71], data_r[72:72], data_r[73:73], data_r[74:74], data_r[75:75], data_r[76:76], data_r[77:77], data_r[78:78], data_r[79:79], data_r[80:80], data_r[81:81], data_r[82:82], data_r[83:83], data_r[84:84], data_r[85:85], data_r[86:86], data_r[87:87], data_r[88:88], data_r[89:89], data_r[90:90], data_r[91:91], data_r[92:92], data_r[93:93], data_r[94:94], data_r[95:95] } : 1'b0;
  assign N14 = N31;
  assign { data_n_3__0_, data_n_3__1_, data_n_3__2_, data_n_3__3_, data_n_3__4_, data_n_3__5_, data_n_3__6_, data_n_3__7_, data_n_3__8_, data_n_3__9_, data_n_3__10_, data_n_3__11_, data_n_3__12_, data_n_3__13_, data_n_3__14_, data_n_3__15_, data_n_3__16_, data_n_3__17_, data_n_3__18_, data_n_3__19_, data_n_3__20_, data_n_3__21_, data_n_3__22_, data_n_3__23_, data_n_3__24_, data_n_3__25_, data_n_3__26_, data_n_3__27_, data_n_3__28_, data_n_3__29_, data_n_3__30_, data_n_3__31_ } = (N15)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = N32;
  assign valid_o[0] = (N16)? N41 : 
                      (N42)? valid_r[0] : 1'b0;
  assign N16 = N37;
  assign valid_o[1] = (N17)? N41 : 
                      (N43)? valid_r[1] : 1'b0;
  assign N17 = N38;
  assign valid_n[2] = (N18)? N41 : 
                      (N44)? valid_r[2] : 1'b0;
  assign N18 = N39;
  assign valid_n[3] = (N19)? N41 : 
                      (N45)? 1'b0 : 1'b0;
  assign N19 = N40;
  assign data_nn[63:32] = (N20)? { data_n_3__31_, data_n_3__30_, data_n_3__29_, data_n_3__28_, data_n_3__27_, data_n_3__26_, data_n_3__25_, data_n_3__24_, data_n_3__23_, data_n_3__22_, data_n_3__21_, data_n_3__20_, data_n_3__19_, data_n_3__18_, data_n_3__17_, data_n_3__16_, data_n_3__15_, data_n_3__14_, data_n_3__13_, data_n_3__12_, data_n_3__11_, data_n_3__10_, data_n_3__9_, data_n_3__8_, data_n_3__7_, data_n_3__6_, data_n_3__5_, data_n_3__4_, data_n_3__3_, data_n_3__2_, data_n_3__1_, data_n_3__0_ } : 
                          (N21)? { data_n_2__31_, data_n_2__30_, data_n_2__29_, data_n_2__28_, data_n_2__27_, data_n_2__26_, data_n_2__25_, data_n_2__24_, data_n_2__23_, data_n_2__22_, data_n_2__21_, data_n_2__20_, data_n_2__19_, data_n_2__18_, data_n_2__17_, data_n_2__16_, data_n_2__15_, data_n_2__14_, data_n_2__13_, data_n_2__12_, data_n_2__11_, data_n_2__10_, data_n_2__9_, data_n_2__8_, data_n_2__7_, data_n_2__6_, data_n_2__5_, data_n_2__4_, data_n_2__3_, data_n_2__2_, data_n_2__1_, data_n_2__0_ } : 
                          (N22)? data_o[63:32] : 1'b0;
  assign N20 = N55;
  assign N21 = N54;
  assign N22 = N53;
  assign data_nn[95:64] = (N21)? { data_n_3__31_, data_n_3__30_, data_n_3__29_, data_n_3__28_, data_n_3__27_, data_n_3__26_, data_n_3__25_, data_n_3__24_, data_n_3__23_, data_n_3__22_, data_n_3__21_, data_n_3__20_, data_n_3__19_, data_n_3__18_, data_n_3__17_, data_n_3__16_, data_n_3__15_, data_n_3__14_, data_n_3__13_, data_n_3__12_, data_n_3__11_, data_n_3__10_, data_n_3__9_, data_n_3__8_, data_n_3__7_, data_n_3__6_, data_n_3__5_, data_n_3__4_, data_n_3__3_, data_n_3__2_, data_n_3__1_, data_n_3__0_ } : 
                          (N22)? { data_n_2__31_, data_n_2__30_, data_n_2__29_, data_n_2__28_, data_n_2__27_, data_n_2__26_, data_n_2__25_, data_n_2__24_, data_n_2__23_, data_n_2__22_, data_n_2__21_, data_n_2__20_, data_n_2__19_, data_n_2__18_, data_n_2__17_, data_n_2__16_, data_n_2__15_, data_n_2__14_, data_n_2__13_, data_n_2__12_, data_n_2__11_, data_n_2__10_, data_n_2__9_, data_n_2__8_, data_n_2__7_, data_n_2__6_, data_n_2__5_, data_n_2__4_, data_n_2__3_, data_n_2__2_, data_n_2__1_, data_n_2__0_ } : 1'b0;
  assign { N59, N58, N57, N56 } = (N23)? { 1'b0, 1'b0, valid_n } : 
                                  (N47)? { valid_n, valid_o } : 1'b0;
  assign N23 = yumi_cnt_i[1];
  assign valid_nn = (N24)? { N59, N58, N57 } : 
                    (N46)? { N58, N57, N56 } : 1'b0;
  assign N24 = yumi_cnt_i[0];
  assign data_nn[31] = (N48)? data_o[31] : 
                       (N50)? data_o[63] : 
                       (N49)? data_n_2__31_ : 
                       (N51)? data_n_3__31_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign N25 = 1'b0;
  assign data_nn[30] = (N48)? data_o[30] : 
                       (N50)? data_o[62] : 
                       (N49)? data_n_2__30_ : 
                       (N51)? data_n_3__30_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[29] = (N48)? data_o[29] : 
                       (N50)? data_o[61] : 
                       (N49)? data_n_2__29_ : 
                       (N51)? data_n_3__29_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[28] = (N48)? data_o[28] : 
                       (N50)? data_o[60] : 
                       (N49)? data_n_2__28_ : 
                       (N51)? data_n_3__28_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[27] = (N48)? data_o[27] : 
                       (N50)? data_o[59] : 
                       (N49)? data_n_2__27_ : 
                       (N51)? data_n_3__27_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[26] = (N48)? data_o[26] : 
                       (N50)? data_o[58] : 
                       (N49)? data_n_2__26_ : 
                       (N51)? data_n_3__26_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[25] = (N48)? data_o[25] : 
                       (N50)? data_o[57] : 
                       (N49)? data_n_2__25_ : 
                       (N51)? data_n_3__25_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[24] = (N48)? data_o[24] : 
                       (N50)? data_o[56] : 
                       (N49)? data_n_2__24_ : 
                       (N51)? data_n_3__24_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[23] = (N48)? data_o[23] : 
                       (N50)? data_o[55] : 
                       (N49)? data_n_2__23_ : 
                       (N51)? data_n_3__23_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[22] = (N48)? data_o[22] : 
                       (N50)? data_o[54] : 
                       (N49)? data_n_2__22_ : 
                       (N51)? data_n_3__22_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[21] = (N48)? data_o[21] : 
                       (N50)? data_o[53] : 
                       (N49)? data_n_2__21_ : 
                       (N51)? data_n_3__21_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[20] = (N48)? data_o[20] : 
                       (N50)? data_o[52] : 
                       (N49)? data_n_2__20_ : 
                       (N51)? data_n_3__20_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[19] = (N48)? data_o[19] : 
                       (N50)? data_o[51] : 
                       (N49)? data_n_2__19_ : 
                       (N51)? data_n_3__19_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[18] = (N48)? data_o[18] : 
                       (N50)? data_o[50] : 
                       (N49)? data_n_2__18_ : 
                       (N51)? data_n_3__18_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[17] = (N48)? data_o[17] : 
                       (N50)? data_o[49] : 
                       (N49)? data_n_2__17_ : 
                       (N51)? data_n_3__17_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[16] = (N48)? data_o[16] : 
                       (N50)? data_o[48] : 
                       (N49)? data_n_2__16_ : 
                       (N51)? data_n_3__16_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[15] = (N48)? data_o[15] : 
                       (N50)? data_o[47] : 
                       (N49)? data_n_2__15_ : 
                       (N51)? data_n_3__15_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[14] = (N48)? data_o[14] : 
                       (N50)? data_o[46] : 
                       (N49)? data_n_2__14_ : 
                       (N51)? data_n_3__14_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[13] = (N48)? data_o[13] : 
                       (N50)? data_o[45] : 
                       (N49)? data_n_2__13_ : 
                       (N51)? data_n_3__13_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[12] = (N48)? data_o[12] : 
                       (N50)? data_o[44] : 
                       (N49)? data_n_2__12_ : 
                       (N51)? data_n_3__12_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[11] = (N48)? data_o[11] : 
                       (N50)? data_o[43] : 
                       (N49)? data_n_2__11_ : 
                       (N51)? data_n_3__11_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[10] = (N48)? data_o[10] : 
                       (N50)? data_o[42] : 
                       (N49)? data_n_2__10_ : 
                       (N51)? data_n_3__10_ : 
                       (N25)? 1'b0 : 
                       (N25)? 1'b0 : 1'b0;
  assign data_nn[9] = (N48)? data_o[9] : 
                      (N50)? data_o[41] : 
                      (N49)? data_n_2__9_ : 
                      (N51)? data_n_3__9_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[8] = (N48)? data_o[8] : 
                      (N50)? data_o[40] : 
                      (N49)? data_n_2__8_ : 
                      (N51)? data_n_3__8_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[7] = (N48)? data_o[7] : 
                      (N50)? data_o[39] : 
                      (N49)? data_n_2__7_ : 
                      (N51)? data_n_3__7_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[6] = (N48)? data_o[6] : 
                      (N50)? data_o[38] : 
                      (N49)? data_n_2__6_ : 
                      (N51)? data_n_3__6_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[5] = (N48)? data_o[5] : 
                      (N50)? data_o[37] : 
                      (N49)? data_n_2__5_ : 
                      (N51)? data_n_3__5_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[4] = (N48)? data_o[4] : 
                      (N50)? data_o[36] : 
                      (N49)? data_n_2__4_ : 
                      (N51)? data_n_3__4_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[3] = (N48)? data_o[3] : 
                      (N50)? data_o[35] : 
                      (N49)? data_n_2__3_ : 
                      (N51)? data_n_3__3_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[2] = (N48)? data_o[2] : 
                      (N50)? data_o[34] : 
                      (N49)? data_n_2__2_ : 
                      (N51)? data_n_3__2_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[1] = (N48)? data_o[1] : 
                      (N50)? data_o[33] : 
                      (N49)? data_n_2__1_ : 
                      (N51)? data_n_3__1_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign data_nn[0] = (N48)? data_o[0] : 
                      (N50)? data_o[32] : 
                      (N49)? data_n_2__0_ : 
                      (N51)? data_n_3__0_ : 
                      (N25)? 1'b0 : 
                      (N25)? 1'b0 : 1'b0;
  assign ready_o = ~valid_r[2];
  assign N26 = valid_i & ready_o;
  assign N33 = ~N29;
  assign N34 = ~N30;
  assign N35 = ~N31;
  assign N36 = ~N32;
  assign N41 = valid_i & ready_o;
  assign N42 = ~N37;
  assign N43 = ~N38;
  assign N44 = ~N39;
  assign N45 = ~N40;
  assign N46 = ~yumi_cnt_i[0];
  assign N47 = ~yumi_cnt_i[1];
  assign N48 = N46 & N47;
  assign N49 = N46 & yumi_cnt_i[1];
  assign N50 = yumi_cnt_i[0] & N47;
  assign N51 = yumi_cnt_i[0] & yumi_cnt_i[1];

  always @(posedge clk_i) begin
    if(reset_i) begin
      valid_r_2_sv2v_reg <= 1'b0;
      valid_r_1_sv2v_reg <= 1'b0;
      valid_r_0_sv2v_reg <= 1'b0;
      num_els_r_1_sv2v_reg <= 1'b0;
      num_els_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      valid_r_2_sv2v_reg <= valid_nn[2];
      valid_r_1_sv2v_reg <= valid_nn[1];
      valid_r_0_sv2v_reg <= valid_nn[0];
      num_els_r_1_sv2v_reg <= num_els_n[1];
      num_els_r_0_sv2v_reg <= num_els_n[0];
    end 
    if(N60) begin
      data_r_95_sv2v_reg <= 1'b0;
      data_r_94_sv2v_reg <= 1'b0;
      data_r_93_sv2v_reg <= 1'b0;
      data_r_92_sv2v_reg <= 1'b0;
      data_r_91_sv2v_reg <= 1'b0;
      data_r_90_sv2v_reg <= 1'b0;
      data_r_89_sv2v_reg <= 1'b0;
      data_r_88_sv2v_reg <= 1'b0;
      data_r_87_sv2v_reg <= 1'b0;
      data_r_86_sv2v_reg <= 1'b0;
      data_r_85_sv2v_reg <= 1'b0;
      data_r_84_sv2v_reg <= 1'b0;
      data_r_83_sv2v_reg <= 1'b0;
      data_r_82_sv2v_reg <= 1'b0;
      data_r_81_sv2v_reg <= 1'b0;
      data_r_80_sv2v_reg <= 1'b0;
      data_r_79_sv2v_reg <= 1'b0;
      data_r_78_sv2v_reg <= 1'b0;
      data_r_77_sv2v_reg <= 1'b0;
      data_r_76_sv2v_reg <= 1'b0;
      data_r_75_sv2v_reg <= 1'b0;
      data_r_74_sv2v_reg <= 1'b0;
      data_r_73_sv2v_reg <= 1'b0;
      data_r_72_sv2v_reg <= 1'b0;
      data_r_71_sv2v_reg <= 1'b0;
      data_r_70_sv2v_reg <= 1'b0;
      data_r_69_sv2v_reg <= 1'b0;
      data_r_68_sv2v_reg <= 1'b0;
      data_r_67_sv2v_reg <= 1'b0;
      data_r_66_sv2v_reg <= 1'b0;
      data_r_65_sv2v_reg <= 1'b0;
      data_r_64_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_r_95_sv2v_reg <= data_nn[95];
      data_r_94_sv2v_reg <= data_nn[94];
      data_r_93_sv2v_reg <= data_nn[93];
      data_r_92_sv2v_reg <= data_nn[92];
      data_r_91_sv2v_reg <= data_nn[91];
      data_r_90_sv2v_reg <= data_nn[90];
      data_r_89_sv2v_reg <= data_nn[89];
      data_r_88_sv2v_reg <= data_nn[88];
      data_r_87_sv2v_reg <= data_nn[87];
      data_r_86_sv2v_reg <= data_nn[86];
      data_r_85_sv2v_reg <= data_nn[85];
      data_r_84_sv2v_reg <= data_nn[84];
      data_r_83_sv2v_reg <= data_nn[83];
      data_r_82_sv2v_reg <= data_nn[82];
      data_r_81_sv2v_reg <= data_nn[81];
      data_r_80_sv2v_reg <= data_nn[80];
      data_r_79_sv2v_reg <= data_nn[79];
      data_r_78_sv2v_reg <= data_nn[78];
      data_r_77_sv2v_reg <= data_nn[77];
      data_r_76_sv2v_reg <= data_nn[76];
      data_r_75_sv2v_reg <= data_nn[75];
      data_r_74_sv2v_reg <= data_nn[74];
      data_r_73_sv2v_reg <= data_nn[73];
      data_r_72_sv2v_reg <= data_nn[72];
      data_r_71_sv2v_reg <= data_nn[71];
      data_r_70_sv2v_reg <= data_nn[70];
      data_r_69_sv2v_reg <= data_nn[69];
      data_r_68_sv2v_reg <= data_nn[68];
      data_r_67_sv2v_reg <= data_nn[67];
      data_r_66_sv2v_reg <= data_nn[66];
      data_r_65_sv2v_reg <= data_nn[65];
      data_r_64_sv2v_reg <= data_nn[64];
    end 
    if(N52) begin
      data_r_63_sv2v_reg <= 1'b0;
      data_r_62_sv2v_reg <= 1'b0;
      data_r_61_sv2v_reg <= 1'b0;
      data_r_60_sv2v_reg <= 1'b0;
      data_r_59_sv2v_reg <= 1'b0;
      data_r_58_sv2v_reg <= 1'b0;
      data_r_57_sv2v_reg <= 1'b0;
      data_r_56_sv2v_reg <= 1'b0;
      data_r_55_sv2v_reg <= 1'b0;
      data_r_54_sv2v_reg <= 1'b0;
      data_r_53_sv2v_reg <= 1'b0;
      data_r_52_sv2v_reg <= 1'b0;
      data_r_51_sv2v_reg <= 1'b0;
      data_r_50_sv2v_reg <= 1'b0;
      data_r_49_sv2v_reg <= 1'b0;
      data_r_48_sv2v_reg <= 1'b0;
      data_r_47_sv2v_reg <= 1'b0;
      data_r_46_sv2v_reg <= 1'b0;
      data_r_45_sv2v_reg <= 1'b0;
      data_r_44_sv2v_reg <= 1'b0;
      data_r_43_sv2v_reg <= 1'b0;
      data_r_42_sv2v_reg <= 1'b0;
      data_r_41_sv2v_reg <= 1'b0;
      data_r_40_sv2v_reg <= 1'b0;
      data_r_39_sv2v_reg <= 1'b0;
      data_r_38_sv2v_reg <= 1'b0;
      data_r_37_sv2v_reg <= 1'b0;
      data_r_36_sv2v_reg <= 1'b0;
      data_r_35_sv2v_reg <= 1'b0;
      data_r_34_sv2v_reg <= 1'b0;
      data_r_33_sv2v_reg <= 1'b0;
      data_r_32_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_r_63_sv2v_reg <= data_nn[63];
      data_r_62_sv2v_reg <= data_nn[62];
      data_r_61_sv2v_reg <= data_nn[61];
      data_r_60_sv2v_reg <= data_nn[60];
      data_r_59_sv2v_reg <= data_nn[59];
      data_r_58_sv2v_reg <= data_nn[58];
      data_r_57_sv2v_reg <= data_nn[57];
      data_r_56_sv2v_reg <= data_nn[56];
      data_r_55_sv2v_reg <= data_nn[55];
      data_r_54_sv2v_reg <= data_nn[54];
      data_r_53_sv2v_reg <= data_nn[53];
      data_r_52_sv2v_reg <= data_nn[52];
      data_r_51_sv2v_reg <= data_nn[51];
      data_r_50_sv2v_reg <= data_nn[50];
      data_r_49_sv2v_reg <= data_nn[49];
      data_r_48_sv2v_reg <= data_nn[48];
      data_r_47_sv2v_reg <= data_nn[47];
      data_r_46_sv2v_reg <= data_nn[46];
      data_r_45_sv2v_reg <= data_nn[45];
      data_r_44_sv2v_reg <= data_nn[44];
      data_r_43_sv2v_reg <= data_nn[43];
      data_r_42_sv2v_reg <= data_nn[42];
      data_r_41_sv2v_reg <= data_nn[41];
      data_r_40_sv2v_reg <= data_nn[40];
      data_r_39_sv2v_reg <= data_nn[39];
      data_r_38_sv2v_reg <= data_nn[38];
      data_r_37_sv2v_reg <= data_nn[37];
      data_r_36_sv2v_reg <= data_nn[36];
      data_r_35_sv2v_reg <= data_nn[35];
      data_r_34_sv2v_reg <= data_nn[34];
      data_r_33_sv2v_reg <= data_nn[33];
      data_r_32_sv2v_reg <= data_nn[32];
    end 
    if(1'b1) begin
      data_r_31_sv2v_reg <= data_nn[31];
      data_r_30_sv2v_reg <= data_nn[30];
      data_r_29_sv2v_reg <= data_nn[29];
      data_r_28_sv2v_reg <= data_nn[28];
      data_r_27_sv2v_reg <= data_nn[27];
      data_r_26_sv2v_reg <= data_nn[26];
      data_r_25_sv2v_reg <= data_nn[25];
      data_r_24_sv2v_reg <= data_nn[24];
      data_r_23_sv2v_reg <= data_nn[23];
      data_r_22_sv2v_reg <= data_nn[22];
      data_r_21_sv2v_reg <= data_nn[21];
      data_r_20_sv2v_reg <= data_nn[20];
      data_r_19_sv2v_reg <= data_nn[19];
      data_r_18_sv2v_reg <= data_nn[18];
      data_r_17_sv2v_reg <= data_nn[17];
      data_r_16_sv2v_reg <= data_nn[16];
      data_r_15_sv2v_reg <= data_nn[15];
      data_r_14_sv2v_reg <= data_nn[14];
      data_r_13_sv2v_reg <= data_nn[13];
      data_r_12_sv2v_reg <= data_nn[12];
      data_r_11_sv2v_reg <= data_nn[11];
      data_r_10_sv2v_reg <= data_nn[10];
      data_r_9_sv2v_reg <= data_nn[9];
      data_r_8_sv2v_reg <= data_nn[8];
      data_r_7_sv2v_reg <= data_nn[7];
      data_r_6_sv2v_reg <= data_nn[6];
      data_r_5_sv2v_reg <= data_nn[5];
      data_r_4_sv2v_reg <= data_nn[4];
      data_r_3_sv2v_reg <= data_nn[3];
      data_r_2_sv2v_reg <= data_nn[2];
      data_r_1_sv2v_reg <= data_nn[1];
      data_r_0_sv2v_reg <= data_nn[0];
    end 
  end


endmodule



module bsg_circular_ptr_slots_p16_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [3:0] o;
  output [3:0] n_o;
  input clk;
  input reset_i;
  wire [3:0] o,n_o,\genblk1.genblk1.ptr_r_p1 ;
  wire N0,N1,N2;
  reg o_3_sv2v_reg,o_2_sv2v_reg,o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[3] = o_3_sv2v_reg;
  assign o[2] = o_2_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign \genblk1.genblk1.ptr_r_p1  = o + 1'b1;
  assign n_o = (N0)? \genblk1.genblk1.ptr_r_p1  : 
               (N1)? o : 1'b0;
  assign N0 = add_i[0];
  assign N1 = N2;
  assign N2 = ~add_i[0];

  always @(posedge clk) begin
    if(reset_i) begin
      o_3_sv2v_reg <= 1'b0;
      o_2_sv2v_reg <= 1'b0;
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_3_sv2v_reg <= n_o[3];
      o_2_sv2v_reg <= n_o[2];
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_synth_width_p64_els_p16_latch_last_read_p0_verbose_p1
(
  clk_i,
  v_i,
  reset_i,
  data_i,
  addr_i,
  w_i,
  data_o
);

  input [63:0] data_i;
  input [3:0] addr_i;
  output [63:0] data_o;
  input clk_i;
  input v_i;
  input reset_i;
  input w_i;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82;
  wire [3:0] \nz.addr_r ;
  wire [1023:0] \nz.mem ;
  reg \nz.addr_r_3_sv2v_reg ,\nz.addr_r_2_sv2v_reg ,\nz.addr_r_1_sv2v_reg ,
  \nz.addr_r_0_sv2v_reg ,\nz.mem_1023_sv2v_reg ,\nz.mem_1022_sv2v_reg ,
  \nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,\nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,
  \nz.mem_1017_sv2v_reg ,\nz.mem_1016_sv2v_reg ,\nz.mem_1015_sv2v_reg ,
  \nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,\nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,
  \nz.mem_1010_sv2v_reg ,\nz.mem_1009_sv2v_reg ,\nz.mem_1008_sv2v_reg ,
  \nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,\nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,
  \nz.mem_1003_sv2v_reg ,\nz.mem_1002_sv2v_reg ,\nz.mem_1001_sv2v_reg ,
  \nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,\nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,
  \nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,\nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,
  \nz.mem_992_sv2v_reg ,\nz.mem_991_sv2v_reg ,\nz.mem_990_sv2v_reg ,
  \nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,\nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,
  \nz.mem_985_sv2v_reg ,\nz.mem_984_sv2v_reg ,\nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,
  \nz.mem_981_sv2v_reg ,\nz.mem_980_sv2v_reg ,\nz.mem_979_sv2v_reg ,
  \nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,\nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,
  \nz.mem_974_sv2v_reg ,\nz.mem_973_sv2v_reg ,\nz.mem_972_sv2v_reg ,
  \nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,\nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,
  \nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,\nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,
  \nz.mem_963_sv2v_reg ,\nz.mem_962_sv2v_reg ,\nz.mem_961_sv2v_reg ,
  \nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,\nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,
  \nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,\nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,
  \nz.mem_952_sv2v_reg ,\nz.mem_951_sv2v_reg ,\nz.mem_950_sv2v_reg ,
  \nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,\nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,
  \nz.mem_945_sv2v_reg ,\nz.mem_944_sv2v_reg ,\nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,
  \nz.mem_941_sv2v_reg ,\nz.mem_940_sv2v_reg ,\nz.mem_939_sv2v_reg ,
  \nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,\nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,
  \nz.mem_934_sv2v_reg ,\nz.mem_933_sv2v_reg ,\nz.mem_932_sv2v_reg ,
  \nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,\nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,
  \nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,\nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,
  \nz.mem_923_sv2v_reg ,\nz.mem_922_sv2v_reg ,\nz.mem_921_sv2v_reg ,
  \nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,\nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,
  \nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,\nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,
  \nz.mem_912_sv2v_reg ,\nz.mem_911_sv2v_reg ,\nz.mem_910_sv2v_reg ,
  \nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,\nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,
  \nz.mem_905_sv2v_reg ,\nz.mem_904_sv2v_reg ,\nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,
  \nz.mem_901_sv2v_reg ,\nz.mem_900_sv2v_reg ,\nz.mem_899_sv2v_reg ,
  \nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,\nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,
  \nz.mem_894_sv2v_reg ,\nz.mem_893_sv2v_reg ,\nz.mem_892_sv2v_reg ,
  \nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,\nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,
  \nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,\nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,
  \nz.mem_883_sv2v_reg ,\nz.mem_882_sv2v_reg ,\nz.mem_881_sv2v_reg ,
  \nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,\nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,
  \nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,\nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,
  \nz.mem_872_sv2v_reg ,\nz.mem_871_sv2v_reg ,\nz.mem_870_sv2v_reg ,
  \nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,\nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,
  \nz.mem_865_sv2v_reg ,\nz.mem_864_sv2v_reg ,\nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,
  \nz.mem_861_sv2v_reg ,\nz.mem_860_sv2v_reg ,\nz.mem_859_sv2v_reg ,
  \nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,\nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,
  \nz.mem_854_sv2v_reg ,\nz.mem_853_sv2v_reg ,\nz.mem_852_sv2v_reg ,
  \nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,\nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,
  \nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,\nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,
  \nz.mem_843_sv2v_reg ,\nz.mem_842_sv2v_reg ,\nz.mem_841_sv2v_reg ,
  \nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,\nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,
  \nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,\nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,
  \nz.mem_832_sv2v_reg ,\nz.mem_831_sv2v_reg ,\nz.mem_830_sv2v_reg ,
  \nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,\nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,
  \nz.mem_825_sv2v_reg ,\nz.mem_824_sv2v_reg ,\nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,
  \nz.mem_821_sv2v_reg ,\nz.mem_820_sv2v_reg ,\nz.mem_819_sv2v_reg ,
  \nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,\nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,
  \nz.mem_814_sv2v_reg ,\nz.mem_813_sv2v_reg ,\nz.mem_812_sv2v_reg ,
  \nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,\nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,
  \nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,\nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,
  \nz.mem_803_sv2v_reg ,\nz.mem_802_sv2v_reg ,\nz.mem_801_sv2v_reg ,
  \nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,\nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,
  \nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,\nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,
  \nz.mem_792_sv2v_reg ,\nz.mem_791_sv2v_reg ,\nz.mem_790_sv2v_reg ,
  \nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,\nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,
  \nz.mem_785_sv2v_reg ,\nz.mem_784_sv2v_reg ,\nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,
  \nz.mem_781_sv2v_reg ,\nz.mem_780_sv2v_reg ,\nz.mem_779_sv2v_reg ,
  \nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,\nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,
  \nz.mem_774_sv2v_reg ,\nz.mem_773_sv2v_reg ,\nz.mem_772_sv2v_reg ,
  \nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,\nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,
  \nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,\nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,
  \nz.mem_763_sv2v_reg ,\nz.mem_762_sv2v_reg ,\nz.mem_761_sv2v_reg ,
  \nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,\nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,
  \nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,\nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,
  \nz.mem_752_sv2v_reg ,\nz.mem_751_sv2v_reg ,\nz.mem_750_sv2v_reg ,
  \nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,\nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,
  \nz.mem_745_sv2v_reg ,\nz.mem_744_sv2v_reg ,\nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,
  \nz.mem_741_sv2v_reg ,\nz.mem_740_sv2v_reg ,\nz.mem_739_sv2v_reg ,
  \nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,\nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,
  \nz.mem_734_sv2v_reg ,\nz.mem_733_sv2v_reg ,\nz.mem_732_sv2v_reg ,
  \nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,\nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,
  \nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,\nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,
  \nz.mem_723_sv2v_reg ,\nz.mem_722_sv2v_reg ,\nz.mem_721_sv2v_reg ,
  \nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,\nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,
  \nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,\nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,
  \nz.mem_712_sv2v_reg ,\nz.mem_711_sv2v_reg ,\nz.mem_710_sv2v_reg ,
  \nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,\nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,
  \nz.mem_705_sv2v_reg ,\nz.mem_704_sv2v_reg ,\nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,
  \nz.mem_701_sv2v_reg ,\nz.mem_700_sv2v_reg ,\nz.mem_699_sv2v_reg ,
  \nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,\nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,
  \nz.mem_694_sv2v_reg ,\nz.mem_693_sv2v_reg ,\nz.mem_692_sv2v_reg ,
  \nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,\nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,
  \nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,\nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,
  \nz.mem_683_sv2v_reg ,\nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,
  \nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,\nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,
  \nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,\nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,
  \nz.mem_672_sv2v_reg ,\nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,
  \nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,\nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,
  \nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,\nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,
  \nz.mem_661_sv2v_reg ,\nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,
  \nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,\nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,
  \nz.mem_654_sv2v_reg ,\nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,
  \nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,\nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,
  \nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,\nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,
  \nz.mem_643_sv2v_reg ,\nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,
  \nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,\nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,
  \nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,\nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,
  \nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,
  \nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,\nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,
  \nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,
  \nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,
  \nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,\nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,
  \nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,
  \nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,\nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,
  \nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,\nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,
  \nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,
  \nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,\nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,
  \nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,\nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,
  \nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,
  \nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,\nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,
  \nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,
  \nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,
  \nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,\nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,
  \nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,
  \nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,\nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,
  \nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,\nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,
  \nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,
  \nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,\nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,
  \nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,\nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,
  \nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,
  \nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,\nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,
  \nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,
  \nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,
  \nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,\nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,
  \nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,
  \nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,\nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,
  \nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,\nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,
  \nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,
  \nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,\nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,
  \nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,\nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,
  \nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,
  \nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,\nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,
  \nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,
  \nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,
  \nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,\nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,
  \nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,
  \nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,\nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,
  \nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,\nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,
  \nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,
  \nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,\nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,
  \nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,\nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,
  \nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,
  \nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,\nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,
  \nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,
  \nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,
  \nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,\nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,
  \nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,
  \nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,\nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,
  \nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,
  \nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,
  \nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,\nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,
  \nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,
  \nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,
  \nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,\nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,
  \nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,
  \nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,
  \nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,
  \nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,
  \nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,\nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,
  \nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,
  \nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,
  \nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,\nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,
  \nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,
  \nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,
  \nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,\nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,
  \nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,
  \nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,
  \nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,
  \nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,
  \nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,\nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,
  \nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,
  \nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,
  \nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,\nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,
  \nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,
  \nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,
  \nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,\nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,
  \nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,
  \nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,
  \nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,
  \nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,
  \nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,\nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,
  \nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,
  \nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,
  \nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,\nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,
  \nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,
  \nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,
  \nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,\nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,
  \nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,
  \nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,
  \nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,
  \nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,
  \nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,
  \nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,
  \nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,
  \nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,
  \nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,
  \nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,
  \nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,
  \nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,
  \nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,
  \nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,
  \nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,
  \nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,
  \nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,
  \nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,
  \nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,
  \nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,
  \nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,
  \nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,
  \nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,
  \nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,
  \nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,
  \nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,
  \nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,
  \nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,
  \nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,
  \nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,
  \nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,
  \nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,
  \nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,
  \nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,
  \nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,
  \nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,
  \nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,
  \nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,
  \nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,
  \nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,
  \nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,
  \nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,
  \nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,
  \nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,
  \nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,
  \nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,
  \nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,
  \nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,
  \nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,
  \nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,
  \nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,
  \nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,
  \nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,
  \nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,
  \nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,
  \nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,
  \nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,
  \nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,
  \nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,
  \nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,
  \nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,
  \nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,
  \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign data_o[63] = (N25)? \nz.mem [63] : 
                      (N27)? \nz.mem [127] : 
                      (N29)? \nz.mem [191] : 
                      (N31)? \nz.mem [255] : 
                      (N33)? \nz.mem [319] : 
                      (N35)? \nz.mem [383] : 
                      (N37)? \nz.mem [447] : 
                      (N39)? \nz.mem [511] : 
                      (N26)? \nz.mem [575] : 
                      (N28)? \nz.mem [639] : 
                      (N30)? \nz.mem [703] : 
                      (N32)? \nz.mem [767] : 
                      (N34)? \nz.mem [831] : 
                      (N36)? \nz.mem [895] : 
                      (N38)? \nz.mem [959] : 
                      (N40)? \nz.mem [1023] : 1'b0;
  assign data_o[62] = (N25)? \nz.mem [62] : 
                      (N27)? \nz.mem [126] : 
                      (N29)? \nz.mem [190] : 
                      (N31)? \nz.mem [254] : 
                      (N33)? \nz.mem [318] : 
                      (N35)? \nz.mem [382] : 
                      (N37)? \nz.mem [446] : 
                      (N39)? \nz.mem [510] : 
                      (N26)? \nz.mem [574] : 
                      (N28)? \nz.mem [638] : 
                      (N30)? \nz.mem [702] : 
                      (N32)? \nz.mem [766] : 
                      (N34)? \nz.mem [830] : 
                      (N36)? \nz.mem [894] : 
                      (N38)? \nz.mem [958] : 
                      (N40)? \nz.mem [1022] : 1'b0;
  assign data_o[61] = (N25)? \nz.mem [61] : 
                      (N27)? \nz.mem [125] : 
                      (N29)? \nz.mem [189] : 
                      (N31)? \nz.mem [253] : 
                      (N33)? \nz.mem [317] : 
                      (N35)? \nz.mem [381] : 
                      (N37)? \nz.mem [445] : 
                      (N39)? \nz.mem [509] : 
                      (N26)? \nz.mem [573] : 
                      (N28)? \nz.mem [637] : 
                      (N30)? \nz.mem [701] : 
                      (N32)? \nz.mem [765] : 
                      (N34)? \nz.mem [829] : 
                      (N36)? \nz.mem [893] : 
                      (N38)? \nz.mem [957] : 
                      (N40)? \nz.mem [1021] : 1'b0;
  assign data_o[60] = (N25)? \nz.mem [60] : 
                      (N27)? \nz.mem [124] : 
                      (N29)? \nz.mem [188] : 
                      (N31)? \nz.mem [252] : 
                      (N33)? \nz.mem [316] : 
                      (N35)? \nz.mem [380] : 
                      (N37)? \nz.mem [444] : 
                      (N39)? \nz.mem [508] : 
                      (N26)? \nz.mem [572] : 
                      (N28)? \nz.mem [636] : 
                      (N30)? \nz.mem [700] : 
                      (N32)? \nz.mem [764] : 
                      (N34)? \nz.mem [828] : 
                      (N36)? \nz.mem [892] : 
                      (N38)? \nz.mem [956] : 
                      (N40)? \nz.mem [1020] : 1'b0;
  assign data_o[59] = (N25)? \nz.mem [59] : 
                      (N27)? \nz.mem [123] : 
                      (N29)? \nz.mem [187] : 
                      (N31)? \nz.mem [251] : 
                      (N33)? \nz.mem [315] : 
                      (N35)? \nz.mem [379] : 
                      (N37)? \nz.mem [443] : 
                      (N39)? \nz.mem [507] : 
                      (N26)? \nz.mem [571] : 
                      (N28)? \nz.mem [635] : 
                      (N30)? \nz.mem [699] : 
                      (N32)? \nz.mem [763] : 
                      (N34)? \nz.mem [827] : 
                      (N36)? \nz.mem [891] : 
                      (N38)? \nz.mem [955] : 
                      (N40)? \nz.mem [1019] : 1'b0;
  assign data_o[58] = (N25)? \nz.mem [58] : 
                      (N27)? \nz.mem [122] : 
                      (N29)? \nz.mem [186] : 
                      (N31)? \nz.mem [250] : 
                      (N33)? \nz.mem [314] : 
                      (N35)? \nz.mem [378] : 
                      (N37)? \nz.mem [442] : 
                      (N39)? \nz.mem [506] : 
                      (N26)? \nz.mem [570] : 
                      (N28)? \nz.mem [634] : 
                      (N30)? \nz.mem [698] : 
                      (N32)? \nz.mem [762] : 
                      (N34)? \nz.mem [826] : 
                      (N36)? \nz.mem [890] : 
                      (N38)? \nz.mem [954] : 
                      (N40)? \nz.mem [1018] : 1'b0;
  assign data_o[57] = (N25)? \nz.mem [57] : 
                      (N27)? \nz.mem [121] : 
                      (N29)? \nz.mem [185] : 
                      (N31)? \nz.mem [249] : 
                      (N33)? \nz.mem [313] : 
                      (N35)? \nz.mem [377] : 
                      (N37)? \nz.mem [441] : 
                      (N39)? \nz.mem [505] : 
                      (N26)? \nz.mem [569] : 
                      (N28)? \nz.mem [633] : 
                      (N30)? \nz.mem [697] : 
                      (N32)? \nz.mem [761] : 
                      (N34)? \nz.mem [825] : 
                      (N36)? \nz.mem [889] : 
                      (N38)? \nz.mem [953] : 
                      (N40)? \nz.mem [1017] : 1'b0;
  assign data_o[56] = (N25)? \nz.mem [56] : 
                      (N27)? \nz.mem [120] : 
                      (N29)? \nz.mem [184] : 
                      (N31)? \nz.mem [248] : 
                      (N33)? \nz.mem [312] : 
                      (N35)? \nz.mem [376] : 
                      (N37)? \nz.mem [440] : 
                      (N39)? \nz.mem [504] : 
                      (N26)? \nz.mem [568] : 
                      (N28)? \nz.mem [632] : 
                      (N30)? \nz.mem [696] : 
                      (N32)? \nz.mem [760] : 
                      (N34)? \nz.mem [824] : 
                      (N36)? \nz.mem [888] : 
                      (N38)? \nz.mem [952] : 
                      (N40)? \nz.mem [1016] : 1'b0;
  assign data_o[55] = (N25)? \nz.mem [55] : 
                      (N27)? \nz.mem [119] : 
                      (N29)? \nz.mem [183] : 
                      (N31)? \nz.mem [247] : 
                      (N33)? \nz.mem [311] : 
                      (N35)? \nz.mem [375] : 
                      (N37)? \nz.mem [439] : 
                      (N39)? \nz.mem [503] : 
                      (N26)? \nz.mem [567] : 
                      (N28)? \nz.mem [631] : 
                      (N30)? \nz.mem [695] : 
                      (N32)? \nz.mem [759] : 
                      (N34)? \nz.mem [823] : 
                      (N36)? \nz.mem [887] : 
                      (N38)? \nz.mem [951] : 
                      (N40)? \nz.mem [1015] : 1'b0;
  assign data_o[54] = (N25)? \nz.mem [54] : 
                      (N27)? \nz.mem [118] : 
                      (N29)? \nz.mem [182] : 
                      (N31)? \nz.mem [246] : 
                      (N33)? \nz.mem [310] : 
                      (N35)? \nz.mem [374] : 
                      (N37)? \nz.mem [438] : 
                      (N39)? \nz.mem [502] : 
                      (N26)? \nz.mem [566] : 
                      (N28)? \nz.mem [630] : 
                      (N30)? \nz.mem [694] : 
                      (N32)? \nz.mem [758] : 
                      (N34)? \nz.mem [822] : 
                      (N36)? \nz.mem [886] : 
                      (N38)? \nz.mem [950] : 
                      (N40)? \nz.mem [1014] : 1'b0;
  assign data_o[53] = (N25)? \nz.mem [53] : 
                      (N27)? \nz.mem [117] : 
                      (N29)? \nz.mem [181] : 
                      (N31)? \nz.mem [245] : 
                      (N33)? \nz.mem [309] : 
                      (N35)? \nz.mem [373] : 
                      (N37)? \nz.mem [437] : 
                      (N39)? \nz.mem [501] : 
                      (N26)? \nz.mem [565] : 
                      (N28)? \nz.mem [629] : 
                      (N30)? \nz.mem [693] : 
                      (N32)? \nz.mem [757] : 
                      (N34)? \nz.mem [821] : 
                      (N36)? \nz.mem [885] : 
                      (N38)? \nz.mem [949] : 
                      (N40)? \nz.mem [1013] : 1'b0;
  assign data_o[52] = (N25)? \nz.mem [52] : 
                      (N27)? \nz.mem [116] : 
                      (N29)? \nz.mem [180] : 
                      (N31)? \nz.mem [244] : 
                      (N33)? \nz.mem [308] : 
                      (N35)? \nz.mem [372] : 
                      (N37)? \nz.mem [436] : 
                      (N39)? \nz.mem [500] : 
                      (N26)? \nz.mem [564] : 
                      (N28)? \nz.mem [628] : 
                      (N30)? \nz.mem [692] : 
                      (N32)? \nz.mem [756] : 
                      (N34)? \nz.mem [820] : 
                      (N36)? \nz.mem [884] : 
                      (N38)? \nz.mem [948] : 
                      (N40)? \nz.mem [1012] : 1'b0;
  assign data_o[51] = (N25)? \nz.mem [51] : 
                      (N27)? \nz.mem [115] : 
                      (N29)? \nz.mem [179] : 
                      (N31)? \nz.mem [243] : 
                      (N33)? \nz.mem [307] : 
                      (N35)? \nz.mem [371] : 
                      (N37)? \nz.mem [435] : 
                      (N39)? \nz.mem [499] : 
                      (N26)? \nz.mem [563] : 
                      (N28)? \nz.mem [627] : 
                      (N30)? \nz.mem [691] : 
                      (N32)? \nz.mem [755] : 
                      (N34)? \nz.mem [819] : 
                      (N36)? \nz.mem [883] : 
                      (N38)? \nz.mem [947] : 
                      (N40)? \nz.mem [1011] : 1'b0;
  assign data_o[50] = (N25)? \nz.mem [50] : 
                      (N27)? \nz.mem [114] : 
                      (N29)? \nz.mem [178] : 
                      (N31)? \nz.mem [242] : 
                      (N33)? \nz.mem [306] : 
                      (N35)? \nz.mem [370] : 
                      (N37)? \nz.mem [434] : 
                      (N39)? \nz.mem [498] : 
                      (N26)? \nz.mem [562] : 
                      (N28)? \nz.mem [626] : 
                      (N30)? \nz.mem [690] : 
                      (N32)? \nz.mem [754] : 
                      (N34)? \nz.mem [818] : 
                      (N36)? \nz.mem [882] : 
                      (N38)? \nz.mem [946] : 
                      (N40)? \nz.mem [1010] : 1'b0;
  assign data_o[49] = (N25)? \nz.mem [49] : 
                      (N27)? \nz.mem [113] : 
                      (N29)? \nz.mem [177] : 
                      (N31)? \nz.mem [241] : 
                      (N33)? \nz.mem [305] : 
                      (N35)? \nz.mem [369] : 
                      (N37)? \nz.mem [433] : 
                      (N39)? \nz.mem [497] : 
                      (N26)? \nz.mem [561] : 
                      (N28)? \nz.mem [625] : 
                      (N30)? \nz.mem [689] : 
                      (N32)? \nz.mem [753] : 
                      (N34)? \nz.mem [817] : 
                      (N36)? \nz.mem [881] : 
                      (N38)? \nz.mem [945] : 
                      (N40)? \nz.mem [1009] : 1'b0;
  assign data_o[48] = (N25)? \nz.mem [48] : 
                      (N27)? \nz.mem [112] : 
                      (N29)? \nz.mem [176] : 
                      (N31)? \nz.mem [240] : 
                      (N33)? \nz.mem [304] : 
                      (N35)? \nz.mem [368] : 
                      (N37)? \nz.mem [432] : 
                      (N39)? \nz.mem [496] : 
                      (N26)? \nz.mem [560] : 
                      (N28)? \nz.mem [624] : 
                      (N30)? \nz.mem [688] : 
                      (N32)? \nz.mem [752] : 
                      (N34)? \nz.mem [816] : 
                      (N36)? \nz.mem [880] : 
                      (N38)? \nz.mem [944] : 
                      (N40)? \nz.mem [1008] : 1'b0;
  assign data_o[47] = (N25)? \nz.mem [47] : 
                      (N27)? \nz.mem [111] : 
                      (N29)? \nz.mem [175] : 
                      (N31)? \nz.mem [239] : 
                      (N33)? \nz.mem [303] : 
                      (N35)? \nz.mem [367] : 
                      (N37)? \nz.mem [431] : 
                      (N39)? \nz.mem [495] : 
                      (N26)? \nz.mem [559] : 
                      (N28)? \nz.mem [623] : 
                      (N30)? \nz.mem [687] : 
                      (N32)? \nz.mem [751] : 
                      (N34)? \nz.mem [815] : 
                      (N36)? \nz.mem [879] : 
                      (N38)? \nz.mem [943] : 
                      (N40)? \nz.mem [1007] : 1'b0;
  assign data_o[46] = (N25)? \nz.mem [46] : 
                      (N27)? \nz.mem [110] : 
                      (N29)? \nz.mem [174] : 
                      (N31)? \nz.mem [238] : 
                      (N33)? \nz.mem [302] : 
                      (N35)? \nz.mem [366] : 
                      (N37)? \nz.mem [430] : 
                      (N39)? \nz.mem [494] : 
                      (N26)? \nz.mem [558] : 
                      (N28)? \nz.mem [622] : 
                      (N30)? \nz.mem [686] : 
                      (N32)? \nz.mem [750] : 
                      (N34)? \nz.mem [814] : 
                      (N36)? \nz.mem [878] : 
                      (N38)? \nz.mem [942] : 
                      (N40)? \nz.mem [1006] : 1'b0;
  assign data_o[45] = (N25)? \nz.mem [45] : 
                      (N27)? \nz.mem [109] : 
                      (N29)? \nz.mem [173] : 
                      (N31)? \nz.mem [237] : 
                      (N33)? \nz.mem [301] : 
                      (N35)? \nz.mem [365] : 
                      (N37)? \nz.mem [429] : 
                      (N39)? \nz.mem [493] : 
                      (N26)? \nz.mem [557] : 
                      (N28)? \nz.mem [621] : 
                      (N30)? \nz.mem [685] : 
                      (N32)? \nz.mem [749] : 
                      (N34)? \nz.mem [813] : 
                      (N36)? \nz.mem [877] : 
                      (N38)? \nz.mem [941] : 
                      (N40)? \nz.mem [1005] : 1'b0;
  assign data_o[44] = (N25)? \nz.mem [44] : 
                      (N27)? \nz.mem [108] : 
                      (N29)? \nz.mem [172] : 
                      (N31)? \nz.mem [236] : 
                      (N33)? \nz.mem [300] : 
                      (N35)? \nz.mem [364] : 
                      (N37)? \nz.mem [428] : 
                      (N39)? \nz.mem [492] : 
                      (N26)? \nz.mem [556] : 
                      (N28)? \nz.mem [620] : 
                      (N30)? \nz.mem [684] : 
                      (N32)? \nz.mem [748] : 
                      (N34)? \nz.mem [812] : 
                      (N36)? \nz.mem [876] : 
                      (N38)? \nz.mem [940] : 
                      (N40)? \nz.mem [1004] : 1'b0;
  assign data_o[43] = (N25)? \nz.mem [43] : 
                      (N27)? \nz.mem [107] : 
                      (N29)? \nz.mem [171] : 
                      (N31)? \nz.mem [235] : 
                      (N33)? \nz.mem [299] : 
                      (N35)? \nz.mem [363] : 
                      (N37)? \nz.mem [427] : 
                      (N39)? \nz.mem [491] : 
                      (N26)? \nz.mem [555] : 
                      (N28)? \nz.mem [619] : 
                      (N30)? \nz.mem [683] : 
                      (N32)? \nz.mem [747] : 
                      (N34)? \nz.mem [811] : 
                      (N36)? \nz.mem [875] : 
                      (N38)? \nz.mem [939] : 
                      (N40)? \nz.mem [1003] : 1'b0;
  assign data_o[42] = (N25)? \nz.mem [42] : 
                      (N27)? \nz.mem [106] : 
                      (N29)? \nz.mem [170] : 
                      (N31)? \nz.mem [234] : 
                      (N33)? \nz.mem [298] : 
                      (N35)? \nz.mem [362] : 
                      (N37)? \nz.mem [426] : 
                      (N39)? \nz.mem [490] : 
                      (N26)? \nz.mem [554] : 
                      (N28)? \nz.mem [618] : 
                      (N30)? \nz.mem [682] : 
                      (N32)? \nz.mem [746] : 
                      (N34)? \nz.mem [810] : 
                      (N36)? \nz.mem [874] : 
                      (N38)? \nz.mem [938] : 
                      (N40)? \nz.mem [1002] : 1'b0;
  assign data_o[41] = (N25)? \nz.mem [41] : 
                      (N27)? \nz.mem [105] : 
                      (N29)? \nz.mem [169] : 
                      (N31)? \nz.mem [233] : 
                      (N33)? \nz.mem [297] : 
                      (N35)? \nz.mem [361] : 
                      (N37)? \nz.mem [425] : 
                      (N39)? \nz.mem [489] : 
                      (N26)? \nz.mem [553] : 
                      (N28)? \nz.mem [617] : 
                      (N30)? \nz.mem [681] : 
                      (N32)? \nz.mem [745] : 
                      (N34)? \nz.mem [809] : 
                      (N36)? \nz.mem [873] : 
                      (N38)? \nz.mem [937] : 
                      (N40)? \nz.mem [1001] : 1'b0;
  assign data_o[40] = (N25)? \nz.mem [40] : 
                      (N27)? \nz.mem [104] : 
                      (N29)? \nz.mem [168] : 
                      (N31)? \nz.mem [232] : 
                      (N33)? \nz.mem [296] : 
                      (N35)? \nz.mem [360] : 
                      (N37)? \nz.mem [424] : 
                      (N39)? \nz.mem [488] : 
                      (N26)? \nz.mem [552] : 
                      (N28)? \nz.mem [616] : 
                      (N30)? \nz.mem [680] : 
                      (N32)? \nz.mem [744] : 
                      (N34)? \nz.mem [808] : 
                      (N36)? \nz.mem [872] : 
                      (N38)? \nz.mem [936] : 
                      (N40)? \nz.mem [1000] : 1'b0;
  assign data_o[39] = (N25)? \nz.mem [39] : 
                      (N27)? \nz.mem [103] : 
                      (N29)? \nz.mem [167] : 
                      (N31)? \nz.mem [231] : 
                      (N33)? \nz.mem [295] : 
                      (N35)? \nz.mem [359] : 
                      (N37)? \nz.mem [423] : 
                      (N39)? \nz.mem [487] : 
                      (N26)? \nz.mem [551] : 
                      (N28)? \nz.mem [615] : 
                      (N30)? \nz.mem [679] : 
                      (N32)? \nz.mem [743] : 
                      (N34)? \nz.mem [807] : 
                      (N36)? \nz.mem [871] : 
                      (N38)? \nz.mem [935] : 
                      (N40)? \nz.mem [999] : 1'b0;
  assign data_o[38] = (N25)? \nz.mem [38] : 
                      (N27)? \nz.mem [102] : 
                      (N29)? \nz.mem [166] : 
                      (N31)? \nz.mem [230] : 
                      (N33)? \nz.mem [294] : 
                      (N35)? \nz.mem [358] : 
                      (N37)? \nz.mem [422] : 
                      (N39)? \nz.mem [486] : 
                      (N26)? \nz.mem [550] : 
                      (N28)? \nz.mem [614] : 
                      (N30)? \nz.mem [678] : 
                      (N32)? \nz.mem [742] : 
                      (N34)? \nz.mem [806] : 
                      (N36)? \nz.mem [870] : 
                      (N38)? \nz.mem [934] : 
                      (N40)? \nz.mem [998] : 1'b0;
  assign data_o[37] = (N25)? \nz.mem [37] : 
                      (N27)? \nz.mem [101] : 
                      (N29)? \nz.mem [165] : 
                      (N31)? \nz.mem [229] : 
                      (N33)? \nz.mem [293] : 
                      (N35)? \nz.mem [357] : 
                      (N37)? \nz.mem [421] : 
                      (N39)? \nz.mem [485] : 
                      (N26)? \nz.mem [549] : 
                      (N28)? \nz.mem [613] : 
                      (N30)? \nz.mem [677] : 
                      (N32)? \nz.mem [741] : 
                      (N34)? \nz.mem [805] : 
                      (N36)? \nz.mem [869] : 
                      (N38)? \nz.mem [933] : 
                      (N40)? \nz.mem [997] : 1'b0;
  assign data_o[36] = (N25)? \nz.mem [36] : 
                      (N27)? \nz.mem [100] : 
                      (N29)? \nz.mem [164] : 
                      (N31)? \nz.mem [228] : 
                      (N33)? \nz.mem [292] : 
                      (N35)? \nz.mem [356] : 
                      (N37)? \nz.mem [420] : 
                      (N39)? \nz.mem [484] : 
                      (N26)? \nz.mem [548] : 
                      (N28)? \nz.mem [612] : 
                      (N30)? \nz.mem [676] : 
                      (N32)? \nz.mem [740] : 
                      (N34)? \nz.mem [804] : 
                      (N36)? \nz.mem [868] : 
                      (N38)? \nz.mem [932] : 
                      (N40)? \nz.mem [996] : 1'b0;
  assign data_o[35] = (N25)? \nz.mem [35] : 
                      (N27)? \nz.mem [99] : 
                      (N29)? \nz.mem [163] : 
                      (N31)? \nz.mem [227] : 
                      (N33)? \nz.mem [291] : 
                      (N35)? \nz.mem [355] : 
                      (N37)? \nz.mem [419] : 
                      (N39)? \nz.mem [483] : 
                      (N26)? \nz.mem [547] : 
                      (N28)? \nz.mem [611] : 
                      (N30)? \nz.mem [675] : 
                      (N32)? \nz.mem [739] : 
                      (N34)? \nz.mem [803] : 
                      (N36)? \nz.mem [867] : 
                      (N38)? \nz.mem [931] : 
                      (N40)? \nz.mem [995] : 1'b0;
  assign data_o[34] = (N25)? \nz.mem [34] : 
                      (N27)? \nz.mem [98] : 
                      (N29)? \nz.mem [162] : 
                      (N31)? \nz.mem [226] : 
                      (N33)? \nz.mem [290] : 
                      (N35)? \nz.mem [354] : 
                      (N37)? \nz.mem [418] : 
                      (N39)? \nz.mem [482] : 
                      (N26)? \nz.mem [546] : 
                      (N28)? \nz.mem [610] : 
                      (N30)? \nz.mem [674] : 
                      (N32)? \nz.mem [738] : 
                      (N34)? \nz.mem [802] : 
                      (N36)? \nz.mem [866] : 
                      (N38)? \nz.mem [930] : 
                      (N40)? \nz.mem [994] : 1'b0;
  assign data_o[33] = (N25)? \nz.mem [33] : 
                      (N27)? \nz.mem [97] : 
                      (N29)? \nz.mem [161] : 
                      (N31)? \nz.mem [225] : 
                      (N33)? \nz.mem [289] : 
                      (N35)? \nz.mem [353] : 
                      (N37)? \nz.mem [417] : 
                      (N39)? \nz.mem [481] : 
                      (N26)? \nz.mem [545] : 
                      (N28)? \nz.mem [609] : 
                      (N30)? \nz.mem [673] : 
                      (N32)? \nz.mem [737] : 
                      (N34)? \nz.mem [801] : 
                      (N36)? \nz.mem [865] : 
                      (N38)? \nz.mem [929] : 
                      (N40)? \nz.mem [993] : 1'b0;
  assign data_o[32] = (N25)? \nz.mem [32] : 
                      (N27)? \nz.mem [96] : 
                      (N29)? \nz.mem [160] : 
                      (N31)? \nz.mem [224] : 
                      (N33)? \nz.mem [288] : 
                      (N35)? \nz.mem [352] : 
                      (N37)? \nz.mem [416] : 
                      (N39)? \nz.mem [480] : 
                      (N26)? \nz.mem [544] : 
                      (N28)? \nz.mem [608] : 
                      (N30)? \nz.mem [672] : 
                      (N32)? \nz.mem [736] : 
                      (N34)? \nz.mem [800] : 
                      (N36)? \nz.mem [864] : 
                      (N38)? \nz.mem [928] : 
                      (N40)? \nz.mem [992] : 1'b0;
  assign data_o[31] = (N25)? \nz.mem [31] : 
                      (N27)? \nz.mem [95] : 
                      (N29)? \nz.mem [159] : 
                      (N31)? \nz.mem [223] : 
                      (N33)? \nz.mem [287] : 
                      (N35)? \nz.mem [351] : 
                      (N37)? \nz.mem [415] : 
                      (N39)? \nz.mem [479] : 
                      (N26)? \nz.mem [543] : 
                      (N28)? \nz.mem [607] : 
                      (N30)? \nz.mem [671] : 
                      (N32)? \nz.mem [735] : 
                      (N34)? \nz.mem [799] : 
                      (N36)? \nz.mem [863] : 
                      (N38)? \nz.mem [927] : 
                      (N40)? \nz.mem [991] : 1'b0;
  assign data_o[30] = (N25)? \nz.mem [30] : 
                      (N27)? \nz.mem [94] : 
                      (N29)? \nz.mem [158] : 
                      (N31)? \nz.mem [222] : 
                      (N33)? \nz.mem [286] : 
                      (N35)? \nz.mem [350] : 
                      (N37)? \nz.mem [414] : 
                      (N39)? \nz.mem [478] : 
                      (N26)? \nz.mem [542] : 
                      (N28)? \nz.mem [606] : 
                      (N30)? \nz.mem [670] : 
                      (N32)? \nz.mem [734] : 
                      (N34)? \nz.mem [798] : 
                      (N36)? \nz.mem [862] : 
                      (N38)? \nz.mem [926] : 
                      (N40)? \nz.mem [990] : 1'b0;
  assign data_o[29] = (N25)? \nz.mem [29] : 
                      (N27)? \nz.mem [93] : 
                      (N29)? \nz.mem [157] : 
                      (N31)? \nz.mem [221] : 
                      (N33)? \nz.mem [285] : 
                      (N35)? \nz.mem [349] : 
                      (N37)? \nz.mem [413] : 
                      (N39)? \nz.mem [477] : 
                      (N26)? \nz.mem [541] : 
                      (N28)? \nz.mem [605] : 
                      (N30)? \nz.mem [669] : 
                      (N32)? \nz.mem [733] : 
                      (N34)? \nz.mem [797] : 
                      (N36)? \nz.mem [861] : 
                      (N38)? \nz.mem [925] : 
                      (N40)? \nz.mem [989] : 1'b0;
  assign data_o[28] = (N25)? \nz.mem [28] : 
                      (N27)? \nz.mem [92] : 
                      (N29)? \nz.mem [156] : 
                      (N31)? \nz.mem [220] : 
                      (N33)? \nz.mem [284] : 
                      (N35)? \nz.mem [348] : 
                      (N37)? \nz.mem [412] : 
                      (N39)? \nz.mem [476] : 
                      (N26)? \nz.mem [540] : 
                      (N28)? \nz.mem [604] : 
                      (N30)? \nz.mem [668] : 
                      (N32)? \nz.mem [732] : 
                      (N34)? \nz.mem [796] : 
                      (N36)? \nz.mem [860] : 
                      (N38)? \nz.mem [924] : 
                      (N40)? \nz.mem [988] : 1'b0;
  assign data_o[27] = (N25)? \nz.mem [27] : 
                      (N27)? \nz.mem [91] : 
                      (N29)? \nz.mem [155] : 
                      (N31)? \nz.mem [219] : 
                      (N33)? \nz.mem [283] : 
                      (N35)? \nz.mem [347] : 
                      (N37)? \nz.mem [411] : 
                      (N39)? \nz.mem [475] : 
                      (N26)? \nz.mem [539] : 
                      (N28)? \nz.mem [603] : 
                      (N30)? \nz.mem [667] : 
                      (N32)? \nz.mem [731] : 
                      (N34)? \nz.mem [795] : 
                      (N36)? \nz.mem [859] : 
                      (N38)? \nz.mem [923] : 
                      (N40)? \nz.mem [987] : 1'b0;
  assign data_o[26] = (N25)? \nz.mem [26] : 
                      (N27)? \nz.mem [90] : 
                      (N29)? \nz.mem [154] : 
                      (N31)? \nz.mem [218] : 
                      (N33)? \nz.mem [282] : 
                      (N35)? \nz.mem [346] : 
                      (N37)? \nz.mem [410] : 
                      (N39)? \nz.mem [474] : 
                      (N26)? \nz.mem [538] : 
                      (N28)? \nz.mem [602] : 
                      (N30)? \nz.mem [666] : 
                      (N32)? \nz.mem [730] : 
                      (N34)? \nz.mem [794] : 
                      (N36)? \nz.mem [858] : 
                      (N38)? \nz.mem [922] : 
                      (N40)? \nz.mem [986] : 1'b0;
  assign data_o[25] = (N25)? \nz.mem [25] : 
                      (N27)? \nz.mem [89] : 
                      (N29)? \nz.mem [153] : 
                      (N31)? \nz.mem [217] : 
                      (N33)? \nz.mem [281] : 
                      (N35)? \nz.mem [345] : 
                      (N37)? \nz.mem [409] : 
                      (N39)? \nz.mem [473] : 
                      (N26)? \nz.mem [537] : 
                      (N28)? \nz.mem [601] : 
                      (N30)? \nz.mem [665] : 
                      (N32)? \nz.mem [729] : 
                      (N34)? \nz.mem [793] : 
                      (N36)? \nz.mem [857] : 
                      (N38)? \nz.mem [921] : 
                      (N40)? \nz.mem [985] : 1'b0;
  assign data_o[24] = (N25)? \nz.mem [24] : 
                      (N27)? \nz.mem [88] : 
                      (N29)? \nz.mem [152] : 
                      (N31)? \nz.mem [216] : 
                      (N33)? \nz.mem [280] : 
                      (N35)? \nz.mem [344] : 
                      (N37)? \nz.mem [408] : 
                      (N39)? \nz.mem [472] : 
                      (N26)? \nz.mem [536] : 
                      (N28)? \nz.mem [600] : 
                      (N30)? \nz.mem [664] : 
                      (N32)? \nz.mem [728] : 
                      (N34)? \nz.mem [792] : 
                      (N36)? \nz.mem [856] : 
                      (N38)? \nz.mem [920] : 
                      (N40)? \nz.mem [984] : 1'b0;
  assign data_o[23] = (N25)? \nz.mem [23] : 
                      (N27)? \nz.mem [87] : 
                      (N29)? \nz.mem [151] : 
                      (N31)? \nz.mem [215] : 
                      (N33)? \nz.mem [279] : 
                      (N35)? \nz.mem [343] : 
                      (N37)? \nz.mem [407] : 
                      (N39)? \nz.mem [471] : 
                      (N26)? \nz.mem [535] : 
                      (N28)? \nz.mem [599] : 
                      (N30)? \nz.mem [663] : 
                      (N32)? \nz.mem [727] : 
                      (N34)? \nz.mem [791] : 
                      (N36)? \nz.mem [855] : 
                      (N38)? \nz.mem [919] : 
                      (N40)? \nz.mem [983] : 1'b0;
  assign data_o[22] = (N25)? \nz.mem [22] : 
                      (N27)? \nz.mem [86] : 
                      (N29)? \nz.mem [150] : 
                      (N31)? \nz.mem [214] : 
                      (N33)? \nz.mem [278] : 
                      (N35)? \nz.mem [342] : 
                      (N37)? \nz.mem [406] : 
                      (N39)? \nz.mem [470] : 
                      (N26)? \nz.mem [534] : 
                      (N28)? \nz.mem [598] : 
                      (N30)? \nz.mem [662] : 
                      (N32)? \nz.mem [726] : 
                      (N34)? \nz.mem [790] : 
                      (N36)? \nz.mem [854] : 
                      (N38)? \nz.mem [918] : 
                      (N40)? \nz.mem [982] : 1'b0;
  assign data_o[21] = (N25)? \nz.mem [21] : 
                      (N27)? \nz.mem [85] : 
                      (N29)? \nz.mem [149] : 
                      (N31)? \nz.mem [213] : 
                      (N33)? \nz.mem [277] : 
                      (N35)? \nz.mem [341] : 
                      (N37)? \nz.mem [405] : 
                      (N39)? \nz.mem [469] : 
                      (N26)? \nz.mem [533] : 
                      (N28)? \nz.mem [597] : 
                      (N30)? \nz.mem [661] : 
                      (N32)? \nz.mem [725] : 
                      (N34)? \nz.mem [789] : 
                      (N36)? \nz.mem [853] : 
                      (N38)? \nz.mem [917] : 
                      (N40)? \nz.mem [981] : 1'b0;
  assign data_o[20] = (N25)? \nz.mem [20] : 
                      (N27)? \nz.mem [84] : 
                      (N29)? \nz.mem [148] : 
                      (N31)? \nz.mem [212] : 
                      (N33)? \nz.mem [276] : 
                      (N35)? \nz.mem [340] : 
                      (N37)? \nz.mem [404] : 
                      (N39)? \nz.mem [468] : 
                      (N26)? \nz.mem [532] : 
                      (N28)? \nz.mem [596] : 
                      (N30)? \nz.mem [660] : 
                      (N32)? \nz.mem [724] : 
                      (N34)? \nz.mem [788] : 
                      (N36)? \nz.mem [852] : 
                      (N38)? \nz.mem [916] : 
                      (N40)? \nz.mem [980] : 1'b0;
  assign data_o[19] = (N25)? \nz.mem [19] : 
                      (N27)? \nz.mem [83] : 
                      (N29)? \nz.mem [147] : 
                      (N31)? \nz.mem [211] : 
                      (N33)? \nz.mem [275] : 
                      (N35)? \nz.mem [339] : 
                      (N37)? \nz.mem [403] : 
                      (N39)? \nz.mem [467] : 
                      (N26)? \nz.mem [531] : 
                      (N28)? \nz.mem [595] : 
                      (N30)? \nz.mem [659] : 
                      (N32)? \nz.mem [723] : 
                      (N34)? \nz.mem [787] : 
                      (N36)? \nz.mem [851] : 
                      (N38)? \nz.mem [915] : 
                      (N40)? \nz.mem [979] : 1'b0;
  assign data_o[18] = (N25)? \nz.mem [18] : 
                      (N27)? \nz.mem [82] : 
                      (N29)? \nz.mem [146] : 
                      (N31)? \nz.mem [210] : 
                      (N33)? \nz.mem [274] : 
                      (N35)? \nz.mem [338] : 
                      (N37)? \nz.mem [402] : 
                      (N39)? \nz.mem [466] : 
                      (N26)? \nz.mem [530] : 
                      (N28)? \nz.mem [594] : 
                      (N30)? \nz.mem [658] : 
                      (N32)? \nz.mem [722] : 
                      (N34)? \nz.mem [786] : 
                      (N36)? \nz.mem [850] : 
                      (N38)? \nz.mem [914] : 
                      (N40)? \nz.mem [978] : 1'b0;
  assign data_o[17] = (N25)? \nz.mem [17] : 
                      (N27)? \nz.mem [81] : 
                      (N29)? \nz.mem [145] : 
                      (N31)? \nz.mem [209] : 
                      (N33)? \nz.mem [273] : 
                      (N35)? \nz.mem [337] : 
                      (N37)? \nz.mem [401] : 
                      (N39)? \nz.mem [465] : 
                      (N26)? \nz.mem [529] : 
                      (N28)? \nz.mem [593] : 
                      (N30)? \nz.mem [657] : 
                      (N32)? \nz.mem [721] : 
                      (N34)? \nz.mem [785] : 
                      (N36)? \nz.mem [849] : 
                      (N38)? \nz.mem [913] : 
                      (N40)? \nz.mem [977] : 1'b0;
  assign data_o[16] = (N25)? \nz.mem [16] : 
                      (N27)? \nz.mem [80] : 
                      (N29)? \nz.mem [144] : 
                      (N31)? \nz.mem [208] : 
                      (N33)? \nz.mem [272] : 
                      (N35)? \nz.mem [336] : 
                      (N37)? \nz.mem [400] : 
                      (N39)? \nz.mem [464] : 
                      (N26)? \nz.mem [528] : 
                      (N28)? \nz.mem [592] : 
                      (N30)? \nz.mem [656] : 
                      (N32)? \nz.mem [720] : 
                      (N34)? \nz.mem [784] : 
                      (N36)? \nz.mem [848] : 
                      (N38)? \nz.mem [912] : 
                      (N40)? \nz.mem [976] : 1'b0;
  assign data_o[15] = (N25)? \nz.mem [15] : 
                      (N27)? \nz.mem [79] : 
                      (N29)? \nz.mem [143] : 
                      (N31)? \nz.mem [207] : 
                      (N33)? \nz.mem [271] : 
                      (N35)? \nz.mem [335] : 
                      (N37)? \nz.mem [399] : 
                      (N39)? \nz.mem [463] : 
                      (N26)? \nz.mem [527] : 
                      (N28)? \nz.mem [591] : 
                      (N30)? \nz.mem [655] : 
                      (N32)? \nz.mem [719] : 
                      (N34)? \nz.mem [783] : 
                      (N36)? \nz.mem [847] : 
                      (N38)? \nz.mem [911] : 
                      (N40)? \nz.mem [975] : 1'b0;
  assign data_o[14] = (N25)? \nz.mem [14] : 
                      (N27)? \nz.mem [78] : 
                      (N29)? \nz.mem [142] : 
                      (N31)? \nz.mem [206] : 
                      (N33)? \nz.mem [270] : 
                      (N35)? \nz.mem [334] : 
                      (N37)? \nz.mem [398] : 
                      (N39)? \nz.mem [462] : 
                      (N26)? \nz.mem [526] : 
                      (N28)? \nz.mem [590] : 
                      (N30)? \nz.mem [654] : 
                      (N32)? \nz.mem [718] : 
                      (N34)? \nz.mem [782] : 
                      (N36)? \nz.mem [846] : 
                      (N38)? \nz.mem [910] : 
                      (N40)? \nz.mem [974] : 1'b0;
  assign data_o[13] = (N25)? \nz.mem [13] : 
                      (N27)? \nz.mem [77] : 
                      (N29)? \nz.mem [141] : 
                      (N31)? \nz.mem [205] : 
                      (N33)? \nz.mem [269] : 
                      (N35)? \nz.mem [333] : 
                      (N37)? \nz.mem [397] : 
                      (N39)? \nz.mem [461] : 
                      (N26)? \nz.mem [525] : 
                      (N28)? \nz.mem [589] : 
                      (N30)? \nz.mem [653] : 
                      (N32)? \nz.mem [717] : 
                      (N34)? \nz.mem [781] : 
                      (N36)? \nz.mem [845] : 
                      (N38)? \nz.mem [909] : 
                      (N40)? \nz.mem [973] : 1'b0;
  assign data_o[12] = (N25)? \nz.mem [12] : 
                      (N27)? \nz.mem [76] : 
                      (N29)? \nz.mem [140] : 
                      (N31)? \nz.mem [204] : 
                      (N33)? \nz.mem [268] : 
                      (N35)? \nz.mem [332] : 
                      (N37)? \nz.mem [396] : 
                      (N39)? \nz.mem [460] : 
                      (N26)? \nz.mem [524] : 
                      (N28)? \nz.mem [588] : 
                      (N30)? \nz.mem [652] : 
                      (N32)? \nz.mem [716] : 
                      (N34)? \nz.mem [780] : 
                      (N36)? \nz.mem [844] : 
                      (N38)? \nz.mem [908] : 
                      (N40)? \nz.mem [972] : 1'b0;
  assign data_o[11] = (N25)? \nz.mem [11] : 
                      (N27)? \nz.mem [75] : 
                      (N29)? \nz.mem [139] : 
                      (N31)? \nz.mem [203] : 
                      (N33)? \nz.mem [267] : 
                      (N35)? \nz.mem [331] : 
                      (N37)? \nz.mem [395] : 
                      (N39)? \nz.mem [459] : 
                      (N26)? \nz.mem [523] : 
                      (N28)? \nz.mem [587] : 
                      (N30)? \nz.mem [651] : 
                      (N32)? \nz.mem [715] : 
                      (N34)? \nz.mem [779] : 
                      (N36)? \nz.mem [843] : 
                      (N38)? \nz.mem [907] : 
                      (N40)? \nz.mem [971] : 1'b0;
  assign data_o[10] = (N25)? \nz.mem [10] : 
                      (N27)? \nz.mem [74] : 
                      (N29)? \nz.mem [138] : 
                      (N31)? \nz.mem [202] : 
                      (N33)? \nz.mem [266] : 
                      (N35)? \nz.mem [330] : 
                      (N37)? \nz.mem [394] : 
                      (N39)? \nz.mem [458] : 
                      (N26)? \nz.mem [522] : 
                      (N28)? \nz.mem [586] : 
                      (N30)? \nz.mem [650] : 
                      (N32)? \nz.mem [714] : 
                      (N34)? \nz.mem [778] : 
                      (N36)? \nz.mem [842] : 
                      (N38)? \nz.mem [906] : 
                      (N40)? \nz.mem [970] : 1'b0;
  assign data_o[9] = (N25)? \nz.mem [9] : 
                     (N27)? \nz.mem [73] : 
                     (N29)? \nz.mem [137] : 
                     (N31)? \nz.mem [201] : 
                     (N33)? \nz.mem [265] : 
                     (N35)? \nz.mem [329] : 
                     (N37)? \nz.mem [393] : 
                     (N39)? \nz.mem [457] : 
                     (N26)? \nz.mem [521] : 
                     (N28)? \nz.mem [585] : 
                     (N30)? \nz.mem [649] : 
                     (N32)? \nz.mem [713] : 
                     (N34)? \nz.mem [777] : 
                     (N36)? \nz.mem [841] : 
                     (N38)? \nz.mem [905] : 
                     (N40)? \nz.mem [969] : 1'b0;
  assign data_o[8] = (N25)? \nz.mem [8] : 
                     (N27)? \nz.mem [72] : 
                     (N29)? \nz.mem [136] : 
                     (N31)? \nz.mem [200] : 
                     (N33)? \nz.mem [264] : 
                     (N35)? \nz.mem [328] : 
                     (N37)? \nz.mem [392] : 
                     (N39)? \nz.mem [456] : 
                     (N26)? \nz.mem [520] : 
                     (N28)? \nz.mem [584] : 
                     (N30)? \nz.mem [648] : 
                     (N32)? \nz.mem [712] : 
                     (N34)? \nz.mem [776] : 
                     (N36)? \nz.mem [840] : 
                     (N38)? \nz.mem [904] : 
                     (N40)? \nz.mem [968] : 1'b0;
  assign data_o[7] = (N25)? \nz.mem [7] : 
                     (N27)? \nz.mem [71] : 
                     (N29)? \nz.mem [135] : 
                     (N31)? \nz.mem [199] : 
                     (N33)? \nz.mem [263] : 
                     (N35)? \nz.mem [327] : 
                     (N37)? \nz.mem [391] : 
                     (N39)? \nz.mem [455] : 
                     (N26)? \nz.mem [519] : 
                     (N28)? \nz.mem [583] : 
                     (N30)? \nz.mem [647] : 
                     (N32)? \nz.mem [711] : 
                     (N34)? \nz.mem [775] : 
                     (N36)? \nz.mem [839] : 
                     (N38)? \nz.mem [903] : 
                     (N40)? \nz.mem [967] : 1'b0;
  assign data_o[6] = (N25)? \nz.mem [6] : 
                     (N27)? \nz.mem [70] : 
                     (N29)? \nz.mem [134] : 
                     (N31)? \nz.mem [198] : 
                     (N33)? \nz.mem [262] : 
                     (N35)? \nz.mem [326] : 
                     (N37)? \nz.mem [390] : 
                     (N39)? \nz.mem [454] : 
                     (N26)? \nz.mem [518] : 
                     (N28)? \nz.mem [582] : 
                     (N30)? \nz.mem [646] : 
                     (N32)? \nz.mem [710] : 
                     (N34)? \nz.mem [774] : 
                     (N36)? \nz.mem [838] : 
                     (N38)? \nz.mem [902] : 
                     (N40)? \nz.mem [966] : 1'b0;
  assign data_o[5] = (N25)? \nz.mem [5] : 
                     (N27)? \nz.mem [69] : 
                     (N29)? \nz.mem [133] : 
                     (N31)? \nz.mem [197] : 
                     (N33)? \nz.mem [261] : 
                     (N35)? \nz.mem [325] : 
                     (N37)? \nz.mem [389] : 
                     (N39)? \nz.mem [453] : 
                     (N26)? \nz.mem [517] : 
                     (N28)? \nz.mem [581] : 
                     (N30)? \nz.mem [645] : 
                     (N32)? \nz.mem [709] : 
                     (N34)? \nz.mem [773] : 
                     (N36)? \nz.mem [837] : 
                     (N38)? \nz.mem [901] : 
                     (N40)? \nz.mem [965] : 1'b0;
  assign data_o[4] = (N25)? \nz.mem [4] : 
                     (N27)? \nz.mem [68] : 
                     (N29)? \nz.mem [132] : 
                     (N31)? \nz.mem [196] : 
                     (N33)? \nz.mem [260] : 
                     (N35)? \nz.mem [324] : 
                     (N37)? \nz.mem [388] : 
                     (N39)? \nz.mem [452] : 
                     (N26)? \nz.mem [516] : 
                     (N28)? \nz.mem [580] : 
                     (N30)? \nz.mem [644] : 
                     (N32)? \nz.mem [708] : 
                     (N34)? \nz.mem [772] : 
                     (N36)? \nz.mem [836] : 
                     (N38)? \nz.mem [900] : 
                     (N40)? \nz.mem [964] : 1'b0;
  assign data_o[3] = (N25)? \nz.mem [3] : 
                     (N27)? \nz.mem [67] : 
                     (N29)? \nz.mem [131] : 
                     (N31)? \nz.mem [195] : 
                     (N33)? \nz.mem [259] : 
                     (N35)? \nz.mem [323] : 
                     (N37)? \nz.mem [387] : 
                     (N39)? \nz.mem [451] : 
                     (N26)? \nz.mem [515] : 
                     (N28)? \nz.mem [579] : 
                     (N30)? \nz.mem [643] : 
                     (N32)? \nz.mem [707] : 
                     (N34)? \nz.mem [771] : 
                     (N36)? \nz.mem [835] : 
                     (N38)? \nz.mem [899] : 
                     (N40)? \nz.mem [963] : 1'b0;
  assign data_o[2] = (N25)? \nz.mem [2] : 
                     (N27)? \nz.mem [66] : 
                     (N29)? \nz.mem [130] : 
                     (N31)? \nz.mem [194] : 
                     (N33)? \nz.mem [258] : 
                     (N35)? \nz.mem [322] : 
                     (N37)? \nz.mem [386] : 
                     (N39)? \nz.mem [450] : 
                     (N26)? \nz.mem [514] : 
                     (N28)? \nz.mem [578] : 
                     (N30)? \nz.mem [642] : 
                     (N32)? \nz.mem [706] : 
                     (N34)? \nz.mem [770] : 
                     (N36)? \nz.mem [834] : 
                     (N38)? \nz.mem [898] : 
                     (N40)? \nz.mem [962] : 1'b0;
  assign data_o[1] = (N25)? \nz.mem [1] : 
                     (N27)? \nz.mem [65] : 
                     (N29)? \nz.mem [129] : 
                     (N31)? \nz.mem [193] : 
                     (N33)? \nz.mem [257] : 
                     (N35)? \nz.mem [321] : 
                     (N37)? \nz.mem [385] : 
                     (N39)? \nz.mem [449] : 
                     (N26)? \nz.mem [513] : 
                     (N28)? \nz.mem [577] : 
                     (N30)? \nz.mem [641] : 
                     (N32)? \nz.mem [705] : 
                     (N34)? \nz.mem [769] : 
                     (N36)? \nz.mem [833] : 
                     (N38)? \nz.mem [897] : 
                     (N40)? \nz.mem [961] : 1'b0;
  assign data_o[0] = (N25)? \nz.mem [0] : 
                     (N27)? \nz.mem [64] : 
                     (N29)? \nz.mem [128] : 
                     (N31)? \nz.mem [192] : 
                     (N33)? \nz.mem [256] : 
                     (N35)? \nz.mem [320] : 
                     (N37)? \nz.mem [384] : 
                     (N39)? \nz.mem [448] : 
                     (N26)? \nz.mem [512] : 
                     (N28)? \nz.mem [576] : 
                     (N30)? \nz.mem [640] : 
                     (N32)? \nz.mem [704] : 
                     (N34)? \nz.mem [768] : 
                     (N36)? \nz.mem [832] : 
                     (N38)? \nz.mem [896] : 
                     (N40)? \nz.mem [960] : 1'b0;
  assign N75 = addr_i[2] & addr_i[3];
  assign N76 = N0 & addr_i[3];
  assign N0 = ~addr_i[2];
  assign N77 = addr_i[2] & N1;
  assign N1 = ~addr_i[3];
  assign N78 = N2 & N3;
  assign N2 = ~addr_i[2];
  assign N3 = ~addr_i[3];
  assign N79 = addr_i[0] & addr_i[1];
  assign N80 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N81 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N82 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N58 = N75 & N79;
  assign N57 = N75 & N80;
  assign N56 = N75 & N81;
  assign N55 = N75 & N82;
  assign N54 = N76 & N79;
  assign N53 = N76 & N80;
  assign N52 = N76 & N81;
  assign N51 = N76 & N82;
  assign N50 = N77 & N79;
  assign N49 = N77 & N80;
  assign N48 = N77 & N81;
  assign N47 = N77 & N82;
  assign N46 = N78 & N79;
  assign N45 = N78 & N80;
  assign N44 = N78 & N81;
  assign N43 = N78 & N82;
  assign { N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59 } = (N8)? { N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43 } : 
                                                                                              (N42)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N41;
  assign N9 = ~\nz.addr_r [0];
  assign N10 = ~\nz.addr_r [1];
  assign N11 = N9 & N10;
  assign N12 = N9 & \nz.addr_r [1];
  assign N13 = \nz.addr_r [0] & N10;
  assign N14 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N15 = ~\nz.addr_r [2];
  assign N16 = N11 & N15;
  assign N17 = N11 & \nz.addr_r [2];
  assign N18 = N13 & N15;
  assign N19 = N13 & \nz.addr_r [2];
  assign N20 = N12 & N15;
  assign N21 = N12 & \nz.addr_r [2];
  assign N22 = N14 & N15;
  assign N23 = N14 & \nz.addr_r [2];
  assign N24 = ~\nz.addr_r [3];
  assign N25 = N16 & N24;
  assign N26 = N16 & \nz.addr_r [3];
  assign N27 = N18 & N24;
  assign N28 = N18 & \nz.addr_r [3];
  assign N29 = N20 & N24;
  assign N30 = N20 & \nz.addr_r [3];
  assign N31 = N22 & N24;
  assign N32 = N22 & \nz.addr_r [3];
  assign N33 = N17 & N24;
  assign N34 = N17 & \nz.addr_r [3];
  assign N35 = N19 & N24;
  assign N36 = N19 & \nz.addr_r [3];
  assign N37 = N21 & N24;
  assign N38 = N21 & \nz.addr_r [3];
  assign N39 = N23 & N24;
  assign N40 = N23 & \nz.addr_r [3];
  assign N41 = v_i & w_i;
  assign N42 = ~N41;

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N74) begin
      \nz.mem_1023_sv2v_reg  <= data_i[63];
      \nz.mem_1022_sv2v_reg  <= data_i[62];
      \nz.mem_1021_sv2v_reg  <= data_i[61];
      \nz.mem_1020_sv2v_reg  <= data_i[60];
      \nz.mem_1019_sv2v_reg  <= data_i[59];
      \nz.mem_1018_sv2v_reg  <= data_i[58];
      \nz.mem_1017_sv2v_reg  <= data_i[57];
      \nz.mem_1016_sv2v_reg  <= data_i[56];
      \nz.mem_1015_sv2v_reg  <= data_i[55];
      \nz.mem_1014_sv2v_reg  <= data_i[54];
      \nz.mem_1013_sv2v_reg  <= data_i[53];
      \nz.mem_1012_sv2v_reg  <= data_i[52];
      \nz.mem_1011_sv2v_reg  <= data_i[51];
      \nz.mem_1010_sv2v_reg  <= data_i[50];
      \nz.mem_1009_sv2v_reg  <= data_i[49];
      \nz.mem_1008_sv2v_reg  <= data_i[48];
      \nz.mem_1007_sv2v_reg  <= data_i[47];
      \nz.mem_1006_sv2v_reg  <= data_i[46];
      \nz.mem_1005_sv2v_reg  <= data_i[45];
      \nz.mem_1004_sv2v_reg  <= data_i[44];
      \nz.mem_1003_sv2v_reg  <= data_i[43];
      \nz.mem_1002_sv2v_reg  <= data_i[42];
      \nz.mem_1001_sv2v_reg  <= data_i[41];
      \nz.mem_1000_sv2v_reg  <= data_i[40];
      \nz.mem_999_sv2v_reg  <= data_i[39];
      \nz.mem_998_sv2v_reg  <= data_i[38];
      \nz.mem_997_sv2v_reg  <= data_i[37];
      \nz.mem_996_sv2v_reg  <= data_i[36];
      \nz.mem_995_sv2v_reg  <= data_i[35];
      \nz.mem_994_sv2v_reg  <= data_i[34];
      \nz.mem_993_sv2v_reg  <= data_i[33];
      \nz.mem_992_sv2v_reg  <= data_i[32];
      \nz.mem_991_sv2v_reg  <= data_i[31];
      \nz.mem_990_sv2v_reg  <= data_i[30];
      \nz.mem_989_sv2v_reg  <= data_i[29];
      \nz.mem_988_sv2v_reg  <= data_i[28];
      \nz.mem_987_sv2v_reg  <= data_i[27];
      \nz.mem_986_sv2v_reg  <= data_i[26];
      \nz.mem_985_sv2v_reg  <= data_i[25];
      \nz.mem_984_sv2v_reg  <= data_i[24];
      \nz.mem_983_sv2v_reg  <= data_i[23];
      \nz.mem_982_sv2v_reg  <= data_i[22];
      \nz.mem_981_sv2v_reg  <= data_i[21];
      \nz.mem_980_sv2v_reg  <= data_i[20];
      \nz.mem_979_sv2v_reg  <= data_i[19];
      \nz.mem_978_sv2v_reg  <= data_i[18];
      \nz.mem_977_sv2v_reg  <= data_i[17];
      \nz.mem_976_sv2v_reg  <= data_i[16];
      \nz.mem_975_sv2v_reg  <= data_i[15];
      \nz.mem_974_sv2v_reg  <= data_i[14];
      \nz.mem_973_sv2v_reg  <= data_i[13];
      \nz.mem_972_sv2v_reg  <= data_i[12];
      \nz.mem_971_sv2v_reg  <= data_i[11];
      \nz.mem_970_sv2v_reg  <= data_i[10];
      \nz.mem_969_sv2v_reg  <= data_i[9];
      \nz.mem_968_sv2v_reg  <= data_i[8];
      \nz.mem_967_sv2v_reg  <= data_i[7];
      \nz.mem_966_sv2v_reg  <= data_i[6];
      \nz.mem_965_sv2v_reg  <= data_i[5];
      \nz.mem_964_sv2v_reg  <= data_i[4];
      \nz.mem_963_sv2v_reg  <= data_i[3];
      \nz.mem_962_sv2v_reg  <= data_i[2];
      \nz.mem_961_sv2v_reg  <= data_i[1];
      \nz.mem_960_sv2v_reg  <= data_i[0];
    end 
    if(N73) begin
      \nz.mem_959_sv2v_reg  <= data_i[63];
      \nz.mem_958_sv2v_reg  <= data_i[62];
      \nz.mem_957_sv2v_reg  <= data_i[61];
      \nz.mem_956_sv2v_reg  <= data_i[60];
      \nz.mem_955_sv2v_reg  <= data_i[59];
      \nz.mem_954_sv2v_reg  <= data_i[58];
      \nz.mem_953_sv2v_reg  <= data_i[57];
      \nz.mem_952_sv2v_reg  <= data_i[56];
      \nz.mem_951_sv2v_reg  <= data_i[55];
      \nz.mem_950_sv2v_reg  <= data_i[54];
      \nz.mem_949_sv2v_reg  <= data_i[53];
      \nz.mem_948_sv2v_reg  <= data_i[52];
      \nz.mem_947_sv2v_reg  <= data_i[51];
      \nz.mem_946_sv2v_reg  <= data_i[50];
      \nz.mem_945_sv2v_reg  <= data_i[49];
      \nz.mem_944_sv2v_reg  <= data_i[48];
      \nz.mem_943_sv2v_reg  <= data_i[47];
      \nz.mem_942_sv2v_reg  <= data_i[46];
      \nz.mem_941_sv2v_reg  <= data_i[45];
      \nz.mem_940_sv2v_reg  <= data_i[44];
      \nz.mem_939_sv2v_reg  <= data_i[43];
      \nz.mem_938_sv2v_reg  <= data_i[42];
      \nz.mem_937_sv2v_reg  <= data_i[41];
      \nz.mem_936_sv2v_reg  <= data_i[40];
      \nz.mem_935_sv2v_reg  <= data_i[39];
      \nz.mem_934_sv2v_reg  <= data_i[38];
      \nz.mem_933_sv2v_reg  <= data_i[37];
      \nz.mem_932_sv2v_reg  <= data_i[36];
      \nz.mem_931_sv2v_reg  <= data_i[35];
      \nz.mem_930_sv2v_reg  <= data_i[34];
      \nz.mem_929_sv2v_reg  <= data_i[33];
      \nz.mem_928_sv2v_reg  <= data_i[32];
      \nz.mem_927_sv2v_reg  <= data_i[31];
      \nz.mem_926_sv2v_reg  <= data_i[30];
      \nz.mem_925_sv2v_reg  <= data_i[29];
      \nz.mem_924_sv2v_reg  <= data_i[28];
      \nz.mem_923_sv2v_reg  <= data_i[27];
      \nz.mem_922_sv2v_reg  <= data_i[26];
      \nz.mem_921_sv2v_reg  <= data_i[25];
      \nz.mem_920_sv2v_reg  <= data_i[24];
      \nz.mem_919_sv2v_reg  <= data_i[23];
      \nz.mem_918_sv2v_reg  <= data_i[22];
      \nz.mem_917_sv2v_reg  <= data_i[21];
      \nz.mem_916_sv2v_reg  <= data_i[20];
      \nz.mem_915_sv2v_reg  <= data_i[19];
      \nz.mem_914_sv2v_reg  <= data_i[18];
      \nz.mem_913_sv2v_reg  <= data_i[17];
      \nz.mem_912_sv2v_reg  <= data_i[16];
      \nz.mem_911_sv2v_reg  <= data_i[15];
      \nz.mem_910_sv2v_reg  <= data_i[14];
      \nz.mem_909_sv2v_reg  <= data_i[13];
      \nz.mem_908_sv2v_reg  <= data_i[12];
      \nz.mem_907_sv2v_reg  <= data_i[11];
      \nz.mem_906_sv2v_reg  <= data_i[10];
      \nz.mem_905_sv2v_reg  <= data_i[9];
      \nz.mem_904_sv2v_reg  <= data_i[8];
      \nz.mem_903_sv2v_reg  <= data_i[7];
      \nz.mem_902_sv2v_reg  <= data_i[6];
      \nz.mem_901_sv2v_reg  <= data_i[5];
      \nz.mem_900_sv2v_reg  <= data_i[4];
      \nz.mem_899_sv2v_reg  <= data_i[3];
      \nz.mem_898_sv2v_reg  <= data_i[2];
      \nz.mem_897_sv2v_reg  <= data_i[1];
      \nz.mem_896_sv2v_reg  <= data_i[0];
    end 
    if(N72) begin
      \nz.mem_895_sv2v_reg  <= data_i[63];
      \nz.mem_894_sv2v_reg  <= data_i[62];
      \nz.mem_893_sv2v_reg  <= data_i[61];
      \nz.mem_892_sv2v_reg  <= data_i[60];
      \nz.mem_891_sv2v_reg  <= data_i[59];
      \nz.mem_890_sv2v_reg  <= data_i[58];
      \nz.mem_889_sv2v_reg  <= data_i[57];
      \nz.mem_888_sv2v_reg  <= data_i[56];
      \nz.mem_887_sv2v_reg  <= data_i[55];
      \nz.mem_886_sv2v_reg  <= data_i[54];
      \nz.mem_885_sv2v_reg  <= data_i[53];
      \nz.mem_884_sv2v_reg  <= data_i[52];
      \nz.mem_883_sv2v_reg  <= data_i[51];
      \nz.mem_882_sv2v_reg  <= data_i[50];
      \nz.mem_881_sv2v_reg  <= data_i[49];
      \nz.mem_880_sv2v_reg  <= data_i[48];
      \nz.mem_879_sv2v_reg  <= data_i[47];
      \nz.mem_878_sv2v_reg  <= data_i[46];
      \nz.mem_877_sv2v_reg  <= data_i[45];
      \nz.mem_876_sv2v_reg  <= data_i[44];
      \nz.mem_875_sv2v_reg  <= data_i[43];
      \nz.mem_874_sv2v_reg  <= data_i[42];
      \nz.mem_873_sv2v_reg  <= data_i[41];
      \nz.mem_872_sv2v_reg  <= data_i[40];
      \nz.mem_871_sv2v_reg  <= data_i[39];
      \nz.mem_870_sv2v_reg  <= data_i[38];
      \nz.mem_869_sv2v_reg  <= data_i[37];
      \nz.mem_868_sv2v_reg  <= data_i[36];
      \nz.mem_867_sv2v_reg  <= data_i[35];
      \nz.mem_866_sv2v_reg  <= data_i[34];
      \nz.mem_865_sv2v_reg  <= data_i[33];
      \nz.mem_864_sv2v_reg  <= data_i[32];
      \nz.mem_863_sv2v_reg  <= data_i[31];
      \nz.mem_862_sv2v_reg  <= data_i[30];
      \nz.mem_861_sv2v_reg  <= data_i[29];
      \nz.mem_860_sv2v_reg  <= data_i[28];
      \nz.mem_859_sv2v_reg  <= data_i[27];
      \nz.mem_858_sv2v_reg  <= data_i[26];
      \nz.mem_857_sv2v_reg  <= data_i[25];
      \nz.mem_856_sv2v_reg  <= data_i[24];
      \nz.mem_855_sv2v_reg  <= data_i[23];
      \nz.mem_854_sv2v_reg  <= data_i[22];
      \nz.mem_853_sv2v_reg  <= data_i[21];
      \nz.mem_852_sv2v_reg  <= data_i[20];
      \nz.mem_851_sv2v_reg  <= data_i[19];
      \nz.mem_850_sv2v_reg  <= data_i[18];
      \nz.mem_849_sv2v_reg  <= data_i[17];
      \nz.mem_848_sv2v_reg  <= data_i[16];
      \nz.mem_847_sv2v_reg  <= data_i[15];
      \nz.mem_846_sv2v_reg  <= data_i[14];
      \nz.mem_845_sv2v_reg  <= data_i[13];
      \nz.mem_844_sv2v_reg  <= data_i[12];
      \nz.mem_843_sv2v_reg  <= data_i[11];
      \nz.mem_842_sv2v_reg  <= data_i[10];
      \nz.mem_841_sv2v_reg  <= data_i[9];
      \nz.mem_840_sv2v_reg  <= data_i[8];
      \nz.mem_839_sv2v_reg  <= data_i[7];
      \nz.mem_838_sv2v_reg  <= data_i[6];
      \nz.mem_837_sv2v_reg  <= data_i[5];
      \nz.mem_836_sv2v_reg  <= data_i[4];
      \nz.mem_835_sv2v_reg  <= data_i[3];
      \nz.mem_834_sv2v_reg  <= data_i[2];
      \nz.mem_833_sv2v_reg  <= data_i[1];
      \nz.mem_832_sv2v_reg  <= data_i[0];
    end 
    if(N71) begin
      \nz.mem_831_sv2v_reg  <= data_i[63];
      \nz.mem_830_sv2v_reg  <= data_i[62];
      \nz.mem_829_sv2v_reg  <= data_i[61];
      \nz.mem_828_sv2v_reg  <= data_i[60];
      \nz.mem_827_sv2v_reg  <= data_i[59];
      \nz.mem_826_sv2v_reg  <= data_i[58];
      \nz.mem_825_sv2v_reg  <= data_i[57];
      \nz.mem_824_sv2v_reg  <= data_i[56];
      \nz.mem_823_sv2v_reg  <= data_i[55];
      \nz.mem_822_sv2v_reg  <= data_i[54];
      \nz.mem_821_sv2v_reg  <= data_i[53];
      \nz.mem_820_sv2v_reg  <= data_i[52];
      \nz.mem_819_sv2v_reg  <= data_i[51];
      \nz.mem_818_sv2v_reg  <= data_i[50];
      \nz.mem_817_sv2v_reg  <= data_i[49];
      \nz.mem_816_sv2v_reg  <= data_i[48];
      \nz.mem_815_sv2v_reg  <= data_i[47];
      \nz.mem_814_sv2v_reg  <= data_i[46];
      \nz.mem_813_sv2v_reg  <= data_i[45];
      \nz.mem_812_sv2v_reg  <= data_i[44];
      \nz.mem_811_sv2v_reg  <= data_i[43];
      \nz.mem_810_sv2v_reg  <= data_i[42];
      \nz.mem_809_sv2v_reg  <= data_i[41];
      \nz.mem_808_sv2v_reg  <= data_i[40];
      \nz.mem_807_sv2v_reg  <= data_i[39];
      \nz.mem_806_sv2v_reg  <= data_i[38];
      \nz.mem_805_sv2v_reg  <= data_i[37];
      \nz.mem_804_sv2v_reg  <= data_i[36];
      \nz.mem_803_sv2v_reg  <= data_i[35];
      \nz.mem_802_sv2v_reg  <= data_i[34];
      \nz.mem_801_sv2v_reg  <= data_i[33];
      \nz.mem_800_sv2v_reg  <= data_i[32];
      \nz.mem_799_sv2v_reg  <= data_i[31];
      \nz.mem_798_sv2v_reg  <= data_i[30];
      \nz.mem_797_sv2v_reg  <= data_i[29];
      \nz.mem_796_sv2v_reg  <= data_i[28];
      \nz.mem_795_sv2v_reg  <= data_i[27];
      \nz.mem_794_sv2v_reg  <= data_i[26];
      \nz.mem_793_sv2v_reg  <= data_i[25];
      \nz.mem_792_sv2v_reg  <= data_i[24];
      \nz.mem_791_sv2v_reg  <= data_i[23];
      \nz.mem_790_sv2v_reg  <= data_i[22];
      \nz.mem_789_sv2v_reg  <= data_i[21];
      \nz.mem_788_sv2v_reg  <= data_i[20];
      \nz.mem_787_sv2v_reg  <= data_i[19];
      \nz.mem_786_sv2v_reg  <= data_i[18];
      \nz.mem_785_sv2v_reg  <= data_i[17];
      \nz.mem_784_sv2v_reg  <= data_i[16];
      \nz.mem_783_sv2v_reg  <= data_i[15];
      \nz.mem_782_sv2v_reg  <= data_i[14];
      \nz.mem_781_sv2v_reg  <= data_i[13];
      \nz.mem_780_sv2v_reg  <= data_i[12];
      \nz.mem_779_sv2v_reg  <= data_i[11];
      \nz.mem_778_sv2v_reg  <= data_i[10];
      \nz.mem_777_sv2v_reg  <= data_i[9];
      \nz.mem_776_sv2v_reg  <= data_i[8];
      \nz.mem_775_sv2v_reg  <= data_i[7];
      \nz.mem_774_sv2v_reg  <= data_i[6];
      \nz.mem_773_sv2v_reg  <= data_i[5];
      \nz.mem_772_sv2v_reg  <= data_i[4];
      \nz.mem_771_sv2v_reg  <= data_i[3];
      \nz.mem_770_sv2v_reg  <= data_i[2];
      \nz.mem_769_sv2v_reg  <= data_i[1];
      \nz.mem_768_sv2v_reg  <= data_i[0];
    end 
    if(N70) begin
      \nz.mem_767_sv2v_reg  <= data_i[63];
      \nz.mem_766_sv2v_reg  <= data_i[62];
      \nz.mem_765_sv2v_reg  <= data_i[61];
      \nz.mem_764_sv2v_reg  <= data_i[60];
      \nz.mem_763_sv2v_reg  <= data_i[59];
      \nz.mem_762_sv2v_reg  <= data_i[58];
      \nz.mem_761_sv2v_reg  <= data_i[57];
      \nz.mem_760_sv2v_reg  <= data_i[56];
      \nz.mem_759_sv2v_reg  <= data_i[55];
      \nz.mem_758_sv2v_reg  <= data_i[54];
      \nz.mem_757_sv2v_reg  <= data_i[53];
      \nz.mem_756_sv2v_reg  <= data_i[52];
      \nz.mem_755_sv2v_reg  <= data_i[51];
      \nz.mem_754_sv2v_reg  <= data_i[50];
      \nz.mem_753_sv2v_reg  <= data_i[49];
      \nz.mem_752_sv2v_reg  <= data_i[48];
      \nz.mem_751_sv2v_reg  <= data_i[47];
      \nz.mem_750_sv2v_reg  <= data_i[46];
      \nz.mem_749_sv2v_reg  <= data_i[45];
      \nz.mem_748_sv2v_reg  <= data_i[44];
      \nz.mem_747_sv2v_reg  <= data_i[43];
      \nz.mem_746_sv2v_reg  <= data_i[42];
      \nz.mem_745_sv2v_reg  <= data_i[41];
      \nz.mem_744_sv2v_reg  <= data_i[40];
      \nz.mem_743_sv2v_reg  <= data_i[39];
      \nz.mem_742_sv2v_reg  <= data_i[38];
      \nz.mem_741_sv2v_reg  <= data_i[37];
      \nz.mem_740_sv2v_reg  <= data_i[36];
      \nz.mem_739_sv2v_reg  <= data_i[35];
      \nz.mem_738_sv2v_reg  <= data_i[34];
      \nz.mem_737_sv2v_reg  <= data_i[33];
      \nz.mem_736_sv2v_reg  <= data_i[32];
      \nz.mem_735_sv2v_reg  <= data_i[31];
      \nz.mem_734_sv2v_reg  <= data_i[30];
      \nz.mem_733_sv2v_reg  <= data_i[29];
      \nz.mem_732_sv2v_reg  <= data_i[28];
      \nz.mem_731_sv2v_reg  <= data_i[27];
      \nz.mem_730_sv2v_reg  <= data_i[26];
      \nz.mem_729_sv2v_reg  <= data_i[25];
      \nz.mem_728_sv2v_reg  <= data_i[24];
      \nz.mem_727_sv2v_reg  <= data_i[23];
      \nz.mem_726_sv2v_reg  <= data_i[22];
      \nz.mem_725_sv2v_reg  <= data_i[21];
      \nz.mem_724_sv2v_reg  <= data_i[20];
      \nz.mem_723_sv2v_reg  <= data_i[19];
      \nz.mem_722_sv2v_reg  <= data_i[18];
      \nz.mem_721_sv2v_reg  <= data_i[17];
      \nz.mem_720_sv2v_reg  <= data_i[16];
      \nz.mem_719_sv2v_reg  <= data_i[15];
      \nz.mem_718_sv2v_reg  <= data_i[14];
      \nz.mem_717_sv2v_reg  <= data_i[13];
      \nz.mem_716_sv2v_reg  <= data_i[12];
      \nz.mem_715_sv2v_reg  <= data_i[11];
      \nz.mem_714_sv2v_reg  <= data_i[10];
      \nz.mem_713_sv2v_reg  <= data_i[9];
      \nz.mem_712_sv2v_reg  <= data_i[8];
      \nz.mem_711_sv2v_reg  <= data_i[7];
      \nz.mem_710_sv2v_reg  <= data_i[6];
      \nz.mem_709_sv2v_reg  <= data_i[5];
      \nz.mem_708_sv2v_reg  <= data_i[4];
      \nz.mem_707_sv2v_reg  <= data_i[3];
      \nz.mem_706_sv2v_reg  <= data_i[2];
      \nz.mem_705_sv2v_reg  <= data_i[1];
      \nz.mem_704_sv2v_reg  <= data_i[0];
    end 
    if(N69) begin
      \nz.mem_703_sv2v_reg  <= data_i[63];
      \nz.mem_702_sv2v_reg  <= data_i[62];
      \nz.mem_701_sv2v_reg  <= data_i[61];
      \nz.mem_700_sv2v_reg  <= data_i[60];
      \nz.mem_699_sv2v_reg  <= data_i[59];
      \nz.mem_698_sv2v_reg  <= data_i[58];
      \nz.mem_697_sv2v_reg  <= data_i[57];
      \nz.mem_696_sv2v_reg  <= data_i[56];
      \nz.mem_695_sv2v_reg  <= data_i[55];
      \nz.mem_694_sv2v_reg  <= data_i[54];
      \nz.mem_693_sv2v_reg  <= data_i[53];
      \nz.mem_692_sv2v_reg  <= data_i[52];
      \nz.mem_691_sv2v_reg  <= data_i[51];
      \nz.mem_690_sv2v_reg  <= data_i[50];
      \nz.mem_689_sv2v_reg  <= data_i[49];
      \nz.mem_688_sv2v_reg  <= data_i[48];
      \nz.mem_687_sv2v_reg  <= data_i[47];
      \nz.mem_686_sv2v_reg  <= data_i[46];
      \nz.mem_685_sv2v_reg  <= data_i[45];
      \nz.mem_684_sv2v_reg  <= data_i[44];
      \nz.mem_683_sv2v_reg  <= data_i[43];
      \nz.mem_682_sv2v_reg  <= data_i[42];
      \nz.mem_681_sv2v_reg  <= data_i[41];
      \nz.mem_680_sv2v_reg  <= data_i[40];
      \nz.mem_679_sv2v_reg  <= data_i[39];
      \nz.mem_678_sv2v_reg  <= data_i[38];
      \nz.mem_677_sv2v_reg  <= data_i[37];
      \nz.mem_676_sv2v_reg  <= data_i[36];
      \nz.mem_675_sv2v_reg  <= data_i[35];
      \nz.mem_674_sv2v_reg  <= data_i[34];
      \nz.mem_673_sv2v_reg  <= data_i[33];
      \nz.mem_672_sv2v_reg  <= data_i[32];
      \nz.mem_671_sv2v_reg  <= data_i[31];
      \nz.mem_670_sv2v_reg  <= data_i[30];
      \nz.mem_669_sv2v_reg  <= data_i[29];
      \nz.mem_668_sv2v_reg  <= data_i[28];
      \nz.mem_667_sv2v_reg  <= data_i[27];
      \nz.mem_666_sv2v_reg  <= data_i[26];
      \nz.mem_665_sv2v_reg  <= data_i[25];
      \nz.mem_664_sv2v_reg  <= data_i[24];
      \nz.mem_663_sv2v_reg  <= data_i[23];
      \nz.mem_662_sv2v_reg  <= data_i[22];
      \nz.mem_661_sv2v_reg  <= data_i[21];
      \nz.mem_660_sv2v_reg  <= data_i[20];
      \nz.mem_659_sv2v_reg  <= data_i[19];
      \nz.mem_658_sv2v_reg  <= data_i[18];
      \nz.mem_657_sv2v_reg  <= data_i[17];
      \nz.mem_656_sv2v_reg  <= data_i[16];
      \nz.mem_655_sv2v_reg  <= data_i[15];
      \nz.mem_654_sv2v_reg  <= data_i[14];
      \nz.mem_653_sv2v_reg  <= data_i[13];
      \nz.mem_652_sv2v_reg  <= data_i[12];
      \nz.mem_651_sv2v_reg  <= data_i[11];
      \nz.mem_650_sv2v_reg  <= data_i[10];
      \nz.mem_649_sv2v_reg  <= data_i[9];
      \nz.mem_648_sv2v_reg  <= data_i[8];
      \nz.mem_647_sv2v_reg  <= data_i[7];
      \nz.mem_646_sv2v_reg  <= data_i[6];
      \nz.mem_645_sv2v_reg  <= data_i[5];
      \nz.mem_644_sv2v_reg  <= data_i[4];
      \nz.mem_643_sv2v_reg  <= data_i[3];
      \nz.mem_642_sv2v_reg  <= data_i[2];
      \nz.mem_641_sv2v_reg  <= data_i[1];
      \nz.mem_640_sv2v_reg  <= data_i[0];
    end 
    if(N68) begin
      \nz.mem_639_sv2v_reg  <= data_i[63];
      \nz.mem_638_sv2v_reg  <= data_i[62];
      \nz.mem_637_sv2v_reg  <= data_i[61];
      \nz.mem_636_sv2v_reg  <= data_i[60];
      \nz.mem_635_sv2v_reg  <= data_i[59];
      \nz.mem_634_sv2v_reg  <= data_i[58];
      \nz.mem_633_sv2v_reg  <= data_i[57];
      \nz.mem_632_sv2v_reg  <= data_i[56];
      \nz.mem_631_sv2v_reg  <= data_i[55];
      \nz.mem_630_sv2v_reg  <= data_i[54];
      \nz.mem_629_sv2v_reg  <= data_i[53];
      \nz.mem_628_sv2v_reg  <= data_i[52];
      \nz.mem_627_sv2v_reg  <= data_i[51];
      \nz.mem_626_sv2v_reg  <= data_i[50];
      \nz.mem_625_sv2v_reg  <= data_i[49];
      \nz.mem_624_sv2v_reg  <= data_i[48];
      \nz.mem_623_sv2v_reg  <= data_i[47];
      \nz.mem_622_sv2v_reg  <= data_i[46];
      \nz.mem_621_sv2v_reg  <= data_i[45];
      \nz.mem_620_sv2v_reg  <= data_i[44];
      \nz.mem_619_sv2v_reg  <= data_i[43];
      \nz.mem_618_sv2v_reg  <= data_i[42];
      \nz.mem_617_sv2v_reg  <= data_i[41];
      \nz.mem_616_sv2v_reg  <= data_i[40];
      \nz.mem_615_sv2v_reg  <= data_i[39];
      \nz.mem_614_sv2v_reg  <= data_i[38];
      \nz.mem_613_sv2v_reg  <= data_i[37];
      \nz.mem_612_sv2v_reg  <= data_i[36];
      \nz.mem_611_sv2v_reg  <= data_i[35];
      \nz.mem_610_sv2v_reg  <= data_i[34];
      \nz.mem_609_sv2v_reg  <= data_i[33];
      \nz.mem_608_sv2v_reg  <= data_i[32];
      \nz.mem_607_sv2v_reg  <= data_i[31];
      \nz.mem_606_sv2v_reg  <= data_i[30];
      \nz.mem_605_sv2v_reg  <= data_i[29];
      \nz.mem_604_sv2v_reg  <= data_i[28];
      \nz.mem_603_sv2v_reg  <= data_i[27];
      \nz.mem_602_sv2v_reg  <= data_i[26];
      \nz.mem_601_sv2v_reg  <= data_i[25];
      \nz.mem_600_sv2v_reg  <= data_i[24];
      \nz.mem_599_sv2v_reg  <= data_i[23];
      \nz.mem_598_sv2v_reg  <= data_i[22];
      \nz.mem_597_sv2v_reg  <= data_i[21];
      \nz.mem_596_sv2v_reg  <= data_i[20];
      \nz.mem_595_sv2v_reg  <= data_i[19];
      \nz.mem_594_sv2v_reg  <= data_i[18];
      \nz.mem_593_sv2v_reg  <= data_i[17];
      \nz.mem_592_sv2v_reg  <= data_i[16];
      \nz.mem_591_sv2v_reg  <= data_i[15];
      \nz.mem_590_sv2v_reg  <= data_i[14];
      \nz.mem_589_sv2v_reg  <= data_i[13];
      \nz.mem_588_sv2v_reg  <= data_i[12];
      \nz.mem_587_sv2v_reg  <= data_i[11];
      \nz.mem_586_sv2v_reg  <= data_i[10];
      \nz.mem_585_sv2v_reg  <= data_i[9];
      \nz.mem_584_sv2v_reg  <= data_i[8];
      \nz.mem_583_sv2v_reg  <= data_i[7];
      \nz.mem_582_sv2v_reg  <= data_i[6];
      \nz.mem_581_sv2v_reg  <= data_i[5];
      \nz.mem_580_sv2v_reg  <= data_i[4];
      \nz.mem_579_sv2v_reg  <= data_i[3];
      \nz.mem_578_sv2v_reg  <= data_i[2];
      \nz.mem_577_sv2v_reg  <= data_i[1];
      \nz.mem_576_sv2v_reg  <= data_i[0];
    end 
    if(N67) begin
      \nz.mem_575_sv2v_reg  <= data_i[63];
      \nz.mem_574_sv2v_reg  <= data_i[62];
      \nz.mem_573_sv2v_reg  <= data_i[61];
      \nz.mem_572_sv2v_reg  <= data_i[60];
      \nz.mem_571_sv2v_reg  <= data_i[59];
      \nz.mem_570_sv2v_reg  <= data_i[58];
      \nz.mem_569_sv2v_reg  <= data_i[57];
      \nz.mem_568_sv2v_reg  <= data_i[56];
      \nz.mem_567_sv2v_reg  <= data_i[55];
      \nz.mem_566_sv2v_reg  <= data_i[54];
      \nz.mem_565_sv2v_reg  <= data_i[53];
      \nz.mem_564_sv2v_reg  <= data_i[52];
      \nz.mem_563_sv2v_reg  <= data_i[51];
      \nz.mem_562_sv2v_reg  <= data_i[50];
      \nz.mem_561_sv2v_reg  <= data_i[49];
      \nz.mem_560_sv2v_reg  <= data_i[48];
      \nz.mem_559_sv2v_reg  <= data_i[47];
      \nz.mem_558_sv2v_reg  <= data_i[46];
      \nz.mem_557_sv2v_reg  <= data_i[45];
      \nz.mem_556_sv2v_reg  <= data_i[44];
      \nz.mem_555_sv2v_reg  <= data_i[43];
      \nz.mem_554_sv2v_reg  <= data_i[42];
      \nz.mem_553_sv2v_reg  <= data_i[41];
      \nz.mem_552_sv2v_reg  <= data_i[40];
      \nz.mem_551_sv2v_reg  <= data_i[39];
      \nz.mem_550_sv2v_reg  <= data_i[38];
      \nz.mem_549_sv2v_reg  <= data_i[37];
      \nz.mem_548_sv2v_reg  <= data_i[36];
      \nz.mem_547_sv2v_reg  <= data_i[35];
      \nz.mem_546_sv2v_reg  <= data_i[34];
      \nz.mem_545_sv2v_reg  <= data_i[33];
      \nz.mem_544_sv2v_reg  <= data_i[32];
      \nz.mem_543_sv2v_reg  <= data_i[31];
      \nz.mem_542_sv2v_reg  <= data_i[30];
      \nz.mem_541_sv2v_reg  <= data_i[29];
      \nz.mem_540_sv2v_reg  <= data_i[28];
      \nz.mem_539_sv2v_reg  <= data_i[27];
      \nz.mem_538_sv2v_reg  <= data_i[26];
      \nz.mem_537_sv2v_reg  <= data_i[25];
      \nz.mem_536_sv2v_reg  <= data_i[24];
      \nz.mem_535_sv2v_reg  <= data_i[23];
      \nz.mem_534_sv2v_reg  <= data_i[22];
      \nz.mem_533_sv2v_reg  <= data_i[21];
      \nz.mem_532_sv2v_reg  <= data_i[20];
      \nz.mem_531_sv2v_reg  <= data_i[19];
      \nz.mem_530_sv2v_reg  <= data_i[18];
      \nz.mem_529_sv2v_reg  <= data_i[17];
      \nz.mem_528_sv2v_reg  <= data_i[16];
      \nz.mem_527_sv2v_reg  <= data_i[15];
      \nz.mem_526_sv2v_reg  <= data_i[14];
      \nz.mem_525_sv2v_reg  <= data_i[13];
      \nz.mem_524_sv2v_reg  <= data_i[12];
      \nz.mem_523_sv2v_reg  <= data_i[11];
      \nz.mem_522_sv2v_reg  <= data_i[10];
      \nz.mem_521_sv2v_reg  <= data_i[9];
      \nz.mem_520_sv2v_reg  <= data_i[8];
      \nz.mem_519_sv2v_reg  <= data_i[7];
      \nz.mem_518_sv2v_reg  <= data_i[6];
      \nz.mem_517_sv2v_reg  <= data_i[5];
      \nz.mem_516_sv2v_reg  <= data_i[4];
      \nz.mem_515_sv2v_reg  <= data_i[3];
      \nz.mem_514_sv2v_reg  <= data_i[2];
      \nz.mem_513_sv2v_reg  <= data_i[1];
      \nz.mem_512_sv2v_reg  <= data_i[0];
    end 
    if(N66) begin
      \nz.mem_511_sv2v_reg  <= data_i[63];
      \nz.mem_510_sv2v_reg  <= data_i[62];
      \nz.mem_509_sv2v_reg  <= data_i[61];
      \nz.mem_508_sv2v_reg  <= data_i[60];
      \nz.mem_507_sv2v_reg  <= data_i[59];
      \nz.mem_506_sv2v_reg  <= data_i[58];
      \nz.mem_505_sv2v_reg  <= data_i[57];
      \nz.mem_504_sv2v_reg  <= data_i[56];
      \nz.mem_503_sv2v_reg  <= data_i[55];
      \nz.mem_502_sv2v_reg  <= data_i[54];
      \nz.mem_501_sv2v_reg  <= data_i[53];
      \nz.mem_500_sv2v_reg  <= data_i[52];
      \nz.mem_499_sv2v_reg  <= data_i[51];
      \nz.mem_498_sv2v_reg  <= data_i[50];
      \nz.mem_497_sv2v_reg  <= data_i[49];
      \nz.mem_496_sv2v_reg  <= data_i[48];
      \nz.mem_495_sv2v_reg  <= data_i[47];
      \nz.mem_494_sv2v_reg  <= data_i[46];
      \nz.mem_493_sv2v_reg  <= data_i[45];
      \nz.mem_492_sv2v_reg  <= data_i[44];
      \nz.mem_491_sv2v_reg  <= data_i[43];
      \nz.mem_490_sv2v_reg  <= data_i[42];
      \nz.mem_489_sv2v_reg  <= data_i[41];
      \nz.mem_488_sv2v_reg  <= data_i[40];
      \nz.mem_487_sv2v_reg  <= data_i[39];
      \nz.mem_486_sv2v_reg  <= data_i[38];
      \nz.mem_485_sv2v_reg  <= data_i[37];
      \nz.mem_484_sv2v_reg  <= data_i[36];
      \nz.mem_483_sv2v_reg  <= data_i[35];
      \nz.mem_482_sv2v_reg  <= data_i[34];
      \nz.mem_481_sv2v_reg  <= data_i[33];
      \nz.mem_480_sv2v_reg  <= data_i[32];
      \nz.mem_479_sv2v_reg  <= data_i[31];
      \nz.mem_478_sv2v_reg  <= data_i[30];
      \nz.mem_477_sv2v_reg  <= data_i[29];
      \nz.mem_476_sv2v_reg  <= data_i[28];
      \nz.mem_475_sv2v_reg  <= data_i[27];
      \nz.mem_474_sv2v_reg  <= data_i[26];
      \nz.mem_473_sv2v_reg  <= data_i[25];
      \nz.mem_472_sv2v_reg  <= data_i[24];
      \nz.mem_471_sv2v_reg  <= data_i[23];
      \nz.mem_470_sv2v_reg  <= data_i[22];
      \nz.mem_469_sv2v_reg  <= data_i[21];
      \nz.mem_468_sv2v_reg  <= data_i[20];
      \nz.mem_467_sv2v_reg  <= data_i[19];
      \nz.mem_466_sv2v_reg  <= data_i[18];
      \nz.mem_465_sv2v_reg  <= data_i[17];
      \nz.mem_464_sv2v_reg  <= data_i[16];
      \nz.mem_463_sv2v_reg  <= data_i[15];
      \nz.mem_462_sv2v_reg  <= data_i[14];
      \nz.mem_461_sv2v_reg  <= data_i[13];
      \nz.mem_460_sv2v_reg  <= data_i[12];
      \nz.mem_459_sv2v_reg  <= data_i[11];
      \nz.mem_458_sv2v_reg  <= data_i[10];
      \nz.mem_457_sv2v_reg  <= data_i[9];
      \nz.mem_456_sv2v_reg  <= data_i[8];
      \nz.mem_455_sv2v_reg  <= data_i[7];
      \nz.mem_454_sv2v_reg  <= data_i[6];
      \nz.mem_453_sv2v_reg  <= data_i[5];
      \nz.mem_452_sv2v_reg  <= data_i[4];
      \nz.mem_451_sv2v_reg  <= data_i[3];
      \nz.mem_450_sv2v_reg  <= data_i[2];
      \nz.mem_449_sv2v_reg  <= data_i[1];
      \nz.mem_448_sv2v_reg  <= data_i[0];
    end 
    if(N65) begin
      \nz.mem_447_sv2v_reg  <= data_i[63];
      \nz.mem_446_sv2v_reg  <= data_i[62];
      \nz.mem_445_sv2v_reg  <= data_i[61];
      \nz.mem_444_sv2v_reg  <= data_i[60];
      \nz.mem_443_sv2v_reg  <= data_i[59];
      \nz.mem_442_sv2v_reg  <= data_i[58];
      \nz.mem_441_sv2v_reg  <= data_i[57];
      \nz.mem_440_sv2v_reg  <= data_i[56];
      \nz.mem_439_sv2v_reg  <= data_i[55];
      \nz.mem_438_sv2v_reg  <= data_i[54];
      \nz.mem_437_sv2v_reg  <= data_i[53];
      \nz.mem_436_sv2v_reg  <= data_i[52];
      \nz.mem_435_sv2v_reg  <= data_i[51];
      \nz.mem_434_sv2v_reg  <= data_i[50];
      \nz.mem_433_sv2v_reg  <= data_i[49];
      \nz.mem_432_sv2v_reg  <= data_i[48];
      \nz.mem_431_sv2v_reg  <= data_i[47];
      \nz.mem_430_sv2v_reg  <= data_i[46];
      \nz.mem_429_sv2v_reg  <= data_i[45];
      \nz.mem_428_sv2v_reg  <= data_i[44];
      \nz.mem_427_sv2v_reg  <= data_i[43];
      \nz.mem_426_sv2v_reg  <= data_i[42];
      \nz.mem_425_sv2v_reg  <= data_i[41];
      \nz.mem_424_sv2v_reg  <= data_i[40];
      \nz.mem_423_sv2v_reg  <= data_i[39];
      \nz.mem_422_sv2v_reg  <= data_i[38];
      \nz.mem_421_sv2v_reg  <= data_i[37];
      \nz.mem_420_sv2v_reg  <= data_i[36];
      \nz.mem_419_sv2v_reg  <= data_i[35];
      \nz.mem_418_sv2v_reg  <= data_i[34];
      \nz.mem_417_sv2v_reg  <= data_i[33];
      \nz.mem_416_sv2v_reg  <= data_i[32];
      \nz.mem_415_sv2v_reg  <= data_i[31];
      \nz.mem_414_sv2v_reg  <= data_i[30];
      \nz.mem_413_sv2v_reg  <= data_i[29];
      \nz.mem_412_sv2v_reg  <= data_i[28];
      \nz.mem_411_sv2v_reg  <= data_i[27];
      \nz.mem_410_sv2v_reg  <= data_i[26];
      \nz.mem_409_sv2v_reg  <= data_i[25];
      \nz.mem_408_sv2v_reg  <= data_i[24];
      \nz.mem_407_sv2v_reg  <= data_i[23];
      \nz.mem_406_sv2v_reg  <= data_i[22];
      \nz.mem_405_sv2v_reg  <= data_i[21];
      \nz.mem_404_sv2v_reg  <= data_i[20];
      \nz.mem_403_sv2v_reg  <= data_i[19];
      \nz.mem_402_sv2v_reg  <= data_i[18];
      \nz.mem_401_sv2v_reg  <= data_i[17];
      \nz.mem_400_sv2v_reg  <= data_i[16];
      \nz.mem_399_sv2v_reg  <= data_i[15];
      \nz.mem_398_sv2v_reg  <= data_i[14];
      \nz.mem_397_sv2v_reg  <= data_i[13];
      \nz.mem_396_sv2v_reg  <= data_i[12];
      \nz.mem_395_sv2v_reg  <= data_i[11];
      \nz.mem_394_sv2v_reg  <= data_i[10];
      \nz.mem_393_sv2v_reg  <= data_i[9];
      \nz.mem_392_sv2v_reg  <= data_i[8];
      \nz.mem_391_sv2v_reg  <= data_i[7];
      \nz.mem_390_sv2v_reg  <= data_i[6];
      \nz.mem_389_sv2v_reg  <= data_i[5];
      \nz.mem_388_sv2v_reg  <= data_i[4];
      \nz.mem_387_sv2v_reg  <= data_i[3];
      \nz.mem_386_sv2v_reg  <= data_i[2];
      \nz.mem_385_sv2v_reg  <= data_i[1];
      \nz.mem_384_sv2v_reg  <= data_i[0];
    end 
    if(N64) begin
      \nz.mem_383_sv2v_reg  <= data_i[63];
      \nz.mem_382_sv2v_reg  <= data_i[62];
      \nz.mem_381_sv2v_reg  <= data_i[61];
      \nz.mem_380_sv2v_reg  <= data_i[60];
      \nz.mem_379_sv2v_reg  <= data_i[59];
      \nz.mem_378_sv2v_reg  <= data_i[58];
      \nz.mem_377_sv2v_reg  <= data_i[57];
      \nz.mem_376_sv2v_reg  <= data_i[56];
      \nz.mem_375_sv2v_reg  <= data_i[55];
      \nz.mem_374_sv2v_reg  <= data_i[54];
      \nz.mem_373_sv2v_reg  <= data_i[53];
      \nz.mem_372_sv2v_reg  <= data_i[52];
      \nz.mem_371_sv2v_reg  <= data_i[51];
      \nz.mem_370_sv2v_reg  <= data_i[50];
      \nz.mem_369_sv2v_reg  <= data_i[49];
      \nz.mem_368_sv2v_reg  <= data_i[48];
      \nz.mem_367_sv2v_reg  <= data_i[47];
      \nz.mem_366_sv2v_reg  <= data_i[46];
      \nz.mem_365_sv2v_reg  <= data_i[45];
      \nz.mem_364_sv2v_reg  <= data_i[44];
      \nz.mem_363_sv2v_reg  <= data_i[43];
      \nz.mem_362_sv2v_reg  <= data_i[42];
      \nz.mem_361_sv2v_reg  <= data_i[41];
      \nz.mem_360_sv2v_reg  <= data_i[40];
      \nz.mem_359_sv2v_reg  <= data_i[39];
      \nz.mem_358_sv2v_reg  <= data_i[38];
      \nz.mem_357_sv2v_reg  <= data_i[37];
      \nz.mem_356_sv2v_reg  <= data_i[36];
      \nz.mem_355_sv2v_reg  <= data_i[35];
      \nz.mem_354_sv2v_reg  <= data_i[34];
      \nz.mem_353_sv2v_reg  <= data_i[33];
      \nz.mem_352_sv2v_reg  <= data_i[32];
      \nz.mem_351_sv2v_reg  <= data_i[31];
      \nz.mem_350_sv2v_reg  <= data_i[30];
      \nz.mem_349_sv2v_reg  <= data_i[29];
      \nz.mem_348_sv2v_reg  <= data_i[28];
      \nz.mem_347_sv2v_reg  <= data_i[27];
      \nz.mem_346_sv2v_reg  <= data_i[26];
      \nz.mem_345_sv2v_reg  <= data_i[25];
      \nz.mem_344_sv2v_reg  <= data_i[24];
      \nz.mem_343_sv2v_reg  <= data_i[23];
      \nz.mem_342_sv2v_reg  <= data_i[22];
      \nz.mem_341_sv2v_reg  <= data_i[21];
      \nz.mem_340_sv2v_reg  <= data_i[20];
      \nz.mem_339_sv2v_reg  <= data_i[19];
      \nz.mem_338_sv2v_reg  <= data_i[18];
      \nz.mem_337_sv2v_reg  <= data_i[17];
      \nz.mem_336_sv2v_reg  <= data_i[16];
      \nz.mem_335_sv2v_reg  <= data_i[15];
      \nz.mem_334_sv2v_reg  <= data_i[14];
      \nz.mem_333_sv2v_reg  <= data_i[13];
      \nz.mem_332_sv2v_reg  <= data_i[12];
      \nz.mem_331_sv2v_reg  <= data_i[11];
      \nz.mem_330_sv2v_reg  <= data_i[10];
      \nz.mem_329_sv2v_reg  <= data_i[9];
      \nz.mem_328_sv2v_reg  <= data_i[8];
      \nz.mem_327_sv2v_reg  <= data_i[7];
      \nz.mem_326_sv2v_reg  <= data_i[6];
      \nz.mem_325_sv2v_reg  <= data_i[5];
      \nz.mem_324_sv2v_reg  <= data_i[4];
      \nz.mem_323_sv2v_reg  <= data_i[3];
      \nz.mem_322_sv2v_reg  <= data_i[2];
      \nz.mem_321_sv2v_reg  <= data_i[1];
      \nz.mem_320_sv2v_reg  <= data_i[0];
    end 
    if(N63) begin
      \nz.mem_319_sv2v_reg  <= data_i[63];
      \nz.mem_318_sv2v_reg  <= data_i[62];
      \nz.mem_317_sv2v_reg  <= data_i[61];
      \nz.mem_316_sv2v_reg  <= data_i[60];
      \nz.mem_315_sv2v_reg  <= data_i[59];
      \nz.mem_314_sv2v_reg  <= data_i[58];
      \nz.mem_313_sv2v_reg  <= data_i[57];
      \nz.mem_312_sv2v_reg  <= data_i[56];
      \nz.mem_311_sv2v_reg  <= data_i[55];
      \nz.mem_310_sv2v_reg  <= data_i[54];
      \nz.mem_309_sv2v_reg  <= data_i[53];
      \nz.mem_308_sv2v_reg  <= data_i[52];
      \nz.mem_307_sv2v_reg  <= data_i[51];
      \nz.mem_306_sv2v_reg  <= data_i[50];
      \nz.mem_305_sv2v_reg  <= data_i[49];
      \nz.mem_304_sv2v_reg  <= data_i[48];
      \nz.mem_303_sv2v_reg  <= data_i[47];
      \nz.mem_302_sv2v_reg  <= data_i[46];
      \nz.mem_301_sv2v_reg  <= data_i[45];
      \nz.mem_300_sv2v_reg  <= data_i[44];
      \nz.mem_299_sv2v_reg  <= data_i[43];
      \nz.mem_298_sv2v_reg  <= data_i[42];
      \nz.mem_297_sv2v_reg  <= data_i[41];
      \nz.mem_296_sv2v_reg  <= data_i[40];
      \nz.mem_295_sv2v_reg  <= data_i[39];
      \nz.mem_294_sv2v_reg  <= data_i[38];
      \nz.mem_293_sv2v_reg  <= data_i[37];
      \nz.mem_292_sv2v_reg  <= data_i[36];
      \nz.mem_291_sv2v_reg  <= data_i[35];
      \nz.mem_290_sv2v_reg  <= data_i[34];
      \nz.mem_289_sv2v_reg  <= data_i[33];
      \nz.mem_288_sv2v_reg  <= data_i[32];
      \nz.mem_287_sv2v_reg  <= data_i[31];
      \nz.mem_286_sv2v_reg  <= data_i[30];
      \nz.mem_285_sv2v_reg  <= data_i[29];
      \nz.mem_284_sv2v_reg  <= data_i[28];
      \nz.mem_283_sv2v_reg  <= data_i[27];
      \nz.mem_282_sv2v_reg  <= data_i[26];
      \nz.mem_281_sv2v_reg  <= data_i[25];
      \nz.mem_280_sv2v_reg  <= data_i[24];
      \nz.mem_279_sv2v_reg  <= data_i[23];
      \nz.mem_278_sv2v_reg  <= data_i[22];
      \nz.mem_277_sv2v_reg  <= data_i[21];
      \nz.mem_276_sv2v_reg  <= data_i[20];
      \nz.mem_275_sv2v_reg  <= data_i[19];
      \nz.mem_274_sv2v_reg  <= data_i[18];
      \nz.mem_273_sv2v_reg  <= data_i[17];
      \nz.mem_272_sv2v_reg  <= data_i[16];
      \nz.mem_271_sv2v_reg  <= data_i[15];
      \nz.mem_270_sv2v_reg  <= data_i[14];
      \nz.mem_269_sv2v_reg  <= data_i[13];
      \nz.mem_268_sv2v_reg  <= data_i[12];
      \nz.mem_267_sv2v_reg  <= data_i[11];
      \nz.mem_266_sv2v_reg  <= data_i[10];
      \nz.mem_265_sv2v_reg  <= data_i[9];
      \nz.mem_264_sv2v_reg  <= data_i[8];
      \nz.mem_263_sv2v_reg  <= data_i[7];
      \nz.mem_262_sv2v_reg  <= data_i[6];
      \nz.mem_261_sv2v_reg  <= data_i[5];
      \nz.mem_260_sv2v_reg  <= data_i[4];
      \nz.mem_259_sv2v_reg  <= data_i[3];
      \nz.mem_258_sv2v_reg  <= data_i[2];
      \nz.mem_257_sv2v_reg  <= data_i[1];
      \nz.mem_256_sv2v_reg  <= data_i[0];
    end 
    if(N62) begin
      \nz.mem_255_sv2v_reg  <= data_i[63];
      \nz.mem_254_sv2v_reg  <= data_i[62];
      \nz.mem_253_sv2v_reg  <= data_i[61];
      \nz.mem_252_sv2v_reg  <= data_i[60];
      \nz.mem_251_sv2v_reg  <= data_i[59];
      \nz.mem_250_sv2v_reg  <= data_i[58];
      \nz.mem_249_sv2v_reg  <= data_i[57];
      \nz.mem_248_sv2v_reg  <= data_i[56];
      \nz.mem_247_sv2v_reg  <= data_i[55];
      \nz.mem_246_sv2v_reg  <= data_i[54];
      \nz.mem_245_sv2v_reg  <= data_i[53];
      \nz.mem_244_sv2v_reg  <= data_i[52];
      \nz.mem_243_sv2v_reg  <= data_i[51];
      \nz.mem_242_sv2v_reg  <= data_i[50];
      \nz.mem_241_sv2v_reg  <= data_i[49];
      \nz.mem_240_sv2v_reg  <= data_i[48];
      \nz.mem_239_sv2v_reg  <= data_i[47];
      \nz.mem_238_sv2v_reg  <= data_i[46];
      \nz.mem_237_sv2v_reg  <= data_i[45];
      \nz.mem_236_sv2v_reg  <= data_i[44];
      \nz.mem_235_sv2v_reg  <= data_i[43];
      \nz.mem_234_sv2v_reg  <= data_i[42];
      \nz.mem_233_sv2v_reg  <= data_i[41];
      \nz.mem_232_sv2v_reg  <= data_i[40];
      \nz.mem_231_sv2v_reg  <= data_i[39];
      \nz.mem_230_sv2v_reg  <= data_i[38];
      \nz.mem_229_sv2v_reg  <= data_i[37];
      \nz.mem_228_sv2v_reg  <= data_i[36];
      \nz.mem_227_sv2v_reg  <= data_i[35];
      \nz.mem_226_sv2v_reg  <= data_i[34];
      \nz.mem_225_sv2v_reg  <= data_i[33];
      \nz.mem_224_sv2v_reg  <= data_i[32];
      \nz.mem_223_sv2v_reg  <= data_i[31];
      \nz.mem_222_sv2v_reg  <= data_i[30];
      \nz.mem_221_sv2v_reg  <= data_i[29];
      \nz.mem_220_sv2v_reg  <= data_i[28];
      \nz.mem_219_sv2v_reg  <= data_i[27];
      \nz.mem_218_sv2v_reg  <= data_i[26];
      \nz.mem_217_sv2v_reg  <= data_i[25];
      \nz.mem_216_sv2v_reg  <= data_i[24];
      \nz.mem_215_sv2v_reg  <= data_i[23];
      \nz.mem_214_sv2v_reg  <= data_i[22];
      \nz.mem_213_sv2v_reg  <= data_i[21];
      \nz.mem_212_sv2v_reg  <= data_i[20];
      \nz.mem_211_sv2v_reg  <= data_i[19];
      \nz.mem_210_sv2v_reg  <= data_i[18];
      \nz.mem_209_sv2v_reg  <= data_i[17];
      \nz.mem_208_sv2v_reg  <= data_i[16];
      \nz.mem_207_sv2v_reg  <= data_i[15];
      \nz.mem_206_sv2v_reg  <= data_i[14];
      \nz.mem_205_sv2v_reg  <= data_i[13];
      \nz.mem_204_sv2v_reg  <= data_i[12];
      \nz.mem_203_sv2v_reg  <= data_i[11];
      \nz.mem_202_sv2v_reg  <= data_i[10];
      \nz.mem_201_sv2v_reg  <= data_i[9];
      \nz.mem_200_sv2v_reg  <= data_i[8];
      \nz.mem_199_sv2v_reg  <= data_i[7];
      \nz.mem_198_sv2v_reg  <= data_i[6];
      \nz.mem_197_sv2v_reg  <= data_i[5];
      \nz.mem_196_sv2v_reg  <= data_i[4];
      \nz.mem_195_sv2v_reg  <= data_i[3];
      \nz.mem_194_sv2v_reg  <= data_i[2];
      \nz.mem_193_sv2v_reg  <= data_i[1];
      \nz.mem_192_sv2v_reg  <= data_i[0];
    end 
    if(N61) begin
      \nz.mem_191_sv2v_reg  <= data_i[63];
      \nz.mem_190_sv2v_reg  <= data_i[62];
      \nz.mem_189_sv2v_reg  <= data_i[61];
      \nz.mem_188_sv2v_reg  <= data_i[60];
      \nz.mem_187_sv2v_reg  <= data_i[59];
      \nz.mem_186_sv2v_reg  <= data_i[58];
      \nz.mem_185_sv2v_reg  <= data_i[57];
      \nz.mem_184_sv2v_reg  <= data_i[56];
      \nz.mem_183_sv2v_reg  <= data_i[55];
      \nz.mem_182_sv2v_reg  <= data_i[54];
      \nz.mem_181_sv2v_reg  <= data_i[53];
      \nz.mem_180_sv2v_reg  <= data_i[52];
      \nz.mem_179_sv2v_reg  <= data_i[51];
      \nz.mem_178_sv2v_reg  <= data_i[50];
      \nz.mem_177_sv2v_reg  <= data_i[49];
      \nz.mem_176_sv2v_reg  <= data_i[48];
      \nz.mem_175_sv2v_reg  <= data_i[47];
      \nz.mem_174_sv2v_reg  <= data_i[46];
      \nz.mem_173_sv2v_reg  <= data_i[45];
      \nz.mem_172_sv2v_reg  <= data_i[44];
      \nz.mem_171_sv2v_reg  <= data_i[43];
      \nz.mem_170_sv2v_reg  <= data_i[42];
      \nz.mem_169_sv2v_reg  <= data_i[41];
      \nz.mem_168_sv2v_reg  <= data_i[40];
      \nz.mem_167_sv2v_reg  <= data_i[39];
      \nz.mem_166_sv2v_reg  <= data_i[38];
      \nz.mem_165_sv2v_reg  <= data_i[37];
      \nz.mem_164_sv2v_reg  <= data_i[36];
      \nz.mem_163_sv2v_reg  <= data_i[35];
      \nz.mem_162_sv2v_reg  <= data_i[34];
      \nz.mem_161_sv2v_reg  <= data_i[33];
      \nz.mem_160_sv2v_reg  <= data_i[32];
      \nz.mem_159_sv2v_reg  <= data_i[31];
      \nz.mem_158_sv2v_reg  <= data_i[30];
      \nz.mem_157_sv2v_reg  <= data_i[29];
      \nz.mem_156_sv2v_reg  <= data_i[28];
      \nz.mem_155_sv2v_reg  <= data_i[27];
      \nz.mem_154_sv2v_reg  <= data_i[26];
      \nz.mem_153_sv2v_reg  <= data_i[25];
      \nz.mem_152_sv2v_reg  <= data_i[24];
      \nz.mem_151_sv2v_reg  <= data_i[23];
      \nz.mem_150_sv2v_reg  <= data_i[22];
      \nz.mem_149_sv2v_reg  <= data_i[21];
      \nz.mem_148_sv2v_reg  <= data_i[20];
      \nz.mem_147_sv2v_reg  <= data_i[19];
      \nz.mem_146_sv2v_reg  <= data_i[18];
      \nz.mem_145_sv2v_reg  <= data_i[17];
      \nz.mem_144_sv2v_reg  <= data_i[16];
      \nz.mem_143_sv2v_reg  <= data_i[15];
      \nz.mem_142_sv2v_reg  <= data_i[14];
      \nz.mem_141_sv2v_reg  <= data_i[13];
      \nz.mem_140_sv2v_reg  <= data_i[12];
      \nz.mem_139_sv2v_reg  <= data_i[11];
      \nz.mem_138_sv2v_reg  <= data_i[10];
      \nz.mem_137_sv2v_reg  <= data_i[9];
      \nz.mem_136_sv2v_reg  <= data_i[8];
      \nz.mem_135_sv2v_reg  <= data_i[7];
      \nz.mem_134_sv2v_reg  <= data_i[6];
      \nz.mem_133_sv2v_reg  <= data_i[5];
      \nz.mem_132_sv2v_reg  <= data_i[4];
      \nz.mem_131_sv2v_reg  <= data_i[3];
      \nz.mem_130_sv2v_reg  <= data_i[2];
      \nz.mem_129_sv2v_reg  <= data_i[1];
      \nz.mem_128_sv2v_reg  <= data_i[0];
    end 
    if(N60) begin
      \nz.mem_127_sv2v_reg  <= data_i[63];
      \nz.mem_126_sv2v_reg  <= data_i[62];
      \nz.mem_125_sv2v_reg  <= data_i[61];
      \nz.mem_124_sv2v_reg  <= data_i[60];
      \nz.mem_123_sv2v_reg  <= data_i[59];
      \nz.mem_122_sv2v_reg  <= data_i[58];
      \nz.mem_121_sv2v_reg  <= data_i[57];
      \nz.mem_120_sv2v_reg  <= data_i[56];
      \nz.mem_119_sv2v_reg  <= data_i[55];
      \nz.mem_118_sv2v_reg  <= data_i[54];
      \nz.mem_117_sv2v_reg  <= data_i[53];
      \nz.mem_116_sv2v_reg  <= data_i[52];
      \nz.mem_115_sv2v_reg  <= data_i[51];
      \nz.mem_114_sv2v_reg  <= data_i[50];
      \nz.mem_113_sv2v_reg  <= data_i[49];
      \nz.mem_112_sv2v_reg  <= data_i[48];
      \nz.mem_111_sv2v_reg  <= data_i[47];
      \nz.mem_110_sv2v_reg  <= data_i[46];
      \nz.mem_109_sv2v_reg  <= data_i[45];
      \nz.mem_108_sv2v_reg  <= data_i[44];
      \nz.mem_107_sv2v_reg  <= data_i[43];
      \nz.mem_106_sv2v_reg  <= data_i[42];
      \nz.mem_105_sv2v_reg  <= data_i[41];
      \nz.mem_104_sv2v_reg  <= data_i[40];
      \nz.mem_103_sv2v_reg  <= data_i[39];
      \nz.mem_102_sv2v_reg  <= data_i[38];
      \nz.mem_101_sv2v_reg  <= data_i[37];
      \nz.mem_100_sv2v_reg  <= data_i[36];
      \nz.mem_99_sv2v_reg  <= data_i[35];
      \nz.mem_98_sv2v_reg  <= data_i[34];
      \nz.mem_97_sv2v_reg  <= data_i[33];
      \nz.mem_96_sv2v_reg  <= data_i[32];
      \nz.mem_95_sv2v_reg  <= data_i[31];
      \nz.mem_94_sv2v_reg  <= data_i[30];
      \nz.mem_93_sv2v_reg  <= data_i[29];
      \nz.mem_92_sv2v_reg  <= data_i[28];
      \nz.mem_91_sv2v_reg  <= data_i[27];
      \nz.mem_90_sv2v_reg  <= data_i[26];
      \nz.mem_89_sv2v_reg  <= data_i[25];
      \nz.mem_88_sv2v_reg  <= data_i[24];
      \nz.mem_87_sv2v_reg  <= data_i[23];
      \nz.mem_86_sv2v_reg  <= data_i[22];
      \nz.mem_85_sv2v_reg  <= data_i[21];
      \nz.mem_84_sv2v_reg  <= data_i[20];
      \nz.mem_83_sv2v_reg  <= data_i[19];
      \nz.mem_82_sv2v_reg  <= data_i[18];
      \nz.mem_81_sv2v_reg  <= data_i[17];
      \nz.mem_80_sv2v_reg  <= data_i[16];
      \nz.mem_79_sv2v_reg  <= data_i[15];
      \nz.mem_78_sv2v_reg  <= data_i[14];
      \nz.mem_77_sv2v_reg  <= data_i[13];
      \nz.mem_76_sv2v_reg  <= data_i[12];
      \nz.mem_75_sv2v_reg  <= data_i[11];
      \nz.mem_74_sv2v_reg  <= data_i[10];
      \nz.mem_73_sv2v_reg  <= data_i[9];
      \nz.mem_72_sv2v_reg  <= data_i[8];
      \nz.mem_71_sv2v_reg  <= data_i[7];
      \nz.mem_70_sv2v_reg  <= data_i[6];
      \nz.mem_69_sv2v_reg  <= data_i[5];
      \nz.mem_68_sv2v_reg  <= data_i[4];
      \nz.mem_67_sv2v_reg  <= data_i[3];
      \nz.mem_66_sv2v_reg  <= data_i[2];
      \nz.mem_65_sv2v_reg  <= data_i[1];
      \nz.mem_64_sv2v_reg  <= data_i[0];
    end 
    if(N59) begin
      \nz.mem_63_sv2v_reg  <= data_i[63];
      \nz.mem_62_sv2v_reg  <= data_i[62];
      \nz.mem_61_sv2v_reg  <= data_i[61];
      \nz.mem_60_sv2v_reg  <= data_i[60];
      \nz.mem_59_sv2v_reg  <= data_i[59];
      \nz.mem_58_sv2v_reg  <= data_i[58];
      \nz.mem_57_sv2v_reg  <= data_i[57];
      \nz.mem_56_sv2v_reg  <= data_i[56];
      \nz.mem_55_sv2v_reg  <= data_i[55];
      \nz.mem_54_sv2v_reg  <= data_i[54];
      \nz.mem_53_sv2v_reg  <= data_i[53];
      \nz.mem_52_sv2v_reg  <= data_i[52];
      \nz.mem_51_sv2v_reg  <= data_i[51];
      \nz.mem_50_sv2v_reg  <= data_i[50];
      \nz.mem_49_sv2v_reg  <= data_i[49];
      \nz.mem_48_sv2v_reg  <= data_i[48];
      \nz.mem_47_sv2v_reg  <= data_i[47];
      \nz.mem_46_sv2v_reg  <= data_i[46];
      \nz.mem_45_sv2v_reg  <= data_i[45];
      \nz.mem_44_sv2v_reg  <= data_i[44];
      \nz.mem_43_sv2v_reg  <= data_i[43];
      \nz.mem_42_sv2v_reg  <= data_i[42];
      \nz.mem_41_sv2v_reg  <= data_i[41];
      \nz.mem_40_sv2v_reg  <= data_i[40];
      \nz.mem_39_sv2v_reg  <= data_i[39];
      \nz.mem_38_sv2v_reg  <= data_i[38];
      \nz.mem_37_sv2v_reg  <= data_i[37];
      \nz.mem_36_sv2v_reg  <= data_i[36];
      \nz.mem_35_sv2v_reg  <= data_i[35];
      \nz.mem_34_sv2v_reg  <= data_i[34];
      \nz.mem_33_sv2v_reg  <= data_i[33];
      \nz.mem_32_sv2v_reg  <= data_i[32];
      \nz.mem_31_sv2v_reg  <= data_i[31];
      \nz.mem_30_sv2v_reg  <= data_i[30];
      \nz.mem_29_sv2v_reg  <= data_i[29];
      \nz.mem_28_sv2v_reg  <= data_i[28];
      \nz.mem_27_sv2v_reg  <= data_i[27];
      \nz.mem_26_sv2v_reg  <= data_i[26];
      \nz.mem_25_sv2v_reg  <= data_i[25];
      \nz.mem_24_sv2v_reg  <= data_i[24];
      \nz.mem_23_sv2v_reg  <= data_i[23];
      \nz.mem_22_sv2v_reg  <= data_i[22];
      \nz.mem_21_sv2v_reg  <= data_i[21];
      \nz.mem_20_sv2v_reg  <= data_i[20];
      \nz.mem_19_sv2v_reg  <= data_i[19];
      \nz.mem_18_sv2v_reg  <= data_i[18];
      \nz.mem_17_sv2v_reg  <= data_i[17];
      \nz.mem_16_sv2v_reg  <= data_i[16];
      \nz.mem_15_sv2v_reg  <= data_i[15];
      \nz.mem_14_sv2v_reg  <= data_i[14];
      \nz.mem_13_sv2v_reg  <= data_i[13];
      \nz.mem_12_sv2v_reg  <= data_i[12];
      \nz.mem_11_sv2v_reg  <= data_i[11];
      \nz.mem_10_sv2v_reg  <= data_i[10];
      \nz.mem_9_sv2v_reg  <= data_i[9];
      \nz.mem_8_sv2v_reg  <= data_i[8];
      \nz.mem_7_sv2v_reg  <= data_i[7];
      \nz.mem_6_sv2v_reg  <= data_i[6];
      \nz.mem_5_sv2v_reg  <= data_i[5];
      \nz.mem_4_sv2v_reg  <= data_i[4];
      \nz.mem_3_sv2v_reg  <= data_i[3];
      \nz.mem_2_sv2v_reg  <= data_i[2];
      \nz.mem_1_sv2v_reg  <= data_i[1];
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_width_p64_els_p16
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [63:0] data_i;
  input [3:0] addr_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  bsg_mem_1rw_sync_synth_width_p64_els_p16_latch_last_read_p0_verbose_p1
  synth
  (
    .clk_i(clk_i),
    .v_i(v_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_fifo_1rw_large_width_p64_els_p16
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  enq_not_deq_i,
  full_o,
  empty_o,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input enq_not_deq_i;
  output full_o;
  output empty_o;
  wire [63:0] data_o;
  wire full_o,empty_o,N0,N1,N2,mem_we,mem_re,N3,N4,last_op_is_read_r,N5,N6,N7,
  _0_net__3_,_0_net__2_,_0_net__1_,_0_net__0_,N8,N9,N10,N11,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,
  sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8;
  wire [3:0] rd_ptr,wr_ptr;
  reg last_op_is_read_r_sv2v_reg;
  assign last_op_is_read_r = last_op_is_read_r_sv2v_reg;
  assign N6 = rd_ptr == wr_ptr;
  assign N7 = rd_ptr == wr_ptr;

  bsg_circular_ptr_slots_p16_max_add_p1
  rd_circ_ptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(mem_re),
    .o(rd_ptr),
    .n_o({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4 })
  );


  bsg_circular_ptr_slots_p16_max_add_p1
  wr_circ_ptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(mem_we),
    .o(wr_ptr),
    .n_o({ sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8 })
  );


  bsg_mem_1rw_sync_width_p64_els_p16
  mem_1srw
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i({ _0_net__3_, _0_net__2_, _0_net__1_, _0_net__0_ }),
    .v_i(v_i),
    .w_i(mem_we),
    .data_o(data_o)
  );

  assign N5 = (N0)? 1'b1 : 
              (N4)? 1'b0 : 1'b0;
  assign N0 = N3;
  assign { _0_net__3_, _0_net__2_, _0_net__1_, _0_net__0_ } = (N1)? wr_ptr : 
                                                              (N2)? rd_ptr : 1'b0;
  assign N1 = N9;
  assign N2 = N8;
  assign mem_we = enq_not_deq_i & v_i;
  assign mem_re = N10 & v_i;
  assign N10 = ~enq_not_deq_i;
  assign N3 = v_i;
  assign N4 = ~N3;
  assign empty_o = N6 & last_op_is_read_r;
  assign full_o = N7 & N11;
  assign N11 = ~last_op_is_read_r;
  assign N8 = ~mem_we;
  assign N9 = mem_we;

  always @(posedge clk_i) begin
    if(reset_i) begin
      last_op_is_read_r_sv2v_reg <= 1'b1;
    end else if(N5) begin
      last_op_is_read_r_sv2v_reg <= mem_re;
    end 
  end


endmodule



module bsg_thermometer_count_width_p2
(
  i,
  o
);

  input [1:0] i;
  output [1:0] o;
  wire [1:0] o;
  wire o_1_,N0;
  assign o_1_ = i[1];
  assign o[1] = o_1_;
  assign o[0] = i[0] & N0;
  assign N0 = ~o_1_;

endmodule



module bsg_round_robin_2_to_2_width_p32
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  ready_i
);

  input [63:0] data_i;
  input [1:0] v_i;
  output [1:0] ready_o;
  output [63:0] data_o;
  output [1:0] v_o;
  input [1:0] ready_i;
  input clk_i;
  input reset_i;
  wire [1:0] ready_o,v_o;
  wire [63:0] data_o;
  wire N0,N1,head_r,N2,N3,N4,N5,N6;
  reg head_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign data_o = (N0)? { data_i[31:0], data_i[63:32] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = head_r;
  assign N1 = N3;
  assign v_o = (N0)? { v_i[0:0], v_i[1:1] } : 
               (N1)? v_i : 1'b0;
  assign ready_o = (N0)? { ready_i[0:0], ready_i[1:1] } : 
                   (N1)? ready_i : 1'b0;
  assign N2 = N5 ^ N6;
  assign N5 = head_r ^ N4;
  assign N4 = v_i[1] & ready_o[1];
  assign N6 = v_i[0] & ready_o[0];
  assign N3 = ~head_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [63:0] \nz.mem ;
  reg \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [62] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [61] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [60] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [59] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [58] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [57] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [56] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [55] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [54] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [53] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [52] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [51] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [50] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [49] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [48] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [47] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [46] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [45] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [44] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [43] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [42] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [41] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [40] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [39] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [38] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [37] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [36] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [35] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [34] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [33] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_63_sv2v_reg  <= w_data_i[31];
      \nz.mem_62_sv2v_reg  <= w_data_i[30];
      \nz.mem_61_sv2v_reg  <= w_data_i[29];
      \nz.mem_60_sv2v_reg  <= w_data_i[28];
      \nz.mem_59_sv2v_reg  <= w_data_i[27];
      \nz.mem_58_sv2v_reg  <= w_data_i[26];
      \nz.mem_57_sv2v_reg  <= w_data_i[25];
      \nz.mem_56_sv2v_reg  <= w_data_i[24];
      \nz.mem_55_sv2v_reg  <= w_data_i[23];
      \nz.mem_54_sv2v_reg  <= w_data_i[22];
      \nz.mem_53_sv2v_reg  <= w_data_i[21];
      \nz.mem_52_sv2v_reg  <= w_data_i[20];
      \nz.mem_51_sv2v_reg  <= w_data_i[19];
      \nz.mem_50_sv2v_reg  <= w_data_i[18];
      \nz.mem_49_sv2v_reg  <= w_data_i[17];
      \nz.mem_48_sv2v_reg  <= w_data_i[16];
      \nz.mem_47_sv2v_reg  <= w_data_i[15];
      \nz.mem_46_sv2v_reg  <= w_data_i[14];
      \nz.mem_45_sv2v_reg  <= w_data_i[13];
      \nz.mem_44_sv2v_reg  <= w_data_i[12];
      \nz.mem_43_sv2v_reg  <= w_data_i[11];
      \nz.mem_42_sv2v_reg  <= w_data_i[10];
      \nz.mem_41_sv2v_reg  <= w_data_i[9];
      \nz.mem_40_sv2v_reg  <= w_data_i[8];
      \nz.mem_39_sv2v_reg  <= w_data_i[7];
      \nz.mem_38_sv2v_reg  <= w_data_i[6];
      \nz.mem_37_sv2v_reg  <= w_data_i[5];
      \nz.mem_36_sv2v_reg  <= w_data_i[4];
      \nz.mem_35_sv2v_reg  <= w_data_i[3];
      \nz.mem_34_sv2v_reg  <= w_data_i[2];
      \nz.mem_33_sv2v_reg  <= w_data_i[1];
      \nz.mem_32_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_circular_ptr_slots_p2_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [0:0] o;
  output [0:0] n_o;
  input clk;
  input reset_i;
  wire [0:0] o,n_o,\genblk1.genblk1.ptr_r_p1 ;
  wire N0,N1,N2;
  reg o_0_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign \genblk1.genblk1.ptr_r_p1 [0] = o[0] ^ 1'b1;
  assign n_o[0] = (N0)? \genblk1.genblk1.ptr_r_p1 [0] : 
                  (N1)? o[0] : 1'b0;
  assign N0 = add_i[0];
  assign N1 = N2;
  assign N2 = ~add_i[0];

  always @(posedge clk) begin
    if(reset_i) begin
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_round_robin_n_to_1_width_p32_num_in_p2_strict_p1
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  v_o,
  data_o,
  tag_o,
  yumi_i
);

  input [63:0] data_i;
  input [1:0] v_i;
  output [1:0] yumi_o;
  output [31:0] data_o;
  output [0:0] tag_o;
  input clk_i;
  input reset_i;
  input yumi_i;
  output v_o;
  wire [1:0] yumi_o;
  wire [31:0] data_o;
  wire [0:0] tag_o;
  wire v_o,N0,N1,sv2v_dc_1;

  bsg_circular_ptr_slots_p2_max_add_p1
  \strict.circular_ptr 
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(yumi_i),
    .o(tag_o[0]),
    .n_o(sv2v_dc_1)
  );

  assign v_o = (N1)? v_i[0] : 
               (N0)? v_i[1] : 1'b0;
  assign N0 = tag_o[0];
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[63] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[62] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[61] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[60] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[59] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[58] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[57] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[56] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[55] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[54] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[53] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[52] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[51] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[50] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[49] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[48] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[47] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[46] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[45] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[44] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[43] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[42] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[41] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[40] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[39] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[38] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[37] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[36] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[35] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[34] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[33] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[32] : 1'b0;
  assign yumi_o = { 1'b0, yumi_i } << tag_o[0];
  assign N1 = ~tag_o[0];

endmodule



module bsg_fifo_1r1w_large_width_p32_els_p32
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,N0,N1,N2,N3,big_deq_r,big_deq,big_valid,big_full_lo,big_empty_lo,
  bypass_mode,can_spill,emergency,will_spill,N4,N5,N6,_0_net__1_,_0_net__0_,N7,N8,N9,
  N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,sv2v_dc_1;
  wire [1:0] valid_sipo,yumi_cnt_sipo,little_ready,little_ready_rot,valid_int,bypass_vector,
  little_valid,cnt,little_valid_rot,yumi_int;
  wire [63:0] data_sipo,big_data_lo,little_data,little_data_rot,data_int;
  reg big_deq_r_sv2v_reg;
  assign big_deq_r = big_deq_r_sv2v_reg;

  bsg_serial_in_parallel_out_width_p32_els_p3_out_els_p2
  sipo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .valid_i(v_i),
    .data_i(data_i),
    .ready_o(ready_o),
    .valid_o(valid_sipo),
    .data_o(data_sipo),
    .yumi_cnt_i(yumi_cnt_sipo)
  );


  bsg_fifo_1rw_large_width_p64_els_p16
  big1p
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_sipo),
    .v_i(big_valid),
    .enq_not_deq_i(will_spill),
    .full_o(big_full_lo),
    .empty_o(big_empty_lo),
    .data_o(big_data_lo)
  );


  bsg_thermometer_count_width_p2
  thermo
  (
    .i({ _0_net__1_, _0_net__0_ }),
    .o(cnt)
  );


  bsg_round_robin_2_to_2_width_p32
  rr222
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(little_data),
    .v_i(little_valid),
    .ready_o(little_ready),
    .data_o(little_data_rot),
    .v_o(little_valid_rot),
    .ready_i(little_ready_rot)
  );


  bsg_two_fifo_width_p32
  \twofer_0_.little 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(little_ready_rot[0]),
    .data_i(little_data_rot[31:0]),
    .v_i(little_valid_rot[0]),
    .v_o(valid_int[0]),
    .data_o(data_int[31:0]),
    .yumi_i(yumi_int[0])
  );


  bsg_two_fifo_width_p32
  \twofer_1_.little 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(little_ready_rot[1]),
    .data_i(little_data_rot[63:32]),
    .v_i(little_valid_rot[1]),
    .v_o(valid_int[1]),
    .data_o(data_int[63:32]),
    .yumi_i(yumi_int[1])
  );


  bsg_round_robin_n_to_1_width_p32_num_in_p2_strict_p1
  round_robin_n_to_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_int),
    .v_i(valid_int),
    .yumi_o(yumi_int),
    .v_o(v_o),
    .data_o(data_o),
    .tag_o(sv2v_dc_1),
    .yumi_i(yumi_i)
  );

  assign N6 = (N0)? N4 : 
              (N1)? N5 : 1'b0;
  assign N0 = big_deq_r;
  assign N1 = N9;
  assign little_data = (N0)? big_data_lo : 
                       (N1)? data_sipo : 1'b0;
  assign little_valid = (N0)? { 1'b1, 1'b1 } : 
                        (N1)? bypass_vector : 1'b0;
  assign yumi_cnt_sipo = (N2)? { 1'b1, 1'b0 } : 
                         (N3)? cnt : 1'b0;
  assign N2 = N8;
  assign N3 = N7;
  assign bypass_mode = N10 & big_empty_lo;
  assign N10 = N9 & little_ready[0];
  assign N9 = ~big_deq_r;
  assign can_spill = N11 & N12;
  assign N11 = ~big_full_lo;
  assign N12 = ~bypass_mode;
  assign emergency = N15 & N9;
  assign N15 = N13 & N14;
  assign N13 = little_ready_rot[1] & little_ready_rot[0];
  assign N14 = ~big_empty_lo;
  assign will_spill = N17 & N18;
  assign N17 = can_spill & N16;
  assign N16 = valid_sipo[1] & valid_sipo[0];
  assign N18 = ~emergency;
  assign N4 = ~N19;
  assign N19 = valid_int[1] | valid_int[0];
  assign N5 = little_ready_rot[1] & little_ready_rot[0];
  assign big_deq = N21 & N6;
  assign N21 = N20 & N14;
  assign N20 = ~will_spill;
  assign big_valid = will_spill | big_deq;
  assign bypass_vector[1] = valid_sipo[1] & bypass_mode;
  assign bypass_vector[0] = valid_sipo[0] & bypass_mode;
  assign _0_net__1_ = little_ready[1] & bypass_vector[1];
  assign _0_net__0_ = little_ready[0] & bypass_vector[0];
  assign N7 = ~will_spill;
  assign N8 = will_spill;

  always @(posedge clk_i) begin
    if(1'b1) begin
      big_deq_r_sv2v_reg <= big_deq;
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p7_init_val_p0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [2:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [2:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N2,N3,N7,N30,N16;
  reg count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N16 = reset_i | clear_i;
  assign { N8, N6, N5 } = count_o + 1'b1;
  assign N9 = (N0)? 1'b1 : 
              (N7)? 1'b1 : 
              (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N11 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N10 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N15;
  assign N12 = ~reset_i;
  assign N13 = ~clear_i;
  assign N14 = N12 & N13;
  assign N15 = up_i & N14;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N13;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N16) begin
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N11) begin
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N9) begin
      count_o_0_sv2v_reg <= N10;
    end 
  end


endmodule



module bsg_cache_to_dram_ctrl_rx
(
  clk_i,
  reset_i,
  dma_data_o,
  dma_data_v_o,
  dma_data_ready_i,
  app_rd_data_valid_i,
  app_rd_data_end_i,
  app_rd_data_i
);

  output [31:0] dma_data_o;
  input [31:0] app_rd_data_i;
  input clk_i;
  input reset_i;
  input dma_data_ready_i;
  input app_rd_data_valid_i;
  input app_rd_data_end_i;
  output dma_data_v_o;
  wire [31:0] dma_data_o;
  wire dma_data_v_o,N0,fifo_yumi_li,counter_clear_li,counter_up_li,N1,N2,N3;
  wire [2:0] count_lo;

  bsg_fifo_1r1w_large_width_p32_els_p32
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(app_rd_data_i),
    .v_i(app_rd_data_valid_i),
    .v_o(dma_data_v_o),
    .data_o(dma_data_o),
    .yumi_i(fifo_yumi_li)
  );


  bsg_counter_clear_up_max_val_p7_init_val_p0
  counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(counter_clear_li),
    .up_i(counter_up_li),
    .count_o(count_lo)
  );

  assign N2 = count_lo[1] & count_lo[2];
  assign N3 = count_lo[0] & N2;
  assign counter_clear_li = (N0)? fifo_yumi_li : 
                            (N1)? 1'b0 : 1'b0;
  assign N0 = N3;
  assign counter_up_li = (N0)? 1'b0 : 
                         (N1)? fifo_yumi_li : 1'b0;
  assign fifo_yumi_li = dma_data_v_o & dma_data_ready_i;
  assign N1 = ~N3;

endmodule

