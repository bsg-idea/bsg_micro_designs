

module top
(
  en_ls_i,
  clk_i,
  reset_i,
  clk_o,
  reset_o,
  fsb_v_i_o,
  fsb_data_i_o,
  fsb_yumi_o_i,
  fsb_v_o_i,
  fsb_data_o_i,
  fsb_ready_i_o,
  node_v_i_o,
  node_data_i_o,
  node_ready_o_i,
  node_v_o_i,
  node_data_o_i,
  node_yumi_i_o
);

  output [999:0] fsb_data_i_o;
  input [999:0] fsb_data_o_i;
  output [999:0] node_data_i_o;
  input [999:0] node_data_o_i;
  input en_ls_i;
  input clk_i;
  input reset_i;
  input fsb_yumi_o_i;
  input fsb_v_o_i;
  input node_ready_o_i;
  input node_v_o_i;
  output clk_o;
  output reset_o;
  output fsb_v_i_o;
  output fsb_ready_i_o;
  output node_v_i_o;
  output node_yumi_i_o;

  bsg_fsb_node_level_shift_fsb_domain
  wrapper
  (
    .fsb_data_i_o(fsb_data_i_o),
    .fsb_data_o_i(fsb_data_o_i),
    .node_data_i_o(node_data_i_o),
    .node_data_o_i(node_data_o_i),
    .en_ls_i(en_ls_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fsb_yumi_o_i(fsb_yumi_o_i),
    .fsb_v_o_i(fsb_v_o_i),
    .node_ready_o_i(node_ready_o_i),
    .node_v_o_i(node_v_o_i),
    .clk_o(clk_o),
    .reset_o(reset_o),
    .fsb_v_i_o(fsb_v_i_o),
    .fsb_ready_i_o(fsb_ready_i_o),
    .node_v_i_o(node_v_i_o),
    .node_yumi_i_o(node_yumi_i_o)
  );


endmodule



module bsg_level_shift_up_down_source_width_p1
(
  v0_en_i,
  v0_data_i,
  v1_data_o
);

  input [0:0] v0_data_i;
  output [0:0] v1_data_o;
  input v0_en_i;
  wire [0:0] v1_data_o;
  assign v1_data_o[0] = v0_data_i[0] & v0_en_i;

endmodule



module bsg_level_shift_up_down_sink_width_p1
(
  v0_data_i,
  v1_en_i,
  v1_data_o
);

  input [0:0] v0_data_i;
  output [0:0] v1_data_o;
  input v1_en_i;
  wire [0:0] v1_data_o;
  assign v1_data_o[0] = v0_data_i[0] & v1_en_i;

endmodule



module bsg_level_shift_up_down_sink_width_p1000
(
  v0_data_i,
  v1_en_i,
  v1_data_o
);

  input [999:0] v0_data_i;
  output [999:0] v1_data_o;
  input v1_en_i;
  wire [999:0] v1_data_o;
  assign v1_data_o[999] = v0_data_i[999] & v1_en_i;
  assign v1_data_o[998] = v0_data_i[998] & v1_en_i;
  assign v1_data_o[997] = v0_data_i[997] & v1_en_i;
  assign v1_data_o[996] = v0_data_i[996] & v1_en_i;
  assign v1_data_o[995] = v0_data_i[995] & v1_en_i;
  assign v1_data_o[994] = v0_data_i[994] & v1_en_i;
  assign v1_data_o[993] = v0_data_i[993] & v1_en_i;
  assign v1_data_o[992] = v0_data_i[992] & v1_en_i;
  assign v1_data_o[991] = v0_data_i[991] & v1_en_i;
  assign v1_data_o[990] = v0_data_i[990] & v1_en_i;
  assign v1_data_o[989] = v0_data_i[989] & v1_en_i;
  assign v1_data_o[988] = v0_data_i[988] & v1_en_i;
  assign v1_data_o[987] = v0_data_i[987] & v1_en_i;
  assign v1_data_o[986] = v0_data_i[986] & v1_en_i;
  assign v1_data_o[985] = v0_data_i[985] & v1_en_i;
  assign v1_data_o[984] = v0_data_i[984] & v1_en_i;
  assign v1_data_o[983] = v0_data_i[983] & v1_en_i;
  assign v1_data_o[982] = v0_data_i[982] & v1_en_i;
  assign v1_data_o[981] = v0_data_i[981] & v1_en_i;
  assign v1_data_o[980] = v0_data_i[980] & v1_en_i;
  assign v1_data_o[979] = v0_data_i[979] & v1_en_i;
  assign v1_data_o[978] = v0_data_i[978] & v1_en_i;
  assign v1_data_o[977] = v0_data_i[977] & v1_en_i;
  assign v1_data_o[976] = v0_data_i[976] & v1_en_i;
  assign v1_data_o[975] = v0_data_i[975] & v1_en_i;
  assign v1_data_o[974] = v0_data_i[974] & v1_en_i;
  assign v1_data_o[973] = v0_data_i[973] & v1_en_i;
  assign v1_data_o[972] = v0_data_i[972] & v1_en_i;
  assign v1_data_o[971] = v0_data_i[971] & v1_en_i;
  assign v1_data_o[970] = v0_data_i[970] & v1_en_i;
  assign v1_data_o[969] = v0_data_i[969] & v1_en_i;
  assign v1_data_o[968] = v0_data_i[968] & v1_en_i;
  assign v1_data_o[967] = v0_data_i[967] & v1_en_i;
  assign v1_data_o[966] = v0_data_i[966] & v1_en_i;
  assign v1_data_o[965] = v0_data_i[965] & v1_en_i;
  assign v1_data_o[964] = v0_data_i[964] & v1_en_i;
  assign v1_data_o[963] = v0_data_i[963] & v1_en_i;
  assign v1_data_o[962] = v0_data_i[962] & v1_en_i;
  assign v1_data_o[961] = v0_data_i[961] & v1_en_i;
  assign v1_data_o[960] = v0_data_i[960] & v1_en_i;
  assign v1_data_o[959] = v0_data_i[959] & v1_en_i;
  assign v1_data_o[958] = v0_data_i[958] & v1_en_i;
  assign v1_data_o[957] = v0_data_i[957] & v1_en_i;
  assign v1_data_o[956] = v0_data_i[956] & v1_en_i;
  assign v1_data_o[955] = v0_data_i[955] & v1_en_i;
  assign v1_data_o[954] = v0_data_i[954] & v1_en_i;
  assign v1_data_o[953] = v0_data_i[953] & v1_en_i;
  assign v1_data_o[952] = v0_data_i[952] & v1_en_i;
  assign v1_data_o[951] = v0_data_i[951] & v1_en_i;
  assign v1_data_o[950] = v0_data_i[950] & v1_en_i;
  assign v1_data_o[949] = v0_data_i[949] & v1_en_i;
  assign v1_data_o[948] = v0_data_i[948] & v1_en_i;
  assign v1_data_o[947] = v0_data_i[947] & v1_en_i;
  assign v1_data_o[946] = v0_data_i[946] & v1_en_i;
  assign v1_data_o[945] = v0_data_i[945] & v1_en_i;
  assign v1_data_o[944] = v0_data_i[944] & v1_en_i;
  assign v1_data_o[943] = v0_data_i[943] & v1_en_i;
  assign v1_data_o[942] = v0_data_i[942] & v1_en_i;
  assign v1_data_o[941] = v0_data_i[941] & v1_en_i;
  assign v1_data_o[940] = v0_data_i[940] & v1_en_i;
  assign v1_data_o[939] = v0_data_i[939] & v1_en_i;
  assign v1_data_o[938] = v0_data_i[938] & v1_en_i;
  assign v1_data_o[937] = v0_data_i[937] & v1_en_i;
  assign v1_data_o[936] = v0_data_i[936] & v1_en_i;
  assign v1_data_o[935] = v0_data_i[935] & v1_en_i;
  assign v1_data_o[934] = v0_data_i[934] & v1_en_i;
  assign v1_data_o[933] = v0_data_i[933] & v1_en_i;
  assign v1_data_o[932] = v0_data_i[932] & v1_en_i;
  assign v1_data_o[931] = v0_data_i[931] & v1_en_i;
  assign v1_data_o[930] = v0_data_i[930] & v1_en_i;
  assign v1_data_o[929] = v0_data_i[929] & v1_en_i;
  assign v1_data_o[928] = v0_data_i[928] & v1_en_i;
  assign v1_data_o[927] = v0_data_i[927] & v1_en_i;
  assign v1_data_o[926] = v0_data_i[926] & v1_en_i;
  assign v1_data_o[925] = v0_data_i[925] & v1_en_i;
  assign v1_data_o[924] = v0_data_i[924] & v1_en_i;
  assign v1_data_o[923] = v0_data_i[923] & v1_en_i;
  assign v1_data_o[922] = v0_data_i[922] & v1_en_i;
  assign v1_data_o[921] = v0_data_i[921] & v1_en_i;
  assign v1_data_o[920] = v0_data_i[920] & v1_en_i;
  assign v1_data_o[919] = v0_data_i[919] & v1_en_i;
  assign v1_data_o[918] = v0_data_i[918] & v1_en_i;
  assign v1_data_o[917] = v0_data_i[917] & v1_en_i;
  assign v1_data_o[916] = v0_data_i[916] & v1_en_i;
  assign v1_data_o[915] = v0_data_i[915] & v1_en_i;
  assign v1_data_o[914] = v0_data_i[914] & v1_en_i;
  assign v1_data_o[913] = v0_data_i[913] & v1_en_i;
  assign v1_data_o[912] = v0_data_i[912] & v1_en_i;
  assign v1_data_o[911] = v0_data_i[911] & v1_en_i;
  assign v1_data_o[910] = v0_data_i[910] & v1_en_i;
  assign v1_data_o[909] = v0_data_i[909] & v1_en_i;
  assign v1_data_o[908] = v0_data_i[908] & v1_en_i;
  assign v1_data_o[907] = v0_data_i[907] & v1_en_i;
  assign v1_data_o[906] = v0_data_i[906] & v1_en_i;
  assign v1_data_o[905] = v0_data_i[905] & v1_en_i;
  assign v1_data_o[904] = v0_data_i[904] & v1_en_i;
  assign v1_data_o[903] = v0_data_i[903] & v1_en_i;
  assign v1_data_o[902] = v0_data_i[902] & v1_en_i;
  assign v1_data_o[901] = v0_data_i[901] & v1_en_i;
  assign v1_data_o[900] = v0_data_i[900] & v1_en_i;
  assign v1_data_o[899] = v0_data_i[899] & v1_en_i;
  assign v1_data_o[898] = v0_data_i[898] & v1_en_i;
  assign v1_data_o[897] = v0_data_i[897] & v1_en_i;
  assign v1_data_o[896] = v0_data_i[896] & v1_en_i;
  assign v1_data_o[895] = v0_data_i[895] & v1_en_i;
  assign v1_data_o[894] = v0_data_i[894] & v1_en_i;
  assign v1_data_o[893] = v0_data_i[893] & v1_en_i;
  assign v1_data_o[892] = v0_data_i[892] & v1_en_i;
  assign v1_data_o[891] = v0_data_i[891] & v1_en_i;
  assign v1_data_o[890] = v0_data_i[890] & v1_en_i;
  assign v1_data_o[889] = v0_data_i[889] & v1_en_i;
  assign v1_data_o[888] = v0_data_i[888] & v1_en_i;
  assign v1_data_o[887] = v0_data_i[887] & v1_en_i;
  assign v1_data_o[886] = v0_data_i[886] & v1_en_i;
  assign v1_data_o[885] = v0_data_i[885] & v1_en_i;
  assign v1_data_o[884] = v0_data_i[884] & v1_en_i;
  assign v1_data_o[883] = v0_data_i[883] & v1_en_i;
  assign v1_data_o[882] = v0_data_i[882] & v1_en_i;
  assign v1_data_o[881] = v0_data_i[881] & v1_en_i;
  assign v1_data_o[880] = v0_data_i[880] & v1_en_i;
  assign v1_data_o[879] = v0_data_i[879] & v1_en_i;
  assign v1_data_o[878] = v0_data_i[878] & v1_en_i;
  assign v1_data_o[877] = v0_data_i[877] & v1_en_i;
  assign v1_data_o[876] = v0_data_i[876] & v1_en_i;
  assign v1_data_o[875] = v0_data_i[875] & v1_en_i;
  assign v1_data_o[874] = v0_data_i[874] & v1_en_i;
  assign v1_data_o[873] = v0_data_i[873] & v1_en_i;
  assign v1_data_o[872] = v0_data_i[872] & v1_en_i;
  assign v1_data_o[871] = v0_data_i[871] & v1_en_i;
  assign v1_data_o[870] = v0_data_i[870] & v1_en_i;
  assign v1_data_o[869] = v0_data_i[869] & v1_en_i;
  assign v1_data_o[868] = v0_data_i[868] & v1_en_i;
  assign v1_data_o[867] = v0_data_i[867] & v1_en_i;
  assign v1_data_o[866] = v0_data_i[866] & v1_en_i;
  assign v1_data_o[865] = v0_data_i[865] & v1_en_i;
  assign v1_data_o[864] = v0_data_i[864] & v1_en_i;
  assign v1_data_o[863] = v0_data_i[863] & v1_en_i;
  assign v1_data_o[862] = v0_data_i[862] & v1_en_i;
  assign v1_data_o[861] = v0_data_i[861] & v1_en_i;
  assign v1_data_o[860] = v0_data_i[860] & v1_en_i;
  assign v1_data_o[859] = v0_data_i[859] & v1_en_i;
  assign v1_data_o[858] = v0_data_i[858] & v1_en_i;
  assign v1_data_o[857] = v0_data_i[857] & v1_en_i;
  assign v1_data_o[856] = v0_data_i[856] & v1_en_i;
  assign v1_data_o[855] = v0_data_i[855] & v1_en_i;
  assign v1_data_o[854] = v0_data_i[854] & v1_en_i;
  assign v1_data_o[853] = v0_data_i[853] & v1_en_i;
  assign v1_data_o[852] = v0_data_i[852] & v1_en_i;
  assign v1_data_o[851] = v0_data_i[851] & v1_en_i;
  assign v1_data_o[850] = v0_data_i[850] & v1_en_i;
  assign v1_data_o[849] = v0_data_i[849] & v1_en_i;
  assign v1_data_o[848] = v0_data_i[848] & v1_en_i;
  assign v1_data_o[847] = v0_data_i[847] & v1_en_i;
  assign v1_data_o[846] = v0_data_i[846] & v1_en_i;
  assign v1_data_o[845] = v0_data_i[845] & v1_en_i;
  assign v1_data_o[844] = v0_data_i[844] & v1_en_i;
  assign v1_data_o[843] = v0_data_i[843] & v1_en_i;
  assign v1_data_o[842] = v0_data_i[842] & v1_en_i;
  assign v1_data_o[841] = v0_data_i[841] & v1_en_i;
  assign v1_data_o[840] = v0_data_i[840] & v1_en_i;
  assign v1_data_o[839] = v0_data_i[839] & v1_en_i;
  assign v1_data_o[838] = v0_data_i[838] & v1_en_i;
  assign v1_data_o[837] = v0_data_i[837] & v1_en_i;
  assign v1_data_o[836] = v0_data_i[836] & v1_en_i;
  assign v1_data_o[835] = v0_data_i[835] & v1_en_i;
  assign v1_data_o[834] = v0_data_i[834] & v1_en_i;
  assign v1_data_o[833] = v0_data_i[833] & v1_en_i;
  assign v1_data_o[832] = v0_data_i[832] & v1_en_i;
  assign v1_data_o[831] = v0_data_i[831] & v1_en_i;
  assign v1_data_o[830] = v0_data_i[830] & v1_en_i;
  assign v1_data_o[829] = v0_data_i[829] & v1_en_i;
  assign v1_data_o[828] = v0_data_i[828] & v1_en_i;
  assign v1_data_o[827] = v0_data_i[827] & v1_en_i;
  assign v1_data_o[826] = v0_data_i[826] & v1_en_i;
  assign v1_data_o[825] = v0_data_i[825] & v1_en_i;
  assign v1_data_o[824] = v0_data_i[824] & v1_en_i;
  assign v1_data_o[823] = v0_data_i[823] & v1_en_i;
  assign v1_data_o[822] = v0_data_i[822] & v1_en_i;
  assign v1_data_o[821] = v0_data_i[821] & v1_en_i;
  assign v1_data_o[820] = v0_data_i[820] & v1_en_i;
  assign v1_data_o[819] = v0_data_i[819] & v1_en_i;
  assign v1_data_o[818] = v0_data_i[818] & v1_en_i;
  assign v1_data_o[817] = v0_data_i[817] & v1_en_i;
  assign v1_data_o[816] = v0_data_i[816] & v1_en_i;
  assign v1_data_o[815] = v0_data_i[815] & v1_en_i;
  assign v1_data_o[814] = v0_data_i[814] & v1_en_i;
  assign v1_data_o[813] = v0_data_i[813] & v1_en_i;
  assign v1_data_o[812] = v0_data_i[812] & v1_en_i;
  assign v1_data_o[811] = v0_data_i[811] & v1_en_i;
  assign v1_data_o[810] = v0_data_i[810] & v1_en_i;
  assign v1_data_o[809] = v0_data_i[809] & v1_en_i;
  assign v1_data_o[808] = v0_data_i[808] & v1_en_i;
  assign v1_data_o[807] = v0_data_i[807] & v1_en_i;
  assign v1_data_o[806] = v0_data_i[806] & v1_en_i;
  assign v1_data_o[805] = v0_data_i[805] & v1_en_i;
  assign v1_data_o[804] = v0_data_i[804] & v1_en_i;
  assign v1_data_o[803] = v0_data_i[803] & v1_en_i;
  assign v1_data_o[802] = v0_data_i[802] & v1_en_i;
  assign v1_data_o[801] = v0_data_i[801] & v1_en_i;
  assign v1_data_o[800] = v0_data_i[800] & v1_en_i;
  assign v1_data_o[799] = v0_data_i[799] & v1_en_i;
  assign v1_data_o[798] = v0_data_i[798] & v1_en_i;
  assign v1_data_o[797] = v0_data_i[797] & v1_en_i;
  assign v1_data_o[796] = v0_data_i[796] & v1_en_i;
  assign v1_data_o[795] = v0_data_i[795] & v1_en_i;
  assign v1_data_o[794] = v0_data_i[794] & v1_en_i;
  assign v1_data_o[793] = v0_data_i[793] & v1_en_i;
  assign v1_data_o[792] = v0_data_i[792] & v1_en_i;
  assign v1_data_o[791] = v0_data_i[791] & v1_en_i;
  assign v1_data_o[790] = v0_data_i[790] & v1_en_i;
  assign v1_data_o[789] = v0_data_i[789] & v1_en_i;
  assign v1_data_o[788] = v0_data_i[788] & v1_en_i;
  assign v1_data_o[787] = v0_data_i[787] & v1_en_i;
  assign v1_data_o[786] = v0_data_i[786] & v1_en_i;
  assign v1_data_o[785] = v0_data_i[785] & v1_en_i;
  assign v1_data_o[784] = v0_data_i[784] & v1_en_i;
  assign v1_data_o[783] = v0_data_i[783] & v1_en_i;
  assign v1_data_o[782] = v0_data_i[782] & v1_en_i;
  assign v1_data_o[781] = v0_data_i[781] & v1_en_i;
  assign v1_data_o[780] = v0_data_i[780] & v1_en_i;
  assign v1_data_o[779] = v0_data_i[779] & v1_en_i;
  assign v1_data_o[778] = v0_data_i[778] & v1_en_i;
  assign v1_data_o[777] = v0_data_i[777] & v1_en_i;
  assign v1_data_o[776] = v0_data_i[776] & v1_en_i;
  assign v1_data_o[775] = v0_data_i[775] & v1_en_i;
  assign v1_data_o[774] = v0_data_i[774] & v1_en_i;
  assign v1_data_o[773] = v0_data_i[773] & v1_en_i;
  assign v1_data_o[772] = v0_data_i[772] & v1_en_i;
  assign v1_data_o[771] = v0_data_i[771] & v1_en_i;
  assign v1_data_o[770] = v0_data_i[770] & v1_en_i;
  assign v1_data_o[769] = v0_data_i[769] & v1_en_i;
  assign v1_data_o[768] = v0_data_i[768] & v1_en_i;
  assign v1_data_o[767] = v0_data_i[767] & v1_en_i;
  assign v1_data_o[766] = v0_data_i[766] & v1_en_i;
  assign v1_data_o[765] = v0_data_i[765] & v1_en_i;
  assign v1_data_o[764] = v0_data_i[764] & v1_en_i;
  assign v1_data_o[763] = v0_data_i[763] & v1_en_i;
  assign v1_data_o[762] = v0_data_i[762] & v1_en_i;
  assign v1_data_o[761] = v0_data_i[761] & v1_en_i;
  assign v1_data_o[760] = v0_data_i[760] & v1_en_i;
  assign v1_data_o[759] = v0_data_i[759] & v1_en_i;
  assign v1_data_o[758] = v0_data_i[758] & v1_en_i;
  assign v1_data_o[757] = v0_data_i[757] & v1_en_i;
  assign v1_data_o[756] = v0_data_i[756] & v1_en_i;
  assign v1_data_o[755] = v0_data_i[755] & v1_en_i;
  assign v1_data_o[754] = v0_data_i[754] & v1_en_i;
  assign v1_data_o[753] = v0_data_i[753] & v1_en_i;
  assign v1_data_o[752] = v0_data_i[752] & v1_en_i;
  assign v1_data_o[751] = v0_data_i[751] & v1_en_i;
  assign v1_data_o[750] = v0_data_i[750] & v1_en_i;
  assign v1_data_o[749] = v0_data_i[749] & v1_en_i;
  assign v1_data_o[748] = v0_data_i[748] & v1_en_i;
  assign v1_data_o[747] = v0_data_i[747] & v1_en_i;
  assign v1_data_o[746] = v0_data_i[746] & v1_en_i;
  assign v1_data_o[745] = v0_data_i[745] & v1_en_i;
  assign v1_data_o[744] = v0_data_i[744] & v1_en_i;
  assign v1_data_o[743] = v0_data_i[743] & v1_en_i;
  assign v1_data_o[742] = v0_data_i[742] & v1_en_i;
  assign v1_data_o[741] = v0_data_i[741] & v1_en_i;
  assign v1_data_o[740] = v0_data_i[740] & v1_en_i;
  assign v1_data_o[739] = v0_data_i[739] & v1_en_i;
  assign v1_data_o[738] = v0_data_i[738] & v1_en_i;
  assign v1_data_o[737] = v0_data_i[737] & v1_en_i;
  assign v1_data_o[736] = v0_data_i[736] & v1_en_i;
  assign v1_data_o[735] = v0_data_i[735] & v1_en_i;
  assign v1_data_o[734] = v0_data_i[734] & v1_en_i;
  assign v1_data_o[733] = v0_data_i[733] & v1_en_i;
  assign v1_data_o[732] = v0_data_i[732] & v1_en_i;
  assign v1_data_o[731] = v0_data_i[731] & v1_en_i;
  assign v1_data_o[730] = v0_data_i[730] & v1_en_i;
  assign v1_data_o[729] = v0_data_i[729] & v1_en_i;
  assign v1_data_o[728] = v0_data_i[728] & v1_en_i;
  assign v1_data_o[727] = v0_data_i[727] & v1_en_i;
  assign v1_data_o[726] = v0_data_i[726] & v1_en_i;
  assign v1_data_o[725] = v0_data_i[725] & v1_en_i;
  assign v1_data_o[724] = v0_data_i[724] & v1_en_i;
  assign v1_data_o[723] = v0_data_i[723] & v1_en_i;
  assign v1_data_o[722] = v0_data_i[722] & v1_en_i;
  assign v1_data_o[721] = v0_data_i[721] & v1_en_i;
  assign v1_data_o[720] = v0_data_i[720] & v1_en_i;
  assign v1_data_o[719] = v0_data_i[719] & v1_en_i;
  assign v1_data_o[718] = v0_data_i[718] & v1_en_i;
  assign v1_data_o[717] = v0_data_i[717] & v1_en_i;
  assign v1_data_o[716] = v0_data_i[716] & v1_en_i;
  assign v1_data_o[715] = v0_data_i[715] & v1_en_i;
  assign v1_data_o[714] = v0_data_i[714] & v1_en_i;
  assign v1_data_o[713] = v0_data_i[713] & v1_en_i;
  assign v1_data_o[712] = v0_data_i[712] & v1_en_i;
  assign v1_data_o[711] = v0_data_i[711] & v1_en_i;
  assign v1_data_o[710] = v0_data_i[710] & v1_en_i;
  assign v1_data_o[709] = v0_data_i[709] & v1_en_i;
  assign v1_data_o[708] = v0_data_i[708] & v1_en_i;
  assign v1_data_o[707] = v0_data_i[707] & v1_en_i;
  assign v1_data_o[706] = v0_data_i[706] & v1_en_i;
  assign v1_data_o[705] = v0_data_i[705] & v1_en_i;
  assign v1_data_o[704] = v0_data_i[704] & v1_en_i;
  assign v1_data_o[703] = v0_data_i[703] & v1_en_i;
  assign v1_data_o[702] = v0_data_i[702] & v1_en_i;
  assign v1_data_o[701] = v0_data_i[701] & v1_en_i;
  assign v1_data_o[700] = v0_data_i[700] & v1_en_i;
  assign v1_data_o[699] = v0_data_i[699] & v1_en_i;
  assign v1_data_o[698] = v0_data_i[698] & v1_en_i;
  assign v1_data_o[697] = v0_data_i[697] & v1_en_i;
  assign v1_data_o[696] = v0_data_i[696] & v1_en_i;
  assign v1_data_o[695] = v0_data_i[695] & v1_en_i;
  assign v1_data_o[694] = v0_data_i[694] & v1_en_i;
  assign v1_data_o[693] = v0_data_i[693] & v1_en_i;
  assign v1_data_o[692] = v0_data_i[692] & v1_en_i;
  assign v1_data_o[691] = v0_data_i[691] & v1_en_i;
  assign v1_data_o[690] = v0_data_i[690] & v1_en_i;
  assign v1_data_o[689] = v0_data_i[689] & v1_en_i;
  assign v1_data_o[688] = v0_data_i[688] & v1_en_i;
  assign v1_data_o[687] = v0_data_i[687] & v1_en_i;
  assign v1_data_o[686] = v0_data_i[686] & v1_en_i;
  assign v1_data_o[685] = v0_data_i[685] & v1_en_i;
  assign v1_data_o[684] = v0_data_i[684] & v1_en_i;
  assign v1_data_o[683] = v0_data_i[683] & v1_en_i;
  assign v1_data_o[682] = v0_data_i[682] & v1_en_i;
  assign v1_data_o[681] = v0_data_i[681] & v1_en_i;
  assign v1_data_o[680] = v0_data_i[680] & v1_en_i;
  assign v1_data_o[679] = v0_data_i[679] & v1_en_i;
  assign v1_data_o[678] = v0_data_i[678] & v1_en_i;
  assign v1_data_o[677] = v0_data_i[677] & v1_en_i;
  assign v1_data_o[676] = v0_data_i[676] & v1_en_i;
  assign v1_data_o[675] = v0_data_i[675] & v1_en_i;
  assign v1_data_o[674] = v0_data_i[674] & v1_en_i;
  assign v1_data_o[673] = v0_data_i[673] & v1_en_i;
  assign v1_data_o[672] = v0_data_i[672] & v1_en_i;
  assign v1_data_o[671] = v0_data_i[671] & v1_en_i;
  assign v1_data_o[670] = v0_data_i[670] & v1_en_i;
  assign v1_data_o[669] = v0_data_i[669] & v1_en_i;
  assign v1_data_o[668] = v0_data_i[668] & v1_en_i;
  assign v1_data_o[667] = v0_data_i[667] & v1_en_i;
  assign v1_data_o[666] = v0_data_i[666] & v1_en_i;
  assign v1_data_o[665] = v0_data_i[665] & v1_en_i;
  assign v1_data_o[664] = v0_data_i[664] & v1_en_i;
  assign v1_data_o[663] = v0_data_i[663] & v1_en_i;
  assign v1_data_o[662] = v0_data_i[662] & v1_en_i;
  assign v1_data_o[661] = v0_data_i[661] & v1_en_i;
  assign v1_data_o[660] = v0_data_i[660] & v1_en_i;
  assign v1_data_o[659] = v0_data_i[659] & v1_en_i;
  assign v1_data_o[658] = v0_data_i[658] & v1_en_i;
  assign v1_data_o[657] = v0_data_i[657] & v1_en_i;
  assign v1_data_o[656] = v0_data_i[656] & v1_en_i;
  assign v1_data_o[655] = v0_data_i[655] & v1_en_i;
  assign v1_data_o[654] = v0_data_i[654] & v1_en_i;
  assign v1_data_o[653] = v0_data_i[653] & v1_en_i;
  assign v1_data_o[652] = v0_data_i[652] & v1_en_i;
  assign v1_data_o[651] = v0_data_i[651] & v1_en_i;
  assign v1_data_o[650] = v0_data_i[650] & v1_en_i;
  assign v1_data_o[649] = v0_data_i[649] & v1_en_i;
  assign v1_data_o[648] = v0_data_i[648] & v1_en_i;
  assign v1_data_o[647] = v0_data_i[647] & v1_en_i;
  assign v1_data_o[646] = v0_data_i[646] & v1_en_i;
  assign v1_data_o[645] = v0_data_i[645] & v1_en_i;
  assign v1_data_o[644] = v0_data_i[644] & v1_en_i;
  assign v1_data_o[643] = v0_data_i[643] & v1_en_i;
  assign v1_data_o[642] = v0_data_i[642] & v1_en_i;
  assign v1_data_o[641] = v0_data_i[641] & v1_en_i;
  assign v1_data_o[640] = v0_data_i[640] & v1_en_i;
  assign v1_data_o[639] = v0_data_i[639] & v1_en_i;
  assign v1_data_o[638] = v0_data_i[638] & v1_en_i;
  assign v1_data_o[637] = v0_data_i[637] & v1_en_i;
  assign v1_data_o[636] = v0_data_i[636] & v1_en_i;
  assign v1_data_o[635] = v0_data_i[635] & v1_en_i;
  assign v1_data_o[634] = v0_data_i[634] & v1_en_i;
  assign v1_data_o[633] = v0_data_i[633] & v1_en_i;
  assign v1_data_o[632] = v0_data_i[632] & v1_en_i;
  assign v1_data_o[631] = v0_data_i[631] & v1_en_i;
  assign v1_data_o[630] = v0_data_i[630] & v1_en_i;
  assign v1_data_o[629] = v0_data_i[629] & v1_en_i;
  assign v1_data_o[628] = v0_data_i[628] & v1_en_i;
  assign v1_data_o[627] = v0_data_i[627] & v1_en_i;
  assign v1_data_o[626] = v0_data_i[626] & v1_en_i;
  assign v1_data_o[625] = v0_data_i[625] & v1_en_i;
  assign v1_data_o[624] = v0_data_i[624] & v1_en_i;
  assign v1_data_o[623] = v0_data_i[623] & v1_en_i;
  assign v1_data_o[622] = v0_data_i[622] & v1_en_i;
  assign v1_data_o[621] = v0_data_i[621] & v1_en_i;
  assign v1_data_o[620] = v0_data_i[620] & v1_en_i;
  assign v1_data_o[619] = v0_data_i[619] & v1_en_i;
  assign v1_data_o[618] = v0_data_i[618] & v1_en_i;
  assign v1_data_o[617] = v0_data_i[617] & v1_en_i;
  assign v1_data_o[616] = v0_data_i[616] & v1_en_i;
  assign v1_data_o[615] = v0_data_i[615] & v1_en_i;
  assign v1_data_o[614] = v0_data_i[614] & v1_en_i;
  assign v1_data_o[613] = v0_data_i[613] & v1_en_i;
  assign v1_data_o[612] = v0_data_i[612] & v1_en_i;
  assign v1_data_o[611] = v0_data_i[611] & v1_en_i;
  assign v1_data_o[610] = v0_data_i[610] & v1_en_i;
  assign v1_data_o[609] = v0_data_i[609] & v1_en_i;
  assign v1_data_o[608] = v0_data_i[608] & v1_en_i;
  assign v1_data_o[607] = v0_data_i[607] & v1_en_i;
  assign v1_data_o[606] = v0_data_i[606] & v1_en_i;
  assign v1_data_o[605] = v0_data_i[605] & v1_en_i;
  assign v1_data_o[604] = v0_data_i[604] & v1_en_i;
  assign v1_data_o[603] = v0_data_i[603] & v1_en_i;
  assign v1_data_o[602] = v0_data_i[602] & v1_en_i;
  assign v1_data_o[601] = v0_data_i[601] & v1_en_i;
  assign v1_data_o[600] = v0_data_i[600] & v1_en_i;
  assign v1_data_o[599] = v0_data_i[599] & v1_en_i;
  assign v1_data_o[598] = v0_data_i[598] & v1_en_i;
  assign v1_data_o[597] = v0_data_i[597] & v1_en_i;
  assign v1_data_o[596] = v0_data_i[596] & v1_en_i;
  assign v1_data_o[595] = v0_data_i[595] & v1_en_i;
  assign v1_data_o[594] = v0_data_i[594] & v1_en_i;
  assign v1_data_o[593] = v0_data_i[593] & v1_en_i;
  assign v1_data_o[592] = v0_data_i[592] & v1_en_i;
  assign v1_data_o[591] = v0_data_i[591] & v1_en_i;
  assign v1_data_o[590] = v0_data_i[590] & v1_en_i;
  assign v1_data_o[589] = v0_data_i[589] & v1_en_i;
  assign v1_data_o[588] = v0_data_i[588] & v1_en_i;
  assign v1_data_o[587] = v0_data_i[587] & v1_en_i;
  assign v1_data_o[586] = v0_data_i[586] & v1_en_i;
  assign v1_data_o[585] = v0_data_i[585] & v1_en_i;
  assign v1_data_o[584] = v0_data_i[584] & v1_en_i;
  assign v1_data_o[583] = v0_data_i[583] & v1_en_i;
  assign v1_data_o[582] = v0_data_i[582] & v1_en_i;
  assign v1_data_o[581] = v0_data_i[581] & v1_en_i;
  assign v1_data_o[580] = v0_data_i[580] & v1_en_i;
  assign v1_data_o[579] = v0_data_i[579] & v1_en_i;
  assign v1_data_o[578] = v0_data_i[578] & v1_en_i;
  assign v1_data_o[577] = v0_data_i[577] & v1_en_i;
  assign v1_data_o[576] = v0_data_i[576] & v1_en_i;
  assign v1_data_o[575] = v0_data_i[575] & v1_en_i;
  assign v1_data_o[574] = v0_data_i[574] & v1_en_i;
  assign v1_data_o[573] = v0_data_i[573] & v1_en_i;
  assign v1_data_o[572] = v0_data_i[572] & v1_en_i;
  assign v1_data_o[571] = v0_data_i[571] & v1_en_i;
  assign v1_data_o[570] = v0_data_i[570] & v1_en_i;
  assign v1_data_o[569] = v0_data_i[569] & v1_en_i;
  assign v1_data_o[568] = v0_data_i[568] & v1_en_i;
  assign v1_data_o[567] = v0_data_i[567] & v1_en_i;
  assign v1_data_o[566] = v0_data_i[566] & v1_en_i;
  assign v1_data_o[565] = v0_data_i[565] & v1_en_i;
  assign v1_data_o[564] = v0_data_i[564] & v1_en_i;
  assign v1_data_o[563] = v0_data_i[563] & v1_en_i;
  assign v1_data_o[562] = v0_data_i[562] & v1_en_i;
  assign v1_data_o[561] = v0_data_i[561] & v1_en_i;
  assign v1_data_o[560] = v0_data_i[560] & v1_en_i;
  assign v1_data_o[559] = v0_data_i[559] & v1_en_i;
  assign v1_data_o[558] = v0_data_i[558] & v1_en_i;
  assign v1_data_o[557] = v0_data_i[557] & v1_en_i;
  assign v1_data_o[556] = v0_data_i[556] & v1_en_i;
  assign v1_data_o[555] = v0_data_i[555] & v1_en_i;
  assign v1_data_o[554] = v0_data_i[554] & v1_en_i;
  assign v1_data_o[553] = v0_data_i[553] & v1_en_i;
  assign v1_data_o[552] = v0_data_i[552] & v1_en_i;
  assign v1_data_o[551] = v0_data_i[551] & v1_en_i;
  assign v1_data_o[550] = v0_data_i[550] & v1_en_i;
  assign v1_data_o[549] = v0_data_i[549] & v1_en_i;
  assign v1_data_o[548] = v0_data_i[548] & v1_en_i;
  assign v1_data_o[547] = v0_data_i[547] & v1_en_i;
  assign v1_data_o[546] = v0_data_i[546] & v1_en_i;
  assign v1_data_o[545] = v0_data_i[545] & v1_en_i;
  assign v1_data_o[544] = v0_data_i[544] & v1_en_i;
  assign v1_data_o[543] = v0_data_i[543] & v1_en_i;
  assign v1_data_o[542] = v0_data_i[542] & v1_en_i;
  assign v1_data_o[541] = v0_data_i[541] & v1_en_i;
  assign v1_data_o[540] = v0_data_i[540] & v1_en_i;
  assign v1_data_o[539] = v0_data_i[539] & v1_en_i;
  assign v1_data_o[538] = v0_data_i[538] & v1_en_i;
  assign v1_data_o[537] = v0_data_i[537] & v1_en_i;
  assign v1_data_o[536] = v0_data_i[536] & v1_en_i;
  assign v1_data_o[535] = v0_data_i[535] & v1_en_i;
  assign v1_data_o[534] = v0_data_i[534] & v1_en_i;
  assign v1_data_o[533] = v0_data_i[533] & v1_en_i;
  assign v1_data_o[532] = v0_data_i[532] & v1_en_i;
  assign v1_data_o[531] = v0_data_i[531] & v1_en_i;
  assign v1_data_o[530] = v0_data_i[530] & v1_en_i;
  assign v1_data_o[529] = v0_data_i[529] & v1_en_i;
  assign v1_data_o[528] = v0_data_i[528] & v1_en_i;
  assign v1_data_o[527] = v0_data_i[527] & v1_en_i;
  assign v1_data_o[526] = v0_data_i[526] & v1_en_i;
  assign v1_data_o[525] = v0_data_i[525] & v1_en_i;
  assign v1_data_o[524] = v0_data_i[524] & v1_en_i;
  assign v1_data_o[523] = v0_data_i[523] & v1_en_i;
  assign v1_data_o[522] = v0_data_i[522] & v1_en_i;
  assign v1_data_o[521] = v0_data_i[521] & v1_en_i;
  assign v1_data_o[520] = v0_data_i[520] & v1_en_i;
  assign v1_data_o[519] = v0_data_i[519] & v1_en_i;
  assign v1_data_o[518] = v0_data_i[518] & v1_en_i;
  assign v1_data_o[517] = v0_data_i[517] & v1_en_i;
  assign v1_data_o[516] = v0_data_i[516] & v1_en_i;
  assign v1_data_o[515] = v0_data_i[515] & v1_en_i;
  assign v1_data_o[514] = v0_data_i[514] & v1_en_i;
  assign v1_data_o[513] = v0_data_i[513] & v1_en_i;
  assign v1_data_o[512] = v0_data_i[512] & v1_en_i;
  assign v1_data_o[511] = v0_data_i[511] & v1_en_i;
  assign v1_data_o[510] = v0_data_i[510] & v1_en_i;
  assign v1_data_o[509] = v0_data_i[509] & v1_en_i;
  assign v1_data_o[508] = v0_data_i[508] & v1_en_i;
  assign v1_data_o[507] = v0_data_i[507] & v1_en_i;
  assign v1_data_o[506] = v0_data_i[506] & v1_en_i;
  assign v1_data_o[505] = v0_data_i[505] & v1_en_i;
  assign v1_data_o[504] = v0_data_i[504] & v1_en_i;
  assign v1_data_o[503] = v0_data_i[503] & v1_en_i;
  assign v1_data_o[502] = v0_data_i[502] & v1_en_i;
  assign v1_data_o[501] = v0_data_i[501] & v1_en_i;
  assign v1_data_o[500] = v0_data_i[500] & v1_en_i;
  assign v1_data_o[499] = v0_data_i[499] & v1_en_i;
  assign v1_data_o[498] = v0_data_i[498] & v1_en_i;
  assign v1_data_o[497] = v0_data_i[497] & v1_en_i;
  assign v1_data_o[496] = v0_data_i[496] & v1_en_i;
  assign v1_data_o[495] = v0_data_i[495] & v1_en_i;
  assign v1_data_o[494] = v0_data_i[494] & v1_en_i;
  assign v1_data_o[493] = v0_data_i[493] & v1_en_i;
  assign v1_data_o[492] = v0_data_i[492] & v1_en_i;
  assign v1_data_o[491] = v0_data_i[491] & v1_en_i;
  assign v1_data_o[490] = v0_data_i[490] & v1_en_i;
  assign v1_data_o[489] = v0_data_i[489] & v1_en_i;
  assign v1_data_o[488] = v0_data_i[488] & v1_en_i;
  assign v1_data_o[487] = v0_data_i[487] & v1_en_i;
  assign v1_data_o[486] = v0_data_i[486] & v1_en_i;
  assign v1_data_o[485] = v0_data_i[485] & v1_en_i;
  assign v1_data_o[484] = v0_data_i[484] & v1_en_i;
  assign v1_data_o[483] = v0_data_i[483] & v1_en_i;
  assign v1_data_o[482] = v0_data_i[482] & v1_en_i;
  assign v1_data_o[481] = v0_data_i[481] & v1_en_i;
  assign v1_data_o[480] = v0_data_i[480] & v1_en_i;
  assign v1_data_o[479] = v0_data_i[479] & v1_en_i;
  assign v1_data_o[478] = v0_data_i[478] & v1_en_i;
  assign v1_data_o[477] = v0_data_i[477] & v1_en_i;
  assign v1_data_o[476] = v0_data_i[476] & v1_en_i;
  assign v1_data_o[475] = v0_data_i[475] & v1_en_i;
  assign v1_data_o[474] = v0_data_i[474] & v1_en_i;
  assign v1_data_o[473] = v0_data_i[473] & v1_en_i;
  assign v1_data_o[472] = v0_data_i[472] & v1_en_i;
  assign v1_data_o[471] = v0_data_i[471] & v1_en_i;
  assign v1_data_o[470] = v0_data_i[470] & v1_en_i;
  assign v1_data_o[469] = v0_data_i[469] & v1_en_i;
  assign v1_data_o[468] = v0_data_i[468] & v1_en_i;
  assign v1_data_o[467] = v0_data_i[467] & v1_en_i;
  assign v1_data_o[466] = v0_data_i[466] & v1_en_i;
  assign v1_data_o[465] = v0_data_i[465] & v1_en_i;
  assign v1_data_o[464] = v0_data_i[464] & v1_en_i;
  assign v1_data_o[463] = v0_data_i[463] & v1_en_i;
  assign v1_data_o[462] = v0_data_i[462] & v1_en_i;
  assign v1_data_o[461] = v0_data_i[461] & v1_en_i;
  assign v1_data_o[460] = v0_data_i[460] & v1_en_i;
  assign v1_data_o[459] = v0_data_i[459] & v1_en_i;
  assign v1_data_o[458] = v0_data_i[458] & v1_en_i;
  assign v1_data_o[457] = v0_data_i[457] & v1_en_i;
  assign v1_data_o[456] = v0_data_i[456] & v1_en_i;
  assign v1_data_o[455] = v0_data_i[455] & v1_en_i;
  assign v1_data_o[454] = v0_data_i[454] & v1_en_i;
  assign v1_data_o[453] = v0_data_i[453] & v1_en_i;
  assign v1_data_o[452] = v0_data_i[452] & v1_en_i;
  assign v1_data_o[451] = v0_data_i[451] & v1_en_i;
  assign v1_data_o[450] = v0_data_i[450] & v1_en_i;
  assign v1_data_o[449] = v0_data_i[449] & v1_en_i;
  assign v1_data_o[448] = v0_data_i[448] & v1_en_i;
  assign v1_data_o[447] = v0_data_i[447] & v1_en_i;
  assign v1_data_o[446] = v0_data_i[446] & v1_en_i;
  assign v1_data_o[445] = v0_data_i[445] & v1_en_i;
  assign v1_data_o[444] = v0_data_i[444] & v1_en_i;
  assign v1_data_o[443] = v0_data_i[443] & v1_en_i;
  assign v1_data_o[442] = v0_data_i[442] & v1_en_i;
  assign v1_data_o[441] = v0_data_i[441] & v1_en_i;
  assign v1_data_o[440] = v0_data_i[440] & v1_en_i;
  assign v1_data_o[439] = v0_data_i[439] & v1_en_i;
  assign v1_data_o[438] = v0_data_i[438] & v1_en_i;
  assign v1_data_o[437] = v0_data_i[437] & v1_en_i;
  assign v1_data_o[436] = v0_data_i[436] & v1_en_i;
  assign v1_data_o[435] = v0_data_i[435] & v1_en_i;
  assign v1_data_o[434] = v0_data_i[434] & v1_en_i;
  assign v1_data_o[433] = v0_data_i[433] & v1_en_i;
  assign v1_data_o[432] = v0_data_i[432] & v1_en_i;
  assign v1_data_o[431] = v0_data_i[431] & v1_en_i;
  assign v1_data_o[430] = v0_data_i[430] & v1_en_i;
  assign v1_data_o[429] = v0_data_i[429] & v1_en_i;
  assign v1_data_o[428] = v0_data_i[428] & v1_en_i;
  assign v1_data_o[427] = v0_data_i[427] & v1_en_i;
  assign v1_data_o[426] = v0_data_i[426] & v1_en_i;
  assign v1_data_o[425] = v0_data_i[425] & v1_en_i;
  assign v1_data_o[424] = v0_data_i[424] & v1_en_i;
  assign v1_data_o[423] = v0_data_i[423] & v1_en_i;
  assign v1_data_o[422] = v0_data_i[422] & v1_en_i;
  assign v1_data_o[421] = v0_data_i[421] & v1_en_i;
  assign v1_data_o[420] = v0_data_i[420] & v1_en_i;
  assign v1_data_o[419] = v0_data_i[419] & v1_en_i;
  assign v1_data_o[418] = v0_data_i[418] & v1_en_i;
  assign v1_data_o[417] = v0_data_i[417] & v1_en_i;
  assign v1_data_o[416] = v0_data_i[416] & v1_en_i;
  assign v1_data_o[415] = v0_data_i[415] & v1_en_i;
  assign v1_data_o[414] = v0_data_i[414] & v1_en_i;
  assign v1_data_o[413] = v0_data_i[413] & v1_en_i;
  assign v1_data_o[412] = v0_data_i[412] & v1_en_i;
  assign v1_data_o[411] = v0_data_i[411] & v1_en_i;
  assign v1_data_o[410] = v0_data_i[410] & v1_en_i;
  assign v1_data_o[409] = v0_data_i[409] & v1_en_i;
  assign v1_data_o[408] = v0_data_i[408] & v1_en_i;
  assign v1_data_o[407] = v0_data_i[407] & v1_en_i;
  assign v1_data_o[406] = v0_data_i[406] & v1_en_i;
  assign v1_data_o[405] = v0_data_i[405] & v1_en_i;
  assign v1_data_o[404] = v0_data_i[404] & v1_en_i;
  assign v1_data_o[403] = v0_data_i[403] & v1_en_i;
  assign v1_data_o[402] = v0_data_i[402] & v1_en_i;
  assign v1_data_o[401] = v0_data_i[401] & v1_en_i;
  assign v1_data_o[400] = v0_data_i[400] & v1_en_i;
  assign v1_data_o[399] = v0_data_i[399] & v1_en_i;
  assign v1_data_o[398] = v0_data_i[398] & v1_en_i;
  assign v1_data_o[397] = v0_data_i[397] & v1_en_i;
  assign v1_data_o[396] = v0_data_i[396] & v1_en_i;
  assign v1_data_o[395] = v0_data_i[395] & v1_en_i;
  assign v1_data_o[394] = v0_data_i[394] & v1_en_i;
  assign v1_data_o[393] = v0_data_i[393] & v1_en_i;
  assign v1_data_o[392] = v0_data_i[392] & v1_en_i;
  assign v1_data_o[391] = v0_data_i[391] & v1_en_i;
  assign v1_data_o[390] = v0_data_i[390] & v1_en_i;
  assign v1_data_o[389] = v0_data_i[389] & v1_en_i;
  assign v1_data_o[388] = v0_data_i[388] & v1_en_i;
  assign v1_data_o[387] = v0_data_i[387] & v1_en_i;
  assign v1_data_o[386] = v0_data_i[386] & v1_en_i;
  assign v1_data_o[385] = v0_data_i[385] & v1_en_i;
  assign v1_data_o[384] = v0_data_i[384] & v1_en_i;
  assign v1_data_o[383] = v0_data_i[383] & v1_en_i;
  assign v1_data_o[382] = v0_data_i[382] & v1_en_i;
  assign v1_data_o[381] = v0_data_i[381] & v1_en_i;
  assign v1_data_o[380] = v0_data_i[380] & v1_en_i;
  assign v1_data_o[379] = v0_data_i[379] & v1_en_i;
  assign v1_data_o[378] = v0_data_i[378] & v1_en_i;
  assign v1_data_o[377] = v0_data_i[377] & v1_en_i;
  assign v1_data_o[376] = v0_data_i[376] & v1_en_i;
  assign v1_data_o[375] = v0_data_i[375] & v1_en_i;
  assign v1_data_o[374] = v0_data_i[374] & v1_en_i;
  assign v1_data_o[373] = v0_data_i[373] & v1_en_i;
  assign v1_data_o[372] = v0_data_i[372] & v1_en_i;
  assign v1_data_o[371] = v0_data_i[371] & v1_en_i;
  assign v1_data_o[370] = v0_data_i[370] & v1_en_i;
  assign v1_data_o[369] = v0_data_i[369] & v1_en_i;
  assign v1_data_o[368] = v0_data_i[368] & v1_en_i;
  assign v1_data_o[367] = v0_data_i[367] & v1_en_i;
  assign v1_data_o[366] = v0_data_i[366] & v1_en_i;
  assign v1_data_o[365] = v0_data_i[365] & v1_en_i;
  assign v1_data_o[364] = v0_data_i[364] & v1_en_i;
  assign v1_data_o[363] = v0_data_i[363] & v1_en_i;
  assign v1_data_o[362] = v0_data_i[362] & v1_en_i;
  assign v1_data_o[361] = v0_data_i[361] & v1_en_i;
  assign v1_data_o[360] = v0_data_i[360] & v1_en_i;
  assign v1_data_o[359] = v0_data_i[359] & v1_en_i;
  assign v1_data_o[358] = v0_data_i[358] & v1_en_i;
  assign v1_data_o[357] = v0_data_i[357] & v1_en_i;
  assign v1_data_o[356] = v0_data_i[356] & v1_en_i;
  assign v1_data_o[355] = v0_data_i[355] & v1_en_i;
  assign v1_data_o[354] = v0_data_i[354] & v1_en_i;
  assign v1_data_o[353] = v0_data_i[353] & v1_en_i;
  assign v1_data_o[352] = v0_data_i[352] & v1_en_i;
  assign v1_data_o[351] = v0_data_i[351] & v1_en_i;
  assign v1_data_o[350] = v0_data_i[350] & v1_en_i;
  assign v1_data_o[349] = v0_data_i[349] & v1_en_i;
  assign v1_data_o[348] = v0_data_i[348] & v1_en_i;
  assign v1_data_o[347] = v0_data_i[347] & v1_en_i;
  assign v1_data_o[346] = v0_data_i[346] & v1_en_i;
  assign v1_data_o[345] = v0_data_i[345] & v1_en_i;
  assign v1_data_o[344] = v0_data_i[344] & v1_en_i;
  assign v1_data_o[343] = v0_data_i[343] & v1_en_i;
  assign v1_data_o[342] = v0_data_i[342] & v1_en_i;
  assign v1_data_o[341] = v0_data_i[341] & v1_en_i;
  assign v1_data_o[340] = v0_data_i[340] & v1_en_i;
  assign v1_data_o[339] = v0_data_i[339] & v1_en_i;
  assign v1_data_o[338] = v0_data_i[338] & v1_en_i;
  assign v1_data_o[337] = v0_data_i[337] & v1_en_i;
  assign v1_data_o[336] = v0_data_i[336] & v1_en_i;
  assign v1_data_o[335] = v0_data_i[335] & v1_en_i;
  assign v1_data_o[334] = v0_data_i[334] & v1_en_i;
  assign v1_data_o[333] = v0_data_i[333] & v1_en_i;
  assign v1_data_o[332] = v0_data_i[332] & v1_en_i;
  assign v1_data_o[331] = v0_data_i[331] & v1_en_i;
  assign v1_data_o[330] = v0_data_i[330] & v1_en_i;
  assign v1_data_o[329] = v0_data_i[329] & v1_en_i;
  assign v1_data_o[328] = v0_data_i[328] & v1_en_i;
  assign v1_data_o[327] = v0_data_i[327] & v1_en_i;
  assign v1_data_o[326] = v0_data_i[326] & v1_en_i;
  assign v1_data_o[325] = v0_data_i[325] & v1_en_i;
  assign v1_data_o[324] = v0_data_i[324] & v1_en_i;
  assign v1_data_o[323] = v0_data_i[323] & v1_en_i;
  assign v1_data_o[322] = v0_data_i[322] & v1_en_i;
  assign v1_data_o[321] = v0_data_i[321] & v1_en_i;
  assign v1_data_o[320] = v0_data_i[320] & v1_en_i;
  assign v1_data_o[319] = v0_data_i[319] & v1_en_i;
  assign v1_data_o[318] = v0_data_i[318] & v1_en_i;
  assign v1_data_o[317] = v0_data_i[317] & v1_en_i;
  assign v1_data_o[316] = v0_data_i[316] & v1_en_i;
  assign v1_data_o[315] = v0_data_i[315] & v1_en_i;
  assign v1_data_o[314] = v0_data_i[314] & v1_en_i;
  assign v1_data_o[313] = v0_data_i[313] & v1_en_i;
  assign v1_data_o[312] = v0_data_i[312] & v1_en_i;
  assign v1_data_o[311] = v0_data_i[311] & v1_en_i;
  assign v1_data_o[310] = v0_data_i[310] & v1_en_i;
  assign v1_data_o[309] = v0_data_i[309] & v1_en_i;
  assign v1_data_o[308] = v0_data_i[308] & v1_en_i;
  assign v1_data_o[307] = v0_data_i[307] & v1_en_i;
  assign v1_data_o[306] = v0_data_i[306] & v1_en_i;
  assign v1_data_o[305] = v0_data_i[305] & v1_en_i;
  assign v1_data_o[304] = v0_data_i[304] & v1_en_i;
  assign v1_data_o[303] = v0_data_i[303] & v1_en_i;
  assign v1_data_o[302] = v0_data_i[302] & v1_en_i;
  assign v1_data_o[301] = v0_data_i[301] & v1_en_i;
  assign v1_data_o[300] = v0_data_i[300] & v1_en_i;
  assign v1_data_o[299] = v0_data_i[299] & v1_en_i;
  assign v1_data_o[298] = v0_data_i[298] & v1_en_i;
  assign v1_data_o[297] = v0_data_i[297] & v1_en_i;
  assign v1_data_o[296] = v0_data_i[296] & v1_en_i;
  assign v1_data_o[295] = v0_data_i[295] & v1_en_i;
  assign v1_data_o[294] = v0_data_i[294] & v1_en_i;
  assign v1_data_o[293] = v0_data_i[293] & v1_en_i;
  assign v1_data_o[292] = v0_data_i[292] & v1_en_i;
  assign v1_data_o[291] = v0_data_i[291] & v1_en_i;
  assign v1_data_o[290] = v0_data_i[290] & v1_en_i;
  assign v1_data_o[289] = v0_data_i[289] & v1_en_i;
  assign v1_data_o[288] = v0_data_i[288] & v1_en_i;
  assign v1_data_o[287] = v0_data_i[287] & v1_en_i;
  assign v1_data_o[286] = v0_data_i[286] & v1_en_i;
  assign v1_data_o[285] = v0_data_i[285] & v1_en_i;
  assign v1_data_o[284] = v0_data_i[284] & v1_en_i;
  assign v1_data_o[283] = v0_data_i[283] & v1_en_i;
  assign v1_data_o[282] = v0_data_i[282] & v1_en_i;
  assign v1_data_o[281] = v0_data_i[281] & v1_en_i;
  assign v1_data_o[280] = v0_data_i[280] & v1_en_i;
  assign v1_data_o[279] = v0_data_i[279] & v1_en_i;
  assign v1_data_o[278] = v0_data_i[278] & v1_en_i;
  assign v1_data_o[277] = v0_data_i[277] & v1_en_i;
  assign v1_data_o[276] = v0_data_i[276] & v1_en_i;
  assign v1_data_o[275] = v0_data_i[275] & v1_en_i;
  assign v1_data_o[274] = v0_data_i[274] & v1_en_i;
  assign v1_data_o[273] = v0_data_i[273] & v1_en_i;
  assign v1_data_o[272] = v0_data_i[272] & v1_en_i;
  assign v1_data_o[271] = v0_data_i[271] & v1_en_i;
  assign v1_data_o[270] = v0_data_i[270] & v1_en_i;
  assign v1_data_o[269] = v0_data_i[269] & v1_en_i;
  assign v1_data_o[268] = v0_data_i[268] & v1_en_i;
  assign v1_data_o[267] = v0_data_i[267] & v1_en_i;
  assign v1_data_o[266] = v0_data_i[266] & v1_en_i;
  assign v1_data_o[265] = v0_data_i[265] & v1_en_i;
  assign v1_data_o[264] = v0_data_i[264] & v1_en_i;
  assign v1_data_o[263] = v0_data_i[263] & v1_en_i;
  assign v1_data_o[262] = v0_data_i[262] & v1_en_i;
  assign v1_data_o[261] = v0_data_i[261] & v1_en_i;
  assign v1_data_o[260] = v0_data_i[260] & v1_en_i;
  assign v1_data_o[259] = v0_data_i[259] & v1_en_i;
  assign v1_data_o[258] = v0_data_i[258] & v1_en_i;
  assign v1_data_o[257] = v0_data_i[257] & v1_en_i;
  assign v1_data_o[256] = v0_data_i[256] & v1_en_i;
  assign v1_data_o[255] = v0_data_i[255] & v1_en_i;
  assign v1_data_o[254] = v0_data_i[254] & v1_en_i;
  assign v1_data_o[253] = v0_data_i[253] & v1_en_i;
  assign v1_data_o[252] = v0_data_i[252] & v1_en_i;
  assign v1_data_o[251] = v0_data_i[251] & v1_en_i;
  assign v1_data_o[250] = v0_data_i[250] & v1_en_i;
  assign v1_data_o[249] = v0_data_i[249] & v1_en_i;
  assign v1_data_o[248] = v0_data_i[248] & v1_en_i;
  assign v1_data_o[247] = v0_data_i[247] & v1_en_i;
  assign v1_data_o[246] = v0_data_i[246] & v1_en_i;
  assign v1_data_o[245] = v0_data_i[245] & v1_en_i;
  assign v1_data_o[244] = v0_data_i[244] & v1_en_i;
  assign v1_data_o[243] = v0_data_i[243] & v1_en_i;
  assign v1_data_o[242] = v0_data_i[242] & v1_en_i;
  assign v1_data_o[241] = v0_data_i[241] & v1_en_i;
  assign v1_data_o[240] = v0_data_i[240] & v1_en_i;
  assign v1_data_o[239] = v0_data_i[239] & v1_en_i;
  assign v1_data_o[238] = v0_data_i[238] & v1_en_i;
  assign v1_data_o[237] = v0_data_i[237] & v1_en_i;
  assign v1_data_o[236] = v0_data_i[236] & v1_en_i;
  assign v1_data_o[235] = v0_data_i[235] & v1_en_i;
  assign v1_data_o[234] = v0_data_i[234] & v1_en_i;
  assign v1_data_o[233] = v0_data_i[233] & v1_en_i;
  assign v1_data_o[232] = v0_data_i[232] & v1_en_i;
  assign v1_data_o[231] = v0_data_i[231] & v1_en_i;
  assign v1_data_o[230] = v0_data_i[230] & v1_en_i;
  assign v1_data_o[229] = v0_data_i[229] & v1_en_i;
  assign v1_data_o[228] = v0_data_i[228] & v1_en_i;
  assign v1_data_o[227] = v0_data_i[227] & v1_en_i;
  assign v1_data_o[226] = v0_data_i[226] & v1_en_i;
  assign v1_data_o[225] = v0_data_i[225] & v1_en_i;
  assign v1_data_o[224] = v0_data_i[224] & v1_en_i;
  assign v1_data_o[223] = v0_data_i[223] & v1_en_i;
  assign v1_data_o[222] = v0_data_i[222] & v1_en_i;
  assign v1_data_o[221] = v0_data_i[221] & v1_en_i;
  assign v1_data_o[220] = v0_data_i[220] & v1_en_i;
  assign v1_data_o[219] = v0_data_i[219] & v1_en_i;
  assign v1_data_o[218] = v0_data_i[218] & v1_en_i;
  assign v1_data_o[217] = v0_data_i[217] & v1_en_i;
  assign v1_data_o[216] = v0_data_i[216] & v1_en_i;
  assign v1_data_o[215] = v0_data_i[215] & v1_en_i;
  assign v1_data_o[214] = v0_data_i[214] & v1_en_i;
  assign v1_data_o[213] = v0_data_i[213] & v1_en_i;
  assign v1_data_o[212] = v0_data_i[212] & v1_en_i;
  assign v1_data_o[211] = v0_data_i[211] & v1_en_i;
  assign v1_data_o[210] = v0_data_i[210] & v1_en_i;
  assign v1_data_o[209] = v0_data_i[209] & v1_en_i;
  assign v1_data_o[208] = v0_data_i[208] & v1_en_i;
  assign v1_data_o[207] = v0_data_i[207] & v1_en_i;
  assign v1_data_o[206] = v0_data_i[206] & v1_en_i;
  assign v1_data_o[205] = v0_data_i[205] & v1_en_i;
  assign v1_data_o[204] = v0_data_i[204] & v1_en_i;
  assign v1_data_o[203] = v0_data_i[203] & v1_en_i;
  assign v1_data_o[202] = v0_data_i[202] & v1_en_i;
  assign v1_data_o[201] = v0_data_i[201] & v1_en_i;
  assign v1_data_o[200] = v0_data_i[200] & v1_en_i;
  assign v1_data_o[199] = v0_data_i[199] & v1_en_i;
  assign v1_data_o[198] = v0_data_i[198] & v1_en_i;
  assign v1_data_o[197] = v0_data_i[197] & v1_en_i;
  assign v1_data_o[196] = v0_data_i[196] & v1_en_i;
  assign v1_data_o[195] = v0_data_i[195] & v1_en_i;
  assign v1_data_o[194] = v0_data_i[194] & v1_en_i;
  assign v1_data_o[193] = v0_data_i[193] & v1_en_i;
  assign v1_data_o[192] = v0_data_i[192] & v1_en_i;
  assign v1_data_o[191] = v0_data_i[191] & v1_en_i;
  assign v1_data_o[190] = v0_data_i[190] & v1_en_i;
  assign v1_data_o[189] = v0_data_i[189] & v1_en_i;
  assign v1_data_o[188] = v0_data_i[188] & v1_en_i;
  assign v1_data_o[187] = v0_data_i[187] & v1_en_i;
  assign v1_data_o[186] = v0_data_i[186] & v1_en_i;
  assign v1_data_o[185] = v0_data_i[185] & v1_en_i;
  assign v1_data_o[184] = v0_data_i[184] & v1_en_i;
  assign v1_data_o[183] = v0_data_i[183] & v1_en_i;
  assign v1_data_o[182] = v0_data_i[182] & v1_en_i;
  assign v1_data_o[181] = v0_data_i[181] & v1_en_i;
  assign v1_data_o[180] = v0_data_i[180] & v1_en_i;
  assign v1_data_o[179] = v0_data_i[179] & v1_en_i;
  assign v1_data_o[178] = v0_data_i[178] & v1_en_i;
  assign v1_data_o[177] = v0_data_i[177] & v1_en_i;
  assign v1_data_o[176] = v0_data_i[176] & v1_en_i;
  assign v1_data_o[175] = v0_data_i[175] & v1_en_i;
  assign v1_data_o[174] = v0_data_i[174] & v1_en_i;
  assign v1_data_o[173] = v0_data_i[173] & v1_en_i;
  assign v1_data_o[172] = v0_data_i[172] & v1_en_i;
  assign v1_data_o[171] = v0_data_i[171] & v1_en_i;
  assign v1_data_o[170] = v0_data_i[170] & v1_en_i;
  assign v1_data_o[169] = v0_data_i[169] & v1_en_i;
  assign v1_data_o[168] = v0_data_i[168] & v1_en_i;
  assign v1_data_o[167] = v0_data_i[167] & v1_en_i;
  assign v1_data_o[166] = v0_data_i[166] & v1_en_i;
  assign v1_data_o[165] = v0_data_i[165] & v1_en_i;
  assign v1_data_o[164] = v0_data_i[164] & v1_en_i;
  assign v1_data_o[163] = v0_data_i[163] & v1_en_i;
  assign v1_data_o[162] = v0_data_i[162] & v1_en_i;
  assign v1_data_o[161] = v0_data_i[161] & v1_en_i;
  assign v1_data_o[160] = v0_data_i[160] & v1_en_i;
  assign v1_data_o[159] = v0_data_i[159] & v1_en_i;
  assign v1_data_o[158] = v0_data_i[158] & v1_en_i;
  assign v1_data_o[157] = v0_data_i[157] & v1_en_i;
  assign v1_data_o[156] = v0_data_i[156] & v1_en_i;
  assign v1_data_o[155] = v0_data_i[155] & v1_en_i;
  assign v1_data_o[154] = v0_data_i[154] & v1_en_i;
  assign v1_data_o[153] = v0_data_i[153] & v1_en_i;
  assign v1_data_o[152] = v0_data_i[152] & v1_en_i;
  assign v1_data_o[151] = v0_data_i[151] & v1_en_i;
  assign v1_data_o[150] = v0_data_i[150] & v1_en_i;
  assign v1_data_o[149] = v0_data_i[149] & v1_en_i;
  assign v1_data_o[148] = v0_data_i[148] & v1_en_i;
  assign v1_data_o[147] = v0_data_i[147] & v1_en_i;
  assign v1_data_o[146] = v0_data_i[146] & v1_en_i;
  assign v1_data_o[145] = v0_data_i[145] & v1_en_i;
  assign v1_data_o[144] = v0_data_i[144] & v1_en_i;
  assign v1_data_o[143] = v0_data_i[143] & v1_en_i;
  assign v1_data_o[142] = v0_data_i[142] & v1_en_i;
  assign v1_data_o[141] = v0_data_i[141] & v1_en_i;
  assign v1_data_o[140] = v0_data_i[140] & v1_en_i;
  assign v1_data_o[139] = v0_data_i[139] & v1_en_i;
  assign v1_data_o[138] = v0_data_i[138] & v1_en_i;
  assign v1_data_o[137] = v0_data_i[137] & v1_en_i;
  assign v1_data_o[136] = v0_data_i[136] & v1_en_i;
  assign v1_data_o[135] = v0_data_i[135] & v1_en_i;
  assign v1_data_o[134] = v0_data_i[134] & v1_en_i;
  assign v1_data_o[133] = v0_data_i[133] & v1_en_i;
  assign v1_data_o[132] = v0_data_i[132] & v1_en_i;
  assign v1_data_o[131] = v0_data_i[131] & v1_en_i;
  assign v1_data_o[130] = v0_data_i[130] & v1_en_i;
  assign v1_data_o[129] = v0_data_i[129] & v1_en_i;
  assign v1_data_o[128] = v0_data_i[128] & v1_en_i;
  assign v1_data_o[127] = v0_data_i[127] & v1_en_i;
  assign v1_data_o[126] = v0_data_i[126] & v1_en_i;
  assign v1_data_o[125] = v0_data_i[125] & v1_en_i;
  assign v1_data_o[124] = v0_data_i[124] & v1_en_i;
  assign v1_data_o[123] = v0_data_i[123] & v1_en_i;
  assign v1_data_o[122] = v0_data_i[122] & v1_en_i;
  assign v1_data_o[121] = v0_data_i[121] & v1_en_i;
  assign v1_data_o[120] = v0_data_i[120] & v1_en_i;
  assign v1_data_o[119] = v0_data_i[119] & v1_en_i;
  assign v1_data_o[118] = v0_data_i[118] & v1_en_i;
  assign v1_data_o[117] = v0_data_i[117] & v1_en_i;
  assign v1_data_o[116] = v0_data_i[116] & v1_en_i;
  assign v1_data_o[115] = v0_data_i[115] & v1_en_i;
  assign v1_data_o[114] = v0_data_i[114] & v1_en_i;
  assign v1_data_o[113] = v0_data_i[113] & v1_en_i;
  assign v1_data_o[112] = v0_data_i[112] & v1_en_i;
  assign v1_data_o[111] = v0_data_i[111] & v1_en_i;
  assign v1_data_o[110] = v0_data_i[110] & v1_en_i;
  assign v1_data_o[109] = v0_data_i[109] & v1_en_i;
  assign v1_data_o[108] = v0_data_i[108] & v1_en_i;
  assign v1_data_o[107] = v0_data_i[107] & v1_en_i;
  assign v1_data_o[106] = v0_data_i[106] & v1_en_i;
  assign v1_data_o[105] = v0_data_i[105] & v1_en_i;
  assign v1_data_o[104] = v0_data_i[104] & v1_en_i;
  assign v1_data_o[103] = v0_data_i[103] & v1_en_i;
  assign v1_data_o[102] = v0_data_i[102] & v1_en_i;
  assign v1_data_o[101] = v0_data_i[101] & v1_en_i;
  assign v1_data_o[100] = v0_data_i[100] & v1_en_i;
  assign v1_data_o[99] = v0_data_i[99] & v1_en_i;
  assign v1_data_o[98] = v0_data_i[98] & v1_en_i;
  assign v1_data_o[97] = v0_data_i[97] & v1_en_i;
  assign v1_data_o[96] = v0_data_i[96] & v1_en_i;
  assign v1_data_o[95] = v0_data_i[95] & v1_en_i;
  assign v1_data_o[94] = v0_data_i[94] & v1_en_i;
  assign v1_data_o[93] = v0_data_i[93] & v1_en_i;
  assign v1_data_o[92] = v0_data_i[92] & v1_en_i;
  assign v1_data_o[91] = v0_data_i[91] & v1_en_i;
  assign v1_data_o[90] = v0_data_i[90] & v1_en_i;
  assign v1_data_o[89] = v0_data_i[89] & v1_en_i;
  assign v1_data_o[88] = v0_data_i[88] & v1_en_i;
  assign v1_data_o[87] = v0_data_i[87] & v1_en_i;
  assign v1_data_o[86] = v0_data_i[86] & v1_en_i;
  assign v1_data_o[85] = v0_data_i[85] & v1_en_i;
  assign v1_data_o[84] = v0_data_i[84] & v1_en_i;
  assign v1_data_o[83] = v0_data_i[83] & v1_en_i;
  assign v1_data_o[82] = v0_data_i[82] & v1_en_i;
  assign v1_data_o[81] = v0_data_i[81] & v1_en_i;
  assign v1_data_o[80] = v0_data_i[80] & v1_en_i;
  assign v1_data_o[79] = v0_data_i[79] & v1_en_i;
  assign v1_data_o[78] = v0_data_i[78] & v1_en_i;
  assign v1_data_o[77] = v0_data_i[77] & v1_en_i;
  assign v1_data_o[76] = v0_data_i[76] & v1_en_i;
  assign v1_data_o[75] = v0_data_i[75] & v1_en_i;
  assign v1_data_o[74] = v0_data_i[74] & v1_en_i;
  assign v1_data_o[73] = v0_data_i[73] & v1_en_i;
  assign v1_data_o[72] = v0_data_i[72] & v1_en_i;
  assign v1_data_o[71] = v0_data_i[71] & v1_en_i;
  assign v1_data_o[70] = v0_data_i[70] & v1_en_i;
  assign v1_data_o[69] = v0_data_i[69] & v1_en_i;
  assign v1_data_o[68] = v0_data_i[68] & v1_en_i;
  assign v1_data_o[67] = v0_data_i[67] & v1_en_i;
  assign v1_data_o[66] = v0_data_i[66] & v1_en_i;
  assign v1_data_o[65] = v0_data_i[65] & v1_en_i;
  assign v1_data_o[64] = v0_data_i[64] & v1_en_i;
  assign v1_data_o[63] = v0_data_i[63] & v1_en_i;
  assign v1_data_o[62] = v0_data_i[62] & v1_en_i;
  assign v1_data_o[61] = v0_data_i[61] & v1_en_i;
  assign v1_data_o[60] = v0_data_i[60] & v1_en_i;
  assign v1_data_o[59] = v0_data_i[59] & v1_en_i;
  assign v1_data_o[58] = v0_data_i[58] & v1_en_i;
  assign v1_data_o[57] = v0_data_i[57] & v1_en_i;
  assign v1_data_o[56] = v0_data_i[56] & v1_en_i;
  assign v1_data_o[55] = v0_data_i[55] & v1_en_i;
  assign v1_data_o[54] = v0_data_i[54] & v1_en_i;
  assign v1_data_o[53] = v0_data_i[53] & v1_en_i;
  assign v1_data_o[52] = v0_data_i[52] & v1_en_i;
  assign v1_data_o[51] = v0_data_i[51] & v1_en_i;
  assign v1_data_o[50] = v0_data_i[50] & v1_en_i;
  assign v1_data_o[49] = v0_data_i[49] & v1_en_i;
  assign v1_data_o[48] = v0_data_i[48] & v1_en_i;
  assign v1_data_o[47] = v0_data_i[47] & v1_en_i;
  assign v1_data_o[46] = v0_data_i[46] & v1_en_i;
  assign v1_data_o[45] = v0_data_i[45] & v1_en_i;
  assign v1_data_o[44] = v0_data_i[44] & v1_en_i;
  assign v1_data_o[43] = v0_data_i[43] & v1_en_i;
  assign v1_data_o[42] = v0_data_i[42] & v1_en_i;
  assign v1_data_o[41] = v0_data_i[41] & v1_en_i;
  assign v1_data_o[40] = v0_data_i[40] & v1_en_i;
  assign v1_data_o[39] = v0_data_i[39] & v1_en_i;
  assign v1_data_o[38] = v0_data_i[38] & v1_en_i;
  assign v1_data_o[37] = v0_data_i[37] & v1_en_i;
  assign v1_data_o[36] = v0_data_i[36] & v1_en_i;
  assign v1_data_o[35] = v0_data_i[35] & v1_en_i;
  assign v1_data_o[34] = v0_data_i[34] & v1_en_i;
  assign v1_data_o[33] = v0_data_i[33] & v1_en_i;
  assign v1_data_o[32] = v0_data_i[32] & v1_en_i;
  assign v1_data_o[31] = v0_data_i[31] & v1_en_i;
  assign v1_data_o[30] = v0_data_i[30] & v1_en_i;
  assign v1_data_o[29] = v0_data_i[29] & v1_en_i;
  assign v1_data_o[28] = v0_data_i[28] & v1_en_i;
  assign v1_data_o[27] = v0_data_i[27] & v1_en_i;
  assign v1_data_o[26] = v0_data_i[26] & v1_en_i;
  assign v1_data_o[25] = v0_data_i[25] & v1_en_i;
  assign v1_data_o[24] = v0_data_i[24] & v1_en_i;
  assign v1_data_o[23] = v0_data_i[23] & v1_en_i;
  assign v1_data_o[22] = v0_data_i[22] & v1_en_i;
  assign v1_data_o[21] = v0_data_i[21] & v1_en_i;
  assign v1_data_o[20] = v0_data_i[20] & v1_en_i;
  assign v1_data_o[19] = v0_data_i[19] & v1_en_i;
  assign v1_data_o[18] = v0_data_i[18] & v1_en_i;
  assign v1_data_o[17] = v0_data_i[17] & v1_en_i;
  assign v1_data_o[16] = v0_data_i[16] & v1_en_i;
  assign v1_data_o[15] = v0_data_i[15] & v1_en_i;
  assign v1_data_o[14] = v0_data_i[14] & v1_en_i;
  assign v1_data_o[13] = v0_data_i[13] & v1_en_i;
  assign v1_data_o[12] = v0_data_i[12] & v1_en_i;
  assign v1_data_o[11] = v0_data_i[11] & v1_en_i;
  assign v1_data_o[10] = v0_data_i[10] & v1_en_i;
  assign v1_data_o[9] = v0_data_i[9] & v1_en_i;
  assign v1_data_o[8] = v0_data_i[8] & v1_en_i;
  assign v1_data_o[7] = v0_data_i[7] & v1_en_i;
  assign v1_data_o[6] = v0_data_i[6] & v1_en_i;
  assign v1_data_o[5] = v0_data_i[5] & v1_en_i;
  assign v1_data_o[4] = v0_data_i[4] & v1_en_i;
  assign v1_data_o[3] = v0_data_i[3] & v1_en_i;
  assign v1_data_o[2] = v0_data_i[2] & v1_en_i;
  assign v1_data_o[1] = v0_data_i[1] & v1_en_i;
  assign v1_data_o[0] = v0_data_i[0] & v1_en_i;

endmodule



module bsg_level_shift_up_down_source_width_p1000
(
  v0_en_i,
  v0_data_i,
  v1_data_o
);

  input [999:0] v0_data_i;
  output [999:0] v1_data_o;
  input v0_en_i;
  wire [999:0] v1_data_o;
  assign v1_data_o[999] = v0_data_i[999] & v0_en_i;
  assign v1_data_o[998] = v0_data_i[998] & v0_en_i;
  assign v1_data_o[997] = v0_data_i[997] & v0_en_i;
  assign v1_data_o[996] = v0_data_i[996] & v0_en_i;
  assign v1_data_o[995] = v0_data_i[995] & v0_en_i;
  assign v1_data_o[994] = v0_data_i[994] & v0_en_i;
  assign v1_data_o[993] = v0_data_i[993] & v0_en_i;
  assign v1_data_o[992] = v0_data_i[992] & v0_en_i;
  assign v1_data_o[991] = v0_data_i[991] & v0_en_i;
  assign v1_data_o[990] = v0_data_i[990] & v0_en_i;
  assign v1_data_o[989] = v0_data_i[989] & v0_en_i;
  assign v1_data_o[988] = v0_data_i[988] & v0_en_i;
  assign v1_data_o[987] = v0_data_i[987] & v0_en_i;
  assign v1_data_o[986] = v0_data_i[986] & v0_en_i;
  assign v1_data_o[985] = v0_data_i[985] & v0_en_i;
  assign v1_data_o[984] = v0_data_i[984] & v0_en_i;
  assign v1_data_o[983] = v0_data_i[983] & v0_en_i;
  assign v1_data_o[982] = v0_data_i[982] & v0_en_i;
  assign v1_data_o[981] = v0_data_i[981] & v0_en_i;
  assign v1_data_o[980] = v0_data_i[980] & v0_en_i;
  assign v1_data_o[979] = v0_data_i[979] & v0_en_i;
  assign v1_data_o[978] = v0_data_i[978] & v0_en_i;
  assign v1_data_o[977] = v0_data_i[977] & v0_en_i;
  assign v1_data_o[976] = v0_data_i[976] & v0_en_i;
  assign v1_data_o[975] = v0_data_i[975] & v0_en_i;
  assign v1_data_o[974] = v0_data_i[974] & v0_en_i;
  assign v1_data_o[973] = v0_data_i[973] & v0_en_i;
  assign v1_data_o[972] = v0_data_i[972] & v0_en_i;
  assign v1_data_o[971] = v0_data_i[971] & v0_en_i;
  assign v1_data_o[970] = v0_data_i[970] & v0_en_i;
  assign v1_data_o[969] = v0_data_i[969] & v0_en_i;
  assign v1_data_o[968] = v0_data_i[968] & v0_en_i;
  assign v1_data_o[967] = v0_data_i[967] & v0_en_i;
  assign v1_data_o[966] = v0_data_i[966] & v0_en_i;
  assign v1_data_o[965] = v0_data_i[965] & v0_en_i;
  assign v1_data_o[964] = v0_data_i[964] & v0_en_i;
  assign v1_data_o[963] = v0_data_i[963] & v0_en_i;
  assign v1_data_o[962] = v0_data_i[962] & v0_en_i;
  assign v1_data_o[961] = v0_data_i[961] & v0_en_i;
  assign v1_data_o[960] = v0_data_i[960] & v0_en_i;
  assign v1_data_o[959] = v0_data_i[959] & v0_en_i;
  assign v1_data_o[958] = v0_data_i[958] & v0_en_i;
  assign v1_data_o[957] = v0_data_i[957] & v0_en_i;
  assign v1_data_o[956] = v0_data_i[956] & v0_en_i;
  assign v1_data_o[955] = v0_data_i[955] & v0_en_i;
  assign v1_data_o[954] = v0_data_i[954] & v0_en_i;
  assign v1_data_o[953] = v0_data_i[953] & v0_en_i;
  assign v1_data_o[952] = v0_data_i[952] & v0_en_i;
  assign v1_data_o[951] = v0_data_i[951] & v0_en_i;
  assign v1_data_o[950] = v0_data_i[950] & v0_en_i;
  assign v1_data_o[949] = v0_data_i[949] & v0_en_i;
  assign v1_data_o[948] = v0_data_i[948] & v0_en_i;
  assign v1_data_o[947] = v0_data_i[947] & v0_en_i;
  assign v1_data_o[946] = v0_data_i[946] & v0_en_i;
  assign v1_data_o[945] = v0_data_i[945] & v0_en_i;
  assign v1_data_o[944] = v0_data_i[944] & v0_en_i;
  assign v1_data_o[943] = v0_data_i[943] & v0_en_i;
  assign v1_data_o[942] = v0_data_i[942] & v0_en_i;
  assign v1_data_o[941] = v0_data_i[941] & v0_en_i;
  assign v1_data_o[940] = v0_data_i[940] & v0_en_i;
  assign v1_data_o[939] = v0_data_i[939] & v0_en_i;
  assign v1_data_o[938] = v0_data_i[938] & v0_en_i;
  assign v1_data_o[937] = v0_data_i[937] & v0_en_i;
  assign v1_data_o[936] = v0_data_i[936] & v0_en_i;
  assign v1_data_o[935] = v0_data_i[935] & v0_en_i;
  assign v1_data_o[934] = v0_data_i[934] & v0_en_i;
  assign v1_data_o[933] = v0_data_i[933] & v0_en_i;
  assign v1_data_o[932] = v0_data_i[932] & v0_en_i;
  assign v1_data_o[931] = v0_data_i[931] & v0_en_i;
  assign v1_data_o[930] = v0_data_i[930] & v0_en_i;
  assign v1_data_o[929] = v0_data_i[929] & v0_en_i;
  assign v1_data_o[928] = v0_data_i[928] & v0_en_i;
  assign v1_data_o[927] = v0_data_i[927] & v0_en_i;
  assign v1_data_o[926] = v0_data_i[926] & v0_en_i;
  assign v1_data_o[925] = v0_data_i[925] & v0_en_i;
  assign v1_data_o[924] = v0_data_i[924] & v0_en_i;
  assign v1_data_o[923] = v0_data_i[923] & v0_en_i;
  assign v1_data_o[922] = v0_data_i[922] & v0_en_i;
  assign v1_data_o[921] = v0_data_i[921] & v0_en_i;
  assign v1_data_o[920] = v0_data_i[920] & v0_en_i;
  assign v1_data_o[919] = v0_data_i[919] & v0_en_i;
  assign v1_data_o[918] = v0_data_i[918] & v0_en_i;
  assign v1_data_o[917] = v0_data_i[917] & v0_en_i;
  assign v1_data_o[916] = v0_data_i[916] & v0_en_i;
  assign v1_data_o[915] = v0_data_i[915] & v0_en_i;
  assign v1_data_o[914] = v0_data_i[914] & v0_en_i;
  assign v1_data_o[913] = v0_data_i[913] & v0_en_i;
  assign v1_data_o[912] = v0_data_i[912] & v0_en_i;
  assign v1_data_o[911] = v0_data_i[911] & v0_en_i;
  assign v1_data_o[910] = v0_data_i[910] & v0_en_i;
  assign v1_data_o[909] = v0_data_i[909] & v0_en_i;
  assign v1_data_o[908] = v0_data_i[908] & v0_en_i;
  assign v1_data_o[907] = v0_data_i[907] & v0_en_i;
  assign v1_data_o[906] = v0_data_i[906] & v0_en_i;
  assign v1_data_o[905] = v0_data_i[905] & v0_en_i;
  assign v1_data_o[904] = v0_data_i[904] & v0_en_i;
  assign v1_data_o[903] = v0_data_i[903] & v0_en_i;
  assign v1_data_o[902] = v0_data_i[902] & v0_en_i;
  assign v1_data_o[901] = v0_data_i[901] & v0_en_i;
  assign v1_data_o[900] = v0_data_i[900] & v0_en_i;
  assign v1_data_o[899] = v0_data_i[899] & v0_en_i;
  assign v1_data_o[898] = v0_data_i[898] & v0_en_i;
  assign v1_data_o[897] = v0_data_i[897] & v0_en_i;
  assign v1_data_o[896] = v0_data_i[896] & v0_en_i;
  assign v1_data_o[895] = v0_data_i[895] & v0_en_i;
  assign v1_data_o[894] = v0_data_i[894] & v0_en_i;
  assign v1_data_o[893] = v0_data_i[893] & v0_en_i;
  assign v1_data_o[892] = v0_data_i[892] & v0_en_i;
  assign v1_data_o[891] = v0_data_i[891] & v0_en_i;
  assign v1_data_o[890] = v0_data_i[890] & v0_en_i;
  assign v1_data_o[889] = v0_data_i[889] & v0_en_i;
  assign v1_data_o[888] = v0_data_i[888] & v0_en_i;
  assign v1_data_o[887] = v0_data_i[887] & v0_en_i;
  assign v1_data_o[886] = v0_data_i[886] & v0_en_i;
  assign v1_data_o[885] = v0_data_i[885] & v0_en_i;
  assign v1_data_o[884] = v0_data_i[884] & v0_en_i;
  assign v1_data_o[883] = v0_data_i[883] & v0_en_i;
  assign v1_data_o[882] = v0_data_i[882] & v0_en_i;
  assign v1_data_o[881] = v0_data_i[881] & v0_en_i;
  assign v1_data_o[880] = v0_data_i[880] & v0_en_i;
  assign v1_data_o[879] = v0_data_i[879] & v0_en_i;
  assign v1_data_o[878] = v0_data_i[878] & v0_en_i;
  assign v1_data_o[877] = v0_data_i[877] & v0_en_i;
  assign v1_data_o[876] = v0_data_i[876] & v0_en_i;
  assign v1_data_o[875] = v0_data_i[875] & v0_en_i;
  assign v1_data_o[874] = v0_data_i[874] & v0_en_i;
  assign v1_data_o[873] = v0_data_i[873] & v0_en_i;
  assign v1_data_o[872] = v0_data_i[872] & v0_en_i;
  assign v1_data_o[871] = v0_data_i[871] & v0_en_i;
  assign v1_data_o[870] = v0_data_i[870] & v0_en_i;
  assign v1_data_o[869] = v0_data_i[869] & v0_en_i;
  assign v1_data_o[868] = v0_data_i[868] & v0_en_i;
  assign v1_data_o[867] = v0_data_i[867] & v0_en_i;
  assign v1_data_o[866] = v0_data_i[866] & v0_en_i;
  assign v1_data_o[865] = v0_data_i[865] & v0_en_i;
  assign v1_data_o[864] = v0_data_i[864] & v0_en_i;
  assign v1_data_o[863] = v0_data_i[863] & v0_en_i;
  assign v1_data_o[862] = v0_data_i[862] & v0_en_i;
  assign v1_data_o[861] = v0_data_i[861] & v0_en_i;
  assign v1_data_o[860] = v0_data_i[860] & v0_en_i;
  assign v1_data_o[859] = v0_data_i[859] & v0_en_i;
  assign v1_data_o[858] = v0_data_i[858] & v0_en_i;
  assign v1_data_o[857] = v0_data_i[857] & v0_en_i;
  assign v1_data_o[856] = v0_data_i[856] & v0_en_i;
  assign v1_data_o[855] = v0_data_i[855] & v0_en_i;
  assign v1_data_o[854] = v0_data_i[854] & v0_en_i;
  assign v1_data_o[853] = v0_data_i[853] & v0_en_i;
  assign v1_data_o[852] = v0_data_i[852] & v0_en_i;
  assign v1_data_o[851] = v0_data_i[851] & v0_en_i;
  assign v1_data_o[850] = v0_data_i[850] & v0_en_i;
  assign v1_data_o[849] = v0_data_i[849] & v0_en_i;
  assign v1_data_o[848] = v0_data_i[848] & v0_en_i;
  assign v1_data_o[847] = v0_data_i[847] & v0_en_i;
  assign v1_data_o[846] = v0_data_i[846] & v0_en_i;
  assign v1_data_o[845] = v0_data_i[845] & v0_en_i;
  assign v1_data_o[844] = v0_data_i[844] & v0_en_i;
  assign v1_data_o[843] = v0_data_i[843] & v0_en_i;
  assign v1_data_o[842] = v0_data_i[842] & v0_en_i;
  assign v1_data_o[841] = v0_data_i[841] & v0_en_i;
  assign v1_data_o[840] = v0_data_i[840] & v0_en_i;
  assign v1_data_o[839] = v0_data_i[839] & v0_en_i;
  assign v1_data_o[838] = v0_data_i[838] & v0_en_i;
  assign v1_data_o[837] = v0_data_i[837] & v0_en_i;
  assign v1_data_o[836] = v0_data_i[836] & v0_en_i;
  assign v1_data_o[835] = v0_data_i[835] & v0_en_i;
  assign v1_data_o[834] = v0_data_i[834] & v0_en_i;
  assign v1_data_o[833] = v0_data_i[833] & v0_en_i;
  assign v1_data_o[832] = v0_data_i[832] & v0_en_i;
  assign v1_data_o[831] = v0_data_i[831] & v0_en_i;
  assign v1_data_o[830] = v0_data_i[830] & v0_en_i;
  assign v1_data_o[829] = v0_data_i[829] & v0_en_i;
  assign v1_data_o[828] = v0_data_i[828] & v0_en_i;
  assign v1_data_o[827] = v0_data_i[827] & v0_en_i;
  assign v1_data_o[826] = v0_data_i[826] & v0_en_i;
  assign v1_data_o[825] = v0_data_i[825] & v0_en_i;
  assign v1_data_o[824] = v0_data_i[824] & v0_en_i;
  assign v1_data_o[823] = v0_data_i[823] & v0_en_i;
  assign v1_data_o[822] = v0_data_i[822] & v0_en_i;
  assign v1_data_o[821] = v0_data_i[821] & v0_en_i;
  assign v1_data_o[820] = v0_data_i[820] & v0_en_i;
  assign v1_data_o[819] = v0_data_i[819] & v0_en_i;
  assign v1_data_o[818] = v0_data_i[818] & v0_en_i;
  assign v1_data_o[817] = v0_data_i[817] & v0_en_i;
  assign v1_data_o[816] = v0_data_i[816] & v0_en_i;
  assign v1_data_o[815] = v0_data_i[815] & v0_en_i;
  assign v1_data_o[814] = v0_data_i[814] & v0_en_i;
  assign v1_data_o[813] = v0_data_i[813] & v0_en_i;
  assign v1_data_o[812] = v0_data_i[812] & v0_en_i;
  assign v1_data_o[811] = v0_data_i[811] & v0_en_i;
  assign v1_data_o[810] = v0_data_i[810] & v0_en_i;
  assign v1_data_o[809] = v0_data_i[809] & v0_en_i;
  assign v1_data_o[808] = v0_data_i[808] & v0_en_i;
  assign v1_data_o[807] = v0_data_i[807] & v0_en_i;
  assign v1_data_o[806] = v0_data_i[806] & v0_en_i;
  assign v1_data_o[805] = v0_data_i[805] & v0_en_i;
  assign v1_data_o[804] = v0_data_i[804] & v0_en_i;
  assign v1_data_o[803] = v0_data_i[803] & v0_en_i;
  assign v1_data_o[802] = v0_data_i[802] & v0_en_i;
  assign v1_data_o[801] = v0_data_i[801] & v0_en_i;
  assign v1_data_o[800] = v0_data_i[800] & v0_en_i;
  assign v1_data_o[799] = v0_data_i[799] & v0_en_i;
  assign v1_data_o[798] = v0_data_i[798] & v0_en_i;
  assign v1_data_o[797] = v0_data_i[797] & v0_en_i;
  assign v1_data_o[796] = v0_data_i[796] & v0_en_i;
  assign v1_data_o[795] = v0_data_i[795] & v0_en_i;
  assign v1_data_o[794] = v0_data_i[794] & v0_en_i;
  assign v1_data_o[793] = v0_data_i[793] & v0_en_i;
  assign v1_data_o[792] = v0_data_i[792] & v0_en_i;
  assign v1_data_o[791] = v0_data_i[791] & v0_en_i;
  assign v1_data_o[790] = v0_data_i[790] & v0_en_i;
  assign v1_data_o[789] = v0_data_i[789] & v0_en_i;
  assign v1_data_o[788] = v0_data_i[788] & v0_en_i;
  assign v1_data_o[787] = v0_data_i[787] & v0_en_i;
  assign v1_data_o[786] = v0_data_i[786] & v0_en_i;
  assign v1_data_o[785] = v0_data_i[785] & v0_en_i;
  assign v1_data_o[784] = v0_data_i[784] & v0_en_i;
  assign v1_data_o[783] = v0_data_i[783] & v0_en_i;
  assign v1_data_o[782] = v0_data_i[782] & v0_en_i;
  assign v1_data_o[781] = v0_data_i[781] & v0_en_i;
  assign v1_data_o[780] = v0_data_i[780] & v0_en_i;
  assign v1_data_o[779] = v0_data_i[779] & v0_en_i;
  assign v1_data_o[778] = v0_data_i[778] & v0_en_i;
  assign v1_data_o[777] = v0_data_i[777] & v0_en_i;
  assign v1_data_o[776] = v0_data_i[776] & v0_en_i;
  assign v1_data_o[775] = v0_data_i[775] & v0_en_i;
  assign v1_data_o[774] = v0_data_i[774] & v0_en_i;
  assign v1_data_o[773] = v0_data_i[773] & v0_en_i;
  assign v1_data_o[772] = v0_data_i[772] & v0_en_i;
  assign v1_data_o[771] = v0_data_i[771] & v0_en_i;
  assign v1_data_o[770] = v0_data_i[770] & v0_en_i;
  assign v1_data_o[769] = v0_data_i[769] & v0_en_i;
  assign v1_data_o[768] = v0_data_i[768] & v0_en_i;
  assign v1_data_o[767] = v0_data_i[767] & v0_en_i;
  assign v1_data_o[766] = v0_data_i[766] & v0_en_i;
  assign v1_data_o[765] = v0_data_i[765] & v0_en_i;
  assign v1_data_o[764] = v0_data_i[764] & v0_en_i;
  assign v1_data_o[763] = v0_data_i[763] & v0_en_i;
  assign v1_data_o[762] = v0_data_i[762] & v0_en_i;
  assign v1_data_o[761] = v0_data_i[761] & v0_en_i;
  assign v1_data_o[760] = v0_data_i[760] & v0_en_i;
  assign v1_data_o[759] = v0_data_i[759] & v0_en_i;
  assign v1_data_o[758] = v0_data_i[758] & v0_en_i;
  assign v1_data_o[757] = v0_data_i[757] & v0_en_i;
  assign v1_data_o[756] = v0_data_i[756] & v0_en_i;
  assign v1_data_o[755] = v0_data_i[755] & v0_en_i;
  assign v1_data_o[754] = v0_data_i[754] & v0_en_i;
  assign v1_data_o[753] = v0_data_i[753] & v0_en_i;
  assign v1_data_o[752] = v0_data_i[752] & v0_en_i;
  assign v1_data_o[751] = v0_data_i[751] & v0_en_i;
  assign v1_data_o[750] = v0_data_i[750] & v0_en_i;
  assign v1_data_o[749] = v0_data_i[749] & v0_en_i;
  assign v1_data_o[748] = v0_data_i[748] & v0_en_i;
  assign v1_data_o[747] = v0_data_i[747] & v0_en_i;
  assign v1_data_o[746] = v0_data_i[746] & v0_en_i;
  assign v1_data_o[745] = v0_data_i[745] & v0_en_i;
  assign v1_data_o[744] = v0_data_i[744] & v0_en_i;
  assign v1_data_o[743] = v0_data_i[743] & v0_en_i;
  assign v1_data_o[742] = v0_data_i[742] & v0_en_i;
  assign v1_data_o[741] = v0_data_i[741] & v0_en_i;
  assign v1_data_o[740] = v0_data_i[740] & v0_en_i;
  assign v1_data_o[739] = v0_data_i[739] & v0_en_i;
  assign v1_data_o[738] = v0_data_i[738] & v0_en_i;
  assign v1_data_o[737] = v0_data_i[737] & v0_en_i;
  assign v1_data_o[736] = v0_data_i[736] & v0_en_i;
  assign v1_data_o[735] = v0_data_i[735] & v0_en_i;
  assign v1_data_o[734] = v0_data_i[734] & v0_en_i;
  assign v1_data_o[733] = v0_data_i[733] & v0_en_i;
  assign v1_data_o[732] = v0_data_i[732] & v0_en_i;
  assign v1_data_o[731] = v0_data_i[731] & v0_en_i;
  assign v1_data_o[730] = v0_data_i[730] & v0_en_i;
  assign v1_data_o[729] = v0_data_i[729] & v0_en_i;
  assign v1_data_o[728] = v0_data_i[728] & v0_en_i;
  assign v1_data_o[727] = v0_data_i[727] & v0_en_i;
  assign v1_data_o[726] = v0_data_i[726] & v0_en_i;
  assign v1_data_o[725] = v0_data_i[725] & v0_en_i;
  assign v1_data_o[724] = v0_data_i[724] & v0_en_i;
  assign v1_data_o[723] = v0_data_i[723] & v0_en_i;
  assign v1_data_o[722] = v0_data_i[722] & v0_en_i;
  assign v1_data_o[721] = v0_data_i[721] & v0_en_i;
  assign v1_data_o[720] = v0_data_i[720] & v0_en_i;
  assign v1_data_o[719] = v0_data_i[719] & v0_en_i;
  assign v1_data_o[718] = v0_data_i[718] & v0_en_i;
  assign v1_data_o[717] = v0_data_i[717] & v0_en_i;
  assign v1_data_o[716] = v0_data_i[716] & v0_en_i;
  assign v1_data_o[715] = v0_data_i[715] & v0_en_i;
  assign v1_data_o[714] = v0_data_i[714] & v0_en_i;
  assign v1_data_o[713] = v0_data_i[713] & v0_en_i;
  assign v1_data_o[712] = v0_data_i[712] & v0_en_i;
  assign v1_data_o[711] = v0_data_i[711] & v0_en_i;
  assign v1_data_o[710] = v0_data_i[710] & v0_en_i;
  assign v1_data_o[709] = v0_data_i[709] & v0_en_i;
  assign v1_data_o[708] = v0_data_i[708] & v0_en_i;
  assign v1_data_o[707] = v0_data_i[707] & v0_en_i;
  assign v1_data_o[706] = v0_data_i[706] & v0_en_i;
  assign v1_data_o[705] = v0_data_i[705] & v0_en_i;
  assign v1_data_o[704] = v0_data_i[704] & v0_en_i;
  assign v1_data_o[703] = v0_data_i[703] & v0_en_i;
  assign v1_data_o[702] = v0_data_i[702] & v0_en_i;
  assign v1_data_o[701] = v0_data_i[701] & v0_en_i;
  assign v1_data_o[700] = v0_data_i[700] & v0_en_i;
  assign v1_data_o[699] = v0_data_i[699] & v0_en_i;
  assign v1_data_o[698] = v0_data_i[698] & v0_en_i;
  assign v1_data_o[697] = v0_data_i[697] & v0_en_i;
  assign v1_data_o[696] = v0_data_i[696] & v0_en_i;
  assign v1_data_o[695] = v0_data_i[695] & v0_en_i;
  assign v1_data_o[694] = v0_data_i[694] & v0_en_i;
  assign v1_data_o[693] = v0_data_i[693] & v0_en_i;
  assign v1_data_o[692] = v0_data_i[692] & v0_en_i;
  assign v1_data_o[691] = v0_data_i[691] & v0_en_i;
  assign v1_data_o[690] = v0_data_i[690] & v0_en_i;
  assign v1_data_o[689] = v0_data_i[689] & v0_en_i;
  assign v1_data_o[688] = v0_data_i[688] & v0_en_i;
  assign v1_data_o[687] = v0_data_i[687] & v0_en_i;
  assign v1_data_o[686] = v0_data_i[686] & v0_en_i;
  assign v1_data_o[685] = v0_data_i[685] & v0_en_i;
  assign v1_data_o[684] = v0_data_i[684] & v0_en_i;
  assign v1_data_o[683] = v0_data_i[683] & v0_en_i;
  assign v1_data_o[682] = v0_data_i[682] & v0_en_i;
  assign v1_data_o[681] = v0_data_i[681] & v0_en_i;
  assign v1_data_o[680] = v0_data_i[680] & v0_en_i;
  assign v1_data_o[679] = v0_data_i[679] & v0_en_i;
  assign v1_data_o[678] = v0_data_i[678] & v0_en_i;
  assign v1_data_o[677] = v0_data_i[677] & v0_en_i;
  assign v1_data_o[676] = v0_data_i[676] & v0_en_i;
  assign v1_data_o[675] = v0_data_i[675] & v0_en_i;
  assign v1_data_o[674] = v0_data_i[674] & v0_en_i;
  assign v1_data_o[673] = v0_data_i[673] & v0_en_i;
  assign v1_data_o[672] = v0_data_i[672] & v0_en_i;
  assign v1_data_o[671] = v0_data_i[671] & v0_en_i;
  assign v1_data_o[670] = v0_data_i[670] & v0_en_i;
  assign v1_data_o[669] = v0_data_i[669] & v0_en_i;
  assign v1_data_o[668] = v0_data_i[668] & v0_en_i;
  assign v1_data_o[667] = v0_data_i[667] & v0_en_i;
  assign v1_data_o[666] = v0_data_i[666] & v0_en_i;
  assign v1_data_o[665] = v0_data_i[665] & v0_en_i;
  assign v1_data_o[664] = v0_data_i[664] & v0_en_i;
  assign v1_data_o[663] = v0_data_i[663] & v0_en_i;
  assign v1_data_o[662] = v0_data_i[662] & v0_en_i;
  assign v1_data_o[661] = v0_data_i[661] & v0_en_i;
  assign v1_data_o[660] = v0_data_i[660] & v0_en_i;
  assign v1_data_o[659] = v0_data_i[659] & v0_en_i;
  assign v1_data_o[658] = v0_data_i[658] & v0_en_i;
  assign v1_data_o[657] = v0_data_i[657] & v0_en_i;
  assign v1_data_o[656] = v0_data_i[656] & v0_en_i;
  assign v1_data_o[655] = v0_data_i[655] & v0_en_i;
  assign v1_data_o[654] = v0_data_i[654] & v0_en_i;
  assign v1_data_o[653] = v0_data_i[653] & v0_en_i;
  assign v1_data_o[652] = v0_data_i[652] & v0_en_i;
  assign v1_data_o[651] = v0_data_i[651] & v0_en_i;
  assign v1_data_o[650] = v0_data_i[650] & v0_en_i;
  assign v1_data_o[649] = v0_data_i[649] & v0_en_i;
  assign v1_data_o[648] = v0_data_i[648] & v0_en_i;
  assign v1_data_o[647] = v0_data_i[647] & v0_en_i;
  assign v1_data_o[646] = v0_data_i[646] & v0_en_i;
  assign v1_data_o[645] = v0_data_i[645] & v0_en_i;
  assign v1_data_o[644] = v0_data_i[644] & v0_en_i;
  assign v1_data_o[643] = v0_data_i[643] & v0_en_i;
  assign v1_data_o[642] = v0_data_i[642] & v0_en_i;
  assign v1_data_o[641] = v0_data_i[641] & v0_en_i;
  assign v1_data_o[640] = v0_data_i[640] & v0_en_i;
  assign v1_data_o[639] = v0_data_i[639] & v0_en_i;
  assign v1_data_o[638] = v0_data_i[638] & v0_en_i;
  assign v1_data_o[637] = v0_data_i[637] & v0_en_i;
  assign v1_data_o[636] = v0_data_i[636] & v0_en_i;
  assign v1_data_o[635] = v0_data_i[635] & v0_en_i;
  assign v1_data_o[634] = v0_data_i[634] & v0_en_i;
  assign v1_data_o[633] = v0_data_i[633] & v0_en_i;
  assign v1_data_o[632] = v0_data_i[632] & v0_en_i;
  assign v1_data_o[631] = v0_data_i[631] & v0_en_i;
  assign v1_data_o[630] = v0_data_i[630] & v0_en_i;
  assign v1_data_o[629] = v0_data_i[629] & v0_en_i;
  assign v1_data_o[628] = v0_data_i[628] & v0_en_i;
  assign v1_data_o[627] = v0_data_i[627] & v0_en_i;
  assign v1_data_o[626] = v0_data_i[626] & v0_en_i;
  assign v1_data_o[625] = v0_data_i[625] & v0_en_i;
  assign v1_data_o[624] = v0_data_i[624] & v0_en_i;
  assign v1_data_o[623] = v0_data_i[623] & v0_en_i;
  assign v1_data_o[622] = v0_data_i[622] & v0_en_i;
  assign v1_data_o[621] = v0_data_i[621] & v0_en_i;
  assign v1_data_o[620] = v0_data_i[620] & v0_en_i;
  assign v1_data_o[619] = v0_data_i[619] & v0_en_i;
  assign v1_data_o[618] = v0_data_i[618] & v0_en_i;
  assign v1_data_o[617] = v0_data_i[617] & v0_en_i;
  assign v1_data_o[616] = v0_data_i[616] & v0_en_i;
  assign v1_data_o[615] = v0_data_i[615] & v0_en_i;
  assign v1_data_o[614] = v0_data_i[614] & v0_en_i;
  assign v1_data_o[613] = v0_data_i[613] & v0_en_i;
  assign v1_data_o[612] = v0_data_i[612] & v0_en_i;
  assign v1_data_o[611] = v0_data_i[611] & v0_en_i;
  assign v1_data_o[610] = v0_data_i[610] & v0_en_i;
  assign v1_data_o[609] = v0_data_i[609] & v0_en_i;
  assign v1_data_o[608] = v0_data_i[608] & v0_en_i;
  assign v1_data_o[607] = v0_data_i[607] & v0_en_i;
  assign v1_data_o[606] = v0_data_i[606] & v0_en_i;
  assign v1_data_o[605] = v0_data_i[605] & v0_en_i;
  assign v1_data_o[604] = v0_data_i[604] & v0_en_i;
  assign v1_data_o[603] = v0_data_i[603] & v0_en_i;
  assign v1_data_o[602] = v0_data_i[602] & v0_en_i;
  assign v1_data_o[601] = v0_data_i[601] & v0_en_i;
  assign v1_data_o[600] = v0_data_i[600] & v0_en_i;
  assign v1_data_o[599] = v0_data_i[599] & v0_en_i;
  assign v1_data_o[598] = v0_data_i[598] & v0_en_i;
  assign v1_data_o[597] = v0_data_i[597] & v0_en_i;
  assign v1_data_o[596] = v0_data_i[596] & v0_en_i;
  assign v1_data_o[595] = v0_data_i[595] & v0_en_i;
  assign v1_data_o[594] = v0_data_i[594] & v0_en_i;
  assign v1_data_o[593] = v0_data_i[593] & v0_en_i;
  assign v1_data_o[592] = v0_data_i[592] & v0_en_i;
  assign v1_data_o[591] = v0_data_i[591] & v0_en_i;
  assign v1_data_o[590] = v0_data_i[590] & v0_en_i;
  assign v1_data_o[589] = v0_data_i[589] & v0_en_i;
  assign v1_data_o[588] = v0_data_i[588] & v0_en_i;
  assign v1_data_o[587] = v0_data_i[587] & v0_en_i;
  assign v1_data_o[586] = v0_data_i[586] & v0_en_i;
  assign v1_data_o[585] = v0_data_i[585] & v0_en_i;
  assign v1_data_o[584] = v0_data_i[584] & v0_en_i;
  assign v1_data_o[583] = v0_data_i[583] & v0_en_i;
  assign v1_data_o[582] = v0_data_i[582] & v0_en_i;
  assign v1_data_o[581] = v0_data_i[581] & v0_en_i;
  assign v1_data_o[580] = v0_data_i[580] & v0_en_i;
  assign v1_data_o[579] = v0_data_i[579] & v0_en_i;
  assign v1_data_o[578] = v0_data_i[578] & v0_en_i;
  assign v1_data_o[577] = v0_data_i[577] & v0_en_i;
  assign v1_data_o[576] = v0_data_i[576] & v0_en_i;
  assign v1_data_o[575] = v0_data_i[575] & v0_en_i;
  assign v1_data_o[574] = v0_data_i[574] & v0_en_i;
  assign v1_data_o[573] = v0_data_i[573] & v0_en_i;
  assign v1_data_o[572] = v0_data_i[572] & v0_en_i;
  assign v1_data_o[571] = v0_data_i[571] & v0_en_i;
  assign v1_data_o[570] = v0_data_i[570] & v0_en_i;
  assign v1_data_o[569] = v0_data_i[569] & v0_en_i;
  assign v1_data_o[568] = v0_data_i[568] & v0_en_i;
  assign v1_data_o[567] = v0_data_i[567] & v0_en_i;
  assign v1_data_o[566] = v0_data_i[566] & v0_en_i;
  assign v1_data_o[565] = v0_data_i[565] & v0_en_i;
  assign v1_data_o[564] = v0_data_i[564] & v0_en_i;
  assign v1_data_o[563] = v0_data_i[563] & v0_en_i;
  assign v1_data_o[562] = v0_data_i[562] & v0_en_i;
  assign v1_data_o[561] = v0_data_i[561] & v0_en_i;
  assign v1_data_o[560] = v0_data_i[560] & v0_en_i;
  assign v1_data_o[559] = v0_data_i[559] & v0_en_i;
  assign v1_data_o[558] = v0_data_i[558] & v0_en_i;
  assign v1_data_o[557] = v0_data_i[557] & v0_en_i;
  assign v1_data_o[556] = v0_data_i[556] & v0_en_i;
  assign v1_data_o[555] = v0_data_i[555] & v0_en_i;
  assign v1_data_o[554] = v0_data_i[554] & v0_en_i;
  assign v1_data_o[553] = v0_data_i[553] & v0_en_i;
  assign v1_data_o[552] = v0_data_i[552] & v0_en_i;
  assign v1_data_o[551] = v0_data_i[551] & v0_en_i;
  assign v1_data_o[550] = v0_data_i[550] & v0_en_i;
  assign v1_data_o[549] = v0_data_i[549] & v0_en_i;
  assign v1_data_o[548] = v0_data_i[548] & v0_en_i;
  assign v1_data_o[547] = v0_data_i[547] & v0_en_i;
  assign v1_data_o[546] = v0_data_i[546] & v0_en_i;
  assign v1_data_o[545] = v0_data_i[545] & v0_en_i;
  assign v1_data_o[544] = v0_data_i[544] & v0_en_i;
  assign v1_data_o[543] = v0_data_i[543] & v0_en_i;
  assign v1_data_o[542] = v0_data_i[542] & v0_en_i;
  assign v1_data_o[541] = v0_data_i[541] & v0_en_i;
  assign v1_data_o[540] = v0_data_i[540] & v0_en_i;
  assign v1_data_o[539] = v0_data_i[539] & v0_en_i;
  assign v1_data_o[538] = v0_data_i[538] & v0_en_i;
  assign v1_data_o[537] = v0_data_i[537] & v0_en_i;
  assign v1_data_o[536] = v0_data_i[536] & v0_en_i;
  assign v1_data_o[535] = v0_data_i[535] & v0_en_i;
  assign v1_data_o[534] = v0_data_i[534] & v0_en_i;
  assign v1_data_o[533] = v0_data_i[533] & v0_en_i;
  assign v1_data_o[532] = v0_data_i[532] & v0_en_i;
  assign v1_data_o[531] = v0_data_i[531] & v0_en_i;
  assign v1_data_o[530] = v0_data_i[530] & v0_en_i;
  assign v1_data_o[529] = v0_data_i[529] & v0_en_i;
  assign v1_data_o[528] = v0_data_i[528] & v0_en_i;
  assign v1_data_o[527] = v0_data_i[527] & v0_en_i;
  assign v1_data_o[526] = v0_data_i[526] & v0_en_i;
  assign v1_data_o[525] = v0_data_i[525] & v0_en_i;
  assign v1_data_o[524] = v0_data_i[524] & v0_en_i;
  assign v1_data_o[523] = v0_data_i[523] & v0_en_i;
  assign v1_data_o[522] = v0_data_i[522] & v0_en_i;
  assign v1_data_o[521] = v0_data_i[521] & v0_en_i;
  assign v1_data_o[520] = v0_data_i[520] & v0_en_i;
  assign v1_data_o[519] = v0_data_i[519] & v0_en_i;
  assign v1_data_o[518] = v0_data_i[518] & v0_en_i;
  assign v1_data_o[517] = v0_data_i[517] & v0_en_i;
  assign v1_data_o[516] = v0_data_i[516] & v0_en_i;
  assign v1_data_o[515] = v0_data_i[515] & v0_en_i;
  assign v1_data_o[514] = v0_data_i[514] & v0_en_i;
  assign v1_data_o[513] = v0_data_i[513] & v0_en_i;
  assign v1_data_o[512] = v0_data_i[512] & v0_en_i;
  assign v1_data_o[511] = v0_data_i[511] & v0_en_i;
  assign v1_data_o[510] = v0_data_i[510] & v0_en_i;
  assign v1_data_o[509] = v0_data_i[509] & v0_en_i;
  assign v1_data_o[508] = v0_data_i[508] & v0_en_i;
  assign v1_data_o[507] = v0_data_i[507] & v0_en_i;
  assign v1_data_o[506] = v0_data_i[506] & v0_en_i;
  assign v1_data_o[505] = v0_data_i[505] & v0_en_i;
  assign v1_data_o[504] = v0_data_i[504] & v0_en_i;
  assign v1_data_o[503] = v0_data_i[503] & v0_en_i;
  assign v1_data_o[502] = v0_data_i[502] & v0_en_i;
  assign v1_data_o[501] = v0_data_i[501] & v0_en_i;
  assign v1_data_o[500] = v0_data_i[500] & v0_en_i;
  assign v1_data_o[499] = v0_data_i[499] & v0_en_i;
  assign v1_data_o[498] = v0_data_i[498] & v0_en_i;
  assign v1_data_o[497] = v0_data_i[497] & v0_en_i;
  assign v1_data_o[496] = v0_data_i[496] & v0_en_i;
  assign v1_data_o[495] = v0_data_i[495] & v0_en_i;
  assign v1_data_o[494] = v0_data_i[494] & v0_en_i;
  assign v1_data_o[493] = v0_data_i[493] & v0_en_i;
  assign v1_data_o[492] = v0_data_i[492] & v0_en_i;
  assign v1_data_o[491] = v0_data_i[491] & v0_en_i;
  assign v1_data_o[490] = v0_data_i[490] & v0_en_i;
  assign v1_data_o[489] = v0_data_i[489] & v0_en_i;
  assign v1_data_o[488] = v0_data_i[488] & v0_en_i;
  assign v1_data_o[487] = v0_data_i[487] & v0_en_i;
  assign v1_data_o[486] = v0_data_i[486] & v0_en_i;
  assign v1_data_o[485] = v0_data_i[485] & v0_en_i;
  assign v1_data_o[484] = v0_data_i[484] & v0_en_i;
  assign v1_data_o[483] = v0_data_i[483] & v0_en_i;
  assign v1_data_o[482] = v0_data_i[482] & v0_en_i;
  assign v1_data_o[481] = v0_data_i[481] & v0_en_i;
  assign v1_data_o[480] = v0_data_i[480] & v0_en_i;
  assign v1_data_o[479] = v0_data_i[479] & v0_en_i;
  assign v1_data_o[478] = v0_data_i[478] & v0_en_i;
  assign v1_data_o[477] = v0_data_i[477] & v0_en_i;
  assign v1_data_o[476] = v0_data_i[476] & v0_en_i;
  assign v1_data_o[475] = v0_data_i[475] & v0_en_i;
  assign v1_data_o[474] = v0_data_i[474] & v0_en_i;
  assign v1_data_o[473] = v0_data_i[473] & v0_en_i;
  assign v1_data_o[472] = v0_data_i[472] & v0_en_i;
  assign v1_data_o[471] = v0_data_i[471] & v0_en_i;
  assign v1_data_o[470] = v0_data_i[470] & v0_en_i;
  assign v1_data_o[469] = v0_data_i[469] & v0_en_i;
  assign v1_data_o[468] = v0_data_i[468] & v0_en_i;
  assign v1_data_o[467] = v0_data_i[467] & v0_en_i;
  assign v1_data_o[466] = v0_data_i[466] & v0_en_i;
  assign v1_data_o[465] = v0_data_i[465] & v0_en_i;
  assign v1_data_o[464] = v0_data_i[464] & v0_en_i;
  assign v1_data_o[463] = v0_data_i[463] & v0_en_i;
  assign v1_data_o[462] = v0_data_i[462] & v0_en_i;
  assign v1_data_o[461] = v0_data_i[461] & v0_en_i;
  assign v1_data_o[460] = v0_data_i[460] & v0_en_i;
  assign v1_data_o[459] = v0_data_i[459] & v0_en_i;
  assign v1_data_o[458] = v0_data_i[458] & v0_en_i;
  assign v1_data_o[457] = v0_data_i[457] & v0_en_i;
  assign v1_data_o[456] = v0_data_i[456] & v0_en_i;
  assign v1_data_o[455] = v0_data_i[455] & v0_en_i;
  assign v1_data_o[454] = v0_data_i[454] & v0_en_i;
  assign v1_data_o[453] = v0_data_i[453] & v0_en_i;
  assign v1_data_o[452] = v0_data_i[452] & v0_en_i;
  assign v1_data_o[451] = v0_data_i[451] & v0_en_i;
  assign v1_data_o[450] = v0_data_i[450] & v0_en_i;
  assign v1_data_o[449] = v0_data_i[449] & v0_en_i;
  assign v1_data_o[448] = v0_data_i[448] & v0_en_i;
  assign v1_data_o[447] = v0_data_i[447] & v0_en_i;
  assign v1_data_o[446] = v0_data_i[446] & v0_en_i;
  assign v1_data_o[445] = v0_data_i[445] & v0_en_i;
  assign v1_data_o[444] = v0_data_i[444] & v0_en_i;
  assign v1_data_o[443] = v0_data_i[443] & v0_en_i;
  assign v1_data_o[442] = v0_data_i[442] & v0_en_i;
  assign v1_data_o[441] = v0_data_i[441] & v0_en_i;
  assign v1_data_o[440] = v0_data_i[440] & v0_en_i;
  assign v1_data_o[439] = v0_data_i[439] & v0_en_i;
  assign v1_data_o[438] = v0_data_i[438] & v0_en_i;
  assign v1_data_o[437] = v0_data_i[437] & v0_en_i;
  assign v1_data_o[436] = v0_data_i[436] & v0_en_i;
  assign v1_data_o[435] = v0_data_i[435] & v0_en_i;
  assign v1_data_o[434] = v0_data_i[434] & v0_en_i;
  assign v1_data_o[433] = v0_data_i[433] & v0_en_i;
  assign v1_data_o[432] = v0_data_i[432] & v0_en_i;
  assign v1_data_o[431] = v0_data_i[431] & v0_en_i;
  assign v1_data_o[430] = v0_data_i[430] & v0_en_i;
  assign v1_data_o[429] = v0_data_i[429] & v0_en_i;
  assign v1_data_o[428] = v0_data_i[428] & v0_en_i;
  assign v1_data_o[427] = v0_data_i[427] & v0_en_i;
  assign v1_data_o[426] = v0_data_i[426] & v0_en_i;
  assign v1_data_o[425] = v0_data_i[425] & v0_en_i;
  assign v1_data_o[424] = v0_data_i[424] & v0_en_i;
  assign v1_data_o[423] = v0_data_i[423] & v0_en_i;
  assign v1_data_o[422] = v0_data_i[422] & v0_en_i;
  assign v1_data_o[421] = v0_data_i[421] & v0_en_i;
  assign v1_data_o[420] = v0_data_i[420] & v0_en_i;
  assign v1_data_o[419] = v0_data_i[419] & v0_en_i;
  assign v1_data_o[418] = v0_data_i[418] & v0_en_i;
  assign v1_data_o[417] = v0_data_i[417] & v0_en_i;
  assign v1_data_o[416] = v0_data_i[416] & v0_en_i;
  assign v1_data_o[415] = v0_data_i[415] & v0_en_i;
  assign v1_data_o[414] = v0_data_i[414] & v0_en_i;
  assign v1_data_o[413] = v0_data_i[413] & v0_en_i;
  assign v1_data_o[412] = v0_data_i[412] & v0_en_i;
  assign v1_data_o[411] = v0_data_i[411] & v0_en_i;
  assign v1_data_o[410] = v0_data_i[410] & v0_en_i;
  assign v1_data_o[409] = v0_data_i[409] & v0_en_i;
  assign v1_data_o[408] = v0_data_i[408] & v0_en_i;
  assign v1_data_o[407] = v0_data_i[407] & v0_en_i;
  assign v1_data_o[406] = v0_data_i[406] & v0_en_i;
  assign v1_data_o[405] = v0_data_i[405] & v0_en_i;
  assign v1_data_o[404] = v0_data_i[404] & v0_en_i;
  assign v1_data_o[403] = v0_data_i[403] & v0_en_i;
  assign v1_data_o[402] = v0_data_i[402] & v0_en_i;
  assign v1_data_o[401] = v0_data_i[401] & v0_en_i;
  assign v1_data_o[400] = v0_data_i[400] & v0_en_i;
  assign v1_data_o[399] = v0_data_i[399] & v0_en_i;
  assign v1_data_o[398] = v0_data_i[398] & v0_en_i;
  assign v1_data_o[397] = v0_data_i[397] & v0_en_i;
  assign v1_data_o[396] = v0_data_i[396] & v0_en_i;
  assign v1_data_o[395] = v0_data_i[395] & v0_en_i;
  assign v1_data_o[394] = v0_data_i[394] & v0_en_i;
  assign v1_data_o[393] = v0_data_i[393] & v0_en_i;
  assign v1_data_o[392] = v0_data_i[392] & v0_en_i;
  assign v1_data_o[391] = v0_data_i[391] & v0_en_i;
  assign v1_data_o[390] = v0_data_i[390] & v0_en_i;
  assign v1_data_o[389] = v0_data_i[389] & v0_en_i;
  assign v1_data_o[388] = v0_data_i[388] & v0_en_i;
  assign v1_data_o[387] = v0_data_i[387] & v0_en_i;
  assign v1_data_o[386] = v0_data_i[386] & v0_en_i;
  assign v1_data_o[385] = v0_data_i[385] & v0_en_i;
  assign v1_data_o[384] = v0_data_i[384] & v0_en_i;
  assign v1_data_o[383] = v0_data_i[383] & v0_en_i;
  assign v1_data_o[382] = v0_data_i[382] & v0_en_i;
  assign v1_data_o[381] = v0_data_i[381] & v0_en_i;
  assign v1_data_o[380] = v0_data_i[380] & v0_en_i;
  assign v1_data_o[379] = v0_data_i[379] & v0_en_i;
  assign v1_data_o[378] = v0_data_i[378] & v0_en_i;
  assign v1_data_o[377] = v0_data_i[377] & v0_en_i;
  assign v1_data_o[376] = v0_data_i[376] & v0_en_i;
  assign v1_data_o[375] = v0_data_i[375] & v0_en_i;
  assign v1_data_o[374] = v0_data_i[374] & v0_en_i;
  assign v1_data_o[373] = v0_data_i[373] & v0_en_i;
  assign v1_data_o[372] = v0_data_i[372] & v0_en_i;
  assign v1_data_o[371] = v0_data_i[371] & v0_en_i;
  assign v1_data_o[370] = v0_data_i[370] & v0_en_i;
  assign v1_data_o[369] = v0_data_i[369] & v0_en_i;
  assign v1_data_o[368] = v0_data_i[368] & v0_en_i;
  assign v1_data_o[367] = v0_data_i[367] & v0_en_i;
  assign v1_data_o[366] = v0_data_i[366] & v0_en_i;
  assign v1_data_o[365] = v0_data_i[365] & v0_en_i;
  assign v1_data_o[364] = v0_data_i[364] & v0_en_i;
  assign v1_data_o[363] = v0_data_i[363] & v0_en_i;
  assign v1_data_o[362] = v0_data_i[362] & v0_en_i;
  assign v1_data_o[361] = v0_data_i[361] & v0_en_i;
  assign v1_data_o[360] = v0_data_i[360] & v0_en_i;
  assign v1_data_o[359] = v0_data_i[359] & v0_en_i;
  assign v1_data_o[358] = v0_data_i[358] & v0_en_i;
  assign v1_data_o[357] = v0_data_i[357] & v0_en_i;
  assign v1_data_o[356] = v0_data_i[356] & v0_en_i;
  assign v1_data_o[355] = v0_data_i[355] & v0_en_i;
  assign v1_data_o[354] = v0_data_i[354] & v0_en_i;
  assign v1_data_o[353] = v0_data_i[353] & v0_en_i;
  assign v1_data_o[352] = v0_data_i[352] & v0_en_i;
  assign v1_data_o[351] = v0_data_i[351] & v0_en_i;
  assign v1_data_o[350] = v0_data_i[350] & v0_en_i;
  assign v1_data_o[349] = v0_data_i[349] & v0_en_i;
  assign v1_data_o[348] = v0_data_i[348] & v0_en_i;
  assign v1_data_o[347] = v0_data_i[347] & v0_en_i;
  assign v1_data_o[346] = v0_data_i[346] & v0_en_i;
  assign v1_data_o[345] = v0_data_i[345] & v0_en_i;
  assign v1_data_o[344] = v0_data_i[344] & v0_en_i;
  assign v1_data_o[343] = v0_data_i[343] & v0_en_i;
  assign v1_data_o[342] = v0_data_i[342] & v0_en_i;
  assign v1_data_o[341] = v0_data_i[341] & v0_en_i;
  assign v1_data_o[340] = v0_data_i[340] & v0_en_i;
  assign v1_data_o[339] = v0_data_i[339] & v0_en_i;
  assign v1_data_o[338] = v0_data_i[338] & v0_en_i;
  assign v1_data_o[337] = v0_data_i[337] & v0_en_i;
  assign v1_data_o[336] = v0_data_i[336] & v0_en_i;
  assign v1_data_o[335] = v0_data_i[335] & v0_en_i;
  assign v1_data_o[334] = v0_data_i[334] & v0_en_i;
  assign v1_data_o[333] = v0_data_i[333] & v0_en_i;
  assign v1_data_o[332] = v0_data_i[332] & v0_en_i;
  assign v1_data_o[331] = v0_data_i[331] & v0_en_i;
  assign v1_data_o[330] = v0_data_i[330] & v0_en_i;
  assign v1_data_o[329] = v0_data_i[329] & v0_en_i;
  assign v1_data_o[328] = v0_data_i[328] & v0_en_i;
  assign v1_data_o[327] = v0_data_i[327] & v0_en_i;
  assign v1_data_o[326] = v0_data_i[326] & v0_en_i;
  assign v1_data_o[325] = v0_data_i[325] & v0_en_i;
  assign v1_data_o[324] = v0_data_i[324] & v0_en_i;
  assign v1_data_o[323] = v0_data_i[323] & v0_en_i;
  assign v1_data_o[322] = v0_data_i[322] & v0_en_i;
  assign v1_data_o[321] = v0_data_i[321] & v0_en_i;
  assign v1_data_o[320] = v0_data_i[320] & v0_en_i;
  assign v1_data_o[319] = v0_data_i[319] & v0_en_i;
  assign v1_data_o[318] = v0_data_i[318] & v0_en_i;
  assign v1_data_o[317] = v0_data_i[317] & v0_en_i;
  assign v1_data_o[316] = v0_data_i[316] & v0_en_i;
  assign v1_data_o[315] = v0_data_i[315] & v0_en_i;
  assign v1_data_o[314] = v0_data_i[314] & v0_en_i;
  assign v1_data_o[313] = v0_data_i[313] & v0_en_i;
  assign v1_data_o[312] = v0_data_i[312] & v0_en_i;
  assign v1_data_o[311] = v0_data_i[311] & v0_en_i;
  assign v1_data_o[310] = v0_data_i[310] & v0_en_i;
  assign v1_data_o[309] = v0_data_i[309] & v0_en_i;
  assign v1_data_o[308] = v0_data_i[308] & v0_en_i;
  assign v1_data_o[307] = v0_data_i[307] & v0_en_i;
  assign v1_data_o[306] = v0_data_i[306] & v0_en_i;
  assign v1_data_o[305] = v0_data_i[305] & v0_en_i;
  assign v1_data_o[304] = v0_data_i[304] & v0_en_i;
  assign v1_data_o[303] = v0_data_i[303] & v0_en_i;
  assign v1_data_o[302] = v0_data_i[302] & v0_en_i;
  assign v1_data_o[301] = v0_data_i[301] & v0_en_i;
  assign v1_data_o[300] = v0_data_i[300] & v0_en_i;
  assign v1_data_o[299] = v0_data_i[299] & v0_en_i;
  assign v1_data_o[298] = v0_data_i[298] & v0_en_i;
  assign v1_data_o[297] = v0_data_i[297] & v0_en_i;
  assign v1_data_o[296] = v0_data_i[296] & v0_en_i;
  assign v1_data_o[295] = v0_data_i[295] & v0_en_i;
  assign v1_data_o[294] = v0_data_i[294] & v0_en_i;
  assign v1_data_o[293] = v0_data_i[293] & v0_en_i;
  assign v1_data_o[292] = v0_data_i[292] & v0_en_i;
  assign v1_data_o[291] = v0_data_i[291] & v0_en_i;
  assign v1_data_o[290] = v0_data_i[290] & v0_en_i;
  assign v1_data_o[289] = v0_data_i[289] & v0_en_i;
  assign v1_data_o[288] = v0_data_i[288] & v0_en_i;
  assign v1_data_o[287] = v0_data_i[287] & v0_en_i;
  assign v1_data_o[286] = v0_data_i[286] & v0_en_i;
  assign v1_data_o[285] = v0_data_i[285] & v0_en_i;
  assign v1_data_o[284] = v0_data_i[284] & v0_en_i;
  assign v1_data_o[283] = v0_data_i[283] & v0_en_i;
  assign v1_data_o[282] = v0_data_i[282] & v0_en_i;
  assign v1_data_o[281] = v0_data_i[281] & v0_en_i;
  assign v1_data_o[280] = v0_data_i[280] & v0_en_i;
  assign v1_data_o[279] = v0_data_i[279] & v0_en_i;
  assign v1_data_o[278] = v0_data_i[278] & v0_en_i;
  assign v1_data_o[277] = v0_data_i[277] & v0_en_i;
  assign v1_data_o[276] = v0_data_i[276] & v0_en_i;
  assign v1_data_o[275] = v0_data_i[275] & v0_en_i;
  assign v1_data_o[274] = v0_data_i[274] & v0_en_i;
  assign v1_data_o[273] = v0_data_i[273] & v0_en_i;
  assign v1_data_o[272] = v0_data_i[272] & v0_en_i;
  assign v1_data_o[271] = v0_data_i[271] & v0_en_i;
  assign v1_data_o[270] = v0_data_i[270] & v0_en_i;
  assign v1_data_o[269] = v0_data_i[269] & v0_en_i;
  assign v1_data_o[268] = v0_data_i[268] & v0_en_i;
  assign v1_data_o[267] = v0_data_i[267] & v0_en_i;
  assign v1_data_o[266] = v0_data_i[266] & v0_en_i;
  assign v1_data_o[265] = v0_data_i[265] & v0_en_i;
  assign v1_data_o[264] = v0_data_i[264] & v0_en_i;
  assign v1_data_o[263] = v0_data_i[263] & v0_en_i;
  assign v1_data_o[262] = v0_data_i[262] & v0_en_i;
  assign v1_data_o[261] = v0_data_i[261] & v0_en_i;
  assign v1_data_o[260] = v0_data_i[260] & v0_en_i;
  assign v1_data_o[259] = v0_data_i[259] & v0_en_i;
  assign v1_data_o[258] = v0_data_i[258] & v0_en_i;
  assign v1_data_o[257] = v0_data_i[257] & v0_en_i;
  assign v1_data_o[256] = v0_data_i[256] & v0_en_i;
  assign v1_data_o[255] = v0_data_i[255] & v0_en_i;
  assign v1_data_o[254] = v0_data_i[254] & v0_en_i;
  assign v1_data_o[253] = v0_data_i[253] & v0_en_i;
  assign v1_data_o[252] = v0_data_i[252] & v0_en_i;
  assign v1_data_o[251] = v0_data_i[251] & v0_en_i;
  assign v1_data_o[250] = v0_data_i[250] & v0_en_i;
  assign v1_data_o[249] = v0_data_i[249] & v0_en_i;
  assign v1_data_o[248] = v0_data_i[248] & v0_en_i;
  assign v1_data_o[247] = v0_data_i[247] & v0_en_i;
  assign v1_data_o[246] = v0_data_i[246] & v0_en_i;
  assign v1_data_o[245] = v0_data_i[245] & v0_en_i;
  assign v1_data_o[244] = v0_data_i[244] & v0_en_i;
  assign v1_data_o[243] = v0_data_i[243] & v0_en_i;
  assign v1_data_o[242] = v0_data_i[242] & v0_en_i;
  assign v1_data_o[241] = v0_data_i[241] & v0_en_i;
  assign v1_data_o[240] = v0_data_i[240] & v0_en_i;
  assign v1_data_o[239] = v0_data_i[239] & v0_en_i;
  assign v1_data_o[238] = v0_data_i[238] & v0_en_i;
  assign v1_data_o[237] = v0_data_i[237] & v0_en_i;
  assign v1_data_o[236] = v0_data_i[236] & v0_en_i;
  assign v1_data_o[235] = v0_data_i[235] & v0_en_i;
  assign v1_data_o[234] = v0_data_i[234] & v0_en_i;
  assign v1_data_o[233] = v0_data_i[233] & v0_en_i;
  assign v1_data_o[232] = v0_data_i[232] & v0_en_i;
  assign v1_data_o[231] = v0_data_i[231] & v0_en_i;
  assign v1_data_o[230] = v0_data_i[230] & v0_en_i;
  assign v1_data_o[229] = v0_data_i[229] & v0_en_i;
  assign v1_data_o[228] = v0_data_i[228] & v0_en_i;
  assign v1_data_o[227] = v0_data_i[227] & v0_en_i;
  assign v1_data_o[226] = v0_data_i[226] & v0_en_i;
  assign v1_data_o[225] = v0_data_i[225] & v0_en_i;
  assign v1_data_o[224] = v0_data_i[224] & v0_en_i;
  assign v1_data_o[223] = v0_data_i[223] & v0_en_i;
  assign v1_data_o[222] = v0_data_i[222] & v0_en_i;
  assign v1_data_o[221] = v0_data_i[221] & v0_en_i;
  assign v1_data_o[220] = v0_data_i[220] & v0_en_i;
  assign v1_data_o[219] = v0_data_i[219] & v0_en_i;
  assign v1_data_o[218] = v0_data_i[218] & v0_en_i;
  assign v1_data_o[217] = v0_data_i[217] & v0_en_i;
  assign v1_data_o[216] = v0_data_i[216] & v0_en_i;
  assign v1_data_o[215] = v0_data_i[215] & v0_en_i;
  assign v1_data_o[214] = v0_data_i[214] & v0_en_i;
  assign v1_data_o[213] = v0_data_i[213] & v0_en_i;
  assign v1_data_o[212] = v0_data_i[212] & v0_en_i;
  assign v1_data_o[211] = v0_data_i[211] & v0_en_i;
  assign v1_data_o[210] = v0_data_i[210] & v0_en_i;
  assign v1_data_o[209] = v0_data_i[209] & v0_en_i;
  assign v1_data_o[208] = v0_data_i[208] & v0_en_i;
  assign v1_data_o[207] = v0_data_i[207] & v0_en_i;
  assign v1_data_o[206] = v0_data_i[206] & v0_en_i;
  assign v1_data_o[205] = v0_data_i[205] & v0_en_i;
  assign v1_data_o[204] = v0_data_i[204] & v0_en_i;
  assign v1_data_o[203] = v0_data_i[203] & v0_en_i;
  assign v1_data_o[202] = v0_data_i[202] & v0_en_i;
  assign v1_data_o[201] = v0_data_i[201] & v0_en_i;
  assign v1_data_o[200] = v0_data_i[200] & v0_en_i;
  assign v1_data_o[199] = v0_data_i[199] & v0_en_i;
  assign v1_data_o[198] = v0_data_i[198] & v0_en_i;
  assign v1_data_o[197] = v0_data_i[197] & v0_en_i;
  assign v1_data_o[196] = v0_data_i[196] & v0_en_i;
  assign v1_data_o[195] = v0_data_i[195] & v0_en_i;
  assign v1_data_o[194] = v0_data_i[194] & v0_en_i;
  assign v1_data_o[193] = v0_data_i[193] & v0_en_i;
  assign v1_data_o[192] = v0_data_i[192] & v0_en_i;
  assign v1_data_o[191] = v0_data_i[191] & v0_en_i;
  assign v1_data_o[190] = v0_data_i[190] & v0_en_i;
  assign v1_data_o[189] = v0_data_i[189] & v0_en_i;
  assign v1_data_o[188] = v0_data_i[188] & v0_en_i;
  assign v1_data_o[187] = v0_data_i[187] & v0_en_i;
  assign v1_data_o[186] = v0_data_i[186] & v0_en_i;
  assign v1_data_o[185] = v0_data_i[185] & v0_en_i;
  assign v1_data_o[184] = v0_data_i[184] & v0_en_i;
  assign v1_data_o[183] = v0_data_i[183] & v0_en_i;
  assign v1_data_o[182] = v0_data_i[182] & v0_en_i;
  assign v1_data_o[181] = v0_data_i[181] & v0_en_i;
  assign v1_data_o[180] = v0_data_i[180] & v0_en_i;
  assign v1_data_o[179] = v0_data_i[179] & v0_en_i;
  assign v1_data_o[178] = v0_data_i[178] & v0_en_i;
  assign v1_data_o[177] = v0_data_i[177] & v0_en_i;
  assign v1_data_o[176] = v0_data_i[176] & v0_en_i;
  assign v1_data_o[175] = v0_data_i[175] & v0_en_i;
  assign v1_data_o[174] = v0_data_i[174] & v0_en_i;
  assign v1_data_o[173] = v0_data_i[173] & v0_en_i;
  assign v1_data_o[172] = v0_data_i[172] & v0_en_i;
  assign v1_data_o[171] = v0_data_i[171] & v0_en_i;
  assign v1_data_o[170] = v0_data_i[170] & v0_en_i;
  assign v1_data_o[169] = v0_data_i[169] & v0_en_i;
  assign v1_data_o[168] = v0_data_i[168] & v0_en_i;
  assign v1_data_o[167] = v0_data_i[167] & v0_en_i;
  assign v1_data_o[166] = v0_data_i[166] & v0_en_i;
  assign v1_data_o[165] = v0_data_i[165] & v0_en_i;
  assign v1_data_o[164] = v0_data_i[164] & v0_en_i;
  assign v1_data_o[163] = v0_data_i[163] & v0_en_i;
  assign v1_data_o[162] = v0_data_i[162] & v0_en_i;
  assign v1_data_o[161] = v0_data_i[161] & v0_en_i;
  assign v1_data_o[160] = v0_data_i[160] & v0_en_i;
  assign v1_data_o[159] = v0_data_i[159] & v0_en_i;
  assign v1_data_o[158] = v0_data_i[158] & v0_en_i;
  assign v1_data_o[157] = v0_data_i[157] & v0_en_i;
  assign v1_data_o[156] = v0_data_i[156] & v0_en_i;
  assign v1_data_o[155] = v0_data_i[155] & v0_en_i;
  assign v1_data_o[154] = v0_data_i[154] & v0_en_i;
  assign v1_data_o[153] = v0_data_i[153] & v0_en_i;
  assign v1_data_o[152] = v0_data_i[152] & v0_en_i;
  assign v1_data_o[151] = v0_data_i[151] & v0_en_i;
  assign v1_data_o[150] = v0_data_i[150] & v0_en_i;
  assign v1_data_o[149] = v0_data_i[149] & v0_en_i;
  assign v1_data_o[148] = v0_data_i[148] & v0_en_i;
  assign v1_data_o[147] = v0_data_i[147] & v0_en_i;
  assign v1_data_o[146] = v0_data_i[146] & v0_en_i;
  assign v1_data_o[145] = v0_data_i[145] & v0_en_i;
  assign v1_data_o[144] = v0_data_i[144] & v0_en_i;
  assign v1_data_o[143] = v0_data_i[143] & v0_en_i;
  assign v1_data_o[142] = v0_data_i[142] & v0_en_i;
  assign v1_data_o[141] = v0_data_i[141] & v0_en_i;
  assign v1_data_o[140] = v0_data_i[140] & v0_en_i;
  assign v1_data_o[139] = v0_data_i[139] & v0_en_i;
  assign v1_data_o[138] = v0_data_i[138] & v0_en_i;
  assign v1_data_o[137] = v0_data_i[137] & v0_en_i;
  assign v1_data_o[136] = v0_data_i[136] & v0_en_i;
  assign v1_data_o[135] = v0_data_i[135] & v0_en_i;
  assign v1_data_o[134] = v0_data_i[134] & v0_en_i;
  assign v1_data_o[133] = v0_data_i[133] & v0_en_i;
  assign v1_data_o[132] = v0_data_i[132] & v0_en_i;
  assign v1_data_o[131] = v0_data_i[131] & v0_en_i;
  assign v1_data_o[130] = v0_data_i[130] & v0_en_i;
  assign v1_data_o[129] = v0_data_i[129] & v0_en_i;
  assign v1_data_o[128] = v0_data_i[128] & v0_en_i;
  assign v1_data_o[127] = v0_data_i[127] & v0_en_i;
  assign v1_data_o[126] = v0_data_i[126] & v0_en_i;
  assign v1_data_o[125] = v0_data_i[125] & v0_en_i;
  assign v1_data_o[124] = v0_data_i[124] & v0_en_i;
  assign v1_data_o[123] = v0_data_i[123] & v0_en_i;
  assign v1_data_o[122] = v0_data_i[122] & v0_en_i;
  assign v1_data_o[121] = v0_data_i[121] & v0_en_i;
  assign v1_data_o[120] = v0_data_i[120] & v0_en_i;
  assign v1_data_o[119] = v0_data_i[119] & v0_en_i;
  assign v1_data_o[118] = v0_data_i[118] & v0_en_i;
  assign v1_data_o[117] = v0_data_i[117] & v0_en_i;
  assign v1_data_o[116] = v0_data_i[116] & v0_en_i;
  assign v1_data_o[115] = v0_data_i[115] & v0_en_i;
  assign v1_data_o[114] = v0_data_i[114] & v0_en_i;
  assign v1_data_o[113] = v0_data_i[113] & v0_en_i;
  assign v1_data_o[112] = v0_data_i[112] & v0_en_i;
  assign v1_data_o[111] = v0_data_i[111] & v0_en_i;
  assign v1_data_o[110] = v0_data_i[110] & v0_en_i;
  assign v1_data_o[109] = v0_data_i[109] & v0_en_i;
  assign v1_data_o[108] = v0_data_i[108] & v0_en_i;
  assign v1_data_o[107] = v0_data_i[107] & v0_en_i;
  assign v1_data_o[106] = v0_data_i[106] & v0_en_i;
  assign v1_data_o[105] = v0_data_i[105] & v0_en_i;
  assign v1_data_o[104] = v0_data_i[104] & v0_en_i;
  assign v1_data_o[103] = v0_data_i[103] & v0_en_i;
  assign v1_data_o[102] = v0_data_i[102] & v0_en_i;
  assign v1_data_o[101] = v0_data_i[101] & v0_en_i;
  assign v1_data_o[100] = v0_data_i[100] & v0_en_i;
  assign v1_data_o[99] = v0_data_i[99] & v0_en_i;
  assign v1_data_o[98] = v0_data_i[98] & v0_en_i;
  assign v1_data_o[97] = v0_data_i[97] & v0_en_i;
  assign v1_data_o[96] = v0_data_i[96] & v0_en_i;
  assign v1_data_o[95] = v0_data_i[95] & v0_en_i;
  assign v1_data_o[94] = v0_data_i[94] & v0_en_i;
  assign v1_data_o[93] = v0_data_i[93] & v0_en_i;
  assign v1_data_o[92] = v0_data_i[92] & v0_en_i;
  assign v1_data_o[91] = v0_data_i[91] & v0_en_i;
  assign v1_data_o[90] = v0_data_i[90] & v0_en_i;
  assign v1_data_o[89] = v0_data_i[89] & v0_en_i;
  assign v1_data_o[88] = v0_data_i[88] & v0_en_i;
  assign v1_data_o[87] = v0_data_i[87] & v0_en_i;
  assign v1_data_o[86] = v0_data_i[86] & v0_en_i;
  assign v1_data_o[85] = v0_data_i[85] & v0_en_i;
  assign v1_data_o[84] = v0_data_i[84] & v0_en_i;
  assign v1_data_o[83] = v0_data_i[83] & v0_en_i;
  assign v1_data_o[82] = v0_data_i[82] & v0_en_i;
  assign v1_data_o[81] = v0_data_i[81] & v0_en_i;
  assign v1_data_o[80] = v0_data_i[80] & v0_en_i;
  assign v1_data_o[79] = v0_data_i[79] & v0_en_i;
  assign v1_data_o[78] = v0_data_i[78] & v0_en_i;
  assign v1_data_o[77] = v0_data_i[77] & v0_en_i;
  assign v1_data_o[76] = v0_data_i[76] & v0_en_i;
  assign v1_data_o[75] = v0_data_i[75] & v0_en_i;
  assign v1_data_o[74] = v0_data_i[74] & v0_en_i;
  assign v1_data_o[73] = v0_data_i[73] & v0_en_i;
  assign v1_data_o[72] = v0_data_i[72] & v0_en_i;
  assign v1_data_o[71] = v0_data_i[71] & v0_en_i;
  assign v1_data_o[70] = v0_data_i[70] & v0_en_i;
  assign v1_data_o[69] = v0_data_i[69] & v0_en_i;
  assign v1_data_o[68] = v0_data_i[68] & v0_en_i;
  assign v1_data_o[67] = v0_data_i[67] & v0_en_i;
  assign v1_data_o[66] = v0_data_i[66] & v0_en_i;
  assign v1_data_o[65] = v0_data_i[65] & v0_en_i;
  assign v1_data_o[64] = v0_data_i[64] & v0_en_i;
  assign v1_data_o[63] = v0_data_i[63] & v0_en_i;
  assign v1_data_o[62] = v0_data_i[62] & v0_en_i;
  assign v1_data_o[61] = v0_data_i[61] & v0_en_i;
  assign v1_data_o[60] = v0_data_i[60] & v0_en_i;
  assign v1_data_o[59] = v0_data_i[59] & v0_en_i;
  assign v1_data_o[58] = v0_data_i[58] & v0_en_i;
  assign v1_data_o[57] = v0_data_i[57] & v0_en_i;
  assign v1_data_o[56] = v0_data_i[56] & v0_en_i;
  assign v1_data_o[55] = v0_data_i[55] & v0_en_i;
  assign v1_data_o[54] = v0_data_i[54] & v0_en_i;
  assign v1_data_o[53] = v0_data_i[53] & v0_en_i;
  assign v1_data_o[52] = v0_data_i[52] & v0_en_i;
  assign v1_data_o[51] = v0_data_i[51] & v0_en_i;
  assign v1_data_o[50] = v0_data_i[50] & v0_en_i;
  assign v1_data_o[49] = v0_data_i[49] & v0_en_i;
  assign v1_data_o[48] = v0_data_i[48] & v0_en_i;
  assign v1_data_o[47] = v0_data_i[47] & v0_en_i;
  assign v1_data_o[46] = v0_data_i[46] & v0_en_i;
  assign v1_data_o[45] = v0_data_i[45] & v0_en_i;
  assign v1_data_o[44] = v0_data_i[44] & v0_en_i;
  assign v1_data_o[43] = v0_data_i[43] & v0_en_i;
  assign v1_data_o[42] = v0_data_i[42] & v0_en_i;
  assign v1_data_o[41] = v0_data_i[41] & v0_en_i;
  assign v1_data_o[40] = v0_data_i[40] & v0_en_i;
  assign v1_data_o[39] = v0_data_i[39] & v0_en_i;
  assign v1_data_o[38] = v0_data_i[38] & v0_en_i;
  assign v1_data_o[37] = v0_data_i[37] & v0_en_i;
  assign v1_data_o[36] = v0_data_i[36] & v0_en_i;
  assign v1_data_o[35] = v0_data_i[35] & v0_en_i;
  assign v1_data_o[34] = v0_data_i[34] & v0_en_i;
  assign v1_data_o[33] = v0_data_i[33] & v0_en_i;
  assign v1_data_o[32] = v0_data_i[32] & v0_en_i;
  assign v1_data_o[31] = v0_data_i[31] & v0_en_i;
  assign v1_data_o[30] = v0_data_i[30] & v0_en_i;
  assign v1_data_o[29] = v0_data_i[29] & v0_en_i;
  assign v1_data_o[28] = v0_data_i[28] & v0_en_i;
  assign v1_data_o[27] = v0_data_i[27] & v0_en_i;
  assign v1_data_o[26] = v0_data_i[26] & v0_en_i;
  assign v1_data_o[25] = v0_data_i[25] & v0_en_i;
  assign v1_data_o[24] = v0_data_i[24] & v0_en_i;
  assign v1_data_o[23] = v0_data_i[23] & v0_en_i;
  assign v1_data_o[22] = v0_data_i[22] & v0_en_i;
  assign v1_data_o[21] = v0_data_i[21] & v0_en_i;
  assign v1_data_o[20] = v0_data_i[20] & v0_en_i;
  assign v1_data_o[19] = v0_data_i[19] & v0_en_i;
  assign v1_data_o[18] = v0_data_i[18] & v0_en_i;
  assign v1_data_o[17] = v0_data_i[17] & v0_en_i;
  assign v1_data_o[16] = v0_data_i[16] & v0_en_i;
  assign v1_data_o[15] = v0_data_i[15] & v0_en_i;
  assign v1_data_o[14] = v0_data_i[14] & v0_en_i;
  assign v1_data_o[13] = v0_data_i[13] & v0_en_i;
  assign v1_data_o[12] = v0_data_i[12] & v0_en_i;
  assign v1_data_o[11] = v0_data_i[11] & v0_en_i;
  assign v1_data_o[10] = v0_data_i[10] & v0_en_i;
  assign v1_data_o[9] = v0_data_i[9] & v0_en_i;
  assign v1_data_o[8] = v0_data_i[8] & v0_en_i;
  assign v1_data_o[7] = v0_data_i[7] & v0_en_i;
  assign v1_data_o[6] = v0_data_i[6] & v0_en_i;
  assign v1_data_o[5] = v0_data_i[5] & v0_en_i;
  assign v1_data_o[4] = v0_data_i[4] & v0_en_i;
  assign v1_data_o[3] = v0_data_i[3] & v0_en_i;
  assign v1_data_o[2] = v0_data_i[2] & v0_en_i;
  assign v1_data_o[1] = v0_data_i[1] & v0_en_i;
  assign v1_data_o[0] = v0_data_i[0] & v0_en_i;

endmodule



module bsg_fsb_node_level_shift_fsb_domain
(
  en_ls_i,
  clk_i,
  reset_i,
  clk_o,
  reset_o,
  fsb_v_i_o,
  fsb_data_i_o,
  fsb_yumi_o_i,
  fsb_v_o_i,
  fsb_data_o_i,
  fsb_ready_i_o,
  node_v_i_o,
  node_data_i_o,
  node_ready_o_i,
  node_v_o_i,
  node_data_o_i,
  node_yumi_i_o
);

  output [999:0] fsb_data_i_o;
  input [999:0] fsb_data_o_i;
  output [999:0] node_data_i_o;
  input [999:0] node_data_o_i;
  input en_ls_i;
  input clk_i;
  input reset_i;
  input fsb_yumi_o_i;
  input fsb_v_o_i;
  input node_ready_o_i;
  input node_v_o_i;
  output clk_o;
  output reset_o;
  output fsb_v_i_o;
  output fsb_ready_i_o;
  output node_v_i_o;
  output node_yumi_i_o;
  wire [999:0] fsb_data_i_o,node_data_i_o;
  wire clk_o,reset_o,fsb_v_i_o,fsb_ready_i_o,node_v_i_o,node_yumi_i_o;

  bsg_level_shift_up_down_source_width_p1
  clk_ls_inst
  (
    .v0_en_i(1'b1),
    .v0_data_i(clk_i),
    .v1_data_o(clk_o)
  );


  bsg_level_shift_up_down_source_width_p1
  reset_ls_inst
  (
    .v0_en_i(1'b1),
    .v0_data_i(reset_i),
    .v1_data_o(reset_o)
  );


  bsg_level_shift_up_down_sink_width_p1
  n2f_v_ls_inst
  (
    .v0_data_i(node_v_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(fsb_v_i_o)
  );


  bsg_level_shift_up_down_sink_width_p1000
  n2f_data_ls_inst
  (
    .v0_data_i(node_data_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(fsb_data_i_o)
  );


  bsg_level_shift_up_down_source_width_p1
  f2n_yumi_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(fsb_yumi_o_i),
    .v1_data_o(node_yumi_i_o)
  );


  bsg_level_shift_up_down_source_width_p1
  f2n_v_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(fsb_v_o_i),
    .v1_data_o(node_v_i_o)
  );


  bsg_level_shift_up_down_source_width_p1000
  f2n_data_ls_inst
  (
    .v0_en_i(en_ls_i),
    .v0_data_i(fsb_data_o_i),
    .v1_data_o(node_data_i_o)
  );


  bsg_level_shift_up_down_sink_width_p1
  n2f_ready_ls_inst
  (
    .v0_data_i(node_ready_o_i),
    .v1_en_i(en_ls_i),
    .v1_data_o(fsb_ready_i_o)
  );


endmodule

