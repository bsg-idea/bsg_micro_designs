

module top
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_cnt_i
);

  input [31:0] data_i;
  output [63:0] valid_o;
  output [2047:0] data_o;
  input [6:0] yumi_cnt_i;
  input clk_i;
  input reset_i;
  input valid_i;
  output ready_o;

  bsg_serial_in_parallel_out
  wrapper
  (
    .data_i(data_i),
    .valid_o(valid_o),
    .data_o(data_o),
    .yumi_cnt_i(yumi_cnt_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .valid_i(valid_i),
    .ready_o(ready_o)
  );


endmodule



module bsg_serial_in_parallel_out
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_cnt_i
);

  input [31:0] data_i;
  output [63:0] valid_o;
  output [2047:0] data_o;
  input [6:0] yumi_cnt_i;
  input clk_i;
  input reset_i;
  input valid_i;
  output ready_o;
  wire [63:0] valid_o,valid_r,valid_nn;
  wire [2047:0] data_o,data_r,data_nn;
  wire ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,
  N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
  N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,
  N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,
  N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,
  N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,
  N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,
  N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
  N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,
  N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,
  N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
  N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,
  N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,
  N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,
  N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,
  N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,
  N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,
  N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,
  N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,
  N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,
  N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,
  N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,
  N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,
  N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,
  N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
  N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,
  N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,
  N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,
  N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,
  N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,
  N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,
  N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,
  N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,
  N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,
  N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,
  N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
  N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,
  N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,
  N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,
  N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,
  N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,
  N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,
  N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,
  N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,
  N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,
  N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,
  N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,
  N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,
  N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,
  N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,
  N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,
  N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,
  N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,
  N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,
  N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,
  N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,
  N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,
  N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,
  N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,
  N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,
  N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,
  N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,
  N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,
  N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,
  N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,
  N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,
  N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,
  N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,
  N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,
  N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,
  N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,
  N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,
  N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,
  N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,
  N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,
  N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,
  N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,
  N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,
  N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,
  N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,
  N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,
  N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,
  N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,
  N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,
  N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,
  N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,
  N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,
  N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,
  N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,
  N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,
  N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,
  N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,
  N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,
  N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,
  N2237,data_n_127__31_,data_n_127__30_,data_n_127__29_,data_n_127__28_,
  data_n_127__27_,data_n_127__26_,data_n_127__25_,data_n_127__24_,data_n_127__23_,
  data_n_127__22_,data_n_127__21_,data_n_127__20_,data_n_127__19_,data_n_127__18_,
  data_n_127__17_,data_n_127__16_,data_n_127__15_,data_n_127__14_,data_n_127__13_,
  data_n_127__12_,data_n_127__11_,data_n_127__10_,data_n_127__9_,data_n_127__8_,
  data_n_127__7_,data_n_127__6_,data_n_127__5_,data_n_127__4_,data_n_127__3_,data_n_127__2_,
  data_n_127__1_,data_n_127__0_,data_n_126__31_,data_n_126__30_,data_n_126__29_,
  data_n_126__28_,data_n_126__27_,data_n_126__26_,data_n_126__25_,data_n_126__24_,
  data_n_126__23_,data_n_126__22_,data_n_126__21_,data_n_126__20_,data_n_126__19_,
  data_n_126__18_,data_n_126__17_,data_n_126__16_,data_n_126__15_,data_n_126__14_,
  data_n_126__13_,data_n_126__12_,data_n_126__11_,data_n_126__10_,data_n_126__9_,
  data_n_126__8_,data_n_126__7_,data_n_126__6_,data_n_126__5_,data_n_126__4_,
  data_n_126__3_,data_n_126__2_,data_n_126__1_,data_n_126__0_,data_n_125__31_,
  data_n_125__30_,data_n_125__29_,data_n_125__28_,data_n_125__27_,data_n_125__26_,
  data_n_125__25_,data_n_125__24_,data_n_125__23_,data_n_125__22_,data_n_125__21_,
  data_n_125__20_,data_n_125__19_,data_n_125__18_,data_n_125__17_,data_n_125__16_,
  data_n_125__15_,data_n_125__14_,data_n_125__13_,data_n_125__12_,data_n_125__11_,
  data_n_125__10_,data_n_125__9_,data_n_125__8_,data_n_125__7_,data_n_125__6_,data_n_125__5_,
  data_n_125__4_,data_n_125__3_,data_n_125__2_,data_n_125__1_,data_n_125__0_,
  data_n_124__31_,data_n_124__30_,data_n_124__29_,data_n_124__28_,data_n_124__27_,
  data_n_124__26_,data_n_124__25_,data_n_124__24_,data_n_124__23_,data_n_124__22_,
  data_n_124__21_,data_n_124__20_,data_n_124__19_,data_n_124__18_,data_n_124__17_,
  data_n_124__16_,data_n_124__15_,data_n_124__14_,data_n_124__13_,data_n_124__12_,
  data_n_124__11_,data_n_124__10_,data_n_124__9_,data_n_124__8_,data_n_124__7_,
  data_n_124__6_,data_n_124__5_,data_n_124__4_,data_n_124__3_,data_n_124__2_,data_n_124__1_,
  data_n_124__0_,data_n_123__31_,data_n_123__30_,data_n_123__29_,data_n_123__28_,
  data_n_123__27_,data_n_123__26_,data_n_123__25_,data_n_123__24_,data_n_123__23_,
  data_n_123__22_,data_n_123__21_,data_n_123__20_,data_n_123__19_,data_n_123__18_,
  data_n_123__17_,data_n_123__16_,data_n_123__15_,data_n_123__14_,data_n_123__13_,
  data_n_123__12_,data_n_123__11_,data_n_123__10_,data_n_123__9_,data_n_123__8_,
  data_n_123__7_,data_n_123__6_,data_n_123__5_,data_n_123__4_,data_n_123__3_,
  data_n_123__2_,data_n_123__1_,data_n_123__0_,data_n_122__31_,data_n_122__30_,
  data_n_122__29_,data_n_122__28_,data_n_122__27_,data_n_122__26_,data_n_122__25_,
  data_n_122__24_,data_n_122__23_,data_n_122__22_,data_n_122__21_,data_n_122__20_,
  data_n_122__19_,data_n_122__18_,data_n_122__17_,data_n_122__16_,data_n_122__15_,
  data_n_122__14_,data_n_122__13_,data_n_122__12_,data_n_122__11_,data_n_122__10_,
  data_n_122__9_,data_n_122__8_,data_n_122__7_,data_n_122__6_,data_n_122__5_,data_n_122__4_,
  data_n_122__3_,data_n_122__2_,data_n_122__1_,data_n_122__0_,data_n_121__31_,
  data_n_121__30_,data_n_121__29_,data_n_121__28_,data_n_121__27_,data_n_121__26_,
  data_n_121__25_,data_n_121__24_,data_n_121__23_,data_n_121__22_,data_n_121__21_,
  data_n_121__20_,data_n_121__19_,data_n_121__18_,data_n_121__17_,data_n_121__16_,
  data_n_121__15_,data_n_121__14_,data_n_121__13_,data_n_121__12_,data_n_121__11_,
  data_n_121__10_,data_n_121__9_,data_n_121__8_,data_n_121__7_,data_n_121__6_,
  data_n_121__5_,data_n_121__4_,data_n_121__3_,data_n_121__2_,data_n_121__1_,data_n_121__0_,
  data_n_120__31_,data_n_120__30_,data_n_120__29_,data_n_120__28_,data_n_120__27_,
  data_n_120__26_,data_n_120__25_,data_n_120__24_,data_n_120__23_,data_n_120__22_,
  data_n_120__21_,data_n_120__20_,data_n_120__19_,data_n_120__18_,data_n_120__17_,
  data_n_120__16_,data_n_120__15_,data_n_120__14_,data_n_120__13_,data_n_120__12_,
  data_n_120__11_,data_n_120__10_,data_n_120__9_,data_n_120__8_,data_n_120__7_,
  data_n_120__6_,data_n_120__5_,data_n_120__4_,data_n_120__3_,data_n_120__2_,
  data_n_120__1_,data_n_120__0_,data_n_119__31_,data_n_119__30_,data_n_119__29_,
  data_n_119__28_,data_n_119__27_,data_n_119__26_,data_n_119__25_,data_n_119__24_,
  data_n_119__23_,data_n_119__22_,data_n_119__21_,data_n_119__20_,data_n_119__19_,
  data_n_119__18_,data_n_119__17_,data_n_119__16_,data_n_119__15_,data_n_119__14_,
  data_n_119__13_,data_n_119__12_,data_n_119__11_,data_n_119__10_,data_n_119__9_,
  data_n_119__8_,data_n_119__7_,data_n_119__6_,data_n_119__5_,data_n_119__4_,data_n_119__3_,
  data_n_119__2_,data_n_119__1_,data_n_119__0_,data_n_118__31_,data_n_118__30_,
  data_n_118__29_,data_n_118__28_,data_n_118__27_,data_n_118__26_,data_n_118__25_,
  data_n_118__24_,data_n_118__23_,data_n_118__22_,data_n_118__21_,data_n_118__20_,
  data_n_118__19_,data_n_118__18_,data_n_118__17_,data_n_118__16_,data_n_118__15_,
  data_n_118__14_,data_n_118__13_,data_n_118__12_,data_n_118__11_,data_n_118__10_,
  data_n_118__9_,data_n_118__8_,data_n_118__7_,data_n_118__6_,data_n_118__5_,
  data_n_118__4_,data_n_118__3_,data_n_118__2_,data_n_118__1_,data_n_118__0_,
  data_n_117__31_,data_n_117__30_,data_n_117__29_,data_n_117__28_,data_n_117__27_,
  data_n_117__26_,data_n_117__25_,data_n_117__24_,data_n_117__23_,data_n_117__22_,
  data_n_117__21_,data_n_117__20_,data_n_117__19_,data_n_117__18_,data_n_117__17_,
  data_n_117__16_,data_n_117__15_,data_n_117__14_,data_n_117__13_,data_n_117__12_,
  data_n_117__11_,data_n_117__10_,data_n_117__9_,data_n_117__8_,data_n_117__7_,data_n_117__6_,
  data_n_117__5_,data_n_117__4_,data_n_117__3_,data_n_117__2_,data_n_117__1_,
  data_n_117__0_,data_n_116__31_,data_n_116__30_,data_n_116__29_,data_n_116__28_,
  data_n_116__27_,data_n_116__26_,data_n_116__25_,data_n_116__24_,data_n_116__23_,
  data_n_116__22_,data_n_116__21_,data_n_116__20_,data_n_116__19_,data_n_116__18_,
  data_n_116__17_,data_n_116__16_,data_n_116__15_,data_n_116__14_,data_n_116__13_,
  data_n_116__12_,data_n_116__11_,data_n_116__10_,data_n_116__9_,data_n_116__8_,
  data_n_116__7_,data_n_116__6_,data_n_116__5_,data_n_116__4_,data_n_116__3_,data_n_116__2_,
  data_n_116__1_,data_n_116__0_,data_n_115__31_,data_n_115__30_,data_n_115__29_,
  data_n_115__28_,data_n_115__27_,data_n_115__26_,data_n_115__25_,data_n_115__24_,
  data_n_115__23_,data_n_115__22_,data_n_115__21_,data_n_115__20_,data_n_115__19_,
  data_n_115__18_,data_n_115__17_,data_n_115__16_,data_n_115__15_,data_n_115__14_,
  data_n_115__13_,data_n_115__12_,data_n_115__11_,data_n_115__10_,data_n_115__9_,
  data_n_115__8_,data_n_115__7_,data_n_115__6_,data_n_115__5_,data_n_115__4_,
  data_n_115__3_,data_n_115__2_,data_n_115__1_,data_n_115__0_,data_n_114__31_,
  data_n_114__30_,data_n_114__29_,data_n_114__28_,data_n_114__27_,data_n_114__26_,
  data_n_114__25_,data_n_114__24_,data_n_114__23_,data_n_114__22_,data_n_114__21_,
  data_n_114__20_,data_n_114__19_,data_n_114__18_,data_n_114__17_,data_n_114__16_,
  data_n_114__15_,data_n_114__14_,data_n_114__13_,data_n_114__12_,data_n_114__11_,
  data_n_114__10_,data_n_114__9_,data_n_114__8_,data_n_114__7_,data_n_114__6_,data_n_114__5_,
  data_n_114__4_,data_n_114__3_,data_n_114__2_,data_n_114__1_,data_n_114__0_,
  data_n_113__31_,data_n_113__30_,data_n_113__29_,data_n_113__28_,data_n_113__27_,
  data_n_113__26_,data_n_113__25_,data_n_113__24_,data_n_113__23_,data_n_113__22_,
  data_n_113__21_,data_n_113__20_,data_n_113__19_,data_n_113__18_,data_n_113__17_,
  data_n_113__16_,data_n_113__15_,data_n_113__14_,data_n_113__13_,data_n_113__12_,
  data_n_113__11_,data_n_113__10_,data_n_113__9_,data_n_113__8_,data_n_113__7_,
  data_n_113__6_,data_n_113__5_,data_n_113__4_,data_n_113__3_,data_n_113__2_,
  data_n_113__1_,data_n_113__0_,data_n_112__31_,data_n_112__30_,data_n_112__29_,data_n_112__28_,
  data_n_112__27_,data_n_112__26_,data_n_112__25_,data_n_112__24_,data_n_112__23_,
  data_n_112__22_,data_n_112__21_,data_n_112__20_,data_n_112__19_,data_n_112__18_,
  data_n_112__17_,data_n_112__16_,data_n_112__15_,data_n_112__14_,data_n_112__13_,
  data_n_112__12_,data_n_112__11_,data_n_112__10_,data_n_112__9_,data_n_112__8_,
  data_n_112__7_,data_n_112__6_,data_n_112__5_,data_n_112__4_,data_n_112__3_,
  data_n_112__2_,data_n_112__1_,data_n_112__0_,data_n_111__31_,data_n_111__30_,
  data_n_111__29_,data_n_111__28_,data_n_111__27_,data_n_111__26_,data_n_111__25_,
  data_n_111__24_,data_n_111__23_,data_n_111__22_,data_n_111__21_,data_n_111__20_,
  data_n_111__19_,data_n_111__18_,data_n_111__17_,data_n_111__16_,data_n_111__15_,
  data_n_111__14_,data_n_111__13_,data_n_111__12_,data_n_111__11_,data_n_111__10_,
  data_n_111__9_,data_n_111__8_,data_n_111__7_,data_n_111__6_,data_n_111__5_,data_n_111__4_,
  data_n_111__3_,data_n_111__2_,data_n_111__1_,data_n_111__0_,data_n_110__31_,
  data_n_110__30_,data_n_110__29_,data_n_110__28_,data_n_110__27_,data_n_110__26_,
  data_n_110__25_,data_n_110__24_,data_n_110__23_,data_n_110__22_,data_n_110__21_,
  data_n_110__20_,data_n_110__19_,data_n_110__18_,data_n_110__17_,data_n_110__16_,
  data_n_110__15_,data_n_110__14_,data_n_110__13_,data_n_110__12_,data_n_110__11_,
  data_n_110__10_,data_n_110__9_,data_n_110__8_,data_n_110__7_,data_n_110__6_,
  data_n_110__5_,data_n_110__4_,data_n_110__3_,data_n_110__2_,data_n_110__1_,
  data_n_110__0_,data_n_109__31_,data_n_109__30_,data_n_109__29_,data_n_109__28_,
  data_n_109__27_,data_n_109__26_,data_n_109__25_,data_n_109__24_,data_n_109__23_,
  data_n_109__22_,data_n_109__21_,data_n_109__20_,data_n_109__19_,data_n_109__18_,
  data_n_109__17_,data_n_109__16_,data_n_109__15_,data_n_109__14_,data_n_109__13_,
  data_n_109__12_,data_n_109__11_,data_n_109__10_,data_n_109__9_,data_n_109__8_,data_n_109__7_,
  data_n_109__6_,data_n_109__5_,data_n_109__4_,data_n_109__3_,data_n_109__2_,
  data_n_109__1_,data_n_109__0_,data_n_108__31_,data_n_108__30_,data_n_108__29_,
  data_n_108__28_,data_n_108__27_,data_n_108__26_,data_n_108__25_,data_n_108__24_,
  data_n_108__23_,data_n_108__22_,data_n_108__21_,data_n_108__20_,data_n_108__19_,
  data_n_108__18_,data_n_108__17_,data_n_108__16_,data_n_108__15_,data_n_108__14_,
  data_n_108__13_,data_n_108__12_,data_n_108__11_,data_n_108__10_,data_n_108__9_,
  data_n_108__8_,data_n_108__7_,data_n_108__6_,data_n_108__5_,data_n_108__4_,
  data_n_108__3_,data_n_108__2_,data_n_108__1_,data_n_108__0_,data_n_107__31_,data_n_107__30_,
  data_n_107__29_,data_n_107__28_,data_n_107__27_,data_n_107__26_,data_n_107__25_,
  data_n_107__24_,data_n_107__23_,data_n_107__22_,data_n_107__21_,data_n_107__20_,
  data_n_107__19_,data_n_107__18_,data_n_107__17_,data_n_107__16_,data_n_107__15_,
  data_n_107__14_,data_n_107__13_,data_n_107__12_,data_n_107__11_,data_n_107__10_,
  data_n_107__9_,data_n_107__8_,data_n_107__7_,data_n_107__6_,data_n_107__5_,
  data_n_107__4_,data_n_107__3_,data_n_107__2_,data_n_107__1_,data_n_107__0_,
  data_n_106__31_,data_n_106__30_,data_n_106__29_,data_n_106__28_,data_n_106__27_,
  data_n_106__26_,data_n_106__25_,data_n_106__24_,data_n_106__23_,data_n_106__22_,
  data_n_106__21_,data_n_106__20_,data_n_106__19_,data_n_106__18_,data_n_106__17_,
  data_n_106__16_,data_n_106__15_,data_n_106__14_,data_n_106__13_,data_n_106__12_,
  data_n_106__11_,data_n_106__10_,data_n_106__9_,data_n_106__8_,data_n_106__7_,data_n_106__6_,
  data_n_106__5_,data_n_106__4_,data_n_106__3_,data_n_106__2_,data_n_106__1_,
  data_n_106__0_,data_n_105__31_,data_n_105__30_,data_n_105__29_,data_n_105__28_,
  data_n_105__27_,data_n_105__26_,data_n_105__25_,data_n_105__24_,data_n_105__23_,
  data_n_105__22_,data_n_105__21_,data_n_105__20_,data_n_105__19_,data_n_105__18_,
  data_n_105__17_,data_n_105__16_,data_n_105__15_,data_n_105__14_,data_n_105__13_,
  data_n_105__12_,data_n_105__11_,data_n_105__10_,data_n_105__9_,data_n_105__8_,
  data_n_105__7_,data_n_105__6_,data_n_105__5_,data_n_105__4_,data_n_105__3_,
  data_n_105__2_,data_n_105__1_,data_n_105__0_,data_n_104__31_,data_n_104__30_,data_n_104__29_,
  data_n_104__28_,data_n_104__27_,data_n_104__26_,data_n_104__25_,data_n_104__24_,
  data_n_104__23_,data_n_104__22_,data_n_104__21_,data_n_104__20_,data_n_104__19_,
  data_n_104__18_,data_n_104__17_,data_n_104__16_,data_n_104__15_,data_n_104__14_,
  data_n_104__13_,data_n_104__12_,data_n_104__11_,data_n_104__10_,data_n_104__9_,
  data_n_104__8_,data_n_104__7_,data_n_104__6_,data_n_104__5_,data_n_104__4_,
  data_n_104__3_,data_n_104__2_,data_n_104__1_,data_n_104__0_,data_n_103__31_,
  data_n_103__30_,data_n_103__29_,data_n_103__28_,data_n_103__27_,data_n_103__26_,
  data_n_103__25_,data_n_103__24_,data_n_103__23_,data_n_103__22_,data_n_103__21_,
  data_n_103__20_,data_n_103__19_,data_n_103__18_,data_n_103__17_,data_n_103__16_,
  data_n_103__15_,data_n_103__14_,data_n_103__13_,data_n_103__12_,data_n_103__11_,
  data_n_103__10_,data_n_103__9_,data_n_103__8_,data_n_103__7_,data_n_103__6_,
  data_n_103__5_,data_n_103__4_,data_n_103__3_,data_n_103__2_,data_n_103__1_,data_n_103__0_,
  data_n_102__31_,data_n_102__30_,data_n_102__29_,data_n_102__28_,data_n_102__27_,
  data_n_102__26_,data_n_102__25_,data_n_102__24_,data_n_102__23_,data_n_102__22_,
  data_n_102__21_,data_n_102__20_,data_n_102__19_,data_n_102__18_,data_n_102__17_,
  data_n_102__16_,data_n_102__15_,data_n_102__14_,data_n_102__13_,data_n_102__12_,
  data_n_102__11_,data_n_102__10_,data_n_102__9_,data_n_102__8_,data_n_102__7_,
  data_n_102__6_,data_n_102__5_,data_n_102__4_,data_n_102__3_,data_n_102__2_,
  data_n_102__1_,data_n_102__0_,data_n_101__31_,data_n_101__30_,data_n_101__29_,
  data_n_101__28_,data_n_101__27_,data_n_101__26_,data_n_101__25_,data_n_101__24_,
  data_n_101__23_,data_n_101__22_,data_n_101__21_,data_n_101__20_,data_n_101__19_,
  data_n_101__18_,data_n_101__17_,data_n_101__16_,data_n_101__15_,data_n_101__14_,
  data_n_101__13_,data_n_101__12_,data_n_101__11_,data_n_101__10_,data_n_101__9_,data_n_101__8_,
  data_n_101__7_,data_n_101__6_,data_n_101__5_,data_n_101__4_,data_n_101__3_,
  data_n_101__2_,data_n_101__1_,data_n_101__0_,data_n_100__31_,data_n_100__30_,
  data_n_100__29_,data_n_100__28_,data_n_100__27_,data_n_100__26_,data_n_100__25_,
  data_n_100__24_,data_n_100__23_,data_n_100__22_,data_n_100__21_,data_n_100__20_,
  data_n_100__19_,data_n_100__18_,data_n_100__17_,data_n_100__16_,data_n_100__15_,
  data_n_100__14_,data_n_100__13_,data_n_100__12_,data_n_100__11_,data_n_100__10_,
  data_n_100__9_,data_n_100__8_,data_n_100__7_,data_n_100__6_,data_n_100__5_,
  data_n_100__4_,data_n_100__3_,data_n_100__2_,data_n_100__1_,data_n_100__0_,data_n_99__31_,
  data_n_99__30_,data_n_99__29_,data_n_99__28_,data_n_99__27_,data_n_99__26_,
  data_n_99__25_,data_n_99__24_,data_n_99__23_,data_n_99__22_,data_n_99__21_,
  data_n_99__20_,data_n_99__19_,data_n_99__18_,data_n_99__17_,data_n_99__16_,data_n_99__15_,
  data_n_99__14_,data_n_99__13_,data_n_99__12_,data_n_99__11_,data_n_99__10_,
  data_n_99__9_,data_n_99__8_,data_n_99__7_,data_n_99__6_,data_n_99__5_,data_n_99__4_,
  data_n_99__3_,data_n_99__2_,data_n_99__1_,data_n_99__0_,data_n_98__31_,
  data_n_98__30_,data_n_98__29_,data_n_98__28_,data_n_98__27_,data_n_98__26_,data_n_98__25_,
  data_n_98__24_,data_n_98__23_,data_n_98__22_,data_n_98__21_,data_n_98__20_,
  data_n_98__19_,data_n_98__18_,data_n_98__17_,data_n_98__16_,data_n_98__15_,
  data_n_98__14_,data_n_98__13_,data_n_98__12_,data_n_98__11_,data_n_98__10_,data_n_98__9_,
  data_n_98__8_,data_n_98__7_,data_n_98__6_,data_n_98__5_,data_n_98__4_,data_n_98__3_,
  data_n_98__2_,data_n_98__1_,data_n_98__0_,data_n_97__31_,data_n_97__30_,
  data_n_97__29_,data_n_97__28_,data_n_97__27_,data_n_97__26_,data_n_97__25_,
  data_n_97__24_,data_n_97__23_,data_n_97__22_,data_n_97__21_,data_n_97__20_,data_n_97__19_,
  data_n_97__18_,data_n_97__17_,data_n_97__16_,data_n_97__15_,data_n_97__14_,
  data_n_97__13_,data_n_97__12_,data_n_97__11_,data_n_97__10_,data_n_97__9_,data_n_97__8_,
  data_n_97__7_,data_n_97__6_,data_n_97__5_,data_n_97__4_,data_n_97__3_,
  data_n_97__2_,data_n_97__1_,data_n_97__0_,data_n_96__31_,data_n_96__30_,data_n_96__29_,
  data_n_96__28_,data_n_96__27_,data_n_96__26_,data_n_96__25_,data_n_96__24_,
  data_n_96__23_,data_n_96__22_,data_n_96__21_,data_n_96__20_,data_n_96__19_,
  data_n_96__18_,data_n_96__17_,data_n_96__16_,data_n_96__15_,data_n_96__14_,data_n_96__13_,
  data_n_96__12_,data_n_96__11_,data_n_96__10_,data_n_96__9_,data_n_96__8_,
  data_n_96__7_,data_n_96__6_,data_n_96__5_,data_n_96__4_,data_n_96__3_,data_n_96__2_,
  data_n_96__1_,data_n_96__0_,data_n_95__31_,data_n_95__30_,data_n_95__29_,
  data_n_95__28_,data_n_95__27_,data_n_95__26_,data_n_95__25_,data_n_95__24_,data_n_95__23_,
  data_n_95__22_,data_n_95__21_,data_n_95__20_,data_n_95__19_,data_n_95__18_,
  data_n_95__17_,data_n_95__16_,data_n_95__15_,data_n_95__14_,data_n_95__13_,
  data_n_95__12_,data_n_95__11_,data_n_95__10_,data_n_95__9_,data_n_95__8_,data_n_95__7_,
  data_n_95__6_,data_n_95__5_,data_n_95__4_,data_n_95__3_,data_n_95__2_,data_n_95__1_,
  data_n_95__0_,data_n_94__31_,data_n_94__30_,data_n_94__29_,data_n_94__28_,
  data_n_94__27_,data_n_94__26_,data_n_94__25_,data_n_94__24_,data_n_94__23_,
  data_n_94__22_,data_n_94__21_,data_n_94__20_,data_n_94__19_,data_n_94__18_,data_n_94__17_,
  data_n_94__16_,data_n_94__15_,data_n_94__14_,data_n_94__13_,data_n_94__12_,
  data_n_94__11_,data_n_94__10_,data_n_94__9_,data_n_94__8_,data_n_94__7_,data_n_94__6_,
  data_n_94__5_,data_n_94__4_,data_n_94__3_,data_n_94__2_,data_n_94__1_,
  data_n_94__0_,data_n_93__31_,data_n_93__30_,data_n_93__29_,data_n_93__28_,data_n_93__27_,
  data_n_93__26_,data_n_93__25_,data_n_93__24_,data_n_93__23_,data_n_93__22_,
  data_n_93__21_,data_n_93__20_,data_n_93__19_,data_n_93__18_,data_n_93__17_,
  data_n_93__16_,data_n_93__15_,data_n_93__14_,data_n_93__13_,data_n_93__12_,data_n_93__11_,
  data_n_93__10_,data_n_93__9_,data_n_93__8_,data_n_93__7_,data_n_93__6_,
  data_n_93__5_,data_n_93__4_,data_n_93__3_,data_n_93__2_,data_n_93__1_,data_n_93__0_,
  data_n_92__31_,data_n_92__30_,data_n_92__29_,data_n_92__28_,data_n_92__27_,
  data_n_92__26_,data_n_92__25_,data_n_92__24_,data_n_92__23_,data_n_92__22_,data_n_92__21_,
  data_n_92__20_,data_n_92__19_,data_n_92__18_,data_n_92__17_,data_n_92__16_,
  data_n_92__15_,data_n_92__14_,data_n_92__13_,data_n_92__12_,data_n_92__11_,
  data_n_92__10_,data_n_92__9_,data_n_92__8_,data_n_92__7_,data_n_92__6_,data_n_92__5_,
  data_n_92__4_,data_n_92__3_,data_n_92__2_,data_n_92__1_,data_n_92__0_,data_n_91__31_,
  data_n_91__30_,data_n_91__29_,data_n_91__28_,data_n_91__27_,data_n_91__26_,
  data_n_91__25_,data_n_91__24_,data_n_91__23_,data_n_91__22_,data_n_91__21_,
  data_n_91__20_,data_n_91__19_,data_n_91__18_,data_n_91__17_,data_n_91__16_,data_n_91__15_,
  data_n_91__14_,data_n_91__13_,data_n_91__12_,data_n_91__11_,data_n_91__10_,
  data_n_91__9_,data_n_91__8_,data_n_91__7_,data_n_91__6_,data_n_91__5_,data_n_91__4_,
  data_n_91__3_,data_n_91__2_,data_n_91__1_,data_n_91__0_,data_n_90__31_,
  data_n_90__30_,data_n_90__29_,data_n_90__28_,data_n_90__27_,data_n_90__26_,data_n_90__25_,
  data_n_90__24_,data_n_90__23_,data_n_90__22_,data_n_90__21_,data_n_90__20_,
  data_n_90__19_,data_n_90__18_,data_n_90__17_,data_n_90__16_,data_n_90__15_,
  data_n_90__14_,data_n_90__13_,data_n_90__12_,data_n_90__11_,data_n_90__10_,data_n_90__9_,
  data_n_90__8_,data_n_90__7_,data_n_90__6_,data_n_90__5_,data_n_90__4_,data_n_90__3_,
  data_n_90__2_,data_n_90__1_,data_n_90__0_,data_n_89__31_,data_n_89__30_,
  data_n_89__29_,data_n_89__28_,data_n_89__27_,data_n_89__26_,data_n_89__25_,
  data_n_89__24_,data_n_89__23_,data_n_89__22_,data_n_89__21_,data_n_89__20_,data_n_89__19_,
  data_n_89__18_,data_n_89__17_,data_n_89__16_,data_n_89__15_,data_n_89__14_,
  data_n_89__13_,data_n_89__12_,data_n_89__11_,data_n_89__10_,data_n_89__9_,data_n_89__8_,
  data_n_89__7_,data_n_89__6_,data_n_89__5_,data_n_89__4_,data_n_89__3_,
  data_n_89__2_,data_n_89__1_,data_n_89__0_,data_n_88__31_,data_n_88__30_,data_n_88__29_,
  data_n_88__28_,data_n_88__27_,data_n_88__26_,data_n_88__25_,data_n_88__24_,
  data_n_88__23_,data_n_88__22_,data_n_88__21_,data_n_88__20_,data_n_88__19_,
  data_n_88__18_,data_n_88__17_,data_n_88__16_,data_n_88__15_,data_n_88__14_,data_n_88__13_,
  data_n_88__12_,data_n_88__11_,data_n_88__10_,data_n_88__9_,data_n_88__8_,
  data_n_88__7_,data_n_88__6_,data_n_88__5_,data_n_88__4_,data_n_88__3_,data_n_88__2_,
  data_n_88__1_,data_n_88__0_,data_n_87__31_,data_n_87__30_,data_n_87__29_,
  data_n_87__28_,data_n_87__27_,data_n_87__26_,data_n_87__25_,data_n_87__24_,data_n_87__23_,
  data_n_87__22_,data_n_87__21_,data_n_87__20_,data_n_87__19_,data_n_87__18_,
  data_n_87__17_,data_n_87__16_,data_n_87__15_,data_n_87__14_,data_n_87__13_,
  data_n_87__12_,data_n_87__11_,data_n_87__10_,data_n_87__9_,data_n_87__8_,data_n_87__7_,
  data_n_87__6_,data_n_87__5_,data_n_87__4_,data_n_87__3_,data_n_87__2_,data_n_87__1_,
  data_n_87__0_,data_n_86__31_,data_n_86__30_,data_n_86__29_,data_n_86__28_,
  data_n_86__27_,data_n_86__26_,data_n_86__25_,data_n_86__24_,data_n_86__23_,
  data_n_86__22_,data_n_86__21_,data_n_86__20_,data_n_86__19_,data_n_86__18_,data_n_86__17_,
  data_n_86__16_,data_n_86__15_,data_n_86__14_,data_n_86__13_,data_n_86__12_,
  data_n_86__11_,data_n_86__10_,data_n_86__9_,data_n_86__8_,data_n_86__7_,data_n_86__6_,
  data_n_86__5_,data_n_86__4_,data_n_86__3_,data_n_86__2_,data_n_86__1_,
  data_n_86__0_,data_n_85__31_,data_n_85__30_,data_n_85__29_,data_n_85__28_,data_n_85__27_,
  data_n_85__26_,data_n_85__25_,data_n_85__24_,data_n_85__23_,data_n_85__22_,
  data_n_85__21_,data_n_85__20_,data_n_85__19_,data_n_85__18_,data_n_85__17_,
  data_n_85__16_,data_n_85__15_,data_n_85__14_,data_n_85__13_,data_n_85__12_,data_n_85__11_,
  data_n_85__10_,data_n_85__9_,data_n_85__8_,data_n_85__7_,data_n_85__6_,
  data_n_85__5_,data_n_85__4_,data_n_85__3_,data_n_85__2_,data_n_85__1_,data_n_85__0_,
  data_n_84__31_,data_n_84__30_,data_n_84__29_,data_n_84__28_,data_n_84__27_,
  data_n_84__26_,data_n_84__25_,data_n_84__24_,data_n_84__23_,data_n_84__22_,data_n_84__21_,
  data_n_84__20_,data_n_84__19_,data_n_84__18_,data_n_84__17_,data_n_84__16_,
  data_n_84__15_,data_n_84__14_,data_n_84__13_,data_n_84__12_,data_n_84__11_,
  data_n_84__10_,data_n_84__9_,data_n_84__8_,data_n_84__7_,data_n_84__6_,data_n_84__5_,
  data_n_84__4_,data_n_84__3_,data_n_84__2_,data_n_84__1_,data_n_84__0_,data_n_83__31_,
  data_n_83__30_,data_n_83__29_,data_n_83__28_,data_n_83__27_,data_n_83__26_,
  data_n_83__25_,data_n_83__24_,data_n_83__23_,data_n_83__22_,data_n_83__21_,
  data_n_83__20_,data_n_83__19_,data_n_83__18_,data_n_83__17_,data_n_83__16_,data_n_83__15_,
  data_n_83__14_,data_n_83__13_,data_n_83__12_,data_n_83__11_,data_n_83__10_,
  data_n_83__9_,data_n_83__8_,data_n_83__7_,data_n_83__6_,data_n_83__5_,data_n_83__4_,
  data_n_83__3_,data_n_83__2_,data_n_83__1_,data_n_83__0_,data_n_82__31_,
  data_n_82__30_,data_n_82__29_,data_n_82__28_,data_n_82__27_,data_n_82__26_,data_n_82__25_,
  data_n_82__24_,data_n_82__23_,data_n_82__22_,data_n_82__21_,data_n_82__20_,
  data_n_82__19_,data_n_82__18_,data_n_82__17_,data_n_82__16_,data_n_82__15_,
  data_n_82__14_,data_n_82__13_,data_n_82__12_,data_n_82__11_,data_n_82__10_,data_n_82__9_,
  data_n_82__8_,data_n_82__7_,data_n_82__6_,data_n_82__5_,data_n_82__4_,data_n_82__3_,
  data_n_82__2_,data_n_82__1_,data_n_82__0_,data_n_81__31_,data_n_81__30_,
  data_n_81__29_,data_n_81__28_,data_n_81__27_,data_n_81__26_,data_n_81__25_,
  data_n_81__24_,data_n_81__23_,data_n_81__22_,data_n_81__21_,data_n_81__20_,data_n_81__19_,
  data_n_81__18_,data_n_81__17_,data_n_81__16_,data_n_81__15_,data_n_81__14_,
  data_n_81__13_,data_n_81__12_,data_n_81__11_,data_n_81__10_,data_n_81__9_,data_n_81__8_,
  data_n_81__7_,data_n_81__6_,data_n_81__5_,data_n_81__4_,data_n_81__3_,
  data_n_81__2_,data_n_81__1_,data_n_81__0_,data_n_80__31_,data_n_80__30_,data_n_80__29_,
  data_n_80__28_,data_n_80__27_,data_n_80__26_,data_n_80__25_,data_n_80__24_,
  data_n_80__23_,data_n_80__22_,data_n_80__21_,data_n_80__20_,data_n_80__19_,
  data_n_80__18_,data_n_80__17_,data_n_80__16_,data_n_80__15_,data_n_80__14_,data_n_80__13_,
  data_n_80__12_,data_n_80__11_,data_n_80__10_,data_n_80__9_,data_n_80__8_,
  data_n_80__7_,data_n_80__6_,data_n_80__5_,data_n_80__4_,data_n_80__3_,data_n_80__2_,
  data_n_80__1_,data_n_80__0_,data_n_79__31_,data_n_79__30_,data_n_79__29_,
  data_n_79__28_,data_n_79__27_,data_n_79__26_,data_n_79__25_,data_n_79__24_,data_n_79__23_,
  data_n_79__22_,data_n_79__21_,data_n_79__20_,data_n_79__19_,data_n_79__18_,
  data_n_79__17_,data_n_79__16_,data_n_79__15_,data_n_79__14_,data_n_79__13_,
  data_n_79__12_,data_n_79__11_,data_n_79__10_,data_n_79__9_,data_n_79__8_,data_n_79__7_,
  data_n_79__6_,data_n_79__5_,data_n_79__4_,data_n_79__3_,data_n_79__2_,data_n_79__1_,
  data_n_79__0_,data_n_78__31_,data_n_78__30_,data_n_78__29_,data_n_78__28_,
  data_n_78__27_,data_n_78__26_,data_n_78__25_,data_n_78__24_,data_n_78__23_,
  data_n_78__22_,data_n_78__21_,data_n_78__20_,data_n_78__19_,data_n_78__18_,data_n_78__17_,
  data_n_78__16_,data_n_78__15_,data_n_78__14_,data_n_78__13_,data_n_78__12_,
  data_n_78__11_,data_n_78__10_,data_n_78__9_,data_n_78__8_,data_n_78__7_,data_n_78__6_,
  data_n_78__5_,data_n_78__4_,data_n_78__3_,data_n_78__2_,data_n_78__1_,
  data_n_78__0_,data_n_77__31_,data_n_77__30_,data_n_77__29_,data_n_77__28_,data_n_77__27_,
  data_n_77__26_,data_n_77__25_,data_n_77__24_,data_n_77__23_,data_n_77__22_,
  data_n_77__21_,data_n_77__20_,data_n_77__19_,data_n_77__18_,data_n_77__17_,
  data_n_77__16_,data_n_77__15_,data_n_77__14_,data_n_77__13_,data_n_77__12_,data_n_77__11_,
  data_n_77__10_,data_n_77__9_,data_n_77__8_,data_n_77__7_,data_n_77__6_,
  data_n_77__5_,data_n_77__4_,data_n_77__3_,data_n_77__2_,data_n_77__1_,data_n_77__0_,
  data_n_76__31_,data_n_76__30_,data_n_76__29_,data_n_76__28_,data_n_76__27_,
  data_n_76__26_,data_n_76__25_,data_n_76__24_,data_n_76__23_,data_n_76__22_,data_n_76__21_,
  data_n_76__20_,data_n_76__19_,data_n_76__18_,data_n_76__17_,data_n_76__16_,
  data_n_76__15_,data_n_76__14_,data_n_76__13_,data_n_76__12_,data_n_76__11_,
  data_n_76__10_,data_n_76__9_,data_n_76__8_,data_n_76__7_,data_n_76__6_,data_n_76__5_,
  data_n_76__4_,data_n_76__3_,data_n_76__2_,data_n_76__1_,data_n_76__0_,data_n_75__31_,
  data_n_75__30_,data_n_75__29_,data_n_75__28_,data_n_75__27_,data_n_75__26_,
  data_n_75__25_,data_n_75__24_,data_n_75__23_,data_n_75__22_,data_n_75__21_,
  data_n_75__20_,data_n_75__19_,data_n_75__18_,data_n_75__17_,data_n_75__16_,data_n_75__15_,
  data_n_75__14_,data_n_75__13_,data_n_75__12_,data_n_75__11_,data_n_75__10_,
  data_n_75__9_,data_n_75__8_,data_n_75__7_,data_n_75__6_,data_n_75__5_,data_n_75__4_,
  data_n_75__3_,data_n_75__2_,data_n_75__1_,data_n_75__0_,data_n_74__31_,
  data_n_74__30_,data_n_74__29_,data_n_74__28_,data_n_74__27_,data_n_74__26_,data_n_74__25_,
  data_n_74__24_,data_n_74__23_,data_n_74__22_,data_n_74__21_,data_n_74__20_,
  data_n_74__19_,data_n_74__18_,data_n_74__17_,data_n_74__16_,data_n_74__15_,
  data_n_74__14_,data_n_74__13_,data_n_74__12_,data_n_74__11_,data_n_74__10_,data_n_74__9_,
  data_n_74__8_,data_n_74__7_,data_n_74__6_,data_n_74__5_,data_n_74__4_,data_n_74__3_,
  data_n_74__2_,data_n_74__1_,data_n_74__0_,data_n_73__31_,data_n_73__30_,
  data_n_73__29_,data_n_73__28_,data_n_73__27_,data_n_73__26_,data_n_73__25_,
  data_n_73__24_,data_n_73__23_,data_n_73__22_,data_n_73__21_,data_n_73__20_,data_n_73__19_,
  data_n_73__18_,data_n_73__17_,data_n_73__16_,data_n_73__15_,data_n_73__14_,
  data_n_73__13_,data_n_73__12_,data_n_73__11_,data_n_73__10_,data_n_73__9_,data_n_73__8_,
  data_n_73__7_,data_n_73__6_,data_n_73__5_,data_n_73__4_,data_n_73__3_,
  data_n_73__2_,data_n_73__1_,data_n_73__0_,data_n_72__31_,data_n_72__30_,data_n_72__29_,
  data_n_72__28_,data_n_72__27_,data_n_72__26_,data_n_72__25_,data_n_72__24_,
  data_n_72__23_,data_n_72__22_,data_n_72__21_,data_n_72__20_,data_n_72__19_,
  data_n_72__18_,data_n_72__17_,data_n_72__16_,data_n_72__15_,data_n_72__14_,data_n_72__13_,
  data_n_72__12_,data_n_72__11_,data_n_72__10_,data_n_72__9_,data_n_72__8_,
  data_n_72__7_,data_n_72__6_,data_n_72__5_,data_n_72__4_,data_n_72__3_,data_n_72__2_,
  data_n_72__1_,data_n_72__0_,data_n_71__31_,data_n_71__30_,data_n_71__29_,
  data_n_71__28_,data_n_71__27_,data_n_71__26_,data_n_71__25_,data_n_71__24_,data_n_71__23_,
  data_n_71__22_,data_n_71__21_,data_n_71__20_,data_n_71__19_,data_n_71__18_,
  data_n_71__17_,data_n_71__16_,data_n_71__15_,data_n_71__14_,data_n_71__13_,
  data_n_71__12_,data_n_71__11_,data_n_71__10_,data_n_71__9_,data_n_71__8_,data_n_71__7_,
  data_n_71__6_,data_n_71__5_,data_n_71__4_,data_n_71__3_,data_n_71__2_,data_n_71__1_,
  data_n_71__0_,data_n_70__31_,data_n_70__30_,data_n_70__29_,data_n_70__28_,
  data_n_70__27_,data_n_70__26_,data_n_70__25_,data_n_70__24_,data_n_70__23_,
  data_n_70__22_,data_n_70__21_,data_n_70__20_,data_n_70__19_,data_n_70__18_,data_n_70__17_,
  data_n_70__16_,data_n_70__15_,data_n_70__14_,data_n_70__13_,data_n_70__12_,
  data_n_70__11_,data_n_70__10_,data_n_70__9_,data_n_70__8_,data_n_70__7_,data_n_70__6_,
  data_n_70__5_,data_n_70__4_,data_n_70__3_,data_n_70__2_,data_n_70__1_,
  data_n_70__0_,data_n_69__31_,data_n_69__30_,data_n_69__29_,data_n_69__28_,data_n_69__27_,
  data_n_69__26_,data_n_69__25_,data_n_69__24_,data_n_69__23_,data_n_69__22_,
  data_n_69__21_,data_n_69__20_,data_n_69__19_,data_n_69__18_,data_n_69__17_,
  data_n_69__16_,data_n_69__15_,data_n_69__14_,data_n_69__13_,data_n_69__12_,data_n_69__11_,
  data_n_69__10_,data_n_69__9_,data_n_69__8_,data_n_69__7_,data_n_69__6_,
  data_n_69__5_,data_n_69__4_,data_n_69__3_,data_n_69__2_,data_n_69__1_,data_n_69__0_,
  data_n_68__31_,data_n_68__30_,data_n_68__29_,data_n_68__28_,data_n_68__27_,
  data_n_68__26_,data_n_68__25_,data_n_68__24_,data_n_68__23_,data_n_68__22_,data_n_68__21_,
  data_n_68__20_,data_n_68__19_,data_n_68__18_,data_n_68__17_,data_n_68__16_,
  data_n_68__15_,data_n_68__14_,data_n_68__13_,data_n_68__12_,data_n_68__11_,
  data_n_68__10_,data_n_68__9_,data_n_68__8_,data_n_68__7_,data_n_68__6_,data_n_68__5_,
  data_n_68__4_,data_n_68__3_,data_n_68__2_,data_n_68__1_,data_n_68__0_,data_n_67__31_,
  data_n_67__30_,data_n_67__29_,data_n_67__28_,data_n_67__27_,data_n_67__26_,
  data_n_67__25_,data_n_67__24_,data_n_67__23_,data_n_67__22_,data_n_67__21_,
  data_n_67__20_,data_n_67__19_,data_n_67__18_,data_n_67__17_,data_n_67__16_,data_n_67__15_,
  data_n_67__14_,data_n_67__13_,data_n_67__12_,data_n_67__11_,data_n_67__10_,
  data_n_67__9_,data_n_67__8_,data_n_67__7_,data_n_67__6_,data_n_67__5_,data_n_67__4_,
  data_n_67__3_,data_n_67__2_,data_n_67__1_,data_n_67__0_,data_n_66__31_,
  data_n_66__30_,data_n_66__29_,data_n_66__28_,data_n_66__27_,data_n_66__26_,data_n_66__25_,
  data_n_66__24_,data_n_66__23_,data_n_66__22_,data_n_66__21_,data_n_66__20_,
  data_n_66__19_,data_n_66__18_,data_n_66__17_,data_n_66__16_,data_n_66__15_,
  data_n_66__14_,data_n_66__13_,data_n_66__12_,data_n_66__11_,data_n_66__10_,data_n_66__9_,
  data_n_66__8_,data_n_66__7_,data_n_66__6_,data_n_66__5_,data_n_66__4_,data_n_66__3_,
  data_n_66__2_,data_n_66__1_,data_n_66__0_,data_n_65__31_,data_n_65__30_,
  data_n_65__29_,data_n_65__28_,data_n_65__27_,data_n_65__26_,data_n_65__25_,
  data_n_65__24_,data_n_65__23_,data_n_65__22_,data_n_65__21_,data_n_65__20_,data_n_65__19_,
  data_n_65__18_,data_n_65__17_,data_n_65__16_,data_n_65__15_,data_n_65__14_,
  data_n_65__13_,data_n_65__12_,data_n_65__11_,data_n_65__10_,data_n_65__9_,data_n_65__8_,
  data_n_65__7_,data_n_65__6_,data_n_65__5_,data_n_65__4_,data_n_65__3_,
  data_n_65__2_,data_n_65__1_,data_n_65__0_,data_n_64__31_,data_n_64__30_,data_n_64__29_,
  data_n_64__28_,data_n_64__27_,data_n_64__26_,data_n_64__25_,data_n_64__24_,
  data_n_64__23_,data_n_64__22_,data_n_64__21_,data_n_64__20_,data_n_64__19_,
  data_n_64__18_,data_n_64__17_,data_n_64__16_,data_n_64__15_,data_n_64__14_,data_n_64__13_,
  data_n_64__12_,data_n_64__11_,data_n_64__10_,data_n_64__9_,data_n_64__8_,
  data_n_64__7_,data_n_64__6_,data_n_64__5_,data_n_64__4_,data_n_64__3_,data_n_64__2_,
  data_n_64__1_,data_n_64__0_,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,
  N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,
  N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,
  N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,
  N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,
  N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,
  N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,
  N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,
  N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,
  N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
  N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,
  N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,
  N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,
  N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,
  N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,
  N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,
  N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,
  N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,
  N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,
  N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,
  N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,
  N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,
  N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,
  N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,
  N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,
  N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,
  N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,
  N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,
  N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,
  N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,
  N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,
  N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,
  N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,
  N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,
  N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,
  N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,
  N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,
  N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,
  N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,
  N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,
  N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,
  N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,
  N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,
  N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,
  N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,
  N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,
  N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,
  N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,
  N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,
  N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
  N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,
  N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,
  N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,
  N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,
  N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,
  N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,
  N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,
  N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,
  N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,
  N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,
  N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,
  N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,
  N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,
  N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,
  N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,
  N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,
  N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,
  N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,
  N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,
  N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,
  N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,
  N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,
  N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,
  N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,
  N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,
  N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,
  N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,
  N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,
  N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,
  N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,
  N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,
  N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,
  N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,
  N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,
  N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,
  N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,
  N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,
  N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,
  N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,
  N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,
  N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,
  N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,
  N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,
  N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,
  N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,
  N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,
  N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,
  N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,
  N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,
  N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,
  N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,
  N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,
  N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,
  N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,
  N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,
  N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,
  N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,
  N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,
  N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,
  N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,
  N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,
  N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,
  N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,
  N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,
  N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,
  N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,
  N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,
  N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,
  N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,
  N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,
  N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,
  N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,
  N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,
  N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,
  N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,
  N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,
  N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,
  N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,
  N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,
  N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,
  N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,
  N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,
  N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,
  N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,
  N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,
  N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,
  N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,
  N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,
  N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,
  N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,
  N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,
  N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,
  N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,
  N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,
  N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,
  N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,
  N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,
  N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,
  N4207,N4208,N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,
  N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,
  N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,
  N4247,N4248,N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,
  N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,
  N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,
  N4287,N4288,N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,
  N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,
  N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,
  N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,
  N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,
  N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,
  N4367,N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,
  N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,
  N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,
  N4407,N4408,N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,
  N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,
  N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,
  N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,
  N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,
  N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,
  N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,
  N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,
  N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,
  N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,
  N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,
  N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,
  N4567,N4568,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,
  N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,
  N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,
  N4607,N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,
  N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,
  N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,
  N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,
  N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,
  N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,
  N4687,N4688,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,
  N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,
  N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,
  N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,
  N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,
  N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,
  N4767,N4768,N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,
  N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,
  N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,
  N4807,N4808,N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,
  N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,
  N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,
  N4847,N4848,N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,
  N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,
  N4874,N4875,N4876,N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,
  N4887,N4888,N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,N4900,
  N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,
  N4914,N4915,N4916,N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,
  N4927,N4928,N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,
  N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,
  N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,
  N4967,N4968,N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,
  N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,
  N4994,N4995,N4996,N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,
  N5007,N5008,N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,
  N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,
  N5034,N5035,N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,
  N5047,N5048,N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,
  N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,
  N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,
  N5087,N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,
  N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,
  N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,
  N5127,N5128,N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,
  N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,
  N5154,N5155,N5156,N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,
  N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,
  N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,
  N5194,N5195,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,
  N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,
  N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,
  N5234,N5235,N5236,N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,
  N5247,N5248,N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,
  N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,
  N5274,N5275,N5276,N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,
  N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,
  N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,
  N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,
  N5327,N5328,N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,
  N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,
  N5354,N5355,N5356,N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,
  N5367,N5368,N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,
  N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,
  N5394,N5395,N5396,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,
  N5407,N5408,N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,
  N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,
  N5434,N5435,N5436,N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,
  N5447,N5448,N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,
  N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,
  N5474,N5475,N5476,N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,
  N5487,N5488,N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,
  N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,
  N5514,N5515,N5516,N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,
  N5527,N5528,N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,
  N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,
  N5554,N5555,N5556,N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,
  N5567,N5568,N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,
  N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,
  N5594,N5595,N5596,N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,
  N5607,N5608,N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,
  N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,
  N5634,N5635,N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,
  N5647,N5648,N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,
  N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,
  N5674,N5675,N5676,N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,
  N5687,N5688,N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,
  N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,
  N5714,N5715,N5716,N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,
  N5727,N5728,N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,
  N5741,N5742,N5743;
  wire [6:0] num_els_r,num_els_n;
  wire [127:64] valid_n;
  reg valid_r_63_sv2v_reg,valid_r_62_sv2v_reg,valid_r_61_sv2v_reg,valid_r_60_sv2v_reg,
  valid_r_59_sv2v_reg,valid_r_58_sv2v_reg,valid_r_57_sv2v_reg,valid_r_56_sv2v_reg,
  valid_r_55_sv2v_reg,valid_r_54_sv2v_reg,valid_r_53_sv2v_reg,valid_r_52_sv2v_reg,
  valid_r_51_sv2v_reg,valid_r_50_sv2v_reg,valid_r_49_sv2v_reg,valid_r_48_sv2v_reg,
  valid_r_47_sv2v_reg,valid_r_46_sv2v_reg,valid_r_45_sv2v_reg,valid_r_44_sv2v_reg,
  valid_r_43_sv2v_reg,valid_r_42_sv2v_reg,valid_r_41_sv2v_reg,valid_r_40_sv2v_reg,
  valid_r_39_sv2v_reg,valid_r_38_sv2v_reg,valid_r_37_sv2v_reg,valid_r_36_sv2v_reg,
  valid_r_35_sv2v_reg,valid_r_34_sv2v_reg,valid_r_33_sv2v_reg,valid_r_32_sv2v_reg,
  valid_r_31_sv2v_reg,valid_r_30_sv2v_reg,valid_r_29_sv2v_reg,valid_r_28_sv2v_reg,
  valid_r_27_sv2v_reg,valid_r_26_sv2v_reg,valid_r_25_sv2v_reg,valid_r_24_sv2v_reg,
  valid_r_23_sv2v_reg,valid_r_22_sv2v_reg,valid_r_21_sv2v_reg,valid_r_20_sv2v_reg,
  valid_r_19_sv2v_reg,valid_r_18_sv2v_reg,valid_r_17_sv2v_reg,valid_r_16_sv2v_reg,
  valid_r_15_sv2v_reg,valid_r_14_sv2v_reg,valid_r_13_sv2v_reg,valid_r_12_sv2v_reg,
  valid_r_11_sv2v_reg,valid_r_10_sv2v_reg,valid_r_9_sv2v_reg,valid_r_8_sv2v_reg,
  valid_r_7_sv2v_reg,valid_r_6_sv2v_reg,valid_r_5_sv2v_reg,valid_r_4_sv2v_reg,
  valid_r_3_sv2v_reg,valid_r_2_sv2v_reg,valid_r_1_sv2v_reg,valid_r_0_sv2v_reg,
  num_els_r_6_sv2v_reg,num_els_r_5_sv2v_reg,num_els_r_4_sv2v_reg,num_els_r_3_sv2v_reg,
  num_els_r_2_sv2v_reg,num_els_r_1_sv2v_reg,num_els_r_0_sv2v_reg,data_r_2047_sv2v_reg,
  data_r_2046_sv2v_reg,data_r_2045_sv2v_reg,data_r_2044_sv2v_reg,
  data_r_2043_sv2v_reg,data_r_2042_sv2v_reg,data_r_2041_sv2v_reg,data_r_2040_sv2v_reg,
  data_r_2039_sv2v_reg,data_r_2038_sv2v_reg,data_r_2037_sv2v_reg,data_r_2036_sv2v_reg,
  data_r_2035_sv2v_reg,data_r_2034_sv2v_reg,data_r_2033_sv2v_reg,data_r_2032_sv2v_reg,
  data_r_2031_sv2v_reg,data_r_2030_sv2v_reg,data_r_2029_sv2v_reg,data_r_2028_sv2v_reg,
  data_r_2027_sv2v_reg,data_r_2026_sv2v_reg,data_r_2025_sv2v_reg,
  data_r_2024_sv2v_reg,data_r_2023_sv2v_reg,data_r_2022_sv2v_reg,data_r_2021_sv2v_reg,
  data_r_2020_sv2v_reg,data_r_2019_sv2v_reg,data_r_2018_sv2v_reg,data_r_2017_sv2v_reg,
  data_r_2016_sv2v_reg,data_r_2015_sv2v_reg,data_r_2014_sv2v_reg,data_r_2013_sv2v_reg,
  data_r_2012_sv2v_reg,data_r_2011_sv2v_reg,data_r_2010_sv2v_reg,data_r_2009_sv2v_reg,
  data_r_2008_sv2v_reg,data_r_2007_sv2v_reg,data_r_2006_sv2v_reg,data_r_2005_sv2v_reg,
  data_r_2004_sv2v_reg,data_r_2003_sv2v_reg,data_r_2002_sv2v_reg,
  data_r_2001_sv2v_reg,data_r_2000_sv2v_reg,data_r_1999_sv2v_reg,data_r_1998_sv2v_reg,
  data_r_1997_sv2v_reg,data_r_1996_sv2v_reg,data_r_1995_sv2v_reg,data_r_1994_sv2v_reg,
  data_r_1993_sv2v_reg,data_r_1992_sv2v_reg,data_r_1991_sv2v_reg,data_r_1990_sv2v_reg,
  data_r_1989_sv2v_reg,data_r_1988_sv2v_reg,data_r_1987_sv2v_reg,data_r_1986_sv2v_reg,
  data_r_1985_sv2v_reg,data_r_1984_sv2v_reg,data_r_1983_sv2v_reg,
  data_r_1982_sv2v_reg,data_r_1981_sv2v_reg,data_r_1980_sv2v_reg,data_r_1979_sv2v_reg,
  data_r_1978_sv2v_reg,data_r_1977_sv2v_reg,data_r_1976_sv2v_reg,data_r_1975_sv2v_reg,
  data_r_1974_sv2v_reg,data_r_1973_sv2v_reg,data_r_1972_sv2v_reg,data_r_1971_sv2v_reg,
  data_r_1970_sv2v_reg,data_r_1969_sv2v_reg,data_r_1968_sv2v_reg,data_r_1967_sv2v_reg,
  data_r_1966_sv2v_reg,data_r_1965_sv2v_reg,data_r_1964_sv2v_reg,
  data_r_1963_sv2v_reg,data_r_1962_sv2v_reg,data_r_1961_sv2v_reg,data_r_1960_sv2v_reg,
  data_r_1959_sv2v_reg,data_r_1958_sv2v_reg,data_r_1957_sv2v_reg,data_r_1956_sv2v_reg,
  data_r_1955_sv2v_reg,data_r_1954_sv2v_reg,data_r_1953_sv2v_reg,data_r_1952_sv2v_reg,
  data_r_1951_sv2v_reg,data_r_1950_sv2v_reg,data_r_1949_sv2v_reg,data_r_1948_sv2v_reg,
  data_r_1947_sv2v_reg,data_r_1946_sv2v_reg,data_r_1945_sv2v_reg,
  data_r_1944_sv2v_reg,data_r_1943_sv2v_reg,data_r_1942_sv2v_reg,data_r_1941_sv2v_reg,
  data_r_1940_sv2v_reg,data_r_1939_sv2v_reg,data_r_1938_sv2v_reg,data_r_1937_sv2v_reg,
  data_r_1936_sv2v_reg,data_r_1935_sv2v_reg,data_r_1934_sv2v_reg,data_r_1933_sv2v_reg,
  data_r_1932_sv2v_reg,data_r_1931_sv2v_reg,data_r_1930_sv2v_reg,data_r_1929_sv2v_reg,
  data_r_1928_sv2v_reg,data_r_1927_sv2v_reg,data_r_1926_sv2v_reg,data_r_1925_sv2v_reg,
  data_r_1924_sv2v_reg,data_r_1923_sv2v_reg,data_r_1922_sv2v_reg,
  data_r_1921_sv2v_reg,data_r_1920_sv2v_reg,data_r_1919_sv2v_reg,data_r_1918_sv2v_reg,
  data_r_1917_sv2v_reg,data_r_1916_sv2v_reg,data_r_1915_sv2v_reg,data_r_1914_sv2v_reg,
  data_r_1913_sv2v_reg,data_r_1912_sv2v_reg,data_r_1911_sv2v_reg,data_r_1910_sv2v_reg,
  data_r_1909_sv2v_reg,data_r_1908_sv2v_reg,data_r_1907_sv2v_reg,data_r_1906_sv2v_reg,
  data_r_1905_sv2v_reg,data_r_1904_sv2v_reg,data_r_1903_sv2v_reg,
  data_r_1902_sv2v_reg,data_r_1901_sv2v_reg,data_r_1900_sv2v_reg,data_r_1899_sv2v_reg,
  data_r_1898_sv2v_reg,data_r_1897_sv2v_reg,data_r_1896_sv2v_reg,data_r_1895_sv2v_reg,
  data_r_1894_sv2v_reg,data_r_1893_sv2v_reg,data_r_1892_sv2v_reg,data_r_1891_sv2v_reg,
  data_r_1890_sv2v_reg,data_r_1889_sv2v_reg,data_r_1888_sv2v_reg,data_r_1887_sv2v_reg,
  data_r_1886_sv2v_reg,data_r_1885_sv2v_reg,data_r_1884_sv2v_reg,
  data_r_1883_sv2v_reg,data_r_1882_sv2v_reg,data_r_1881_sv2v_reg,data_r_1880_sv2v_reg,
  data_r_1879_sv2v_reg,data_r_1878_sv2v_reg,data_r_1877_sv2v_reg,data_r_1876_sv2v_reg,
  data_r_1875_sv2v_reg,data_r_1874_sv2v_reg,data_r_1873_sv2v_reg,data_r_1872_sv2v_reg,
  data_r_1871_sv2v_reg,data_r_1870_sv2v_reg,data_r_1869_sv2v_reg,data_r_1868_sv2v_reg,
  data_r_1867_sv2v_reg,data_r_1866_sv2v_reg,data_r_1865_sv2v_reg,
  data_r_1864_sv2v_reg,data_r_1863_sv2v_reg,data_r_1862_sv2v_reg,data_r_1861_sv2v_reg,
  data_r_1860_sv2v_reg,data_r_1859_sv2v_reg,data_r_1858_sv2v_reg,data_r_1857_sv2v_reg,
  data_r_1856_sv2v_reg,data_r_1855_sv2v_reg,data_r_1854_sv2v_reg,data_r_1853_sv2v_reg,
  data_r_1852_sv2v_reg,data_r_1851_sv2v_reg,data_r_1850_sv2v_reg,data_r_1849_sv2v_reg,
  data_r_1848_sv2v_reg,data_r_1847_sv2v_reg,data_r_1846_sv2v_reg,data_r_1845_sv2v_reg,
  data_r_1844_sv2v_reg,data_r_1843_sv2v_reg,data_r_1842_sv2v_reg,
  data_r_1841_sv2v_reg,data_r_1840_sv2v_reg,data_r_1839_sv2v_reg,data_r_1838_sv2v_reg,
  data_r_1837_sv2v_reg,data_r_1836_sv2v_reg,data_r_1835_sv2v_reg,data_r_1834_sv2v_reg,
  data_r_1833_sv2v_reg,data_r_1832_sv2v_reg,data_r_1831_sv2v_reg,data_r_1830_sv2v_reg,
  data_r_1829_sv2v_reg,data_r_1828_sv2v_reg,data_r_1827_sv2v_reg,data_r_1826_sv2v_reg,
  data_r_1825_sv2v_reg,data_r_1824_sv2v_reg,data_r_1823_sv2v_reg,
  data_r_1822_sv2v_reg,data_r_1821_sv2v_reg,data_r_1820_sv2v_reg,data_r_1819_sv2v_reg,
  data_r_1818_sv2v_reg,data_r_1817_sv2v_reg,data_r_1816_sv2v_reg,data_r_1815_sv2v_reg,
  data_r_1814_sv2v_reg,data_r_1813_sv2v_reg,data_r_1812_sv2v_reg,data_r_1811_sv2v_reg,
  data_r_1810_sv2v_reg,data_r_1809_sv2v_reg,data_r_1808_sv2v_reg,data_r_1807_sv2v_reg,
  data_r_1806_sv2v_reg,data_r_1805_sv2v_reg,data_r_1804_sv2v_reg,
  data_r_1803_sv2v_reg,data_r_1802_sv2v_reg,data_r_1801_sv2v_reg,data_r_1800_sv2v_reg,
  data_r_1799_sv2v_reg,data_r_1798_sv2v_reg,data_r_1797_sv2v_reg,data_r_1796_sv2v_reg,
  data_r_1795_sv2v_reg,data_r_1794_sv2v_reg,data_r_1793_sv2v_reg,data_r_1792_sv2v_reg,
  data_r_1791_sv2v_reg,data_r_1790_sv2v_reg,data_r_1789_sv2v_reg,data_r_1788_sv2v_reg,
  data_r_1787_sv2v_reg,data_r_1786_sv2v_reg,data_r_1785_sv2v_reg,
  data_r_1784_sv2v_reg,data_r_1783_sv2v_reg,data_r_1782_sv2v_reg,data_r_1781_sv2v_reg,
  data_r_1780_sv2v_reg,data_r_1779_sv2v_reg,data_r_1778_sv2v_reg,data_r_1777_sv2v_reg,
  data_r_1776_sv2v_reg,data_r_1775_sv2v_reg,data_r_1774_sv2v_reg,data_r_1773_sv2v_reg,
  data_r_1772_sv2v_reg,data_r_1771_sv2v_reg,data_r_1770_sv2v_reg,data_r_1769_sv2v_reg,
  data_r_1768_sv2v_reg,data_r_1767_sv2v_reg,data_r_1766_sv2v_reg,data_r_1765_sv2v_reg,
  data_r_1764_sv2v_reg,data_r_1763_sv2v_reg,data_r_1762_sv2v_reg,
  data_r_1761_sv2v_reg,data_r_1760_sv2v_reg,data_r_1759_sv2v_reg,data_r_1758_sv2v_reg,
  data_r_1757_sv2v_reg,data_r_1756_sv2v_reg,data_r_1755_sv2v_reg,data_r_1754_sv2v_reg,
  data_r_1753_sv2v_reg,data_r_1752_sv2v_reg,data_r_1751_sv2v_reg,data_r_1750_sv2v_reg,
  data_r_1749_sv2v_reg,data_r_1748_sv2v_reg,data_r_1747_sv2v_reg,data_r_1746_sv2v_reg,
  data_r_1745_sv2v_reg,data_r_1744_sv2v_reg,data_r_1743_sv2v_reg,
  data_r_1742_sv2v_reg,data_r_1741_sv2v_reg,data_r_1740_sv2v_reg,data_r_1739_sv2v_reg,
  data_r_1738_sv2v_reg,data_r_1737_sv2v_reg,data_r_1736_sv2v_reg,data_r_1735_sv2v_reg,
  data_r_1734_sv2v_reg,data_r_1733_sv2v_reg,data_r_1732_sv2v_reg,data_r_1731_sv2v_reg,
  data_r_1730_sv2v_reg,data_r_1729_sv2v_reg,data_r_1728_sv2v_reg,data_r_1727_sv2v_reg,
  data_r_1726_sv2v_reg,data_r_1725_sv2v_reg,data_r_1724_sv2v_reg,
  data_r_1723_sv2v_reg,data_r_1722_sv2v_reg,data_r_1721_sv2v_reg,data_r_1720_sv2v_reg,
  data_r_1719_sv2v_reg,data_r_1718_sv2v_reg,data_r_1717_sv2v_reg,data_r_1716_sv2v_reg,
  data_r_1715_sv2v_reg,data_r_1714_sv2v_reg,data_r_1713_sv2v_reg,data_r_1712_sv2v_reg,
  data_r_1711_sv2v_reg,data_r_1710_sv2v_reg,data_r_1709_sv2v_reg,data_r_1708_sv2v_reg,
  data_r_1707_sv2v_reg,data_r_1706_sv2v_reg,data_r_1705_sv2v_reg,
  data_r_1704_sv2v_reg,data_r_1703_sv2v_reg,data_r_1702_sv2v_reg,data_r_1701_sv2v_reg,
  data_r_1700_sv2v_reg,data_r_1699_sv2v_reg,data_r_1698_sv2v_reg,data_r_1697_sv2v_reg,
  data_r_1696_sv2v_reg,data_r_1695_sv2v_reg,data_r_1694_sv2v_reg,data_r_1693_sv2v_reg,
  data_r_1692_sv2v_reg,data_r_1691_sv2v_reg,data_r_1690_sv2v_reg,data_r_1689_sv2v_reg,
  data_r_1688_sv2v_reg,data_r_1687_sv2v_reg,data_r_1686_sv2v_reg,data_r_1685_sv2v_reg,
  data_r_1684_sv2v_reg,data_r_1683_sv2v_reg,data_r_1682_sv2v_reg,
  data_r_1681_sv2v_reg,data_r_1680_sv2v_reg,data_r_1679_sv2v_reg,data_r_1678_sv2v_reg,
  data_r_1677_sv2v_reg,data_r_1676_sv2v_reg,data_r_1675_sv2v_reg,data_r_1674_sv2v_reg,
  data_r_1673_sv2v_reg,data_r_1672_sv2v_reg,data_r_1671_sv2v_reg,data_r_1670_sv2v_reg,
  data_r_1669_sv2v_reg,data_r_1668_sv2v_reg,data_r_1667_sv2v_reg,data_r_1666_sv2v_reg,
  data_r_1665_sv2v_reg,data_r_1664_sv2v_reg,data_r_1663_sv2v_reg,
  data_r_1662_sv2v_reg,data_r_1661_sv2v_reg,data_r_1660_sv2v_reg,data_r_1659_sv2v_reg,
  data_r_1658_sv2v_reg,data_r_1657_sv2v_reg,data_r_1656_sv2v_reg,data_r_1655_sv2v_reg,
  data_r_1654_sv2v_reg,data_r_1653_sv2v_reg,data_r_1652_sv2v_reg,data_r_1651_sv2v_reg,
  data_r_1650_sv2v_reg,data_r_1649_sv2v_reg,data_r_1648_sv2v_reg,data_r_1647_sv2v_reg,
  data_r_1646_sv2v_reg,data_r_1645_sv2v_reg,data_r_1644_sv2v_reg,
  data_r_1643_sv2v_reg,data_r_1642_sv2v_reg,data_r_1641_sv2v_reg,data_r_1640_sv2v_reg,
  data_r_1639_sv2v_reg,data_r_1638_sv2v_reg,data_r_1637_sv2v_reg,data_r_1636_sv2v_reg,
  data_r_1635_sv2v_reg,data_r_1634_sv2v_reg,data_r_1633_sv2v_reg,data_r_1632_sv2v_reg,
  data_r_1631_sv2v_reg,data_r_1630_sv2v_reg,data_r_1629_sv2v_reg,data_r_1628_sv2v_reg,
  data_r_1627_sv2v_reg,data_r_1626_sv2v_reg,data_r_1625_sv2v_reg,
  data_r_1624_sv2v_reg,data_r_1623_sv2v_reg,data_r_1622_sv2v_reg,data_r_1621_sv2v_reg,
  data_r_1620_sv2v_reg,data_r_1619_sv2v_reg,data_r_1618_sv2v_reg,data_r_1617_sv2v_reg,
  data_r_1616_sv2v_reg,data_r_1615_sv2v_reg,data_r_1614_sv2v_reg,data_r_1613_sv2v_reg,
  data_r_1612_sv2v_reg,data_r_1611_sv2v_reg,data_r_1610_sv2v_reg,data_r_1609_sv2v_reg,
  data_r_1608_sv2v_reg,data_r_1607_sv2v_reg,data_r_1606_sv2v_reg,data_r_1605_sv2v_reg,
  data_r_1604_sv2v_reg,data_r_1603_sv2v_reg,data_r_1602_sv2v_reg,
  data_r_1601_sv2v_reg,data_r_1600_sv2v_reg,data_r_1599_sv2v_reg,data_r_1598_sv2v_reg,
  data_r_1597_sv2v_reg,data_r_1596_sv2v_reg,data_r_1595_sv2v_reg,data_r_1594_sv2v_reg,
  data_r_1593_sv2v_reg,data_r_1592_sv2v_reg,data_r_1591_sv2v_reg,data_r_1590_sv2v_reg,
  data_r_1589_sv2v_reg,data_r_1588_sv2v_reg,data_r_1587_sv2v_reg,data_r_1586_sv2v_reg,
  data_r_1585_sv2v_reg,data_r_1584_sv2v_reg,data_r_1583_sv2v_reg,
  data_r_1582_sv2v_reg,data_r_1581_sv2v_reg,data_r_1580_sv2v_reg,data_r_1579_sv2v_reg,
  data_r_1578_sv2v_reg,data_r_1577_sv2v_reg,data_r_1576_sv2v_reg,data_r_1575_sv2v_reg,
  data_r_1574_sv2v_reg,data_r_1573_sv2v_reg,data_r_1572_sv2v_reg,data_r_1571_sv2v_reg,
  data_r_1570_sv2v_reg,data_r_1569_sv2v_reg,data_r_1568_sv2v_reg,data_r_1567_sv2v_reg,
  data_r_1566_sv2v_reg,data_r_1565_sv2v_reg,data_r_1564_sv2v_reg,
  data_r_1563_sv2v_reg,data_r_1562_sv2v_reg,data_r_1561_sv2v_reg,data_r_1560_sv2v_reg,
  data_r_1559_sv2v_reg,data_r_1558_sv2v_reg,data_r_1557_sv2v_reg,data_r_1556_sv2v_reg,
  data_r_1555_sv2v_reg,data_r_1554_sv2v_reg,data_r_1553_sv2v_reg,data_r_1552_sv2v_reg,
  data_r_1551_sv2v_reg,data_r_1550_sv2v_reg,data_r_1549_sv2v_reg,data_r_1548_sv2v_reg,
  data_r_1547_sv2v_reg,data_r_1546_sv2v_reg,data_r_1545_sv2v_reg,
  data_r_1544_sv2v_reg,data_r_1543_sv2v_reg,data_r_1542_sv2v_reg,data_r_1541_sv2v_reg,
  data_r_1540_sv2v_reg,data_r_1539_sv2v_reg,data_r_1538_sv2v_reg,data_r_1537_sv2v_reg,
  data_r_1536_sv2v_reg,data_r_1535_sv2v_reg,data_r_1534_sv2v_reg,data_r_1533_sv2v_reg,
  data_r_1532_sv2v_reg,data_r_1531_sv2v_reg,data_r_1530_sv2v_reg,data_r_1529_sv2v_reg,
  data_r_1528_sv2v_reg,data_r_1527_sv2v_reg,data_r_1526_sv2v_reg,data_r_1525_sv2v_reg,
  data_r_1524_sv2v_reg,data_r_1523_sv2v_reg,data_r_1522_sv2v_reg,
  data_r_1521_sv2v_reg,data_r_1520_sv2v_reg,data_r_1519_sv2v_reg,data_r_1518_sv2v_reg,
  data_r_1517_sv2v_reg,data_r_1516_sv2v_reg,data_r_1515_sv2v_reg,data_r_1514_sv2v_reg,
  data_r_1513_sv2v_reg,data_r_1512_sv2v_reg,data_r_1511_sv2v_reg,data_r_1510_sv2v_reg,
  data_r_1509_sv2v_reg,data_r_1508_sv2v_reg,data_r_1507_sv2v_reg,data_r_1506_sv2v_reg,
  data_r_1505_sv2v_reg,data_r_1504_sv2v_reg,data_r_1503_sv2v_reg,
  data_r_1502_sv2v_reg,data_r_1501_sv2v_reg,data_r_1500_sv2v_reg,data_r_1499_sv2v_reg,
  data_r_1498_sv2v_reg,data_r_1497_sv2v_reg,data_r_1496_sv2v_reg,data_r_1495_sv2v_reg,
  data_r_1494_sv2v_reg,data_r_1493_sv2v_reg,data_r_1492_sv2v_reg,data_r_1491_sv2v_reg,
  data_r_1490_sv2v_reg,data_r_1489_sv2v_reg,data_r_1488_sv2v_reg,data_r_1487_sv2v_reg,
  data_r_1486_sv2v_reg,data_r_1485_sv2v_reg,data_r_1484_sv2v_reg,
  data_r_1483_sv2v_reg,data_r_1482_sv2v_reg,data_r_1481_sv2v_reg,data_r_1480_sv2v_reg,
  data_r_1479_sv2v_reg,data_r_1478_sv2v_reg,data_r_1477_sv2v_reg,data_r_1476_sv2v_reg,
  data_r_1475_sv2v_reg,data_r_1474_sv2v_reg,data_r_1473_sv2v_reg,data_r_1472_sv2v_reg,
  data_r_1471_sv2v_reg,data_r_1470_sv2v_reg,data_r_1469_sv2v_reg,data_r_1468_sv2v_reg,
  data_r_1467_sv2v_reg,data_r_1466_sv2v_reg,data_r_1465_sv2v_reg,
  data_r_1464_sv2v_reg,data_r_1463_sv2v_reg,data_r_1462_sv2v_reg,data_r_1461_sv2v_reg,
  data_r_1460_sv2v_reg,data_r_1459_sv2v_reg,data_r_1458_sv2v_reg,data_r_1457_sv2v_reg,
  data_r_1456_sv2v_reg,data_r_1455_sv2v_reg,data_r_1454_sv2v_reg,data_r_1453_sv2v_reg,
  data_r_1452_sv2v_reg,data_r_1451_sv2v_reg,data_r_1450_sv2v_reg,data_r_1449_sv2v_reg,
  data_r_1448_sv2v_reg,data_r_1447_sv2v_reg,data_r_1446_sv2v_reg,data_r_1445_sv2v_reg,
  data_r_1444_sv2v_reg,data_r_1443_sv2v_reg,data_r_1442_sv2v_reg,
  data_r_1441_sv2v_reg,data_r_1440_sv2v_reg,data_r_1439_sv2v_reg,data_r_1438_sv2v_reg,
  data_r_1437_sv2v_reg,data_r_1436_sv2v_reg,data_r_1435_sv2v_reg,data_r_1434_sv2v_reg,
  data_r_1433_sv2v_reg,data_r_1432_sv2v_reg,data_r_1431_sv2v_reg,data_r_1430_sv2v_reg,
  data_r_1429_sv2v_reg,data_r_1428_sv2v_reg,data_r_1427_sv2v_reg,data_r_1426_sv2v_reg,
  data_r_1425_sv2v_reg,data_r_1424_sv2v_reg,data_r_1423_sv2v_reg,
  data_r_1422_sv2v_reg,data_r_1421_sv2v_reg,data_r_1420_sv2v_reg,data_r_1419_sv2v_reg,
  data_r_1418_sv2v_reg,data_r_1417_sv2v_reg,data_r_1416_sv2v_reg,data_r_1415_sv2v_reg,
  data_r_1414_sv2v_reg,data_r_1413_sv2v_reg,data_r_1412_sv2v_reg,data_r_1411_sv2v_reg,
  data_r_1410_sv2v_reg,data_r_1409_sv2v_reg,data_r_1408_sv2v_reg,data_r_1407_sv2v_reg,
  data_r_1406_sv2v_reg,data_r_1405_sv2v_reg,data_r_1404_sv2v_reg,
  data_r_1403_sv2v_reg,data_r_1402_sv2v_reg,data_r_1401_sv2v_reg,data_r_1400_sv2v_reg,
  data_r_1399_sv2v_reg,data_r_1398_sv2v_reg,data_r_1397_sv2v_reg,data_r_1396_sv2v_reg,
  data_r_1395_sv2v_reg,data_r_1394_sv2v_reg,data_r_1393_sv2v_reg,data_r_1392_sv2v_reg,
  data_r_1391_sv2v_reg,data_r_1390_sv2v_reg,data_r_1389_sv2v_reg,data_r_1388_sv2v_reg,
  data_r_1387_sv2v_reg,data_r_1386_sv2v_reg,data_r_1385_sv2v_reg,
  data_r_1384_sv2v_reg,data_r_1383_sv2v_reg,data_r_1382_sv2v_reg,data_r_1381_sv2v_reg,
  data_r_1380_sv2v_reg,data_r_1379_sv2v_reg,data_r_1378_sv2v_reg,data_r_1377_sv2v_reg,
  data_r_1376_sv2v_reg,data_r_1375_sv2v_reg,data_r_1374_sv2v_reg,data_r_1373_sv2v_reg,
  data_r_1372_sv2v_reg,data_r_1371_sv2v_reg,data_r_1370_sv2v_reg,data_r_1369_sv2v_reg,
  data_r_1368_sv2v_reg,data_r_1367_sv2v_reg,data_r_1366_sv2v_reg,data_r_1365_sv2v_reg,
  data_r_1364_sv2v_reg,data_r_1363_sv2v_reg,data_r_1362_sv2v_reg,
  data_r_1361_sv2v_reg,data_r_1360_sv2v_reg,data_r_1359_sv2v_reg,data_r_1358_sv2v_reg,
  data_r_1357_sv2v_reg,data_r_1356_sv2v_reg,data_r_1355_sv2v_reg,data_r_1354_sv2v_reg,
  data_r_1353_sv2v_reg,data_r_1352_sv2v_reg,data_r_1351_sv2v_reg,data_r_1350_sv2v_reg,
  data_r_1349_sv2v_reg,data_r_1348_sv2v_reg,data_r_1347_sv2v_reg,data_r_1346_sv2v_reg,
  data_r_1345_sv2v_reg,data_r_1344_sv2v_reg,data_r_1343_sv2v_reg,
  data_r_1342_sv2v_reg,data_r_1341_sv2v_reg,data_r_1340_sv2v_reg,data_r_1339_sv2v_reg,
  data_r_1338_sv2v_reg,data_r_1337_sv2v_reg,data_r_1336_sv2v_reg,data_r_1335_sv2v_reg,
  data_r_1334_sv2v_reg,data_r_1333_sv2v_reg,data_r_1332_sv2v_reg,data_r_1331_sv2v_reg,
  data_r_1330_sv2v_reg,data_r_1329_sv2v_reg,data_r_1328_sv2v_reg,data_r_1327_sv2v_reg,
  data_r_1326_sv2v_reg,data_r_1325_sv2v_reg,data_r_1324_sv2v_reg,
  data_r_1323_sv2v_reg,data_r_1322_sv2v_reg,data_r_1321_sv2v_reg,data_r_1320_sv2v_reg,
  data_r_1319_sv2v_reg,data_r_1318_sv2v_reg,data_r_1317_sv2v_reg,data_r_1316_sv2v_reg,
  data_r_1315_sv2v_reg,data_r_1314_sv2v_reg,data_r_1313_sv2v_reg,data_r_1312_sv2v_reg,
  data_r_1311_sv2v_reg,data_r_1310_sv2v_reg,data_r_1309_sv2v_reg,data_r_1308_sv2v_reg,
  data_r_1307_sv2v_reg,data_r_1306_sv2v_reg,data_r_1305_sv2v_reg,
  data_r_1304_sv2v_reg,data_r_1303_sv2v_reg,data_r_1302_sv2v_reg,data_r_1301_sv2v_reg,
  data_r_1300_sv2v_reg,data_r_1299_sv2v_reg,data_r_1298_sv2v_reg,data_r_1297_sv2v_reg,
  data_r_1296_sv2v_reg,data_r_1295_sv2v_reg,data_r_1294_sv2v_reg,data_r_1293_sv2v_reg,
  data_r_1292_sv2v_reg,data_r_1291_sv2v_reg,data_r_1290_sv2v_reg,data_r_1289_sv2v_reg,
  data_r_1288_sv2v_reg,data_r_1287_sv2v_reg,data_r_1286_sv2v_reg,data_r_1285_sv2v_reg,
  data_r_1284_sv2v_reg,data_r_1283_sv2v_reg,data_r_1282_sv2v_reg,
  data_r_1281_sv2v_reg,data_r_1280_sv2v_reg,data_r_1279_sv2v_reg,data_r_1278_sv2v_reg,
  data_r_1277_sv2v_reg,data_r_1276_sv2v_reg,data_r_1275_sv2v_reg,data_r_1274_sv2v_reg,
  data_r_1273_sv2v_reg,data_r_1272_sv2v_reg,data_r_1271_sv2v_reg,data_r_1270_sv2v_reg,
  data_r_1269_sv2v_reg,data_r_1268_sv2v_reg,data_r_1267_sv2v_reg,data_r_1266_sv2v_reg,
  data_r_1265_sv2v_reg,data_r_1264_sv2v_reg,data_r_1263_sv2v_reg,
  data_r_1262_sv2v_reg,data_r_1261_sv2v_reg,data_r_1260_sv2v_reg,data_r_1259_sv2v_reg,
  data_r_1258_sv2v_reg,data_r_1257_sv2v_reg,data_r_1256_sv2v_reg,data_r_1255_sv2v_reg,
  data_r_1254_sv2v_reg,data_r_1253_sv2v_reg,data_r_1252_sv2v_reg,data_r_1251_sv2v_reg,
  data_r_1250_sv2v_reg,data_r_1249_sv2v_reg,data_r_1248_sv2v_reg,data_r_1247_sv2v_reg,
  data_r_1246_sv2v_reg,data_r_1245_sv2v_reg,data_r_1244_sv2v_reg,
  data_r_1243_sv2v_reg,data_r_1242_sv2v_reg,data_r_1241_sv2v_reg,data_r_1240_sv2v_reg,
  data_r_1239_sv2v_reg,data_r_1238_sv2v_reg,data_r_1237_sv2v_reg,data_r_1236_sv2v_reg,
  data_r_1235_sv2v_reg,data_r_1234_sv2v_reg,data_r_1233_sv2v_reg,data_r_1232_sv2v_reg,
  data_r_1231_sv2v_reg,data_r_1230_sv2v_reg,data_r_1229_sv2v_reg,data_r_1228_sv2v_reg,
  data_r_1227_sv2v_reg,data_r_1226_sv2v_reg,data_r_1225_sv2v_reg,
  data_r_1224_sv2v_reg,data_r_1223_sv2v_reg,data_r_1222_sv2v_reg,data_r_1221_sv2v_reg,
  data_r_1220_sv2v_reg,data_r_1219_sv2v_reg,data_r_1218_sv2v_reg,data_r_1217_sv2v_reg,
  data_r_1216_sv2v_reg,data_r_1215_sv2v_reg,data_r_1214_sv2v_reg,data_r_1213_sv2v_reg,
  data_r_1212_sv2v_reg,data_r_1211_sv2v_reg,data_r_1210_sv2v_reg,data_r_1209_sv2v_reg,
  data_r_1208_sv2v_reg,data_r_1207_sv2v_reg,data_r_1206_sv2v_reg,data_r_1205_sv2v_reg,
  data_r_1204_sv2v_reg,data_r_1203_sv2v_reg,data_r_1202_sv2v_reg,
  data_r_1201_sv2v_reg,data_r_1200_sv2v_reg,data_r_1199_sv2v_reg,data_r_1198_sv2v_reg,
  data_r_1197_sv2v_reg,data_r_1196_sv2v_reg,data_r_1195_sv2v_reg,data_r_1194_sv2v_reg,
  data_r_1193_sv2v_reg,data_r_1192_sv2v_reg,data_r_1191_sv2v_reg,data_r_1190_sv2v_reg,
  data_r_1189_sv2v_reg,data_r_1188_sv2v_reg,data_r_1187_sv2v_reg,data_r_1186_sv2v_reg,
  data_r_1185_sv2v_reg,data_r_1184_sv2v_reg,data_r_1183_sv2v_reg,
  data_r_1182_sv2v_reg,data_r_1181_sv2v_reg,data_r_1180_sv2v_reg,data_r_1179_sv2v_reg,
  data_r_1178_sv2v_reg,data_r_1177_sv2v_reg,data_r_1176_sv2v_reg,data_r_1175_sv2v_reg,
  data_r_1174_sv2v_reg,data_r_1173_sv2v_reg,data_r_1172_sv2v_reg,data_r_1171_sv2v_reg,
  data_r_1170_sv2v_reg,data_r_1169_sv2v_reg,data_r_1168_sv2v_reg,data_r_1167_sv2v_reg,
  data_r_1166_sv2v_reg,data_r_1165_sv2v_reg,data_r_1164_sv2v_reg,
  data_r_1163_sv2v_reg,data_r_1162_sv2v_reg,data_r_1161_sv2v_reg,data_r_1160_sv2v_reg,
  data_r_1159_sv2v_reg,data_r_1158_sv2v_reg,data_r_1157_sv2v_reg,data_r_1156_sv2v_reg,
  data_r_1155_sv2v_reg,data_r_1154_sv2v_reg,data_r_1153_sv2v_reg,data_r_1152_sv2v_reg,
  data_r_1151_sv2v_reg,data_r_1150_sv2v_reg,data_r_1149_sv2v_reg,data_r_1148_sv2v_reg,
  data_r_1147_sv2v_reg,data_r_1146_sv2v_reg,data_r_1145_sv2v_reg,
  data_r_1144_sv2v_reg,data_r_1143_sv2v_reg,data_r_1142_sv2v_reg,data_r_1141_sv2v_reg,
  data_r_1140_sv2v_reg,data_r_1139_sv2v_reg,data_r_1138_sv2v_reg,data_r_1137_sv2v_reg,
  data_r_1136_sv2v_reg,data_r_1135_sv2v_reg,data_r_1134_sv2v_reg,data_r_1133_sv2v_reg,
  data_r_1132_sv2v_reg,data_r_1131_sv2v_reg,data_r_1130_sv2v_reg,data_r_1129_sv2v_reg,
  data_r_1128_sv2v_reg,data_r_1127_sv2v_reg,data_r_1126_sv2v_reg,data_r_1125_sv2v_reg,
  data_r_1124_sv2v_reg,data_r_1123_sv2v_reg,data_r_1122_sv2v_reg,
  data_r_1121_sv2v_reg,data_r_1120_sv2v_reg,data_r_1119_sv2v_reg,data_r_1118_sv2v_reg,
  data_r_1117_sv2v_reg,data_r_1116_sv2v_reg,data_r_1115_sv2v_reg,data_r_1114_sv2v_reg,
  data_r_1113_sv2v_reg,data_r_1112_sv2v_reg,data_r_1111_sv2v_reg,data_r_1110_sv2v_reg,
  data_r_1109_sv2v_reg,data_r_1108_sv2v_reg,data_r_1107_sv2v_reg,data_r_1106_sv2v_reg,
  data_r_1105_sv2v_reg,data_r_1104_sv2v_reg,data_r_1103_sv2v_reg,
  data_r_1102_sv2v_reg,data_r_1101_sv2v_reg,data_r_1100_sv2v_reg,data_r_1099_sv2v_reg,
  data_r_1098_sv2v_reg,data_r_1097_sv2v_reg,data_r_1096_sv2v_reg,data_r_1095_sv2v_reg,
  data_r_1094_sv2v_reg,data_r_1093_sv2v_reg,data_r_1092_sv2v_reg,data_r_1091_sv2v_reg,
  data_r_1090_sv2v_reg,data_r_1089_sv2v_reg,data_r_1088_sv2v_reg,data_r_1087_sv2v_reg,
  data_r_1086_sv2v_reg,data_r_1085_sv2v_reg,data_r_1084_sv2v_reg,
  data_r_1083_sv2v_reg,data_r_1082_sv2v_reg,data_r_1081_sv2v_reg,data_r_1080_sv2v_reg,
  data_r_1079_sv2v_reg,data_r_1078_sv2v_reg,data_r_1077_sv2v_reg,data_r_1076_sv2v_reg,
  data_r_1075_sv2v_reg,data_r_1074_sv2v_reg,data_r_1073_sv2v_reg,data_r_1072_sv2v_reg,
  data_r_1071_sv2v_reg,data_r_1070_sv2v_reg,data_r_1069_sv2v_reg,data_r_1068_sv2v_reg,
  data_r_1067_sv2v_reg,data_r_1066_sv2v_reg,data_r_1065_sv2v_reg,
  data_r_1064_sv2v_reg,data_r_1063_sv2v_reg,data_r_1062_sv2v_reg,data_r_1061_sv2v_reg,
  data_r_1060_sv2v_reg,data_r_1059_sv2v_reg,data_r_1058_sv2v_reg,data_r_1057_sv2v_reg,
  data_r_1056_sv2v_reg,data_r_1055_sv2v_reg,data_r_1054_sv2v_reg,data_r_1053_sv2v_reg,
  data_r_1052_sv2v_reg,data_r_1051_sv2v_reg,data_r_1050_sv2v_reg,data_r_1049_sv2v_reg,
  data_r_1048_sv2v_reg,data_r_1047_sv2v_reg,data_r_1046_sv2v_reg,data_r_1045_sv2v_reg,
  data_r_1044_sv2v_reg,data_r_1043_sv2v_reg,data_r_1042_sv2v_reg,
  data_r_1041_sv2v_reg,data_r_1040_sv2v_reg,data_r_1039_sv2v_reg,data_r_1038_sv2v_reg,
  data_r_1037_sv2v_reg,data_r_1036_sv2v_reg,data_r_1035_sv2v_reg,data_r_1034_sv2v_reg,
  data_r_1033_sv2v_reg,data_r_1032_sv2v_reg,data_r_1031_sv2v_reg,data_r_1030_sv2v_reg,
  data_r_1029_sv2v_reg,data_r_1028_sv2v_reg,data_r_1027_sv2v_reg,data_r_1026_sv2v_reg,
  data_r_1025_sv2v_reg,data_r_1024_sv2v_reg,data_r_1023_sv2v_reg,
  data_r_1022_sv2v_reg,data_r_1021_sv2v_reg,data_r_1020_sv2v_reg,data_r_1019_sv2v_reg,
  data_r_1018_sv2v_reg,data_r_1017_sv2v_reg,data_r_1016_sv2v_reg,data_r_1015_sv2v_reg,
  data_r_1014_sv2v_reg,data_r_1013_sv2v_reg,data_r_1012_sv2v_reg,data_r_1011_sv2v_reg,
  data_r_1010_sv2v_reg,data_r_1009_sv2v_reg,data_r_1008_sv2v_reg,data_r_1007_sv2v_reg,
  data_r_1006_sv2v_reg,data_r_1005_sv2v_reg,data_r_1004_sv2v_reg,
  data_r_1003_sv2v_reg,data_r_1002_sv2v_reg,data_r_1001_sv2v_reg,data_r_1000_sv2v_reg,
  data_r_999_sv2v_reg,data_r_998_sv2v_reg,data_r_997_sv2v_reg,data_r_996_sv2v_reg,
  data_r_995_sv2v_reg,data_r_994_sv2v_reg,data_r_993_sv2v_reg,data_r_992_sv2v_reg,
  data_r_991_sv2v_reg,data_r_990_sv2v_reg,data_r_989_sv2v_reg,data_r_988_sv2v_reg,
  data_r_987_sv2v_reg,data_r_986_sv2v_reg,data_r_985_sv2v_reg,data_r_984_sv2v_reg,
  data_r_983_sv2v_reg,data_r_982_sv2v_reg,data_r_981_sv2v_reg,data_r_980_sv2v_reg,
  data_r_979_sv2v_reg,data_r_978_sv2v_reg,data_r_977_sv2v_reg,data_r_976_sv2v_reg,
  data_r_975_sv2v_reg,data_r_974_sv2v_reg,data_r_973_sv2v_reg,data_r_972_sv2v_reg,
  data_r_971_sv2v_reg,data_r_970_sv2v_reg,data_r_969_sv2v_reg,data_r_968_sv2v_reg,
  data_r_967_sv2v_reg,data_r_966_sv2v_reg,data_r_965_sv2v_reg,data_r_964_sv2v_reg,
  data_r_963_sv2v_reg,data_r_962_sv2v_reg,data_r_961_sv2v_reg,data_r_960_sv2v_reg,
  data_r_959_sv2v_reg,data_r_958_sv2v_reg,data_r_957_sv2v_reg,data_r_956_sv2v_reg,
  data_r_955_sv2v_reg,data_r_954_sv2v_reg,data_r_953_sv2v_reg,data_r_952_sv2v_reg,
  data_r_951_sv2v_reg,data_r_950_sv2v_reg,data_r_949_sv2v_reg,data_r_948_sv2v_reg,
  data_r_947_sv2v_reg,data_r_946_sv2v_reg,data_r_945_sv2v_reg,data_r_944_sv2v_reg,
  data_r_943_sv2v_reg,data_r_942_sv2v_reg,data_r_941_sv2v_reg,data_r_940_sv2v_reg,
  data_r_939_sv2v_reg,data_r_938_sv2v_reg,data_r_937_sv2v_reg,data_r_936_sv2v_reg,
  data_r_935_sv2v_reg,data_r_934_sv2v_reg,data_r_933_sv2v_reg,data_r_932_sv2v_reg,
  data_r_931_sv2v_reg,data_r_930_sv2v_reg,data_r_929_sv2v_reg,data_r_928_sv2v_reg,
  data_r_927_sv2v_reg,data_r_926_sv2v_reg,data_r_925_sv2v_reg,data_r_924_sv2v_reg,
  data_r_923_sv2v_reg,data_r_922_sv2v_reg,data_r_921_sv2v_reg,data_r_920_sv2v_reg,
  data_r_919_sv2v_reg,data_r_918_sv2v_reg,data_r_917_sv2v_reg,data_r_916_sv2v_reg,
  data_r_915_sv2v_reg,data_r_914_sv2v_reg,data_r_913_sv2v_reg,data_r_912_sv2v_reg,
  data_r_911_sv2v_reg,data_r_910_sv2v_reg,data_r_909_sv2v_reg,data_r_908_sv2v_reg,
  data_r_907_sv2v_reg,data_r_906_sv2v_reg,data_r_905_sv2v_reg,data_r_904_sv2v_reg,
  data_r_903_sv2v_reg,data_r_902_sv2v_reg,data_r_901_sv2v_reg,data_r_900_sv2v_reg,
  data_r_899_sv2v_reg,data_r_898_sv2v_reg,data_r_897_sv2v_reg,data_r_896_sv2v_reg,
  data_r_895_sv2v_reg,data_r_894_sv2v_reg,data_r_893_sv2v_reg,data_r_892_sv2v_reg,
  data_r_891_sv2v_reg,data_r_890_sv2v_reg,data_r_889_sv2v_reg,data_r_888_sv2v_reg,
  data_r_887_sv2v_reg,data_r_886_sv2v_reg,data_r_885_sv2v_reg,data_r_884_sv2v_reg,
  data_r_883_sv2v_reg,data_r_882_sv2v_reg,data_r_881_sv2v_reg,data_r_880_sv2v_reg,
  data_r_879_sv2v_reg,data_r_878_sv2v_reg,data_r_877_sv2v_reg,data_r_876_sv2v_reg,
  data_r_875_sv2v_reg,data_r_874_sv2v_reg,data_r_873_sv2v_reg,data_r_872_sv2v_reg,
  data_r_871_sv2v_reg,data_r_870_sv2v_reg,data_r_869_sv2v_reg,data_r_868_sv2v_reg,
  data_r_867_sv2v_reg,data_r_866_sv2v_reg,data_r_865_sv2v_reg,data_r_864_sv2v_reg,
  data_r_863_sv2v_reg,data_r_862_sv2v_reg,data_r_861_sv2v_reg,data_r_860_sv2v_reg,
  data_r_859_sv2v_reg,data_r_858_sv2v_reg,data_r_857_sv2v_reg,data_r_856_sv2v_reg,
  data_r_855_sv2v_reg,data_r_854_sv2v_reg,data_r_853_sv2v_reg,data_r_852_sv2v_reg,
  data_r_851_sv2v_reg,data_r_850_sv2v_reg,data_r_849_sv2v_reg,data_r_848_sv2v_reg,
  data_r_847_sv2v_reg,data_r_846_sv2v_reg,data_r_845_sv2v_reg,data_r_844_sv2v_reg,
  data_r_843_sv2v_reg,data_r_842_sv2v_reg,data_r_841_sv2v_reg,data_r_840_sv2v_reg,
  data_r_839_sv2v_reg,data_r_838_sv2v_reg,data_r_837_sv2v_reg,data_r_836_sv2v_reg,
  data_r_835_sv2v_reg,data_r_834_sv2v_reg,data_r_833_sv2v_reg,data_r_832_sv2v_reg,
  data_r_831_sv2v_reg,data_r_830_sv2v_reg,data_r_829_sv2v_reg,data_r_828_sv2v_reg,
  data_r_827_sv2v_reg,data_r_826_sv2v_reg,data_r_825_sv2v_reg,data_r_824_sv2v_reg,
  data_r_823_sv2v_reg,data_r_822_sv2v_reg,data_r_821_sv2v_reg,data_r_820_sv2v_reg,
  data_r_819_sv2v_reg,data_r_818_sv2v_reg,data_r_817_sv2v_reg,data_r_816_sv2v_reg,
  data_r_815_sv2v_reg,data_r_814_sv2v_reg,data_r_813_sv2v_reg,data_r_812_sv2v_reg,
  data_r_811_sv2v_reg,data_r_810_sv2v_reg,data_r_809_sv2v_reg,data_r_808_sv2v_reg,
  data_r_807_sv2v_reg,data_r_806_sv2v_reg,data_r_805_sv2v_reg,data_r_804_sv2v_reg,
  data_r_803_sv2v_reg,data_r_802_sv2v_reg,data_r_801_sv2v_reg,data_r_800_sv2v_reg,
  data_r_799_sv2v_reg,data_r_798_sv2v_reg,data_r_797_sv2v_reg,data_r_796_sv2v_reg,
  data_r_795_sv2v_reg,data_r_794_sv2v_reg,data_r_793_sv2v_reg,data_r_792_sv2v_reg,
  data_r_791_sv2v_reg,data_r_790_sv2v_reg,data_r_789_sv2v_reg,data_r_788_sv2v_reg,
  data_r_787_sv2v_reg,data_r_786_sv2v_reg,data_r_785_sv2v_reg,data_r_784_sv2v_reg,
  data_r_783_sv2v_reg,data_r_782_sv2v_reg,data_r_781_sv2v_reg,data_r_780_sv2v_reg,
  data_r_779_sv2v_reg,data_r_778_sv2v_reg,data_r_777_sv2v_reg,data_r_776_sv2v_reg,
  data_r_775_sv2v_reg,data_r_774_sv2v_reg,data_r_773_sv2v_reg,data_r_772_sv2v_reg,
  data_r_771_sv2v_reg,data_r_770_sv2v_reg,data_r_769_sv2v_reg,data_r_768_sv2v_reg,
  data_r_767_sv2v_reg,data_r_766_sv2v_reg,data_r_765_sv2v_reg,data_r_764_sv2v_reg,
  data_r_763_sv2v_reg,data_r_762_sv2v_reg,data_r_761_sv2v_reg,data_r_760_sv2v_reg,
  data_r_759_sv2v_reg,data_r_758_sv2v_reg,data_r_757_sv2v_reg,data_r_756_sv2v_reg,
  data_r_755_sv2v_reg,data_r_754_sv2v_reg,data_r_753_sv2v_reg,data_r_752_sv2v_reg,
  data_r_751_sv2v_reg,data_r_750_sv2v_reg,data_r_749_sv2v_reg,data_r_748_sv2v_reg,
  data_r_747_sv2v_reg,data_r_746_sv2v_reg,data_r_745_sv2v_reg,data_r_744_sv2v_reg,
  data_r_743_sv2v_reg,data_r_742_sv2v_reg,data_r_741_sv2v_reg,data_r_740_sv2v_reg,
  data_r_739_sv2v_reg,data_r_738_sv2v_reg,data_r_737_sv2v_reg,data_r_736_sv2v_reg,
  data_r_735_sv2v_reg,data_r_734_sv2v_reg,data_r_733_sv2v_reg,data_r_732_sv2v_reg,
  data_r_731_sv2v_reg,data_r_730_sv2v_reg,data_r_729_sv2v_reg,data_r_728_sv2v_reg,
  data_r_727_sv2v_reg,data_r_726_sv2v_reg,data_r_725_sv2v_reg,data_r_724_sv2v_reg,
  data_r_723_sv2v_reg,data_r_722_sv2v_reg,data_r_721_sv2v_reg,data_r_720_sv2v_reg,
  data_r_719_sv2v_reg,data_r_718_sv2v_reg,data_r_717_sv2v_reg,data_r_716_sv2v_reg,
  data_r_715_sv2v_reg,data_r_714_sv2v_reg,data_r_713_sv2v_reg,data_r_712_sv2v_reg,
  data_r_711_sv2v_reg,data_r_710_sv2v_reg,data_r_709_sv2v_reg,data_r_708_sv2v_reg,
  data_r_707_sv2v_reg,data_r_706_sv2v_reg,data_r_705_sv2v_reg,data_r_704_sv2v_reg,
  data_r_703_sv2v_reg,data_r_702_sv2v_reg,data_r_701_sv2v_reg,data_r_700_sv2v_reg,
  data_r_699_sv2v_reg,data_r_698_sv2v_reg,data_r_697_sv2v_reg,data_r_696_sv2v_reg,
  data_r_695_sv2v_reg,data_r_694_sv2v_reg,data_r_693_sv2v_reg,data_r_692_sv2v_reg,
  data_r_691_sv2v_reg,data_r_690_sv2v_reg,data_r_689_sv2v_reg,data_r_688_sv2v_reg,
  data_r_687_sv2v_reg,data_r_686_sv2v_reg,data_r_685_sv2v_reg,data_r_684_sv2v_reg,
  data_r_683_sv2v_reg,data_r_682_sv2v_reg,data_r_681_sv2v_reg,data_r_680_sv2v_reg,
  data_r_679_sv2v_reg,data_r_678_sv2v_reg,data_r_677_sv2v_reg,data_r_676_sv2v_reg,
  data_r_675_sv2v_reg,data_r_674_sv2v_reg,data_r_673_sv2v_reg,data_r_672_sv2v_reg,
  data_r_671_sv2v_reg,data_r_670_sv2v_reg,data_r_669_sv2v_reg,data_r_668_sv2v_reg,
  data_r_667_sv2v_reg,data_r_666_sv2v_reg,data_r_665_sv2v_reg,data_r_664_sv2v_reg,
  data_r_663_sv2v_reg,data_r_662_sv2v_reg,data_r_661_sv2v_reg,data_r_660_sv2v_reg,
  data_r_659_sv2v_reg,data_r_658_sv2v_reg,data_r_657_sv2v_reg,data_r_656_sv2v_reg,
  data_r_655_sv2v_reg,data_r_654_sv2v_reg,data_r_653_sv2v_reg,data_r_652_sv2v_reg,
  data_r_651_sv2v_reg,data_r_650_sv2v_reg,data_r_649_sv2v_reg,data_r_648_sv2v_reg,
  data_r_647_sv2v_reg,data_r_646_sv2v_reg,data_r_645_sv2v_reg,data_r_644_sv2v_reg,
  data_r_643_sv2v_reg,data_r_642_sv2v_reg,data_r_641_sv2v_reg,data_r_640_sv2v_reg,
  data_r_639_sv2v_reg,data_r_638_sv2v_reg,data_r_637_sv2v_reg,data_r_636_sv2v_reg,
  data_r_635_sv2v_reg,data_r_634_sv2v_reg,data_r_633_sv2v_reg,data_r_632_sv2v_reg,
  data_r_631_sv2v_reg,data_r_630_sv2v_reg,data_r_629_sv2v_reg,data_r_628_sv2v_reg,
  data_r_627_sv2v_reg,data_r_626_sv2v_reg,data_r_625_sv2v_reg,data_r_624_sv2v_reg,
  data_r_623_sv2v_reg,data_r_622_sv2v_reg,data_r_621_sv2v_reg,data_r_620_sv2v_reg,
  data_r_619_sv2v_reg,data_r_618_sv2v_reg,data_r_617_sv2v_reg,data_r_616_sv2v_reg,
  data_r_615_sv2v_reg,data_r_614_sv2v_reg,data_r_613_sv2v_reg,data_r_612_sv2v_reg,
  data_r_611_sv2v_reg,data_r_610_sv2v_reg,data_r_609_sv2v_reg,data_r_608_sv2v_reg,
  data_r_607_sv2v_reg,data_r_606_sv2v_reg,data_r_605_sv2v_reg,data_r_604_sv2v_reg,
  data_r_603_sv2v_reg,data_r_602_sv2v_reg,data_r_601_sv2v_reg,data_r_600_sv2v_reg,
  data_r_599_sv2v_reg,data_r_598_sv2v_reg,data_r_597_sv2v_reg,data_r_596_sv2v_reg,
  data_r_595_sv2v_reg,data_r_594_sv2v_reg,data_r_593_sv2v_reg,data_r_592_sv2v_reg,
  data_r_591_sv2v_reg,data_r_590_sv2v_reg,data_r_589_sv2v_reg,data_r_588_sv2v_reg,
  data_r_587_sv2v_reg,data_r_586_sv2v_reg,data_r_585_sv2v_reg,data_r_584_sv2v_reg,
  data_r_583_sv2v_reg,data_r_582_sv2v_reg,data_r_581_sv2v_reg,data_r_580_sv2v_reg,
  data_r_579_sv2v_reg,data_r_578_sv2v_reg,data_r_577_sv2v_reg,data_r_576_sv2v_reg,
  data_r_575_sv2v_reg,data_r_574_sv2v_reg,data_r_573_sv2v_reg,data_r_572_sv2v_reg,
  data_r_571_sv2v_reg,data_r_570_sv2v_reg,data_r_569_sv2v_reg,data_r_568_sv2v_reg,
  data_r_567_sv2v_reg,data_r_566_sv2v_reg,data_r_565_sv2v_reg,data_r_564_sv2v_reg,
  data_r_563_sv2v_reg,data_r_562_sv2v_reg,data_r_561_sv2v_reg,data_r_560_sv2v_reg,
  data_r_559_sv2v_reg,data_r_558_sv2v_reg,data_r_557_sv2v_reg,data_r_556_sv2v_reg,
  data_r_555_sv2v_reg,data_r_554_sv2v_reg,data_r_553_sv2v_reg,data_r_552_sv2v_reg,
  data_r_551_sv2v_reg,data_r_550_sv2v_reg,data_r_549_sv2v_reg,data_r_548_sv2v_reg,
  data_r_547_sv2v_reg,data_r_546_sv2v_reg,data_r_545_sv2v_reg,data_r_544_sv2v_reg,
  data_r_543_sv2v_reg,data_r_542_sv2v_reg,data_r_541_sv2v_reg,data_r_540_sv2v_reg,
  data_r_539_sv2v_reg,data_r_538_sv2v_reg,data_r_537_sv2v_reg,data_r_536_sv2v_reg,
  data_r_535_sv2v_reg,data_r_534_sv2v_reg,data_r_533_sv2v_reg,data_r_532_sv2v_reg,
  data_r_531_sv2v_reg,data_r_530_sv2v_reg,data_r_529_sv2v_reg,data_r_528_sv2v_reg,
  data_r_527_sv2v_reg,data_r_526_sv2v_reg,data_r_525_sv2v_reg,data_r_524_sv2v_reg,
  data_r_523_sv2v_reg,data_r_522_sv2v_reg,data_r_521_sv2v_reg,data_r_520_sv2v_reg,
  data_r_519_sv2v_reg,data_r_518_sv2v_reg,data_r_517_sv2v_reg,data_r_516_sv2v_reg,
  data_r_515_sv2v_reg,data_r_514_sv2v_reg,data_r_513_sv2v_reg,data_r_512_sv2v_reg,
  data_r_511_sv2v_reg,data_r_510_sv2v_reg,data_r_509_sv2v_reg,data_r_508_sv2v_reg,
  data_r_507_sv2v_reg,data_r_506_sv2v_reg,data_r_505_sv2v_reg,data_r_504_sv2v_reg,
  data_r_503_sv2v_reg,data_r_502_sv2v_reg,data_r_501_sv2v_reg,data_r_500_sv2v_reg,
  data_r_499_sv2v_reg,data_r_498_sv2v_reg,data_r_497_sv2v_reg,data_r_496_sv2v_reg,
  data_r_495_sv2v_reg,data_r_494_sv2v_reg,data_r_493_sv2v_reg,data_r_492_sv2v_reg,
  data_r_491_sv2v_reg,data_r_490_sv2v_reg,data_r_489_sv2v_reg,data_r_488_sv2v_reg,
  data_r_487_sv2v_reg,data_r_486_sv2v_reg,data_r_485_sv2v_reg,data_r_484_sv2v_reg,
  data_r_483_sv2v_reg,data_r_482_sv2v_reg,data_r_481_sv2v_reg,data_r_480_sv2v_reg,
  data_r_479_sv2v_reg,data_r_478_sv2v_reg,data_r_477_sv2v_reg,data_r_476_sv2v_reg,
  data_r_475_sv2v_reg,data_r_474_sv2v_reg,data_r_473_sv2v_reg,data_r_472_sv2v_reg,
  data_r_471_sv2v_reg,data_r_470_sv2v_reg,data_r_469_sv2v_reg,data_r_468_sv2v_reg,
  data_r_467_sv2v_reg,data_r_466_sv2v_reg,data_r_465_sv2v_reg,data_r_464_sv2v_reg,
  data_r_463_sv2v_reg,data_r_462_sv2v_reg,data_r_461_sv2v_reg,data_r_460_sv2v_reg,
  data_r_459_sv2v_reg,data_r_458_sv2v_reg,data_r_457_sv2v_reg,data_r_456_sv2v_reg,
  data_r_455_sv2v_reg,data_r_454_sv2v_reg,data_r_453_sv2v_reg,data_r_452_sv2v_reg,
  data_r_451_sv2v_reg,data_r_450_sv2v_reg,data_r_449_sv2v_reg,data_r_448_sv2v_reg,
  data_r_447_sv2v_reg,data_r_446_sv2v_reg,data_r_445_sv2v_reg,data_r_444_sv2v_reg,
  data_r_443_sv2v_reg,data_r_442_sv2v_reg,data_r_441_sv2v_reg,data_r_440_sv2v_reg,
  data_r_439_sv2v_reg,data_r_438_sv2v_reg,data_r_437_sv2v_reg,data_r_436_sv2v_reg,
  data_r_435_sv2v_reg,data_r_434_sv2v_reg,data_r_433_sv2v_reg,data_r_432_sv2v_reg,
  data_r_431_sv2v_reg,data_r_430_sv2v_reg,data_r_429_sv2v_reg,data_r_428_sv2v_reg,
  data_r_427_sv2v_reg,data_r_426_sv2v_reg,data_r_425_sv2v_reg,data_r_424_sv2v_reg,
  data_r_423_sv2v_reg,data_r_422_sv2v_reg,data_r_421_sv2v_reg,data_r_420_sv2v_reg,
  data_r_419_sv2v_reg,data_r_418_sv2v_reg,data_r_417_sv2v_reg,data_r_416_sv2v_reg,
  data_r_415_sv2v_reg,data_r_414_sv2v_reg,data_r_413_sv2v_reg,data_r_412_sv2v_reg,
  data_r_411_sv2v_reg,data_r_410_sv2v_reg,data_r_409_sv2v_reg,data_r_408_sv2v_reg,
  data_r_407_sv2v_reg,data_r_406_sv2v_reg,data_r_405_sv2v_reg,data_r_404_sv2v_reg,
  data_r_403_sv2v_reg,data_r_402_sv2v_reg,data_r_401_sv2v_reg,data_r_400_sv2v_reg,
  data_r_399_sv2v_reg,data_r_398_sv2v_reg,data_r_397_sv2v_reg,data_r_396_sv2v_reg,
  data_r_395_sv2v_reg,data_r_394_sv2v_reg,data_r_393_sv2v_reg,data_r_392_sv2v_reg,
  data_r_391_sv2v_reg,data_r_390_sv2v_reg,data_r_389_sv2v_reg,data_r_388_sv2v_reg,
  data_r_387_sv2v_reg,data_r_386_sv2v_reg,data_r_385_sv2v_reg,data_r_384_sv2v_reg,
  data_r_383_sv2v_reg,data_r_382_sv2v_reg,data_r_381_sv2v_reg,data_r_380_sv2v_reg,
  data_r_379_sv2v_reg,data_r_378_sv2v_reg,data_r_377_sv2v_reg,data_r_376_sv2v_reg,
  data_r_375_sv2v_reg,data_r_374_sv2v_reg,data_r_373_sv2v_reg,data_r_372_sv2v_reg,
  data_r_371_sv2v_reg,data_r_370_sv2v_reg,data_r_369_sv2v_reg,data_r_368_sv2v_reg,
  data_r_367_sv2v_reg,data_r_366_sv2v_reg,data_r_365_sv2v_reg,data_r_364_sv2v_reg,
  data_r_363_sv2v_reg,data_r_362_sv2v_reg,data_r_361_sv2v_reg,data_r_360_sv2v_reg,
  data_r_359_sv2v_reg,data_r_358_sv2v_reg,data_r_357_sv2v_reg,data_r_356_sv2v_reg,
  data_r_355_sv2v_reg,data_r_354_sv2v_reg,data_r_353_sv2v_reg,data_r_352_sv2v_reg,
  data_r_351_sv2v_reg,data_r_350_sv2v_reg,data_r_349_sv2v_reg,data_r_348_sv2v_reg,
  data_r_347_sv2v_reg,data_r_346_sv2v_reg,data_r_345_sv2v_reg,data_r_344_sv2v_reg,
  data_r_343_sv2v_reg,data_r_342_sv2v_reg,data_r_341_sv2v_reg,data_r_340_sv2v_reg,
  data_r_339_sv2v_reg,data_r_338_sv2v_reg,data_r_337_sv2v_reg,data_r_336_sv2v_reg,
  data_r_335_sv2v_reg,data_r_334_sv2v_reg,data_r_333_sv2v_reg,data_r_332_sv2v_reg,
  data_r_331_sv2v_reg,data_r_330_sv2v_reg,data_r_329_sv2v_reg,data_r_328_sv2v_reg,
  data_r_327_sv2v_reg,data_r_326_sv2v_reg,data_r_325_sv2v_reg,data_r_324_sv2v_reg,
  data_r_323_sv2v_reg,data_r_322_sv2v_reg,data_r_321_sv2v_reg,data_r_320_sv2v_reg,
  data_r_319_sv2v_reg,data_r_318_sv2v_reg,data_r_317_sv2v_reg,data_r_316_sv2v_reg,
  data_r_315_sv2v_reg,data_r_314_sv2v_reg,data_r_313_sv2v_reg,data_r_312_sv2v_reg,
  data_r_311_sv2v_reg,data_r_310_sv2v_reg,data_r_309_sv2v_reg,data_r_308_sv2v_reg,
  data_r_307_sv2v_reg,data_r_306_sv2v_reg,data_r_305_sv2v_reg,data_r_304_sv2v_reg,
  data_r_303_sv2v_reg,data_r_302_sv2v_reg,data_r_301_sv2v_reg,data_r_300_sv2v_reg,
  data_r_299_sv2v_reg,data_r_298_sv2v_reg,data_r_297_sv2v_reg,data_r_296_sv2v_reg,
  data_r_295_sv2v_reg,data_r_294_sv2v_reg,data_r_293_sv2v_reg,data_r_292_sv2v_reg,
  data_r_291_sv2v_reg,data_r_290_sv2v_reg,data_r_289_sv2v_reg,data_r_288_sv2v_reg,
  data_r_287_sv2v_reg,data_r_286_sv2v_reg,data_r_285_sv2v_reg,data_r_284_sv2v_reg,
  data_r_283_sv2v_reg,data_r_282_sv2v_reg,data_r_281_sv2v_reg,data_r_280_sv2v_reg,
  data_r_279_sv2v_reg,data_r_278_sv2v_reg,data_r_277_sv2v_reg,data_r_276_sv2v_reg,
  data_r_275_sv2v_reg,data_r_274_sv2v_reg,data_r_273_sv2v_reg,data_r_272_sv2v_reg,
  data_r_271_sv2v_reg,data_r_270_sv2v_reg,data_r_269_sv2v_reg,data_r_268_sv2v_reg,
  data_r_267_sv2v_reg,data_r_266_sv2v_reg,data_r_265_sv2v_reg,data_r_264_sv2v_reg,
  data_r_263_sv2v_reg,data_r_262_sv2v_reg,data_r_261_sv2v_reg,data_r_260_sv2v_reg,
  data_r_259_sv2v_reg,data_r_258_sv2v_reg,data_r_257_sv2v_reg,data_r_256_sv2v_reg,
  data_r_255_sv2v_reg,data_r_254_sv2v_reg,data_r_253_sv2v_reg,data_r_252_sv2v_reg,
  data_r_251_sv2v_reg,data_r_250_sv2v_reg,data_r_249_sv2v_reg,data_r_248_sv2v_reg,
  data_r_247_sv2v_reg,data_r_246_sv2v_reg,data_r_245_sv2v_reg,data_r_244_sv2v_reg,
  data_r_243_sv2v_reg,data_r_242_sv2v_reg,data_r_241_sv2v_reg,data_r_240_sv2v_reg,
  data_r_239_sv2v_reg,data_r_238_sv2v_reg,data_r_237_sv2v_reg,data_r_236_sv2v_reg,
  data_r_235_sv2v_reg,data_r_234_sv2v_reg,data_r_233_sv2v_reg,data_r_232_sv2v_reg,
  data_r_231_sv2v_reg,data_r_230_sv2v_reg,data_r_229_sv2v_reg,data_r_228_sv2v_reg,
  data_r_227_sv2v_reg,data_r_226_sv2v_reg,data_r_225_sv2v_reg,data_r_224_sv2v_reg,
  data_r_223_sv2v_reg,data_r_222_sv2v_reg,data_r_221_sv2v_reg,data_r_220_sv2v_reg,
  data_r_219_sv2v_reg,data_r_218_sv2v_reg,data_r_217_sv2v_reg,data_r_216_sv2v_reg,
  data_r_215_sv2v_reg,data_r_214_sv2v_reg,data_r_213_sv2v_reg,data_r_212_sv2v_reg,
  data_r_211_sv2v_reg,data_r_210_sv2v_reg,data_r_209_sv2v_reg,data_r_208_sv2v_reg,
  data_r_207_sv2v_reg,data_r_206_sv2v_reg,data_r_205_sv2v_reg,data_r_204_sv2v_reg,
  data_r_203_sv2v_reg,data_r_202_sv2v_reg,data_r_201_sv2v_reg,data_r_200_sv2v_reg,
  data_r_199_sv2v_reg,data_r_198_sv2v_reg,data_r_197_sv2v_reg,data_r_196_sv2v_reg,
  data_r_195_sv2v_reg,data_r_194_sv2v_reg,data_r_193_sv2v_reg,data_r_192_sv2v_reg,
  data_r_191_sv2v_reg,data_r_190_sv2v_reg,data_r_189_sv2v_reg,data_r_188_sv2v_reg,
  data_r_187_sv2v_reg,data_r_186_sv2v_reg,data_r_185_sv2v_reg,data_r_184_sv2v_reg,
  data_r_183_sv2v_reg,data_r_182_sv2v_reg,data_r_181_sv2v_reg,data_r_180_sv2v_reg,
  data_r_179_sv2v_reg,data_r_178_sv2v_reg,data_r_177_sv2v_reg,data_r_176_sv2v_reg,
  data_r_175_sv2v_reg,data_r_174_sv2v_reg,data_r_173_sv2v_reg,data_r_172_sv2v_reg,
  data_r_171_sv2v_reg,data_r_170_sv2v_reg,data_r_169_sv2v_reg,data_r_168_sv2v_reg,
  data_r_167_sv2v_reg,data_r_166_sv2v_reg,data_r_165_sv2v_reg,data_r_164_sv2v_reg,
  data_r_163_sv2v_reg,data_r_162_sv2v_reg,data_r_161_sv2v_reg,data_r_160_sv2v_reg,
  data_r_159_sv2v_reg,data_r_158_sv2v_reg,data_r_157_sv2v_reg,data_r_156_sv2v_reg,
  data_r_155_sv2v_reg,data_r_154_sv2v_reg,data_r_153_sv2v_reg,data_r_152_sv2v_reg,
  data_r_151_sv2v_reg,data_r_150_sv2v_reg,data_r_149_sv2v_reg,data_r_148_sv2v_reg,
  data_r_147_sv2v_reg,data_r_146_sv2v_reg,data_r_145_sv2v_reg,data_r_144_sv2v_reg,
  data_r_143_sv2v_reg,data_r_142_sv2v_reg,data_r_141_sv2v_reg,data_r_140_sv2v_reg,
  data_r_139_sv2v_reg,data_r_138_sv2v_reg,data_r_137_sv2v_reg,data_r_136_sv2v_reg,
  data_r_135_sv2v_reg,data_r_134_sv2v_reg,data_r_133_sv2v_reg,data_r_132_sv2v_reg,
  data_r_131_sv2v_reg,data_r_130_sv2v_reg,data_r_129_sv2v_reg,data_r_128_sv2v_reg,
  data_r_127_sv2v_reg,data_r_126_sv2v_reg,data_r_125_sv2v_reg,data_r_124_sv2v_reg,
  data_r_123_sv2v_reg,data_r_122_sv2v_reg,data_r_121_sv2v_reg,data_r_120_sv2v_reg,
  data_r_119_sv2v_reg,data_r_118_sv2v_reg,data_r_117_sv2v_reg,data_r_116_sv2v_reg,
  data_r_115_sv2v_reg,data_r_114_sv2v_reg,data_r_113_sv2v_reg,data_r_112_sv2v_reg,
  data_r_111_sv2v_reg,data_r_110_sv2v_reg,data_r_109_sv2v_reg,data_r_108_sv2v_reg,
  data_r_107_sv2v_reg,data_r_106_sv2v_reg,data_r_105_sv2v_reg,data_r_104_sv2v_reg,
  data_r_103_sv2v_reg,data_r_102_sv2v_reg,data_r_101_sv2v_reg,data_r_100_sv2v_reg,
  data_r_99_sv2v_reg,data_r_98_sv2v_reg,data_r_97_sv2v_reg,data_r_96_sv2v_reg,data_r_95_sv2v_reg,
  data_r_94_sv2v_reg,data_r_93_sv2v_reg,data_r_92_sv2v_reg,data_r_91_sv2v_reg,
  data_r_90_sv2v_reg,data_r_89_sv2v_reg,data_r_88_sv2v_reg,data_r_87_sv2v_reg,
  data_r_86_sv2v_reg,data_r_85_sv2v_reg,data_r_84_sv2v_reg,data_r_83_sv2v_reg,
  data_r_82_sv2v_reg,data_r_81_sv2v_reg,data_r_80_sv2v_reg,data_r_79_sv2v_reg,
  data_r_78_sv2v_reg,data_r_77_sv2v_reg,data_r_76_sv2v_reg,data_r_75_sv2v_reg,data_r_74_sv2v_reg,
  data_r_73_sv2v_reg,data_r_72_sv2v_reg,data_r_71_sv2v_reg,data_r_70_sv2v_reg,
  data_r_69_sv2v_reg,data_r_68_sv2v_reg,data_r_67_sv2v_reg,data_r_66_sv2v_reg,
  data_r_65_sv2v_reg,data_r_64_sv2v_reg,data_r_63_sv2v_reg,data_r_62_sv2v_reg,
  data_r_61_sv2v_reg,data_r_60_sv2v_reg,data_r_59_sv2v_reg,data_r_58_sv2v_reg,
  data_r_57_sv2v_reg,data_r_56_sv2v_reg,data_r_55_sv2v_reg,data_r_54_sv2v_reg,data_r_53_sv2v_reg,
  data_r_52_sv2v_reg,data_r_51_sv2v_reg,data_r_50_sv2v_reg,data_r_49_sv2v_reg,
  data_r_48_sv2v_reg,data_r_47_sv2v_reg,data_r_46_sv2v_reg,data_r_45_sv2v_reg,
  data_r_44_sv2v_reg,data_r_43_sv2v_reg,data_r_42_sv2v_reg,data_r_41_sv2v_reg,
  data_r_40_sv2v_reg,data_r_39_sv2v_reg,data_r_38_sv2v_reg,data_r_37_sv2v_reg,
  data_r_36_sv2v_reg,data_r_35_sv2v_reg,data_r_34_sv2v_reg,data_r_33_sv2v_reg,data_r_32_sv2v_reg,
  data_r_31_sv2v_reg,data_r_30_sv2v_reg,data_r_29_sv2v_reg,data_r_28_sv2v_reg,
  data_r_27_sv2v_reg,data_r_26_sv2v_reg,data_r_25_sv2v_reg,data_r_24_sv2v_reg,
  data_r_23_sv2v_reg,data_r_22_sv2v_reg,data_r_21_sv2v_reg,data_r_20_sv2v_reg,
  data_r_19_sv2v_reg,data_r_18_sv2v_reg,data_r_17_sv2v_reg,data_r_16_sv2v_reg,data_r_15_sv2v_reg,
  data_r_14_sv2v_reg,data_r_13_sv2v_reg,data_r_12_sv2v_reg,data_r_11_sv2v_reg,
  data_r_10_sv2v_reg,data_r_9_sv2v_reg,data_r_8_sv2v_reg,data_r_7_sv2v_reg,
  data_r_6_sv2v_reg,data_r_5_sv2v_reg,data_r_4_sv2v_reg,data_r_3_sv2v_reg,data_r_2_sv2v_reg,
  data_r_1_sv2v_reg,data_r_0_sv2v_reg;
  assign valid_r[63] = valid_r_63_sv2v_reg;
  assign valid_r[62] = valid_r_62_sv2v_reg;
  assign valid_r[61] = valid_r_61_sv2v_reg;
  assign valid_r[60] = valid_r_60_sv2v_reg;
  assign valid_r[59] = valid_r_59_sv2v_reg;
  assign valid_r[58] = valid_r_58_sv2v_reg;
  assign valid_r[57] = valid_r_57_sv2v_reg;
  assign valid_r[56] = valid_r_56_sv2v_reg;
  assign valid_r[55] = valid_r_55_sv2v_reg;
  assign valid_r[54] = valid_r_54_sv2v_reg;
  assign valid_r[53] = valid_r_53_sv2v_reg;
  assign valid_r[52] = valid_r_52_sv2v_reg;
  assign valid_r[51] = valid_r_51_sv2v_reg;
  assign valid_r[50] = valid_r_50_sv2v_reg;
  assign valid_r[49] = valid_r_49_sv2v_reg;
  assign valid_r[48] = valid_r_48_sv2v_reg;
  assign valid_r[47] = valid_r_47_sv2v_reg;
  assign valid_r[46] = valid_r_46_sv2v_reg;
  assign valid_r[45] = valid_r_45_sv2v_reg;
  assign valid_r[44] = valid_r_44_sv2v_reg;
  assign valid_r[43] = valid_r_43_sv2v_reg;
  assign valid_r[42] = valid_r_42_sv2v_reg;
  assign valid_r[41] = valid_r_41_sv2v_reg;
  assign valid_r[40] = valid_r_40_sv2v_reg;
  assign valid_r[39] = valid_r_39_sv2v_reg;
  assign valid_r[38] = valid_r_38_sv2v_reg;
  assign valid_r[37] = valid_r_37_sv2v_reg;
  assign valid_r[36] = valid_r_36_sv2v_reg;
  assign valid_r[35] = valid_r_35_sv2v_reg;
  assign valid_r[34] = valid_r_34_sv2v_reg;
  assign valid_r[33] = valid_r_33_sv2v_reg;
  assign valid_r[32] = valid_r_32_sv2v_reg;
  assign valid_r[31] = valid_r_31_sv2v_reg;
  assign valid_r[30] = valid_r_30_sv2v_reg;
  assign valid_r[29] = valid_r_29_sv2v_reg;
  assign valid_r[28] = valid_r_28_sv2v_reg;
  assign valid_r[27] = valid_r_27_sv2v_reg;
  assign valid_r[26] = valid_r_26_sv2v_reg;
  assign valid_r[25] = valid_r_25_sv2v_reg;
  assign valid_r[24] = valid_r_24_sv2v_reg;
  assign valid_r[23] = valid_r_23_sv2v_reg;
  assign valid_r[22] = valid_r_22_sv2v_reg;
  assign valid_r[21] = valid_r_21_sv2v_reg;
  assign valid_r[20] = valid_r_20_sv2v_reg;
  assign valid_r[19] = valid_r_19_sv2v_reg;
  assign valid_r[18] = valid_r_18_sv2v_reg;
  assign valid_r[17] = valid_r_17_sv2v_reg;
  assign valid_r[16] = valid_r_16_sv2v_reg;
  assign valid_r[15] = valid_r_15_sv2v_reg;
  assign valid_r[14] = valid_r_14_sv2v_reg;
  assign valid_r[13] = valid_r_13_sv2v_reg;
  assign valid_r[12] = valid_r_12_sv2v_reg;
  assign valid_r[11] = valid_r_11_sv2v_reg;
  assign valid_r[10] = valid_r_10_sv2v_reg;
  assign valid_r[9] = valid_r_9_sv2v_reg;
  assign valid_r[8] = valid_r_8_sv2v_reg;
  assign valid_r[7] = valid_r_7_sv2v_reg;
  assign valid_r[6] = valid_r_6_sv2v_reg;
  assign valid_r[5] = valid_r_5_sv2v_reg;
  assign valid_r[4] = valid_r_4_sv2v_reg;
  assign valid_r[3] = valid_r_3_sv2v_reg;
  assign valid_r[2] = valid_r_2_sv2v_reg;
  assign valid_r[1] = valid_r_1_sv2v_reg;
  assign valid_r[0] = valid_r_0_sv2v_reg;
  assign num_els_r[6] = num_els_r_6_sv2v_reg;
  assign num_els_r[5] = num_els_r_5_sv2v_reg;
  assign num_els_r[4] = num_els_r_4_sv2v_reg;
  assign num_els_r[3] = num_els_r_3_sv2v_reg;
  assign num_els_r[2] = num_els_r_2_sv2v_reg;
  assign num_els_r[1] = num_els_r_1_sv2v_reg;
  assign num_els_r[0] = num_els_r_0_sv2v_reg;
  assign data_r[2047] = data_r_2047_sv2v_reg;
  assign data_r[2046] = data_r_2046_sv2v_reg;
  assign data_r[2045] = data_r_2045_sv2v_reg;
  assign data_r[2044] = data_r_2044_sv2v_reg;
  assign data_r[2043] = data_r_2043_sv2v_reg;
  assign data_r[2042] = data_r_2042_sv2v_reg;
  assign data_r[2041] = data_r_2041_sv2v_reg;
  assign data_r[2040] = data_r_2040_sv2v_reg;
  assign data_r[2039] = data_r_2039_sv2v_reg;
  assign data_r[2038] = data_r_2038_sv2v_reg;
  assign data_r[2037] = data_r_2037_sv2v_reg;
  assign data_r[2036] = data_r_2036_sv2v_reg;
  assign data_r[2035] = data_r_2035_sv2v_reg;
  assign data_r[2034] = data_r_2034_sv2v_reg;
  assign data_r[2033] = data_r_2033_sv2v_reg;
  assign data_r[2032] = data_r_2032_sv2v_reg;
  assign data_r[2031] = data_r_2031_sv2v_reg;
  assign data_r[2030] = data_r_2030_sv2v_reg;
  assign data_r[2029] = data_r_2029_sv2v_reg;
  assign data_r[2028] = data_r_2028_sv2v_reg;
  assign data_r[2027] = data_r_2027_sv2v_reg;
  assign data_r[2026] = data_r_2026_sv2v_reg;
  assign data_r[2025] = data_r_2025_sv2v_reg;
  assign data_r[2024] = data_r_2024_sv2v_reg;
  assign data_r[2023] = data_r_2023_sv2v_reg;
  assign data_r[2022] = data_r_2022_sv2v_reg;
  assign data_r[2021] = data_r_2021_sv2v_reg;
  assign data_r[2020] = data_r_2020_sv2v_reg;
  assign data_r[2019] = data_r_2019_sv2v_reg;
  assign data_r[2018] = data_r_2018_sv2v_reg;
  assign data_r[2017] = data_r_2017_sv2v_reg;
  assign data_r[2016] = data_r_2016_sv2v_reg;
  assign data_r[2015] = data_r_2015_sv2v_reg;
  assign data_r[2014] = data_r_2014_sv2v_reg;
  assign data_r[2013] = data_r_2013_sv2v_reg;
  assign data_r[2012] = data_r_2012_sv2v_reg;
  assign data_r[2011] = data_r_2011_sv2v_reg;
  assign data_r[2010] = data_r_2010_sv2v_reg;
  assign data_r[2009] = data_r_2009_sv2v_reg;
  assign data_r[2008] = data_r_2008_sv2v_reg;
  assign data_r[2007] = data_r_2007_sv2v_reg;
  assign data_r[2006] = data_r_2006_sv2v_reg;
  assign data_r[2005] = data_r_2005_sv2v_reg;
  assign data_r[2004] = data_r_2004_sv2v_reg;
  assign data_r[2003] = data_r_2003_sv2v_reg;
  assign data_r[2002] = data_r_2002_sv2v_reg;
  assign data_r[2001] = data_r_2001_sv2v_reg;
  assign data_r[2000] = data_r_2000_sv2v_reg;
  assign data_r[1999] = data_r_1999_sv2v_reg;
  assign data_r[1998] = data_r_1998_sv2v_reg;
  assign data_r[1997] = data_r_1997_sv2v_reg;
  assign data_r[1996] = data_r_1996_sv2v_reg;
  assign data_r[1995] = data_r_1995_sv2v_reg;
  assign data_r[1994] = data_r_1994_sv2v_reg;
  assign data_r[1993] = data_r_1993_sv2v_reg;
  assign data_r[1992] = data_r_1992_sv2v_reg;
  assign data_r[1991] = data_r_1991_sv2v_reg;
  assign data_r[1990] = data_r_1990_sv2v_reg;
  assign data_r[1989] = data_r_1989_sv2v_reg;
  assign data_r[1988] = data_r_1988_sv2v_reg;
  assign data_r[1987] = data_r_1987_sv2v_reg;
  assign data_r[1986] = data_r_1986_sv2v_reg;
  assign data_r[1985] = data_r_1985_sv2v_reg;
  assign data_r[1984] = data_r_1984_sv2v_reg;
  assign data_r[1983] = data_r_1983_sv2v_reg;
  assign data_r[1982] = data_r_1982_sv2v_reg;
  assign data_r[1981] = data_r_1981_sv2v_reg;
  assign data_r[1980] = data_r_1980_sv2v_reg;
  assign data_r[1979] = data_r_1979_sv2v_reg;
  assign data_r[1978] = data_r_1978_sv2v_reg;
  assign data_r[1977] = data_r_1977_sv2v_reg;
  assign data_r[1976] = data_r_1976_sv2v_reg;
  assign data_r[1975] = data_r_1975_sv2v_reg;
  assign data_r[1974] = data_r_1974_sv2v_reg;
  assign data_r[1973] = data_r_1973_sv2v_reg;
  assign data_r[1972] = data_r_1972_sv2v_reg;
  assign data_r[1971] = data_r_1971_sv2v_reg;
  assign data_r[1970] = data_r_1970_sv2v_reg;
  assign data_r[1969] = data_r_1969_sv2v_reg;
  assign data_r[1968] = data_r_1968_sv2v_reg;
  assign data_r[1967] = data_r_1967_sv2v_reg;
  assign data_r[1966] = data_r_1966_sv2v_reg;
  assign data_r[1965] = data_r_1965_sv2v_reg;
  assign data_r[1964] = data_r_1964_sv2v_reg;
  assign data_r[1963] = data_r_1963_sv2v_reg;
  assign data_r[1962] = data_r_1962_sv2v_reg;
  assign data_r[1961] = data_r_1961_sv2v_reg;
  assign data_r[1960] = data_r_1960_sv2v_reg;
  assign data_r[1959] = data_r_1959_sv2v_reg;
  assign data_r[1958] = data_r_1958_sv2v_reg;
  assign data_r[1957] = data_r_1957_sv2v_reg;
  assign data_r[1956] = data_r_1956_sv2v_reg;
  assign data_r[1955] = data_r_1955_sv2v_reg;
  assign data_r[1954] = data_r_1954_sv2v_reg;
  assign data_r[1953] = data_r_1953_sv2v_reg;
  assign data_r[1952] = data_r_1952_sv2v_reg;
  assign data_r[1951] = data_r_1951_sv2v_reg;
  assign data_r[1950] = data_r_1950_sv2v_reg;
  assign data_r[1949] = data_r_1949_sv2v_reg;
  assign data_r[1948] = data_r_1948_sv2v_reg;
  assign data_r[1947] = data_r_1947_sv2v_reg;
  assign data_r[1946] = data_r_1946_sv2v_reg;
  assign data_r[1945] = data_r_1945_sv2v_reg;
  assign data_r[1944] = data_r_1944_sv2v_reg;
  assign data_r[1943] = data_r_1943_sv2v_reg;
  assign data_r[1942] = data_r_1942_sv2v_reg;
  assign data_r[1941] = data_r_1941_sv2v_reg;
  assign data_r[1940] = data_r_1940_sv2v_reg;
  assign data_r[1939] = data_r_1939_sv2v_reg;
  assign data_r[1938] = data_r_1938_sv2v_reg;
  assign data_r[1937] = data_r_1937_sv2v_reg;
  assign data_r[1936] = data_r_1936_sv2v_reg;
  assign data_r[1935] = data_r_1935_sv2v_reg;
  assign data_r[1934] = data_r_1934_sv2v_reg;
  assign data_r[1933] = data_r_1933_sv2v_reg;
  assign data_r[1932] = data_r_1932_sv2v_reg;
  assign data_r[1931] = data_r_1931_sv2v_reg;
  assign data_r[1930] = data_r_1930_sv2v_reg;
  assign data_r[1929] = data_r_1929_sv2v_reg;
  assign data_r[1928] = data_r_1928_sv2v_reg;
  assign data_r[1927] = data_r_1927_sv2v_reg;
  assign data_r[1926] = data_r_1926_sv2v_reg;
  assign data_r[1925] = data_r_1925_sv2v_reg;
  assign data_r[1924] = data_r_1924_sv2v_reg;
  assign data_r[1923] = data_r_1923_sv2v_reg;
  assign data_r[1922] = data_r_1922_sv2v_reg;
  assign data_r[1921] = data_r_1921_sv2v_reg;
  assign data_r[1920] = data_r_1920_sv2v_reg;
  assign data_r[1919] = data_r_1919_sv2v_reg;
  assign data_r[1918] = data_r_1918_sv2v_reg;
  assign data_r[1917] = data_r_1917_sv2v_reg;
  assign data_r[1916] = data_r_1916_sv2v_reg;
  assign data_r[1915] = data_r_1915_sv2v_reg;
  assign data_r[1914] = data_r_1914_sv2v_reg;
  assign data_r[1913] = data_r_1913_sv2v_reg;
  assign data_r[1912] = data_r_1912_sv2v_reg;
  assign data_r[1911] = data_r_1911_sv2v_reg;
  assign data_r[1910] = data_r_1910_sv2v_reg;
  assign data_r[1909] = data_r_1909_sv2v_reg;
  assign data_r[1908] = data_r_1908_sv2v_reg;
  assign data_r[1907] = data_r_1907_sv2v_reg;
  assign data_r[1906] = data_r_1906_sv2v_reg;
  assign data_r[1905] = data_r_1905_sv2v_reg;
  assign data_r[1904] = data_r_1904_sv2v_reg;
  assign data_r[1903] = data_r_1903_sv2v_reg;
  assign data_r[1902] = data_r_1902_sv2v_reg;
  assign data_r[1901] = data_r_1901_sv2v_reg;
  assign data_r[1900] = data_r_1900_sv2v_reg;
  assign data_r[1899] = data_r_1899_sv2v_reg;
  assign data_r[1898] = data_r_1898_sv2v_reg;
  assign data_r[1897] = data_r_1897_sv2v_reg;
  assign data_r[1896] = data_r_1896_sv2v_reg;
  assign data_r[1895] = data_r_1895_sv2v_reg;
  assign data_r[1894] = data_r_1894_sv2v_reg;
  assign data_r[1893] = data_r_1893_sv2v_reg;
  assign data_r[1892] = data_r_1892_sv2v_reg;
  assign data_r[1891] = data_r_1891_sv2v_reg;
  assign data_r[1890] = data_r_1890_sv2v_reg;
  assign data_r[1889] = data_r_1889_sv2v_reg;
  assign data_r[1888] = data_r_1888_sv2v_reg;
  assign data_r[1887] = data_r_1887_sv2v_reg;
  assign data_r[1886] = data_r_1886_sv2v_reg;
  assign data_r[1885] = data_r_1885_sv2v_reg;
  assign data_r[1884] = data_r_1884_sv2v_reg;
  assign data_r[1883] = data_r_1883_sv2v_reg;
  assign data_r[1882] = data_r_1882_sv2v_reg;
  assign data_r[1881] = data_r_1881_sv2v_reg;
  assign data_r[1880] = data_r_1880_sv2v_reg;
  assign data_r[1879] = data_r_1879_sv2v_reg;
  assign data_r[1878] = data_r_1878_sv2v_reg;
  assign data_r[1877] = data_r_1877_sv2v_reg;
  assign data_r[1876] = data_r_1876_sv2v_reg;
  assign data_r[1875] = data_r_1875_sv2v_reg;
  assign data_r[1874] = data_r_1874_sv2v_reg;
  assign data_r[1873] = data_r_1873_sv2v_reg;
  assign data_r[1872] = data_r_1872_sv2v_reg;
  assign data_r[1871] = data_r_1871_sv2v_reg;
  assign data_r[1870] = data_r_1870_sv2v_reg;
  assign data_r[1869] = data_r_1869_sv2v_reg;
  assign data_r[1868] = data_r_1868_sv2v_reg;
  assign data_r[1867] = data_r_1867_sv2v_reg;
  assign data_r[1866] = data_r_1866_sv2v_reg;
  assign data_r[1865] = data_r_1865_sv2v_reg;
  assign data_r[1864] = data_r_1864_sv2v_reg;
  assign data_r[1863] = data_r_1863_sv2v_reg;
  assign data_r[1862] = data_r_1862_sv2v_reg;
  assign data_r[1861] = data_r_1861_sv2v_reg;
  assign data_r[1860] = data_r_1860_sv2v_reg;
  assign data_r[1859] = data_r_1859_sv2v_reg;
  assign data_r[1858] = data_r_1858_sv2v_reg;
  assign data_r[1857] = data_r_1857_sv2v_reg;
  assign data_r[1856] = data_r_1856_sv2v_reg;
  assign data_r[1855] = data_r_1855_sv2v_reg;
  assign data_r[1854] = data_r_1854_sv2v_reg;
  assign data_r[1853] = data_r_1853_sv2v_reg;
  assign data_r[1852] = data_r_1852_sv2v_reg;
  assign data_r[1851] = data_r_1851_sv2v_reg;
  assign data_r[1850] = data_r_1850_sv2v_reg;
  assign data_r[1849] = data_r_1849_sv2v_reg;
  assign data_r[1848] = data_r_1848_sv2v_reg;
  assign data_r[1847] = data_r_1847_sv2v_reg;
  assign data_r[1846] = data_r_1846_sv2v_reg;
  assign data_r[1845] = data_r_1845_sv2v_reg;
  assign data_r[1844] = data_r_1844_sv2v_reg;
  assign data_r[1843] = data_r_1843_sv2v_reg;
  assign data_r[1842] = data_r_1842_sv2v_reg;
  assign data_r[1841] = data_r_1841_sv2v_reg;
  assign data_r[1840] = data_r_1840_sv2v_reg;
  assign data_r[1839] = data_r_1839_sv2v_reg;
  assign data_r[1838] = data_r_1838_sv2v_reg;
  assign data_r[1837] = data_r_1837_sv2v_reg;
  assign data_r[1836] = data_r_1836_sv2v_reg;
  assign data_r[1835] = data_r_1835_sv2v_reg;
  assign data_r[1834] = data_r_1834_sv2v_reg;
  assign data_r[1833] = data_r_1833_sv2v_reg;
  assign data_r[1832] = data_r_1832_sv2v_reg;
  assign data_r[1831] = data_r_1831_sv2v_reg;
  assign data_r[1830] = data_r_1830_sv2v_reg;
  assign data_r[1829] = data_r_1829_sv2v_reg;
  assign data_r[1828] = data_r_1828_sv2v_reg;
  assign data_r[1827] = data_r_1827_sv2v_reg;
  assign data_r[1826] = data_r_1826_sv2v_reg;
  assign data_r[1825] = data_r_1825_sv2v_reg;
  assign data_r[1824] = data_r_1824_sv2v_reg;
  assign data_r[1823] = data_r_1823_sv2v_reg;
  assign data_r[1822] = data_r_1822_sv2v_reg;
  assign data_r[1821] = data_r_1821_sv2v_reg;
  assign data_r[1820] = data_r_1820_sv2v_reg;
  assign data_r[1819] = data_r_1819_sv2v_reg;
  assign data_r[1818] = data_r_1818_sv2v_reg;
  assign data_r[1817] = data_r_1817_sv2v_reg;
  assign data_r[1816] = data_r_1816_sv2v_reg;
  assign data_r[1815] = data_r_1815_sv2v_reg;
  assign data_r[1814] = data_r_1814_sv2v_reg;
  assign data_r[1813] = data_r_1813_sv2v_reg;
  assign data_r[1812] = data_r_1812_sv2v_reg;
  assign data_r[1811] = data_r_1811_sv2v_reg;
  assign data_r[1810] = data_r_1810_sv2v_reg;
  assign data_r[1809] = data_r_1809_sv2v_reg;
  assign data_r[1808] = data_r_1808_sv2v_reg;
  assign data_r[1807] = data_r_1807_sv2v_reg;
  assign data_r[1806] = data_r_1806_sv2v_reg;
  assign data_r[1805] = data_r_1805_sv2v_reg;
  assign data_r[1804] = data_r_1804_sv2v_reg;
  assign data_r[1803] = data_r_1803_sv2v_reg;
  assign data_r[1802] = data_r_1802_sv2v_reg;
  assign data_r[1801] = data_r_1801_sv2v_reg;
  assign data_r[1800] = data_r_1800_sv2v_reg;
  assign data_r[1799] = data_r_1799_sv2v_reg;
  assign data_r[1798] = data_r_1798_sv2v_reg;
  assign data_r[1797] = data_r_1797_sv2v_reg;
  assign data_r[1796] = data_r_1796_sv2v_reg;
  assign data_r[1795] = data_r_1795_sv2v_reg;
  assign data_r[1794] = data_r_1794_sv2v_reg;
  assign data_r[1793] = data_r_1793_sv2v_reg;
  assign data_r[1792] = data_r_1792_sv2v_reg;
  assign data_r[1791] = data_r_1791_sv2v_reg;
  assign data_r[1790] = data_r_1790_sv2v_reg;
  assign data_r[1789] = data_r_1789_sv2v_reg;
  assign data_r[1788] = data_r_1788_sv2v_reg;
  assign data_r[1787] = data_r_1787_sv2v_reg;
  assign data_r[1786] = data_r_1786_sv2v_reg;
  assign data_r[1785] = data_r_1785_sv2v_reg;
  assign data_r[1784] = data_r_1784_sv2v_reg;
  assign data_r[1783] = data_r_1783_sv2v_reg;
  assign data_r[1782] = data_r_1782_sv2v_reg;
  assign data_r[1781] = data_r_1781_sv2v_reg;
  assign data_r[1780] = data_r_1780_sv2v_reg;
  assign data_r[1779] = data_r_1779_sv2v_reg;
  assign data_r[1778] = data_r_1778_sv2v_reg;
  assign data_r[1777] = data_r_1777_sv2v_reg;
  assign data_r[1776] = data_r_1776_sv2v_reg;
  assign data_r[1775] = data_r_1775_sv2v_reg;
  assign data_r[1774] = data_r_1774_sv2v_reg;
  assign data_r[1773] = data_r_1773_sv2v_reg;
  assign data_r[1772] = data_r_1772_sv2v_reg;
  assign data_r[1771] = data_r_1771_sv2v_reg;
  assign data_r[1770] = data_r_1770_sv2v_reg;
  assign data_r[1769] = data_r_1769_sv2v_reg;
  assign data_r[1768] = data_r_1768_sv2v_reg;
  assign data_r[1767] = data_r_1767_sv2v_reg;
  assign data_r[1766] = data_r_1766_sv2v_reg;
  assign data_r[1765] = data_r_1765_sv2v_reg;
  assign data_r[1764] = data_r_1764_sv2v_reg;
  assign data_r[1763] = data_r_1763_sv2v_reg;
  assign data_r[1762] = data_r_1762_sv2v_reg;
  assign data_r[1761] = data_r_1761_sv2v_reg;
  assign data_r[1760] = data_r_1760_sv2v_reg;
  assign data_r[1759] = data_r_1759_sv2v_reg;
  assign data_r[1758] = data_r_1758_sv2v_reg;
  assign data_r[1757] = data_r_1757_sv2v_reg;
  assign data_r[1756] = data_r_1756_sv2v_reg;
  assign data_r[1755] = data_r_1755_sv2v_reg;
  assign data_r[1754] = data_r_1754_sv2v_reg;
  assign data_r[1753] = data_r_1753_sv2v_reg;
  assign data_r[1752] = data_r_1752_sv2v_reg;
  assign data_r[1751] = data_r_1751_sv2v_reg;
  assign data_r[1750] = data_r_1750_sv2v_reg;
  assign data_r[1749] = data_r_1749_sv2v_reg;
  assign data_r[1748] = data_r_1748_sv2v_reg;
  assign data_r[1747] = data_r_1747_sv2v_reg;
  assign data_r[1746] = data_r_1746_sv2v_reg;
  assign data_r[1745] = data_r_1745_sv2v_reg;
  assign data_r[1744] = data_r_1744_sv2v_reg;
  assign data_r[1743] = data_r_1743_sv2v_reg;
  assign data_r[1742] = data_r_1742_sv2v_reg;
  assign data_r[1741] = data_r_1741_sv2v_reg;
  assign data_r[1740] = data_r_1740_sv2v_reg;
  assign data_r[1739] = data_r_1739_sv2v_reg;
  assign data_r[1738] = data_r_1738_sv2v_reg;
  assign data_r[1737] = data_r_1737_sv2v_reg;
  assign data_r[1736] = data_r_1736_sv2v_reg;
  assign data_r[1735] = data_r_1735_sv2v_reg;
  assign data_r[1734] = data_r_1734_sv2v_reg;
  assign data_r[1733] = data_r_1733_sv2v_reg;
  assign data_r[1732] = data_r_1732_sv2v_reg;
  assign data_r[1731] = data_r_1731_sv2v_reg;
  assign data_r[1730] = data_r_1730_sv2v_reg;
  assign data_r[1729] = data_r_1729_sv2v_reg;
  assign data_r[1728] = data_r_1728_sv2v_reg;
  assign data_r[1727] = data_r_1727_sv2v_reg;
  assign data_r[1726] = data_r_1726_sv2v_reg;
  assign data_r[1725] = data_r_1725_sv2v_reg;
  assign data_r[1724] = data_r_1724_sv2v_reg;
  assign data_r[1723] = data_r_1723_sv2v_reg;
  assign data_r[1722] = data_r_1722_sv2v_reg;
  assign data_r[1721] = data_r_1721_sv2v_reg;
  assign data_r[1720] = data_r_1720_sv2v_reg;
  assign data_r[1719] = data_r_1719_sv2v_reg;
  assign data_r[1718] = data_r_1718_sv2v_reg;
  assign data_r[1717] = data_r_1717_sv2v_reg;
  assign data_r[1716] = data_r_1716_sv2v_reg;
  assign data_r[1715] = data_r_1715_sv2v_reg;
  assign data_r[1714] = data_r_1714_sv2v_reg;
  assign data_r[1713] = data_r_1713_sv2v_reg;
  assign data_r[1712] = data_r_1712_sv2v_reg;
  assign data_r[1711] = data_r_1711_sv2v_reg;
  assign data_r[1710] = data_r_1710_sv2v_reg;
  assign data_r[1709] = data_r_1709_sv2v_reg;
  assign data_r[1708] = data_r_1708_sv2v_reg;
  assign data_r[1707] = data_r_1707_sv2v_reg;
  assign data_r[1706] = data_r_1706_sv2v_reg;
  assign data_r[1705] = data_r_1705_sv2v_reg;
  assign data_r[1704] = data_r_1704_sv2v_reg;
  assign data_r[1703] = data_r_1703_sv2v_reg;
  assign data_r[1702] = data_r_1702_sv2v_reg;
  assign data_r[1701] = data_r_1701_sv2v_reg;
  assign data_r[1700] = data_r_1700_sv2v_reg;
  assign data_r[1699] = data_r_1699_sv2v_reg;
  assign data_r[1698] = data_r_1698_sv2v_reg;
  assign data_r[1697] = data_r_1697_sv2v_reg;
  assign data_r[1696] = data_r_1696_sv2v_reg;
  assign data_r[1695] = data_r_1695_sv2v_reg;
  assign data_r[1694] = data_r_1694_sv2v_reg;
  assign data_r[1693] = data_r_1693_sv2v_reg;
  assign data_r[1692] = data_r_1692_sv2v_reg;
  assign data_r[1691] = data_r_1691_sv2v_reg;
  assign data_r[1690] = data_r_1690_sv2v_reg;
  assign data_r[1689] = data_r_1689_sv2v_reg;
  assign data_r[1688] = data_r_1688_sv2v_reg;
  assign data_r[1687] = data_r_1687_sv2v_reg;
  assign data_r[1686] = data_r_1686_sv2v_reg;
  assign data_r[1685] = data_r_1685_sv2v_reg;
  assign data_r[1684] = data_r_1684_sv2v_reg;
  assign data_r[1683] = data_r_1683_sv2v_reg;
  assign data_r[1682] = data_r_1682_sv2v_reg;
  assign data_r[1681] = data_r_1681_sv2v_reg;
  assign data_r[1680] = data_r_1680_sv2v_reg;
  assign data_r[1679] = data_r_1679_sv2v_reg;
  assign data_r[1678] = data_r_1678_sv2v_reg;
  assign data_r[1677] = data_r_1677_sv2v_reg;
  assign data_r[1676] = data_r_1676_sv2v_reg;
  assign data_r[1675] = data_r_1675_sv2v_reg;
  assign data_r[1674] = data_r_1674_sv2v_reg;
  assign data_r[1673] = data_r_1673_sv2v_reg;
  assign data_r[1672] = data_r_1672_sv2v_reg;
  assign data_r[1671] = data_r_1671_sv2v_reg;
  assign data_r[1670] = data_r_1670_sv2v_reg;
  assign data_r[1669] = data_r_1669_sv2v_reg;
  assign data_r[1668] = data_r_1668_sv2v_reg;
  assign data_r[1667] = data_r_1667_sv2v_reg;
  assign data_r[1666] = data_r_1666_sv2v_reg;
  assign data_r[1665] = data_r_1665_sv2v_reg;
  assign data_r[1664] = data_r_1664_sv2v_reg;
  assign data_r[1663] = data_r_1663_sv2v_reg;
  assign data_r[1662] = data_r_1662_sv2v_reg;
  assign data_r[1661] = data_r_1661_sv2v_reg;
  assign data_r[1660] = data_r_1660_sv2v_reg;
  assign data_r[1659] = data_r_1659_sv2v_reg;
  assign data_r[1658] = data_r_1658_sv2v_reg;
  assign data_r[1657] = data_r_1657_sv2v_reg;
  assign data_r[1656] = data_r_1656_sv2v_reg;
  assign data_r[1655] = data_r_1655_sv2v_reg;
  assign data_r[1654] = data_r_1654_sv2v_reg;
  assign data_r[1653] = data_r_1653_sv2v_reg;
  assign data_r[1652] = data_r_1652_sv2v_reg;
  assign data_r[1651] = data_r_1651_sv2v_reg;
  assign data_r[1650] = data_r_1650_sv2v_reg;
  assign data_r[1649] = data_r_1649_sv2v_reg;
  assign data_r[1648] = data_r_1648_sv2v_reg;
  assign data_r[1647] = data_r_1647_sv2v_reg;
  assign data_r[1646] = data_r_1646_sv2v_reg;
  assign data_r[1645] = data_r_1645_sv2v_reg;
  assign data_r[1644] = data_r_1644_sv2v_reg;
  assign data_r[1643] = data_r_1643_sv2v_reg;
  assign data_r[1642] = data_r_1642_sv2v_reg;
  assign data_r[1641] = data_r_1641_sv2v_reg;
  assign data_r[1640] = data_r_1640_sv2v_reg;
  assign data_r[1639] = data_r_1639_sv2v_reg;
  assign data_r[1638] = data_r_1638_sv2v_reg;
  assign data_r[1637] = data_r_1637_sv2v_reg;
  assign data_r[1636] = data_r_1636_sv2v_reg;
  assign data_r[1635] = data_r_1635_sv2v_reg;
  assign data_r[1634] = data_r_1634_sv2v_reg;
  assign data_r[1633] = data_r_1633_sv2v_reg;
  assign data_r[1632] = data_r_1632_sv2v_reg;
  assign data_r[1631] = data_r_1631_sv2v_reg;
  assign data_r[1630] = data_r_1630_sv2v_reg;
  assign data_r[1629] = data_r_1629_sv2v_reg;
  assign data_r[1628] = data_r_1628_sv2v_reg;
  assign data_r[1627] = data_r_1627_sv2v_reg;
  assign data_r[1626] = data_r_1626_sv2v_reg;
  assign data_r[1625] = data_r_1625_sv2v_reg;
  assign data_r[1624] = data_r_1624_sv2v_reg;
  assign data_r[1623] = data_r_1623_sv2v_reg;
  assign data_r[1622] = data_r_1622_sv2v_reg;
  assign data_r[1621] = data_r_1621_sv2v_reg;
  assign data_r[1620] = data_r_1620_sv2v_reg;
  assign data_r[1619] = data_r_1619_sv2v_reg;
  assign data_r[1618] = data_r_1618_sv2v_reg;
  assign data_r[1617] = data_r_1617_sv2v_reg;
  assign data_r[1616] = data_r_1616_sv2v_reg;
  assign data_r[1615] = data_r_1615_sv2v_reg;
  assign data_r[1614] = data_r_1614_sv2v_reg;
  assign data_r[1613] = data_r_1613_sv2v_reg;
  assign data_r[1612] = data_r_1612_sv2v_reg;
  assign data_r[1611] = data_r_1611_sv2v_reg;
  assign data_r[1610] = data_r_1610_sv2v_reg;
  assign data_r[1609] = data_r_1609_sv2v_reg;
  assign data_r[1608] = data_r_1608_sv2v_reg;
  assign data_r[1607] = data_r_1607_sv2v_reg;
  assign data_r[1606] = data_r_1606_sv2v_reg;
  assign data_r[1605] = data_r_1605_sv2v_reg;
  assign data_r[1604] = data_r_1604_sv2v_reg;
  assign data_r[1603] = data_r_1603_sv2v_reg;
  assign data_r[1602] = data_r_1602_sv2v_reg;
  assign data_r[1601] = data_r_1601_sv2v_reg;
  assign data_r[1600] = data_r_1600_sv2v_reg;
  assign data_r[1599] = data_r_1599_sv2v_reg;
  assign data_r[1598] = data_r_1598_sv2v_reg;
  assign data_r[1597] = data_r_1597_sv2v_reg;
  assign data_r[1596] = data_r_1596_sv2v_reg;
  assign data_r[1595] = data_r_1595_sv2v_reg;
  assign data_r[1594] = data_r_1594_sv2v_reg;
  assign data_r[1593] = data_r_1593_sv2v_reg;
  assign data_r[1592] = data_r_1592_sv2v_reg;
  assign data_r[1591] = data_r_1591_sv2v_reg;
  assign data_r[1590] = data_r_1590_sv2v_reg;
  assign data_r[1589] = data_r_1589_sv2v_reg;
  assign data_r[1588] = data_r_1588_sv2v_reg;
  assign data_r[1587] = data_r_1587_sv2v_reg;
  assign data_r[1586] = data_r_1586_sv2v_reg;
  assign data_r[1585] = data_r_1585_sv2v_reg;
  assign data_r[1584] = data_r_1584_sv2v_reg;
  assign data_r[1583] = data_r_1583_sv2v_reg;
  assign data_r[1582] = data_r_1582_sv2v_reg;
  assign data_r[1581] = data_r_1581_sv2v_reg;
  assign data_r[1580] = data_r_1580_sv2v_reg;
  assign data_r[1579] = data_r_1579_sv2v_reg;
  assign data_r[1578] = data_r_1578_sv2v_reg;
  assign data_r[1577] = data_r_1577_sv2v_reg;
  assign data_r[1576] = data_r_1576_sv2v_reg;
  assign data_r[1575] = data_r_1575_sv2v_reg;
  assign data_r[1574] = data_r_1574_sv2v_reg;
  assign data_r[1573] = data_r_1573_sv2v_reg;
  assign data_r[1572] = data_r_1572_sv2v_reg;
  assign data_r[1571] = data_r_1571_sv2v_reg;
  assign data_r[1570] = data_r_1570_sv2v_reg;
  assign data_r[1569] = data_r_1569_sv2v_reg;
  assign data_r[1568] = data_r_1568_sv2v_reg;
  assign data_r[1567] = data_r_1567_sv2v_reg;
  assign data_r[1566] = data_r_1566_sv2v_reg;
  assign data_r[1565] = data_r_1565_sv2v_reg;
  assign data_r[1564] = data_r_1564_sv2v_reg;
  assign data_r[1563] = data_r_1563_sv2v_reg;
  assign data_r[1562] = data_r_1562_sv2v_reg;
  assign data_r[1561] = data_r_1561_sv2v_reg;
  assign data_r[1560] = data_r_1560_sv2v_reg;
  assign data_r[1559] = data_r_1559_sv2v_reg;
  assign data_r[1558] = data_r_1558_sv2v_reg;
  assign data_r[1557] = data_r_1557_sv2v_reg;
  assign data_r[1556] = data_r_1556_sv2v_reg;
  assign data_r[1555] = data_r_1555_sv2v_reg;
  assign data_r[1554] = data_r_1554_sv2v_reg;
  assign data_r[1553] = data_r_1553_sv2v_reg;
  assign data_r[1552] = data_r_1552_sv2v_reg;
  assign data_r[1551] = data_r_1551_sv2v_reg;
  assign data_r[1550] = data_r_1550_sv2v_reg;
  assign data_r[1549] = data_r_1549_sv2v_reg;
  assign data_r[1548] = data_r_1548_sv2v_reg;
  assign data_r[1547] = data_r_1547_sv2v_reg;
  assign data_r[1546] = data_r_1546_sv2v_reg;
  assign data_r[1545] = data_r_1545_sv2v_reg;
  assign data_r[1544] = data_r_1544_sv2v_reg;
  assign data_r[1543] = data_r_1543_sv2v_reg;
  assign data_r[1542] = data_r_1542_sv2v_reg;
  assign data_r[1541] = data_r_1541_sv2v_reg;
  assign data_r[1540] = data_r_1540_sv2v_reg;
  assign data_r[1539] = data_r_1539_sv2v_reg;
  assign data_r[1538] = data_r_1538_sv2v_reg;
  assign data_r[1537] = data_r_1537_sv2v_reg;
  assign data_r[1536] = data_r_1536_sv2v_reg;
  assign data_r[1535] = data_r_1535_sv2v_reg;
  assign data_r[1534] = data_r_1534_sv2v_reg;
  assign data_r[1533] = data_r_1533_sv2v_reg;
  assign data_r[1532] = data_r_1532_sv2v_reg;
  assign data_r[1531] = data_r_1531_sv2v_reg;
  assign data_r[1530] = data_r_1530_sv2v_reg;
  assign data_r[1529] = data_r_1529_sv2v_reg;
  assign data_r[1528] = data_r_1528_sv2v_reg;
  assign data_r[1527] = data_r_1527_sv2v_reg;
  assign data_r[1526] = data_r_1526_sv2v_reg;
  assign data_r[1525] = data_r_1525_sv2v_reg;
  assign data_r[1524] = data_r_1524_sv2v_reg;
  assign data_r[1523] = data_r_1523_sv2v_reg;
  assign data_r[1522] = data_r_1522_sv2v_reg;
  assign data_r[1521] = data_r_1521_sv2v_reg;
  assign data_r[1520] = data_r_1520_sv2v_reg;
  assign data_r[1519] = data_r_1519_sv2v_reg;
  assign data_r[1518] = data_r_1518_sv2v_reg;
  assign data_r[1517] = data_r_1517_sv2v_reg;
  assign data_r[1516] = data_r_1516_sv2v_reg;
  assign data_r[1515] = data_r_1515_sv2v_reg;
  assign data_r[1514] = data_r_1514_sv2v_reg;
  assign data_r[1513] = data_r_1513_sv2v_reg;
  assign data_r[1512] = data_r_1512_sv2v_reg;
  assign data_r[1511] = data_r_1511_sv2v_reg;
  assign data_r[1510] = data_r_1510_sv2v_reg;
  assign data_r[1509] = data_r_1509_sv2v_reg;
  assign data_r[1508] = data_r_1508_sv2v_reg;
  assign data_r[1507] = data_r_1507_sv2v_reg;
  assign data_r[1506] = data_r_1506_sv2v_reg;
  assign data_r[1505] = data_r_1505_sv2v_reg;
  assign data_r[1504] = data_r_1504_sv2v_reg;
  assign data_r[1503] = data_r_1503_sv2v_reg;
  assign data_r[1502] = data_r_1502_sv2v_reg;
  assign data_r[1501] = data_r_1501_sv2v_reg;
  assign data_r[1500] = data_r_1500_sv2v_reg;
  assign data_r[1499] = data_r_1499_sv2v_reg;
  assign data_r[1498] = data_r_1498_sv2v_reg;
  assign data_r[1497] = data_r_1497_sv2v_reg;
  assign data_r[1496] = data_r_1496_sv2v_reg;
  assign data_r[1495] = data_r_1495_sv2v_reg;
  assign data_r[1494] = data_r_1494_sv2v_reg;
  assign data_r[1493] = data_r_1493_sv2v_reg;
  assign data_r[1492] = data_r_1492_sv2v_reg;
  assign data_r[1491] = data_r_1491_sv2v_reg;
  assign data_r[1490] = data_r_1490_sv2v_reg;
  assign data_r[1489] = data_r_1489_sv2v_reg;
  assign data_r[1488] = data_r_1488_sv2v_reg;
  assign data_r[1487] = data_r_1487_sv2v_reg;
  assign data_r[1486] = data_r_1486_sv2v_reg;
  assign data_r[1485] = data_r_1485_sv2v_reg;
  assign data_r[1484] = data_r_1484_sv2v_reg;
  assign data_r[1483] = data_r_1483_sv2v_reg;
  assign data_r[1482] = data_r_1482_sv2v_reg;
  assign data_r[1481] = data_r_1481_sv2v_reg;
  assign data_r[1480] = data_r_1480_sv2v_reg;
  assign data_r[1479] = data_r_1479_sv2v_reg;
  assign data_r[1478] = data_r_1478_sv2v_reg;
  assign data_r[1477] = data_r_1477_sv2v_reg;
  assign data_r[1476] = data_r_1476_sv2v_reg;
  assign data_r[1475] = data_r_1475_sv2v_reg;
  assign data_r[1474] = data_r_1474_sv2v_reg;
  assign data_r[1473] = data_r_1473_sv2v_reg;
  assign data_r[1472] = data_r_1472_sv2v_reg;
  assign data_r[1471] = data_r_1471_sv2v_reg;
  assign data_r[1470] = data_r_1470_sv2v_reg;
  assign data_r[1469] = data_r_1469_sv2v_reg;
  assign data_r[1468] = data_r_1468_sv2v_reg;
  assign data_r[1467] = data_r_1467_sv2v_reg;
  assign data_r[1466] = data_r_1466_sv2v_reg;
  assign data_r[1465] = data_r_1465_sv2v_reg;
  assign data_r[1464] = data_r_1464_sv2v_reg;
  assign data_r[1463] = data_r_1463_sv2v_reg;
  assign data_r[1462] = data_r_1462_sv2v_reg;
  assign data_r[1461] = data_r_1461_sv2v_reg;
  assign data_r[1460] = data_r_1460_sv2v_reg;
  assign data_r[1459] = data_r_1459_sv2v_reg;
  assign data_r[1458] = data_r_1458_sv2v_reg;
  assign data_r[1457] = data_r_1457_sv2v_reg;
  assign data_r[1456] = data_r_1456_sv2v_reg;
  assign data_r[1455] = data_r_1455_sv2v_reg;
  assign data_r[1454] = data_r_1454_sv2v_reg;
  assign data_r[1453] = data_r_1453_sv2v_reg;
  assign data_r[1452] = data_r_1452_sv2v_reg;
  assign data_r[1451] = data_r_1451_sv2v_reg;
  assign data_r[1450] = data_r_1450_sv2v_reg;
  assign data_r[1449] = data_r_1449_sv2v_reg;
  assign data_r[1448] = data_r_1448_sv2v_reg;
  assign data_r[1447] = data_r_1447_sv2v_reg;
  assign data_r[1446] = data_r_1446_sv2v_reg;
  assign data_r[1445] = data_r_1445_sv2v_reg;
  assign data_r[1444] = data_r_1444_sv2v_reg;
  assign data_r[1443] = data_r_1443_sv2v_reg;
  assign data_r[1442] = data_r_1442_sv2v_reg;
  assign data_r[1441] = data_r_1441_sv2v_reg;
  assign data_r[1440] = data_r_1440_sv2v_reg;
  assign data_r[1439] = data_r_1439_sv2v_reg;
  assign data_r[1438] = data_r_1438_sv2v_reg;
  assign data_r[1437] = data_r_1437_sv2v_reg;
  assign data_r[1436] = data_r_1436_sv2v_reg;
  assign data_r[1435] = data_r_1435_sv2v_reg;
  assign data_r[1434] = data_r_1434_sv2v_reg;
  assign data_r[1433] = data_r_1433_sv2v_reg;
  assign data_r[1432] = data_r_1432_sv2v_reg;
  assign data_r[1431] = data_r_1431_sv2v_reg;
  assign data_r[1430] = data_r_1430_sv2v_reg;
  assign data_r[1429] = data_r_1429_sv2v_reg;
  assign data_r[1428] = data_r_1428_sv2v_reg;
  assign data_r[1427] = data_r_1427_sv2v_reg;
  assign data_r[1426] = data_r_1426_sv2v_reg;
  assign data_r[1425] = data_r_1425_sv2v_reg;
  assign data_r[1424] = data_r_1424_sv2v_reg;
  assign data_r[1423] = data_r_1423_sv2v_reg;
  assign data_r[1422] = data_r_1422_sv2v_reg;
  assign data_r[1421] = data_r_1421_sv2v_reg;
  assign data_r[1420] = data_r_1420_sv2v_reg;
  assign data_r[1419] = data_r_1419_sv2v_reg;
  assign data_r[1418] = data_r_1418_sv2v_reg;
  assign data_r[1417] = data_r_1417_sv2v_reg;
  assign data_r[1416] = data_r_1416_sv2v_reg;
  assign data_r[1415] = data_r_1415_sv2v_reg;
  assign data_r[1414] = data_r_1414_sv2v_reg;
  assign data_r[1413] = data_r_1413_sv2v_reg;
  assign data_r[1412] = data_r_1412_sv2v_reg;
  assign data_r[1411] = data_r_1411_sv2v_reg;
  assign data_r[1410] = data_r_1410_sv2v_reg;
  assign data_r[1409] = data_r_1409_sv2v_reg;
  assign data_r[1408] = data_r_1408_sv2v_reg;
  assign data_r[1407] = data_r_1407_sv2v_reg;
  assign data_r[1406] = data_r_1406_sv2v_reg;
  assign data_r[1405] = data_r_1405_sv2v_reg;
  assign data_r[1404] = data_r_1404_sv2v_reg;
  assign data_r[1403] = data_r_1403_sv2v_reg;
  assign data_r[1402] = data_r_1402_sv2v_reg;
  assign data_r[1401] = data_r_1401_sv2v_reg;
  assign data_r[1400] = data_r_1400_sv2v_reg;
  assign data_r[1399] = data_r_1399_sv2v_reg;
  assign data_r[1398] = data_r_1398_sv2v_reg;
  assign data_r[1397] = data_r_1397_sv2v_reg;
  assign data_r[1396] = data_r_1396_sv2v_reg;
  assign data_r[1395] = data_r_1395_sv2v_reg;
  assign data_r[1394] = data_r_1394_sv2v_reg;
  assign data_r[1393] = data_r_1393_sv2v_reg;
  assign data_r[1392] = data_r_1392_sv2v_reg;
  assign data_r[1391] = data_r_1391_sv2v_reg;
  assign data_r[1390] = data_r_1390_sv2v_reg;
  assign data_r[1389] = data_r_1389_sv2v_reg;
  assign data_r[1388] = data_r_1388_sv2v_reg;
  assign data_r[1387] = data_r_1387_sv2v_reg;
  assign data_r[1386] = data_r_1386_sv2v_reg;
  assign data_r[1385] = data_r_1385_sv2v_reg;
  assign data_r[1384] = data_r_1384_sv2v_reg;
  assign data_r[1383] = data_r_1383_sv2v_reg;
  assign data_r[1382] = data_r_1382_sv2v_reg;
  assign data_r[1381] = data_r_1381_sv2v_reg;
  assign data_r[1380] = data_r_1380_sv2v_reg;
  assign data_r[1379] = data_r_1379_sv2v_reg;
  assign data_r[1378] = data_r_1378_sv2v_reg;
  assign data_r[1377] = data_r_1377_sv2v_reg;
  assign data_r[1376] = data_r_1376_sv2v_reg;
  assign data_r[1375] = data_r_1375_sv2v_reg;
  assign data_r[1374] = data_r_1374_sv2v_reg;
  assign data_r[1373] = data_r_1373_sv2v_reg;
  assign data_r[1372] = data_r_1372_sv2v_reg;
  assign data_r[1371] = data_r_1371_sv2v_reg;
  assign data_r[1370] = data_r_1370_sv2v_reg;
  assign data_r[1369] = data_r_1369_sv2v_reg;
  assign data_r[1368] = data_r_1368_sv2v_reg;
  assign data_r[1367] = data_r_1367_sv2v_reg;
  assign data_r[1366] = data_r_1366_sv2v_reg;
  assign data_r[1365] = data_r_1365_sv2v_reg;
  assign data_r[1364] = data_r_1364_sv2v_reg;
  assign data_r[1363] = data_r_1363_sv2v_reg;
  assign data_r[1362] = data_r_1362_sv2v_reg;
  assign data_r[1361] = data_r_1361_sv2v_reg;
  assign data_r[1360] = data_r_1360_sv2v_reg;
  assign data_r[1359] = data_r_1359_sv2v_reg;
  assign data_r[1358] = data_r_1358_sv2v_reg;
  assign data_r[1357] = data_r_1357_sv2v_reg;
  assign data_r[1356] = data_r_1356_sv2v_reg;
  assign data_r[1355] = data_r_1355_sv2v_reg;
  assign data_r[1354] = data_r_1354_sv2v_reg;
  assign data_r[1353] = data_r_1353_sv2v_reg;
  assign data_r[1352] = data_r_1352_sv2v_reg;
  assign data_r[1351] = data_r_1351_sv2v_reg;
  assign data_r[1350] = data_r_1350_sv2v_reg;
  assign data_r[1349] = data_r_1349_sv2v_reg;
  assign data_r[1348] = data_r_1348_sv2v_reg;
  assign data_r[1347] = data_r_1347_sv2v_reg;
  assign data_r[1346] = data_r_1346_sv2v_reg;
  assign data_r[1345] = data_r_1345_sv2v_reg;
  assign data_r[1344] = data_r_1344_sv2v_reg;
  assign data_r[1343] = data_r_1343_sv2v_reg;
  assign data_r[1342] = data_r_1342_sv2v_reg;
  assign data_r[1341] = data_r_1341_sv2v_reg;
  assign data_r[1340] = data_r_1340_sv2v_reg;
  assign data_r[1339] = data_r_1339_sv2v_reg;
  assign data_r[1338] = data_r_1338_sv2v_reg;
  assign data_r[1337] = data_r_1337_sv2v_reg;
  assign data_r[1336] = data_r_1336_sv2v_reg;
  assign data_r[1335] = data_r_1335_sv2v_reg;
  assign data_r[1334] = data_r_1334_sv2v_reg;
  assign data_r[1333] = data_r_1333_sv2v_reg;
  assign data_r[1332] = data_r_1332_sv2v_reg;
  assign data_r[1331] = data_r_1331_sv2v_reg;
  assign data_r[1330] = data_r_1330_sv2v_reg;
  assign data_r[1329] = data_r_1329_sv2v_reg;
  assign data_r[1328] = data_r_1328_sv2v_reg;
  assign data_r[1327] = data_r_1327_sv2v_reg;
  assign data_r[1326] = data_r_1326_sv2v_reg;
  assign data_r[1325] = data_r_1325_sv2v_reg;
  assign data_r[1324] = data_r_1324_sv2v_reg;
  assign data_r[1323] = data_r_1323_sv2v_reg;
  assign data_r[1322] = data_r_1322_sv2v_reg;
  assign data_r[1321] = data_r_1321_sv2v_reg;
  assign data_r[1320] = data_r_1320_sv2v_reg;
  assign data_r[1319] = data_r_1319_sv2v_reg;
  assign data_r[1318] = data_r_1318_sv2v_reg;
  assign data_r[1317] = data_r_1317_sv2v_reg;
  assign data_r[1316] = data_r_1316_sv2v_reg;
  assign data_r[1315] = data_r_1315_sv2v_reg;
  assign data_r[1314] = data_r_1314_sv2v_reg;
  assign data_r[1313] = data_r_1313_sv2v_reg;
  assign data_r[1312] = data_r_1312_sv2v_reg;
  assign data_r[1311] = data_r_1311_sv2v_reg;
  assign data_r[1310] = data_r_1310_sv2v_reg;
  assign data_r[1309] = data_r_1309_sv2v_reg;
  assign data_r[1308] = data_r_1308_sv2v_reg;
  assign data_r[1307] = data_r_1307_sv2v_reg;
  assign data_r[1306] = data_r_1306_sv2v_reg;
  assign data_r[1305] = data_r_1305_sv2v_reg;
  assign data_r[1304] = data_r_1304_sv2v_reg;
  assign data_r[1303] = data_r_1303_sv2v_reg;
  assign data_r[1302] = data_r_1302_sv2v_reg;
  assign data_r[1301] = data_r_1301_sv2v_reg;
  assign data_r[1300] = data_r_1300_sv2v_reg;
  assign data_r[1299] = data_r_1299_sv2v_reg;
  assign data_r[1298] = data_r_1298_sv2v_reg;
  assign data_r[1297] = data_r_1297_sv2v_reg;
  assign data_r[1296] = data_r_1296_sv2v_reg;
  assign data_r[1295] = data_r_1295_sv2v_reg;
  assign data_r[1294] = data_r_1294_sv2v_reg;
  assign data_r[1293] = data_r_1293_sv2v_reg;
  assign data_r[1292] = data_r_1292_sv2v_reg;
  assign data_r[1291] = data_r_1291_sv2v_reg;
  assign data_r[1290] = data_r_1290_sv2v_reg;
  assign data_r[1289] = data_r_1289_sv2v_reg;
  assign data_r[1288] = data_r_1288_sv2v_reg;
  assign data_r[1287] = data_r_1287_sv2v_reg;
  assign data_r[1286] = data_r_1286_sv2v_reg;
  assign data_r[1285] = data_r_1285_sv2v_reg;
  assign data_r[1284] = data_r_1284_sv2v_reg;
  assign data_r[1283] = data_r_1283_sv2v_reg;
  assign data_r[1282] = data_r_1282_sv2v_reg;
  assign data_r[1281] = data_r_1281_sv2v_reg;
  assign data_r[1280] = data_r_1280_sv2v_reg;
  assign data_r[1279] = data_r_1279_sv2v_reg;
  assign data_r[1278] = data_r_1278_sv2v_reg;
  assign data_r[1277] = data_r_1277_sv2v_reg;
  assign data_r[1276] = data_r_1276_sv2v_reg;
  assign data_r[1275] = data_r_1275_sv2v_reg;
  assign data_r[1274] = data_r_1274_sv2v_reg;
  assign data_r[1273] = data_r_1273_sv2v_reg;
  assign data_r[1272] = data_r_1272_sv2v_reg;
  assign data_r[1271] = data_r_1271_sv2v_reg;
  assign data_r[1270] = data_r_1270_sv2v_reg;
  assign data_r[1269] = data_r_1269_sv2v_reg;
  assign data_r[1268] = data_r_1268_sv2v_reg;
  assign data_r[1267] = data_r_1267_sv2v_reg;
  assign data_r[1266] = data_r_1266_sv2v_reg;
  assign data_r[1265] = data_r_1265_sv2v_reg;
  assign data_r[1264] = data_r_1264_sv2v_reg;
  assign data_r[1263] = data_r_1263_sv2v_reg;
  assign data_r[1262] = data_r_1262_sv2v_reg;
  assign data_r[1261] = data_r_1261_sv2v_reg;
  assign data_r[1260] = data_r_1260_sv2v_reg;
  assign data_r[1259] = data_r_1259_sv2v_reg;
  assign data_r[1258] = data_r_1258_sv2v_reg;
  assign data_r[1257] = data_r_1257_sv2v_reg;
  assign data_r[1256] = data_r_1256_sv2v_reg;
  assign data_r[1255] = data_r_1255_sv2v_reg;
  assign data_r[1254] = data_r_1254_sv2v_reg;
  assign data_r[1253] = data_r_1253_sv2v_reg;
  assign data_r[1252] = data_r_1252_sv2v_reg;
  assign data_r[1251] = data_r_1251_sv2v_reg;
  assign data_r[1250] = data_r_1250_sv2v_reg;
  assign data_r[1249] = data_r_1249_sv2v_reg;
  assign data_r[1248] = data_r_1248_sv2v_reg;
  assign data_r[1247] = data_r_1247_sv2v_reg;
  assign data_r[1246] = data_r_1246_sv2v_reg;
  assign data_r[1245] = data_r_1245_sv2v_reg;
  assign data_r[1244] = data_r_1244_sv2v_reg;
  assign data_r[1243] = data_r_1243_sv2v_reg;
  assign data_r[1242] = data_r_1242_sv2v_reg;
  assign data_r[1241] = data_r_1241_sv2v_reg;
  assign data_r[1240] = data_r_1240_sv2v_reg;
  assign data_r[1239] = data_r_1239_sv2v_reg;
  assign data_r[1238] = data_r_1238_sv2v_reg;
  assign data_r[1237] = data_r_1237_sv2v_reg;
  assign data_r[1236] = data_r_1236_sv2v_reg;
  assign data_r[1235] = data_r_1235_sv2v_reg;
  assign data_r[1234] = data_r_1234_sv2v_reg;
  assign data_r[1233] = data_r_1233_sv2v_reg;
  assign data_r[1232] = data_r_1232_sv2v_reg;
  assign data_r[1231] = data_r_1231_sv2v_reg;
  assign data_r[1230] = data_r_1230_sv2v_reg;
  assign data_r[1229] = data_r_1229_sv2v_reg;
  assign data_r[1228] = data_r_1228_sv2v_reg;
  assign data_r[1227] = data_r_1227_sv2v_reg;
  assign data_r[1226] = data_r_1226_sv2v_reg;
  assign data_r[1225] = data_r_1225_sv2v_reg;
  assign data_r[1224] = data_r_1224_sv2v_reg;
  assign data_r[1223] = data_r_1223_sv2v_reg;
  assign data_r[1222] = data_r_1222_sv2v_reg;
  assign data_r[1221] = data_r_1221_sv2v_reg;
  assign data_r[1220] = data_r_1220_sv2v_reg;
  assign data_r[1219] = data_r_1219_sv2v_reg;
  assign data_r[1218] = data_r_1218_sv2v_reg;
  assign data_r[1217] = data_r_1217_sv2v_reg;
  assign data_r[1216] = data_r_1216_sv2v_reg;
  assign data_r[1215] = data_r_1215_sv2v_reg;
  assign data_r[1214] = data_r_1214_sv2v_reg;
  assign data_r[1213] = data_r_1213_sv2v_reg;
  assign data_r[1212] = data_r_1212_sv2v_reg;
  assign data_r[1211] = data_r_1211_sv2v_reg;
  assign data_r[1210] = data_r_1210_sv2v_reg;
  assign data_r[1209] = data_r_1209_sv2v_reg;
  assign data_r[1208] = data_r_1208_sv2v_reg;
  assign data_r[1207] = data_r_1207_sv2v_reg;
  assign data_r[1206] = data_r_1206_sv2v_reg;
  assign data_r[1205] = data_r_1205_sv2v_reg;
  assign data_r[1204] = data_r_1204_sv2v_reg;
  assign data_r[1203] = data_r_1203_sv2v_reg;
  assign data_r[1202] = data_r_1202_sv2v_reg;
  assign data_r[1201] = data_r_1201_sv2v_reg;
  assign data_r[1200] = data_r_1200_sv2v_reg;
  assign data_r[1199] = data_r_1199_sv2v_reg;
  assign data_r[1198] = data_r_1198_sv2v_reg;
  assign data_r[1197] = data_r_1197_sv2v_reg;
  assign data_r[1196] = data_r_1196_sv2v_reg;
  assign data_r[1195] = data_r_1195_sv2v_reg;
  assign data_r[1194] = data_r_1194_sv2v_reg;
  assign data_r[1193] = data_r_1193_sv2v_reg;
  assign data_r[1192] = data_r_1192_sv2v_reg;
  assign data_r[1191] = data_r_1191_sv2v_reg;
  assign data_r[1190] = data_r_1190_sv2v_reg;
  assign data_r[1189] = data_r_1189_sv2v_reg;
  assign data_r[1188] = data_r_1188_sv2v_reg;
  assign data_r[1187] = data_r_1187_sv2v_reg;
  assign data_r[1186] = data_r_1186_sv2v_reg;
  assign data_r[1185] = data_r_1185_sv2v_reg;
  assign data_r[1184] = data_r_1184_sv2v_reg;
  assign data_r[1183] = data_r_1183_sv2v_reg;
  assign data_r[1182] = data_r_1182_sv2v_reg;
  assign data_r[1181] = data_r_1181_sv2v_reg;
  assign data_r[1180] = data_r_1180_sv2v_reg;
  assign data_r[1179] = data_r_1179_sv2v_reg;
  assign data_r[1178] = data_r_1178_sv2v_reg;
  assign data_r[1177] = data_r_1177_sv2v_reg;
  assign data_r[1176] = data_r_1176_sv2v_reg;
  assign data_r[1175] = data_r_1175_sv2v_reg;
  assign data_r[1174] = data_r_1174_sv2v_reg;
  assign data_r[1173] = data_r_1173_sv2v_reg;
  assign data_r[1172] = data_r_1172_sv2v_reg;
  assign data_r[1171] = data_r_1171_sv2v_reg;
  assign data_r[1170] = data_r_1170_sv2v_reg;
  assign data_r[1169] = data_r_1169_sv2v_reg;
  assign data_r[1168] = data_r_1168_sv2v_reg;
  assign data_r[1167] = data_r_1167_sv2v_reg;
  assign data_r[1166] = data_r_1166_sv2v_reg;
  assign data_r[1165] = data_r_1165_sv2v_reg;
  assign data_r[1164] = data_r_1164_sv2v_reg;
  assign data_r[1163] = data_r_1163_sv2v_reg;
  assign data_r[1162] = data_r_1162_sv2v_reg;
  assign data_r[1161] = data_r_1161_sv2v_reg;
  assign data_r[1160] = data_r_1160_sv2v_reg;
  assign data_r[1159] = data_r_1159_sv2v_reg;
  assign data_r[1158] = data_r_1158_sv2v_reg;
  assign data_r[1157] = data_r_1157_sv2v_reg;
  assign data_r[1156] = data_r_1156_sv2v_reg;
  assign data_r[1155] = data_r_1155_sv2v_reg;
  assign data_r[1154] = data_r_1154_sv2v_reg;
  assign data_r[1153] = data_r_1153_sv2v_reg;
  assign data_r[1152] = data_r_1152_sv2v_reg;
  assign data_r[1151] = data_r_1151_sv2v_reg;
  assign data_r[1150] = data_r_1150_sv2v_reg;
  assign data_r[1149] = data_r_1149_sv2v_reg;
  assign data_r[1148] = data_r_1148_sv2v_reg;
  assign data_r[1147] = data_r_1147_sv2v_reg;
  assign data_r[1146] = data_r_1146_sv2v_reg;
  assign data_r[1145] = data_r_1145_sv2v_reg;
  assign data_r[1144] = data_r_1144_sv2v_reg;
  assign data_r[1143] = data_r_1143_sv2v_reg;
  assign data_r[1142] = data_r_1142_sv2v_reg;
  assign data_r[1141] = data_r_1141_sv2v_reg;
  assign data_r[1140] = data_r_1140_sv2v_reg;
  assign data_r[1139] = data_r_1139_sv2v_reg;
  assign data_r[1138] = data_r_1138_sv2v_reg;
  assign data_r[1137] = data_r_1137_sv2v_reg;
  assign data_r[1136] = data_r_1136_sv2v_reg;
  assign data_r[1135] = data_r_1135_sv2v_reg;
  assign data_r[1134] = data_r_1134_sv2v_reg;
  assign data_r[1133] = data_r_1133_sv2v_reg;
  assign data_r[1132] = data_r_1132_sv2v_reg;
  assign data_r[1131] = data_r_1131_sv2v_reg;
  assign data_r[1130] = data_r_1130_sv2v_reg;
  assign data_r[1129] = data_r_1129_sv2v_reg;
  assign data_r[1128] = data_r_1128_sv2v_reg;
  assign data_r[1127] = data_r_1127_sv2v_reg;
  assign data_r[1126] = data_r_1126_sv2v_reg;
  assign data_r[1125] = data_r_1125_sv2v_reg;
  assign data_r[1124] = data_r_1124_sv2v_reg;
  assign data_r[1123] = data_r_1123_sv2v_reg;
  assign data_r[1122] = data_r_1122_sv2v_reg;
  assign data_r[1121] = data_r_1121_sv2v_reg;
  assign data_r[1120] = data_r_1120_sv2v_reg;
  assign data_r[1119] = data_r_1119_sv2v_reg;
  assign data_r[1118] = data_r_1118_sv2v_reg;
  assign data_r[1117] = data_r_1117_sv2v_reg;
  assign data_r[1116] = data_r_1116_sv2v_reg;
  assign data_r[1115] = data_r_1115_sv2v_reg;
  assign data_r[1114] = data_r_1114_sv2v_reg;
  assign data_r[1113] = data_r_1113_sv2v_reg;
  assign data_r[1112] = data_r_1112_sv2v_reg;
  assign data_r[1111] = data_r_1111_sv2v_reg;
  assign data_r[1110] = data_r_1110_sv2v_reg;
  assign data_r[1109] = data_r_1109_sv2v_reg;
  assign data_r[1108] = data_r_1108_sv2v_reg;
  assign data_r[1107] = data_r_1107_sv2v_reg;
  assign data_r[1106] = data_r_1106_sv2v_reg;
  assign data_r[1105] = data_r_1105_sv2v_reg;
  assign data_r[1104] = data_r_1104_sv2v_reg;
  assign data_r[1103] = data_r_1103_sv2v_reg;
  assign data_r[1102] = data_r_1102_sv2v_reg;
  assign data_r[1101] = data_r_1101_sv2v_reg;
  assign data_r[1100] = data_r_1100_sv2v_reg;
  assign data_r[1099] = data_r_1099_sv2v_reg;
  assign data_r[1098] = data_r_1098_sv2v_reg;
  assign data_r[1097] = data_r_1097_sv2v_reg;
  assign data_r[1096] = data_r_1096_sv2v_reg;
  assign data_r[1095] = data_r_1095_sv2v_reg;
  assign data_r[1094] = data_r_1094_sv2v_reg;
  assign data_r[1093] = data_r_1093_sv2v_reg;
  assign data_r[1092] = data_r_1092_sv2v_reg;
  assign data_r[1091] = data_r_1091_sv2v_reg;
  assign data_r[1090] = data_r_1090_sv2v_reg;
  assign data_r[1089] = data_r_1089_sv2v_reg;
  assign data_r[1088] = data_r_1088_sv2v_reg;
  assign data_r[1087] = data_r_1087_sv2v_reg;
  assign data_r[1086] = data_r_1086_sv2v_reg;
  assign data_r[1085] = data_r_1085_sv2v_reg;
  assign data_r[1084] = data_r_1084_sv2v_reg;
  assign data_r[1083] = data_r_1083_sv2v_reg;
  assign data_r[1082] = data_r_1082_sv2v_reg;
  assign data_r[1081] = data_r_1081_sv2v_reg;
  assign data_r[1080] = data_r_1080_sv2v_reg;
  assign data_r[1079] = data_r_1079_sv2v_reg;
  assign data_r[1078] = data_r_1078_sv2v_reg;
  assign data_r[1077] = data_r_1077_sv2v_reg;
  assign data_r[1076] = data_r_1076_sv2v_reg;
  assign data_r[1075] = data_r_1075_sv2v_reg;
  assign data_r[1074] = data_r_1074_sv2v_reg;
  assign data_r[1073] = data_r_1073_sv2v_reg;
  assign data_r[1072] = data_r_1072_sv2v_reg;
  assign data_r[1071] = data_r_1071_sv2v_reg;
  assign data_r[1070] = data_r_1070_sv2v_reg;
  assign data_r[1069] = data_r_1069_sv2v_reg;
  assign data_r[1068] = data_r_1068_sv2v_reg;
  assign data_r[1067] = data_r_1067_sv2v_reg;
  assign data_r[1066] = data_r_1066_sv2v_reg;
  assign data_r[1065] = data_r_1065_sv2v_reg;
  assign data_r[1064] = data_r_1064_sv2v_reg;
  assign data_r[1063] = data_r_1063_sv2v_reg;
  assign data_r[1062] = data_r_1062_sv2v_reg;
  assign data_r[1061] = data_r_1061_sv2v_reg;
  assign data_r[1060] = data_r_1060_sv2v_reg;
  assign data_r[1059] = data_r_1059_sv2v_reg;
  assign data_r[1058] = data_r_1058_sv2v_reg;
  assign data_r[1057] = data_r_1057_sv2v_reg;
  assign data_r[1056] = data_r_1056_sv2v_reg;
  assign data_r[1055] = data_r_1055_sv2v_reg;
  assign data_r[1054] = data_r_1054_sv2v_reg;
  assign data_r[1053] = data_r_1053_sv2v_reg;
  assign data_r[1052] = data_r_1052_sv2v_reg;
  assign data_r[1051] = data_r_1051_sv2v_reg;
  assign data_r[1050] = data_r_1050_sv2v_reg;
  assign data_r[1049] = data_r_1049_sv2v_reg;
  assign data_r[1048] = data_r_1048_sv2v_reg;
  assign data_r[1047] = data_r_1047_sv2v_reg;
  assign data_r[1046] = data_r_1046_sv2v_reg;
  assign data_r[1045] = data_r_1045_sv2v_reg;
  assign data_r[1044] = data_r_1044_sv2v_reg;
  assign data_r[1043] = data_r_1043_sv2v_reg;
  assign data_r[1042] = data_r_1042_sv2v_reg;
  assign data_r[1041] = data_r_1041_sv2v_reg;
  assign data_r[1040] = data_r_1040_sv2v_reg;
  assign data_r[1039] = data_r_1039_sv2v_reg;
  assign data_r[1038] = data_r_1038_sv2v_reg;
  assign data_r[1037] = data_r_1037_sv2v_reg;
  assign data_r[1036] = data_r_1036_sv2v_reg;
  assign data_r[1035] = data_r_1035_sv2v_reg;
  assign data_r[1034] = data_r_1034_sv2v_reg;
  assign data_r[1033] = data_r_1033_sv2v_reg;
  assign data_r[1032] = data_r_1032_sv2v_reg;
  assign data_r[1031] = data_r_1031_sv2v_reg;
  assign data_r[1030] = data_r_1030_sv2v_reg;
  assign data_r[1029] = data_r_1029_sv2v_reg;
  assign data_r[1028] = data_r_1028_sv2v_reg;
  assign data_r[1027] = data_r_1027_sv2v_reg;
  assign data_r[1026] = data_r_1026_sv2v_reg;
  assign data_r[1025] = data_r_1025_sv2v_reg;
  assign data_r[1024] = data_r_1024_sv2v_reg;
  assign data_r[1023] = data_r_1023_sv2v_reg;
  assign data_r[1022] = data_r_1022_sv2v_reg;
  assign data_r[1021] = data_r_1021_sv2v_reg;
  assign data_r[1020] = data_r_1020_sv2v_reg;
  assign data_r[1019] = data_r_1019_sv2v_reg;
  assign data_r[1018] = data_r_1018_sv2v_reg;
  assign data_r[1017] = data_r_1017_sv2v_reg;
  assign data_r[1016] = data_r_1016_sv2v_reg;
  assign data_r[1015] = data_r_1015_sv2v_reg;
  assign data_r[1014] = data_r_1014_sv2v_reg;
  assign data_r[1013] = data_r_1013_sv2v_reg;
  assign data_r[1012] = data_r_1012_sv2v_reg;
  assign data_r[1011] = data_r_1011_sv2v_reg;
  assign data_r[1010] = data_r_1010_sv2v_reg;
  assign data_r[1009] = data_r_1009_sv2v_reg;
  assign data_r[1008] = data_r_1008_sv2v_reg;
  assign data_r[1007] = data_r_1007_sv2v_reg;
  assign data_r[1006] = data_r_1006_sv2v_reg;
  assign data_r[1005] = data_r_1005_sv2v_reg;
  assign data_r[1004] = data_r_1004_sv2v_reg;
  assign data_r[1003] = data_r_1003_sv2v_reg;
  assign data_r[1002] = data_r_1002_sv2v_reg;
  assign data_r[1001] = data_r_1001_sv2v_reg;
  assign data_r[1000] = data_r_1000_sv2v_reg;
  assign data_r[999] = data_r_999_sv2v_reg;
  assign data_r[998] = data_r_998_sv2v_reg;
  assign data_r[997] = data_r_997_sv2v_reg;
  assign data_r[996] = data_r_996_sv2v_reg;
  assign data_r[995] = data_r_995_sv2v_reg;
  assign data_r[994] = data_r_994_sv2v_reg;
  assign data_r[993] = data_r_993_sv2v_reg;
  assign data_r[992] = data_r_992_sv2v_reg;
  assign data_r[991] = data_r_991_sv2v_reg;
  assign data_r[990] = data_r_990_sv2v_reg;
  assign data_r[989] = data_r_989_sv2v_reg;
  assign data_r[988] = data_r_988_sv2v_reg;
  assign data_r[987] = data_r_987_sv2v_reg;
  assign data_r[986] = data_r_986_sv2v_reg;
  assign data_r[985] = data_r_985_sv2v_reg;
  assign data_r[984] = data_r_984_sv2v_reg;
  assign data_r[983] = data_r_983_sv2v_reg;
  assign data_r[982] = data_r_982_sv2v_reg;
  assign data_r[981] = data_r_981_sv2v_reg;
  assign data_r[980] = data_r_980_sv2v_reg;
  assign data_r[979] = data_r_979_sv2v_reg;
  assign data_r[978] = data_r_978_sv2v_reg;
  assign data_r[977] = data_r_977_sv2v_reg;
  assign data_r[976] = data_r_976_sv2v_reg;
  assign data_r[975] = data_r_975_sv2v_reg;
  assign data_r[974] = data_r_974_sv2v_reg;
  assign data_r[973] = data_r_973_sv2v_reg;
  assign data_r[972] = data_r_972_sv2v_reg;
  assign data_r[971] = data_r_971_sv2v_reg;
  assign data_r[970] = data_r_970_sv2v_reg;
  assign data_r[969] = data_r_969_sv2v_reg;
  assign data_r[968] = data_r_968_sv2v_reg;
  assign data_r[967] = data_r_967_sv2v_reg;
  assign data_r[966] = data_r_966_sv2v_reg;
  assign data_r[965] = data_r_965_sv2v_reg;
  assign data_r[964] = data_r_964_sv2v_reg;
  assign data_r[963] = data_r_963_sv2v_reg;
  assign data_r[962] = data_r_962_sv2v_reg;
  assign data_r[961] = data_r_961_sv2v_reg;
  assign data_r[960] = data_r_960_sv2v_reg;
  assign data_r[959] = data_r_959_sv2v_reg;
  assign data_r[958] = data_r_958_sv2v_reg;
  assign data_r[957] = data_r_957_sv2v_reg;
  assign data_r[956] = data_r_956_sv2v_reg;
  assign data_r[955] = data_r_955_sv2v_reg;
  assign data_r[954] = data_r_954_sv2v_reg;
  assign data_r[953] = data_r_953_sv2v_reg;
  assign data_r[952] = data_r_952_sv2v_reg;
  assign data_r[951] = data_r_951_sv2v_reg;
  assign data_r[950] = data_r_950_sv2v_reg;
  assign data_r[949] = data_r_949_sv2v_reg;
  assign data_r[948] = data_r_948_sv2v_reg;
  assign data_r[947] = data_r_947_sv2v_reg;
  assign data_r[946] = data_r_946_sv2v_reg;
  assign data_r[945] = data_r_945_sv2v_reg;
  assign data_r[944] = data_r_944_sv2v_reg;
  assign data_r[943] = data_r_943_sv2v_reg;
  assign data_r[942] = data_r_942_sv2v_reg;
  assign data_r[941] = data_r_941_sv2v_reg;
  assign data_r[940] = data_r_940_sv2v_reg;
  assign data_r[939] = data_r_939_sv2v_reg;
  assign data_r[938] = data_r_938_sv2v_reg;
  assign data_r[937] = data_r_937_sv2v_reg;
  assign data_r[936] = data_r_936_sv2v_reg;
  assign data_r[935] = data_r_935_sv2v_reg;
  assign data_r[934] = data_r_934_sv2v_reg;
  assign data_r[933] = data_r_933_sv2v_reg;
  assign data_r[932] = data_r_932_sv2v_reg;
  assign data_r[931] = data_r_931_sv2v_reg;
  assign data_r[930] = data_r_930_sv2v_reg;
  assign data_r[929] = data_r_929_sv2v_reg;
  assign data_r[928] = data_r_928_sv2v_reg;
  assign data_r[927] = data_r_927_sv2v_reg;
  assign data_r[926] = data_r_926_sv2v_reg;
  assign data_r[925] = data_r_925_sv2v_reg;
  assign data_r[924] = data_r_924_sv2v_reg;
  assign data_r[923] = data_r_923_sv2v_reg;
  assign data_r[922] = data_r_922_sv2v_reg;
  assign data_r[921] = data_r_921_sv2v_reg;
  assign data_r[920] = data_r_920_sv2v_reg;
  assign data_r[919] = data_r_919_sv2v_reg;
  assign data_r[918] = data_r_918_sv2v_reg;
  assign data_r[917] = data_r_917_sv2v_reg;
  assign data_r[916] = data_r_916_sv2v_reg;
  assign data_r[915] = data_r_915_sv2v_reg;
  assign data_r[914] = data_r_914_sv2v_reg;
  assign data_r[913] = data_r_913_sv2v_reg;
  assign data_r[912] = data_r_912_sv2v_reg;
  assign data_r[911] = data_r_911_sv2v_reg;
  assign data_r[910] = data_r_910_sv2v_reg;
  assign data_r[909] = data_r_909_sv2v_reg;
  assign data_r[908] = data_r_908_sv2v_reg;
  assign data_r[907] = data_r_907_sv2v_reg;
  assign data_r[906] = data_r_906_sv2v_reg;
  assign data_r[905] = data_r_905_sv2v_reg;
  assign data_r[904] = data_r_904_sv2v_reg;
  assign data_r[903] = data_r_903_sv2v_reg;
  assign data_r[902] = data_r_902_sv2v_reg;
  assign data_r[901] = data_r_901_sv2v_reg;
  assign data_r[900] = data_r_900_sv2v_reg;
  assign data_r[899] = data_r_899_sv2v_reg;
  assign data_r[898] = data_r_898_sv2v_reg;
  assign data_r[897] = data_r_897_sv2v_reg;
  assign data_r[896] = data_r_896_sv2v_reg;
  assign data_r[895] = data_r_895_sv2v_reg;
  assign data_r[894] = data_r_894_sv2v_reg;
  assign data_r[893] = data_r_893_sv2v_reg;
  assign data_r[892] = data_r_892_sv2v_reg;
  assign data_r[891] = data_r_891_sv2v_reg;
  assign data_r[890] = data_r_890_sv2v_reg;
  assign data_r[889] = data_r_889_sv2v_reg;
  assign data_r[888] = data_r_888_sv2v_reg;
  assign data_r[887] = data_r_887_sv2v_reg;
  assign data_r[886] = data_r_886_sv2v_reg;
  assign data_r[885] = data_r_885_sv2v_reg;
  assign data_r[884] = data_r_884_sv2v_reg;
  assign data_r[883] = data_r_883_sv2v_reg;
  assign data_r[882] = data_r_882_sv2v_reg;
  assign data_r[881] = data_r_881_sv2v_reg;
  assign data_r[880] = data_r_880_sv2v_reg;
  assign data_r[879] = data_r_879_sv2v_reg;
  assign data_r[878] = data_r_878_sv2v_reg;
  assign data_r[877] = data_r_877_sv2v_reg;
  assign data_r[876] = data_r_876_sv2v_reg;
  assign data_r[875] = data_r_875_sv2v_reg;
  assign data_r[874] = data_r_874_sv2v_reg;
  assign data_r[873] = data_r_873_sv2v_reg;
  assign data_r[872] = data_r_872_sv2v_reg;
  assign data_r[871] = data_r_871_sv2v_reg;
  assign data_r[870] = data_r_870_sv2v_reg;
  assign data_r[869] = data_r_869_sv2v_reg;
  assign data_r[868] = data_r_868_sv2v_reg;
  assign data_r[867] = data_r_867_sv2v_reg;
  assign data_r[866] = data_r_866_sv2v_reg;
  assign data_r[865] = data_r_865_sv2v_reg;
  assign data_r[864] = data_r_864_sv2v_reg;
  assign data_r[863] = data_r_863_sv2v_reg;
  assign data_r[862] = data_r_862_sv2v_reg;
  assign data_r[861] = data_r_861_sv2v_reg;
  assign data_r[860] = data_r_860_sv2v_reg;
  assign data_r[859] = data_r_859_sv2v_reg;
  assign data_r[858] = data_r_858_sv2v_reg;
  assign data_r[857] = data_r_857_sv2v_reg;
  assign data_r[856] = data_r_856_sv2v_reg;
  assign data_r[855] = data_r_855_sv2v_reg;
  assign data_r[854] = data_r_854_sv2v_reg;
  assign data_r[853] = data_r_853_sv2v_reg;
  assign data_r[852] = data_r_852_sv2v_reg;
  assign data_r[851] = data_r_851_sv2v_reg;
  assign data_r[850] = data_r_850_sv2v_reg;
  assign data_r[849] = data_r_849_sv2v_reg;
  assign data_r[848] = data_r_848_sv2v_reg;
  assign data_r[847] = data_r_847_sv2v_reg;
  assign data_r[846] = data_r_846_sv2v_reg;
  assign data_r[845] = data_r_845_sv2v_reg;
  assign data_r[844] = data_r_844_sv2v_reg;
  assign data_r[843] = data_r_843_sv2v_reg;
  assign data_r[842] = data_r_842_sv2v_reg;
  assign data_r[841] = data_r_841_sv2v_reg;
  assign data_r[840] = data_r_840_sv2v_reg;
  assign data_r[839] = data_r_839_sv2v_reg;
  assign data_r[838] = data_r_838_sv2v_reg;
  assign data_r[837] = data_r_837_sv2v_reg;
  assign data_r[836] = data_r_836_sv2v_reg;
  assign data_r[835] = data_r_835_sv2v_reg;
  assign data_r[834] = data_r_834_sv2v_reg;
  assign data_r[833] = data_r_833_sv2v_reg;
  assign data_r[832] = data_r_832_sv2v_reg;
  assign data_r[831] = data_r_831_sv2v_reg;
  assign data_r[830] = data_r_830_sv2v_reg;
  assign data_r[829] = data_r_829_sv2v_reg;
  assign data_r[828] = data_r_828_sv2v_reg;
  assign data_r[827] = data_r_827_sv2v_reg;
  assign data_r[826] = data_r_826_sv2v_reg;
  assign data_r[825] = data_r_825_sv2v_reg;
  assign data_r[824] = data_r_824_sv2v_reg;
  assign data_r[823] = data_r_823_sv2v_reg;
  assign data_r[822] = data_r_822_sv2v_reg;
  assign data_r[821] = data_r_821_sv2v_reg;
  assign data_r[820] = data_r_820_sv2v_reg;
  assign data_r[819] = data_r_819_sv2v_reg;
  assign data_r[818] = data_r_818_sv2v_reg;
  assign data_r[817] = data_r_817_sv2v_reg;
  assign data_r[816] = data_r_816_sv2v_reg;
  assign data_r[815] = data_r_815_sv2v_reg;
  assign data_r[814] = data_r_814_sv2v_reg;
  assign data_r[813] = data_r_813_sv2v_reg;
  assign data_r[812] = data_r_812_sv2v_reg;
  assign data_r[811] = data_r_811_sv2v_reg;
  assign data_r[810] = data_r_810_sv2v_reg;
  assign data_r[809] = data_r_809_sv2v_reg;
  assign data_r[808] = data_r_808_sv2v_reg;
  assign data_r[807] = data_r_807_sv2v_reg;
  assign data_r[806] = data_r_806_sv2v_reg;
  assign data_r[805] = data_r_805_sv2v_reg;
  assign data_r[804] = data_r_804_sv2v_reg;
  assign data_r[803] = data_r_803_sv2v_reg;
  assign data_r[802] = data_r_802_sv2v_reg;
  assign data_r[801] = data_r_801_sv2v_reg;
  assign data_r[800] = data_r_800_sv2v_reg;
  assign data_r[799] = data_r_799_sv2v_reg;
  assign data_r[798] = data_r_798_sv2v_reg;
  assign data_r[797] = data_r_797_sv2v_reg;
  assign data_r[796] = data_r_796_sv2v_reg;
  assign data_r[795] = data_r_795_sv2v_reg;
  assign data_r[794] = data_r_794_sv2v_reg;
  assign data_r[793] = data_r_793_sv2v_reg;
  assign data_r[792] = data_r_792_sv2v_reg;
  assign data_r[791] = data_r_791_sv2v_reg;
  assign data_r[790] = data_r_790_sv2v_reg;
  assign data_r[789] = data_r_789_sv2v_reg;
  assign data_r[788] = data_r_788_sv2v_reg;
  assign data_r[787] = data_r_787_sv2v_reg;
  assign data_r[786] = data_r_786_sv2v_reg;
  assign data_r[785] = data_r_785_sv2v_reg;
  assign data_r[784] = data_r_784_sv2v_reg;
  assign data_r[783] = data_r_783_sv2v_reg;
  assign data_r[782] = data_r_782_sv2v_reg;
  assign data_r[781] = data_r_781_sv2v_reg;
  assign data_r[780] = data_r_780_sv2v_reg;
  assign data_r[779] = data_r_779_sv2v_reg;
  assign data_r[778] = data_r_778_sv2v_reg;
  assign data_r[777] = data_r_777_sv2v_reg;
  assign data_r[776] = data_r_776_sv2v_reg;
  assign data_r[775] = data_r_775_sv2v_reg;
  assign data_r[774] = data_r_774_sv2v_reg;
  assign data_r[773] = data_r_773_sv2v_reg;
  assign data_r[772] = data_r_772_sv2v_reg;
  assign data_r[771] = data_r_771_sv2v_reg;
  assign data_r[770] = data_r_770_sv2v_reg;
  assign data_r[769] = data_r_769_sv2v_reg;
  assign data_r[768] = data_r_768_sv2v_reg;
  assign data_r[767] = data_r_767_sv2v_reg;
  assign data_r[766] = data_r_766_sv2v_reg;
  assign data_r[765] = data_r_765_sv2v_reg;
  assign data_r[764] = data_r_764_sv2v_reg;
  assign data_r[763] = data_r_763_sv2v_reg;
  assign data_r[762] = data_r_762_sv2v_reg;
  assign data_r[761] = data_r_761_sv2v_reg;
  assign data_r[760] = data_r_760_sv2v_reg;
  assign data_r[759] = data_r_759_sv2v_reg;
  assign data_r[758] = data_r_758_sv2v_reg;
  assign data_r[757] = data_r_757_sv2v_reg;
  assign data_r[756] = data_r_756_sv2v_reg;
  assign data_r[755] = data_r_755_sv2v_reg;
  assign data_r[754] = data_r_754_sv2v_reg;
  assign data_r[753] = data_r_753_sv2v_reg;
  assign data_r[752] = data_r_752_sv2v_reg;
  assign data_r[751] = data_r_751_sv2v_reg;
  assign data_r[750] = data_r_750_sv2v_reg;
  assign data_r[749] = data_r_749_sv2v_reg;
  assign data_r[748] = data_r_748_sv2v_reg;
  assign data_r[747] = data_r_747_sv2v_reg;
  assign data_r[746] = data_r_746_sv2v_reg;
  assign data_r[745] = data_r_745_sv2v_reg;
  assign data_r[744] = data_r_744_sv2v_reg;
  assign data_r[743] = data_r_743_sv2v_reg;
  assign data_r[742] = data_r_742_sv2v_reg;
  assign data_r[741] = data_r_741_sv2v_reg;
  assign data_r[740] = data_r_740_sv2v_reg;
  assign data_r[739] = data_r_739_sv2v_reg;
  assign data_r[738] = data_r_738_sv2v_reg;
  assign data_r[737] = data_r_737_sv2v_reg;
  assign data_r[736] = data_r_736_sv2v_reg;
  assign data_r[735] = data_r_735_sv2v_reg;
  assign data_r[734] = data_r_734_sv2v_reg;
  assign data_r[733] = data_r_733_sv2v_reg;
  assign data_r[732] = data_r_732_sv2v_reg;
  assign data_r[731] = data_r_731_sv2v_reg;
  assign data_r[730] = data_r_730_sv2v_reg;
  assign data_r[729] = data_r_729_sv2v_reg;
  assign data_r[728] = data_r_728_sv2v_reg;
  assign data_r[727] = data_r_727_sv2v_reg;
  assign data_r[726] = data_r_726_sv2v_reg;
  assign data_r[725] = data_r_725_sv2v_reg;
  assign data_r[724] = data_r_724_sv2v_reg;
  assign data_r[723] = data_r_723_sv2v_reg;
  assign data_r[722] = data_r_722_sv2v_reg;
  assign data_r[721] = data_r_721_sv2v_reg;
  assign data_r[720] = data_r_720_sv2v_reg;
  assign data_r[719] = data_r_719_sv2v_reg;
  assign data_r[718] = data_r_718_sv2v_reg;
  assign data_r[717] = data_r_717_sv2v_reg;
  assign data_r[716] = data_r_716_sv2v_reg;
  assign data_r[715] = data_r_715_sv2v_reg;
  assign data_r[714] = data_r_714_sv2v_reg;
  assign data_r[713] = data_r_713_sv2v_reg;
  assign data_r[712] = data_r_712_sv2v_reg;
  assign data_r[711] = data_r_711_sv2v_reg;
  assign data_r[710] = data_r_710_sv2v_reg;
  assign data_r[709] = data_r_709_sv2v_reg;
  assign data_r[708] = data_r_708_sv2v_reg;
  assign data_r[707] = data_r_707_sv2v_reg;
  assign data_r[706] = data_r_706_sv2v_reg;
  assign data_r[705] = data_r_705_sv2v_reg;
  assign data_r[704] = data_r_704_sv2v_reg;
  assign data_r[703] = data_r_703_sv2v_reg;
  assign data_r[702] = data_r_702_sv2v_reg;
  assign data_r[701] = data_r_701_sv2v_reg;
  assign data_r[700] = data_r_700_sv2v_reg;
  assign data_r[699] = data_r_699_sv2v_reg;
  assign data_r[698] = data_r_698_sv2v_reg;
  assign data_r[697] = data_r_697_sv2v_reg;
  assign data_r[696] = data_r_696_sv2v_reg;
  assign data_r[695] = data_r_695_sv2v_reg;
  assign data_r[694] = data_r_694_sv2v_reg;
  assign data_r[693] = data_r_693_sv2v_reg;
  assign data_r[692] = data_r_692_sv2v_reg;
  assign data_r[691] = data_r_691_sv2v_reg;
  assign data_r[690] = data_r_690_sv2v_reg;
  assign data_r[689] = data_r_689_sv2v_reg;
  assign data_r[688] = data_r_688_sv2v_reg;
  assign data_r[687] = data_r_687_sv2v_reg;
  assign data_r[686] = data_r_686_sv2v_reg;
  assign data_r[685] = data_r_685_sv2v_reg;
  assign data_r[684] = data_r_684_sv2v_reg;
  assign data_r[683] = data_r_683_sv2v_reg;
  assign data_r[682] = data_r_682_sv2v_reg;
  assign data_r[681] = data_r_681_sv2v_reg;
  assign data_r[680] = data_r_680_sv2v_reg;
  assign data_r[679] = data_r_679_sv2v_reg;
  assign data_r[678] = data_r_678_sv2v_reg;
  assign data_r[677] = data_r_677_sv2v_reg;
  assign data_r[676] = data_r_676_sv2v_reg;
  assign data_r[675] = data_r_675_sv2v_reg;
  assign data_r[674] = data_r_674_sv2v_reg;
  assign data_r[673] = data_r_673_sv2v_reg;
  assign data_r[672] = data_r_672_sv2v_reg;
  assign data_r[671] = data_r_671_sv2v_reg;
  assign data_r[670] = data_r_670_sv2v_reg;
  assign data_r[669] = data_r_669_sv2v_reg;
  assign data_r[668] = data_r_668_sv2v_reg;
  assign data_r[667] = data_r_667_sv2v_reg;
  assign data_r[666] = data_r_666_sv2v_reg;
  assign data_r[665] = data_r_665_sv2v_reg;
  assign data_r[664] = data_r_664_sv2v_reg;
  assign data_r[663] = data_r_663_sv2v_reg;
  assign data_r[662] = data_r_662_sv2v_reg;
  assign data_r[661] = data_r_661_sv2v_reg;
  assign data_r[660] = data_r_660_sv2v_reg;
  assign data_r[659] = data_r_659_sv2v_reg;
  assign data_r[658] = data_r_658_sv2v_reg;
  assign data_r[657] = data_r_657_sv2v_reg;
  assign data_r[656] = data_r_656_sv2v_reg;
  assign data_r[655] = data_r_655_sv2v_reg;
  assign data_r[654] = data_r_654_sv2v_reg;
  assign data_r[653] = data_r_653_sv2v_reg;
  assign data_r[652] = data_r_652_sv2v_reg;
  assign data_r[651] = data_r_651_sv2v_reg;
  assign data_r[650] = data_r_650_sv2v_reg;
  assign data_r[649] = data_r_649_sv2v_reg;
  assign data_r[648] = data_r_648_sv2v_reg;
  assign data_r[647] = data_r_647_sv2v_reg;
  assign data_r[646] = data_r_646_sv2v_reg;
  assign data_r[645] = data_r_645_sv2v_reg;
  assign data_r[644] = data_r_644_sv2v_reg;
  assign data_r[643] = data_r_643_sv2v_reg;
  assign data_r[642] = data_r_642_sv2v_reg;
  assign data_r[641] = data_r_641_sv2v_reg;
  assign data_r[640] = data_r_640_sv2v_reg;
  assign data_r[639] = data_r_639_sv2v_reg;
  assign data_r[638] = data_r_638_sv2v_reg;
  assign data_r[637] = data_r_637_sv2v_reg;
  assign data_r[636] = data_r_636_sv2v_reg;
  assign data_r[635] = data_r_635_sv2v_reg;
  assign data_r[634] = data_r_634_sv2v_reg;
  assign data_r[633] = data_r_633_sv2v_reg;
  assign data_r[632] = data_r_632_sv2v_reg;
  assign data_r[631] = data_r_631_sv2v_reg;
  assign data_r[630] = data_r_630_sv2v_reg;
  assign data_r[629] = data_r_629_sv2v_reg;
  assign data_r[628] = data_r_628_sv2v_reg;
  assign data_r[627] = data_r_627_sv2v_reg;
  assign data_r[626] = data_r_626_sv2v_reg;
  assign data_r[625] = data_r_625_sv2v_reg;
  assign data_r[624] = data_r_624_sv2v_reg;
  assign data_r[623] = data_r_623_sv2v_reg;
  assign data_r[622] = data_r_622_sv2v_reg;
  assign data_r[621] = data_r_621_sv2v_reg;
  assign data_r[620] = data_r_620_sv2v_reg;
  assign data_r[619] = data_r_619_sv2v_reg;
  assign data_r[618] = data_r_618_sv2v_reg;
  assign data_r[617] = data_r_617_sv2v_reg;
  assign data_r[616] = data_r_616_sv2v_reg;
  assign data_r[615] = data_r_615_sv2v_reg;
  assign data_r[614] = data_r_614_sv2v_reg;
  assign data_r[613] = data_r_613_sv2v_reg;
  assign data_r[612] = data_r_612_sv2v_reg;
  assign data_r[611] = data_r_611_sv2v_reg;
  assign data_r[610] = data_r_610_sv2v_reg;
  assign data_r[609] = data_r_609_sv2v_reg;
  assign data_r[608] = data_r_608_sv2v_reg;
  assign data_r[607] = data_r_607_sv2v_reg;
  assign data_r[606] = data_r_606_sv2v_reg;
  assign data_r[605] = data_r_605_sv2v_reg;
  assign data_r[604] = data_r_604_sv2v_reg;
  assign data_r[603] = data_r_603_sv2v_reg;
  assign data_r[602] = data_r_602_sv2v_reg;
  assign data_r[601] = data_r_601_sv2v_reg;
  assign data_r[600] = data_r_600_sv2v_reg;
  assign data_r[599] = data_r_599_sv2v_reg;
  assign data_r[598] = data_r_598_sv2v_reg;
  assign data_r[597] = data_r_597_sv2v_reg;
  assign data_r[596] = data_r_596_sv2v_reg;
  assign data_r[595] = data_r_595_sv2v_reg;
  assign data_r[594] = data_r_594_sv2v_reg;
  assign data_r[593] = data_r_593_sv2v_reg;
  assign data_r[592] = data_r_592_sv2v_reg;
  assign data_r[591] = data_r_591_sv2v_reg;
  assign data_r[590] = data_r_590_sv2v_reg;
  assign data_r[589] = data_r_589_sv2v_reg;
  assign data_r[588] = data_r_588_sv2v_reg;
  assign data_r[587] = data_r_587_sv2v_reg;
  assign data_r[586] = data_r_586_sv2v_reg;
  assign data_r[585] = data_r_585_sv2v_reg;
  assign data_r[584] = data_r_584_sv2v_reg;
  assign data_r[583] = data_r_583_sv2v_reg;
  assign data_r[582] = data_r_582_sv2v_reg;
  assign data_r[581] = data_r_581_sv2v_reg;
  assign data_r[580] = data_r_580_sv2v_reg;
  assign data_r[579] = data_r_579_sv2v_reg;
  assign data_r[578] = data_r_578_sv2v_reg;
  assign data_r[577] = data_r_577_sv2v_reg;
  assign data_r[576] = data_r_576_sv2v_reg;
  assign data_r[575] = data_r_575_sv2v_reg;
  assign data_r[574] = data_r_574_sv2v_reg;
  assign data_r[573] = data_r_573_sv2v_reg;
  assign data_r[572] = data_r_572_sv2v_reg;
  assign data_r[571] = data_r_571_sv2v_reg;
  assign data_r[570] = data_r_570_sv2v_reg;
  assign data_r[569] = data_r_569_sv2v_reg;
  assign data_r[568] = data_r_568_sv2v_reg;
  assign data_r[567] = data_r_567_sv2v_reg;
  assign data_r[566] = data_r_566_sv2v_reg;
  assign data_r[565] = data_r_565_sv2v_reg;
  assign data_r[564] = data_r_564_sv2v_reg;
  assign data_r[563] = data_r_563_sv2v_reg;
  assign data_r[562] = data_r_562_sv2v_reg;
  assign data_r[561] = data_r_561_sv2v_reg;
  assign data_r[560] = data_r_560_sv2v_reg;
  assign data_r[559] = data_r_559_sv2v_reg;
  assign data_r[558] = data_r_558_sv2v_reg;
  assign data_r[557] = data_r_557_sv2v_reg;
  assign data_r[556] = data_r_556_sv2v_reg;
  assign data_r[555] = data_r_555_sv2v_reg;
  assign data_r[554] = data_r_554_sv2v_reg;
  assign data_r[553] = data_r_553_sv2v_reg;
  assign data_r[552] = data_r_552_sv2v_reg;
  assign data_r[551] = data_r_551_sv2v_reg;
  assign data_r[550] = data_r_550_sv2v_reg;
  assign data_r[549] = data_r_549_sv2v_reg;
  assign data_r[548] = data_r_548_sv2v_reg;
  assign data_r[547] = data_r_547_sv2v_reg;
  assign data_r[546] = data_r_546_sv2v_reg;
  assign data_r[545] = data_r_545_sv2v_reg;
  assign data_r[544] = data_r_544_sv2v_reg;
  assign data_r[543] = data_r_543_sv2v_reg;
  assign data_r[542] = data_r_542_sv2v_reg;
  assign data_r[541] = data_r_541_sv2v_reg;
  assign data_r[540] = data_r_540_sv2v_reg;
  assign data_r[539] = data_r_539_sv2v_reg;
  assign data_r[538] = data_r_538_sv2v_reg;
  assign data_r[537] = data_r_537_sv2v_reg;
  assign data_r[536] = data_r_536_sv2v_reg;
  assign data_r[535] = data_r_535_sv2v_reg;
  assign data_r[534] = data_r_534_sv2v_reg;
  assign data_r[533] = data_r_533_sv2v_reg;
  assign data_r[532] = data_r_532_sv2v_reg;
  assign data_r[531] = data_r_531_sv2v_reg;
  assign data_r[530] = data_r_530_sv2v_reg;
  assign data_r[529] = data_r_529_sv2v_reg;
  assign data_r[528] = data_r_528_sv2v_reg;
  assign data_r[527] = data_r_527_sv2v_reg;
  assign data_r[526] = data_r_526_sv2v_reg;
  assign data_r[525] = data_r_525_sv2v_reg;
  assign data_r[524] = data_r_524_sv2v_reg;
  assign data_r[523] = data_r_523_sv2v_reg;
  assign data_r[522] = data_r_522_sv2v_reg;
  assign data_r[521] = data_r_521_sv2v_reg;
  assign data_r[520] = data_r_520_sv2v_reg;
  assign data_r[519] = data_r_519_sv2v_reg;
  assign data_r[518] = data_r_518_sv2v_reg;
  assign data_r[517] = data_r_517_sv2v_reg;
  assign data_r[516] = data_r_516_sv2v_reg;
  assign data_r[515] = data_r_515_sv2v_reg;
  assign data_r[514] = data_r_514_sv2v_reg;
  assign data_r[513] = data_r_513_sv2v_reg;
  assign data_r[512] = data_r_512_sv2v_reg;
  assign data_r[511] = data_r_511_sv2v_reg;
  assign data_r[510] = data_r_510_sv2v_reg;
  assign data_r[509] = data_r_509_sv2v_reg;
  assign data_r[508] = data_r_508_sv2v_reg;
  assign data_r[507] = data_r_507_sv2v_reg;
  assign data_r[506] = data_r_506_sv2v_reg;
  assign data_r[505] = data_r_505_sv2v_reg;
  assign data_r[504] = data_r_504_sv2v_reg;
  assign data_r[503] = data_r_503_sv2v_reg;
  assign data_r[502] = data_r_502_sv2v_reg;
  assign data_r[501] = data_r_501_sv2v_reg;
  assign data_r[500] = data_r_500_sv2v_reg;
  assign data_r[499] = data_r_499_sv2v_reg;
  assign data_r[498] = data_r_498_sv2v_reg;
  assign data_r[497] = data_r_497_sv2v_reg;
  assign data_r[496] = data_r_496_sv2v_reg;
  assign data_r[495] = data_r_495_sv2v_reg;
  assign data_r[494] = data_r_494_sv2v_reg;
  assign data_r[493] = data_r_493_sv2v_reg;
  assign data_r[492] = data_r_492_sv2v_reg;
  assign data_r[491] = data_r_491_sv2v_reg;
  assign data_r[490] = data_r_490_sv2v_reg;
  assign data_r[489] = data_r_489_sv2v_reg;
  assign data_r[488] = data_r_488_sv2v_reg;
  assign data_r[487] = data_r_487_sv2v_reg;
  assign data_r[486] = data_r_486_sv2v_reg;
  assign data_r[485] = data_r_485_sv2v_reg;
  assign data_r[484] = data_r_484_sv2v_reg;
  assign data_r[483] = data_r_483_sv2v_reg;
  assign data_r[482] = data_r_482_sv2v_reg;
  assign data_r[481] = data_r_481_sv2v_reg;
  assign data_r[480] = data_r_480_sv2v_reg;
  assign data_r[479] = data_r_479_sv2v_reg;
  assign data_r[478] = data_r_478_sv2v_reg;
  assign data_r[477] = data_r_477_sv2v_reg;
  assign data_r[476] = data_r_476_sv2v_reg;
  assign data_r[475] = data_r_475_sv2v_reg;
  assign data_r[474] = data_r_474_sv2v_reg;
  assign data_r[473] = data_r_473_sv2v_reg;
  assign data_r[472] = data_r_472_sv2v_reg;
  assign data_r[471] = data_r_471_sv2v_reg;
  assign data_r[470] = data_r_470_sv2v_reg;
  assign data_r[469] = data_r_469_sv2v_reg;
  assign data_r[468] = data_r_468_sv2v_reg;
  assign data_r[467] = data_r_467_sv2v_reg;
  assign data_r[466] = data_r_466_sv2v_reg;
  assign data_r[465] = data_r_465_sv2v_reg;
  assign data_r[464] = data_r_464_sv2v_reg;
  assign data_r[463] = data_r_463_sv2v_reg;
  assign data_r[462] = data_r_462_sv2v_reg;
  assign data_r[461] = data_r_461_sv2v_reg;
  assign data_r[460] = data_r_460_sv2v_reg;
  assign data_r[459] = data_r_459_sv2v_reg;
  assign data_r[458] = data_r_458_sv2v_reg;
  assign data_r[457] = data_r_457_sv2v_reg;
  assign data_r[456] = data_r_456_sv2v_reg;
  assign data_r[455] = data_r_455_sv2v_reg;
  assign data_r[454] = data_r_454_sv2v_reg;
  assign data_r[453] = data_r_453_sv2v_reg;
  assign data_r[452] = data_r_452_sv2v_reg;
  assign data_r[451] = data_r_451_sv2v_reg;
  assign data_r[450] = data_r_450_sv2v_reg;
  assign data_r[449] = data_r_449_sv2v_reg;
  assign data_r[448] = data_r_448_sv2v_reg;
  assign data_r[447] = data_r_447_sv2v_reg;
  assign data_r[446] = data_r_446_sv2v_reg;
  assign data_r[445] = data_r_445_sv2v_reg;
  assign data_r[444] = data_r_444_sv2v_reg;
  assign data_r[443] = data_r_443_sv2v_reg;
  assign data_r[442] = data_r_442_sv2v_reg;
  assign data_r[441] = data_r_441_sv2v_reg;
  assign data_r[440] = data_r_440_sv2v_reg;
  assign data_r[439] = data_r_439_sv2v_reg;
  assign data_r[438] = data_r_438_sv2v_reg;
  assign data_r[437] = data_r_437_sv2v_reg;
  assign data_r[436] = data_r_436_sv2v_reg;
  assign data_r[435] = data_r_435_sv2v_reg;
  assign data_r[434] = data_r_434_sv2v_reg;
  assign data_r[433] = data_r_433_sv2v_reg;
  assign data_r[432] = data_r_432_sv2v_reg;
  assign data_r[431] = data_r_431_sv2v_reg;
  assign data_r[430] = data_r_430_sv2v_reg;
  assign data_r[429] = data_r_429_sv2v_reg;
  assign data_r[428] = data_r_428_sv2v_reg;
  assign data_r[427] = data_r_427_sv2v_reg;
  assign data_r[426] = data_r_426_sv2v_reg;
  assign data_r[425] = data_r_425_sv2v_reg;
  assign data_r[424] = data_r_424_sv2v_reg;
  assign data_r[423] = data_r_423_sv2v_reg;
  assign data_r[422] = data_r_422_sv2v_reg;
  assign data_r[421] = data_r_421_sv2v_reg;
  assign data_r[420] = data_r_420_sv2v_reg;
  assign data_r[419] = data_r_419_sv2v_reg;
  assign data_r[418] = data_r_418_sv2v_reg;
  assign data_r[417] = data_r_417_sv2v_reg;
  assign data_r[416] = data_r_416_sv2v_reg;
  assign data_r[415] = data_r_415_sv2v_reg;
  assign data_r[414] = data_r_414_sv2v_reg;
  assign data_r[413] = data_r_413_sv2v_reg;
  assign data_r[412] = data_r_412_sv2v_reg;
  assign data_r[411] = data_r_411_sv2v_reg;
  assign data_r[410] = data_r_410_sv2v_reg;
  assign data_r[409] = data_r_409_sv2v_reg;
  assign data_r[408] = data_r_408_sv2v_reg;
  assign data_r[407] = data_r_407_sv2v_reg;
  assign data_r[406] = data_r_406_sv2v_reg;
  assign data_r[405] = data_r_405_sv2v_reg;
  assign data_r[404] = data_r_404_sv2v_reg;
  assign data_r[403] = data_r_403_sv2v_reg;
  assign data_r[402] = data_r_402_sv2v_reg;
  assign data_r[401] = data_r_401_sv2v_reg;
  assign data_r[400] = data_r_400_sv2v_reg;
  assign data_r[399] = data_r_399_sv2v_reg;
  assign data_r[398] = data_r_398_sv2v_reg;
  assign data_r[397] = data_r_397_sv2v_reg;
  assign data_r[396] = data_r_396_sv2v_reg;
  assign data_r[395] = data_r_395_sv2v_reg;
  assign data_r[394] = data_r_394_sv2v_reg;
  assign data_r[393] = data_r_393_sv2v_reg;
  assign data_r[392] = data_r_392_sv2v_reg;
  assign data_r[391] = data_r_391_sv2v_reg;
  assign data_r[390] = data_r_390_sv2v_reg;
  assign data_r[389] = data_r_389_sv2v_reg;
  assign data_r[388] = data_r_388_sv2v_reg;
  assign data_r[387] = data_r_387_sv2v_reg;
  assign data_r[386] = data_r_386_sv2v_reg;
  assign data_r[385] = data_r_385_sv2v_reg;
  assign data_r[384] = data_r_384_sv2v_reg;
  assign data_r[383] = data_r_383_sv2v_reg;
  assign data_r[382] = data_r_382_sv2v_reg;
  assign data_r[381] = data_r_381_sv2v_reg;
  assign data_r[380] = data_r_380_sv2v_reg;
  assign data_r[379] = data_r_379_sv2v_reg;
  assign data_r[378] = data_r_378_sv2v_reg;
  assign data_r[377] = data_r_377_sv2v_reg;
  assign data_r[376] = data_r_376_sv2v_reg;
  assign data_r[375] = data_r_375_sv2v_reg;
  assign data_r[374] = data_r_374_sv2v_reg;
  assign data_r[373] = data_r_373_sv2v_reg;
  assign data_r[372] = data_r_372_sv2v_reg;
  assign data_r[371] = data_r_371_sv2v_reg;
  assign data_r[370] = data_r_370_sv2v_reg;
  assign data_r[369] = data_r_369_sv2v_reg;
  assign data_r[368] = data_r_368_sv2v_reg;
  assign data_r[367] = data_r_367_sv2v_reg;
  assign data_r[366] = data_r_366_sv2v_reg;
  assign data_r[365] = data_r_365_sv2v_reg;
  assign data_r[364] = data_r_364_sv2v_reg;
  assign data_r[363] = data_r_363_sv2v_reg;
  assign data_r[362] = data_r_362_sv2v_reg;
  assign data_r[361] = data_r_361_sv2v_reg;
  assign data_r[360] = data_r_360_sv2v_reg;
  assign data_r[359] = data_r_359_sv2v_reg;
  assign data_r[358] = data_r_358_sv2v_reg;
  assign data_r[357] = data_r_357_sv2v_reg;
  assign data_r[356] = data_r_356_sv2v_reg;
  assign data_r[355] = data_r_355_sv2v_reg;
  assign data_r[354] = data_r_354_sv2v_reg;
  assign data_r[353] = data_r_353_sv2v_reg;
  assign data_r[352] = data_r_352_sv2v_reg;
  assign data_r[351] = data_r_351_sv2v_reg;
  assign data_r[350] = data_r_350_sv2v_reg;
  assign data_r[349] = data_r_349_sv2v_reg;
  assign data_r[348] = data_r_348_sv2v_reg;
  assign data_r[347] = data_r_347_sv2v_reg;
  assign data_r[346] = data_r_346_sv2v_reg;
  assign data_r[345] = data_r_345_sv2v_reg;
  assign data_r[344] = data_r_344_sv2v_reg;
  assign data_r[343] = data_r_343_sv2v_reg;
  assign data_r[342] = data_r_342_sv2v_reg;
  assign data_r[341] = data_r_341_sv2v_reg;
  assign data_r[340] = data_r_340_sv2v_reg;
  assign data_r[339] = data_r_339_sv2v_reg;
  assign data_r[338] = data_r_338_sv2v_reg;
  assign data_r[337] = data_r_337_sv2v_reg;
  assign data_r[336] = data_r_336_sv2v_reg;
  assign data_r[335] = data_r_335_sv2v_reg;
  assign data_r[334] = data_r_334_sv2v_reg;
  assign data_r[333] = data_r_333_sv2v_reg;
  assign data_r[332] = data_r_332_sv2v_reg;
  assign data_r[331] = data_r_331_sv2v_reg;
  assign data_r[330] = data_r_330_sv2v_reg;
  assign data_r[329] = data_r_329_sv2v_reg;
  assign data_r[328] = data_r_328_sv2v_reg;
  assign data_r[327] = data_r_327_sv2v_reg;
  assign data_r[326] = data_r_326_sv2v_reg;
  assign data_r[325] = data_r_325_sv2v_reg;
  assign data_r[324] = data_r_324_sv2v_reg;
  assign data_r[323] = data_r_323_sv2v_reg;
  assign data_r[322] = data_r_322_sv2v_reg;
  assign data_r[321] = data_r_321_sv2v_reg;
  assign data_r[320] = data_r_320_sv2v_reg;
  assign data_r[319] = data_r_319_sv2v_reg;
  assign data_r[318] = data_r_318_sv2v_reg;
  assign data_r[317] = data_r_317_sv2v_reg;
  assign data_r[316] = data_r_316_sv2v_reg;
  assign data_r[315] = data_r_315_sv2v_reg;
  assign data_r[314] = data_r_314_sv2v_reg;
  assign data_r[313] = data_r_313_sv2v_reg;
  assign data_r[312] = data_r_312_sv2v_reg;
  assign data_r[311] = data_r_311_sv2v_reg;
  assign data_r[310] = data_r_310_sv2v_reg;
  assign data_r[309] = data_r_309_sv2v_reg;
  assign data_r[308] = data_r_308_sv2v_reg;
  assign data_r[307] = data_r_307_sv2v_reg;
  assign data_r[306] = data_r_306_sv2v_reg;
  assign data_r[305] = data_r_305_sv2v_reg;
  assign data_r[304] = data_r_304_sv2v_reg;
  assign data_r[303] = data_r_303_sv2v_reg;
  assign data_r[302] = data_r_302_sv2v_reg;
  assign data_r[301] = data_r_301_sv2v_reg;
  assign data_r[300] = data_r_300_sv2v_reg;
  assign data_r[299] = data_r_299_sv2v_reg;
  assign data_r[298] = data_r_298_sv2v_reg;
  assign data_r[297] = data_r_297_sv2v_reg;
  assign data_r[296] = data_r_296_sv2v_reg;
  assign data_r[295] = data_r_295_sv2v_reg;
  assign data_r[294] = data_r_294_sv2v_reg;
  assign data_r[293] = data_r_293_sv2v_reg;
  assign data_r[292] = data_r_292_sv2v_reg;
  assign data_r[291] = data_r_291_sv2v_reg;
  assign data_r[290] = data_r_290_sv2v_reg;
  assign data_r[289] = data_r_289_sv2v_reg;
  assign data_r[288] = data_r_288_sv2v_reg;
  assign data_r[287] = data_r_287_sv2v_reg;
  assign data_r[286] = data_r_286_sv2v_reg;
  assign data_r[285] = data_r_285_sv2v_reg;
  assign data_r[284] = data_r_284_sv2v_reg;
  assign data_r[283] = data_r_283_sv2v_reg;
  assign data_r[282] = data_r_282_sv2v_reg;
  assign data_r[281] = data_r_281_sv2v_reg;
  assign data_r[280] = data_r_280_sv2v_reg;
  assign data_r[279] = data_r_279_sv2v_reg;
  assign data_r[278] = data_r_278_sv2v_reg;
  assign data_r[277] = data_r_277_sv2v_reg;
  assign data_r[276] = data_r_276_sv2v_reg;
  assign data_r[275] = data_r_275_sv2v_reg;
  assign data_r[274] = data_r_274_sv2v_reg;
  assign data_r[273] = data_r_273_sv2v_reg;
  assign data_r[272] = data_r_272_sv2v_reg;
  assign data_r[271] = data_r_271_sv2v_reg;
  assign data_r[270] = data_r_270_sv2v_reg;
  assign data_r[269] = data_r_269_sv2v_reg;
  assign data_r[268] = data_r_268_sv2v_reg;
  assign data_r[267] = data_r_267_sv2v_reg;
  assign data_r[266] = data_r_266_sv2v_reg;
  assign data_r[265] = data_r_265_sv2v_reg;
  assign data_r[264] = data_r_264_sv2v_reg;
  assign data_r[263] = data_r_263_sv2v_reg;
  assign data_r[262] = data_r_262_sv2v_reg;
  assign data_r[261] = data_r_261_sv2v_reg;
  assign data_r[260] = data_r_260_sv2v_reg;
  assign data_r[259] = data_r_259_sv2v_reg;
  assign data_r[258] = data_r_258_sv2v_reg;
  assign data_r[257] = data_r_257_sv2v_reg;
  assign data_r[256] = data_r_256_sv2v_reg;
  assign data_r[255] = data_r_255_sv2v_reg;
  assign data_r[254] = data_r_254_sv2v_reg;
  assign data_r[253] = data_r_253_sv2v_reg;
  assign data_r[252] = data_r_252_sv2v_reg;
  assign data_r[251] = data_r_251_sv2v_reg;
  assign data_r[250] = data_r_250_sv2v_reg;
  assign data_r[249] = data_r_249_sv2v_reg;
  assign data_r[248] = data_r_248_sv2v_reg;
  assign data_r[247] = data_r_247_sv2v_reg;
  assign data_r[246] = data_r_246_sv2v_reg;
  assign data_r[245] = data_r_245_sv2v_reg;
  assign data_r[244] = data_r_244_sv2v_reg;
  assign data_r[243] = data_r_243_sv2v_reg;
  assign data_r[242] = data_r_242_sv2v_reg;
  assign data_r[241] = data_r_241_sv2v_reg;
  assign data_r[240] = data_r_240_sv2v_reg;
  assign data_r[239] = data_r_239_sv2v_reg;
  assign data_r[238] = data_r_238_sv2v_reg;
  assign data_r[237] = data_r_237_sv2v_reg;
  assign data_r[236] = data_r_236_sv2v_reg;
  assign data_r[235] = data_r_235_sv2v_reg;
  assign data_r[234] = data_r_234_sv2v_reg;
  assign data_r[233] = data_r_233_sv2v_reg;
  assign data_r[232] = data_r_232_sv2v_reg;
  assign data_r[231] = data_r_231_sv2v_reg;
  assign data_r[230] = data_r_230_sv2v_reg;
  assign data_r[229] = data_r_229_sv2v_reg;
  assign data_r[228] = data_r_228_sv2v_reg;
  assign data_r[227] = data_r_227_sv2v_reg;
  assign data_r[226] = data_r_226_sv2v_reg;
  assign data_r[225] = data_r_225_sv2v_reg;
  assign data_r[224] = data_r_224_sv2v_reg;
  assign data_r[223] = data_r_223_sv2v_reg;
  assign data_r[222] = data_r_222_sv2v_reg;
  assign data_r[221] = data_r_221_sv2v_reg;
  assign data_r[220] = data_r_220_sv2v_reg;
  assign data_r[219] = data_r_219_sv2v_reg;
  assign data_r[218] = data_r_218_sv2v_reg;
  assign data_r[217] = data_r_217_sv2v_reg;
  assign data_r[216] = data_r_216_sv2v_reg;
  assign data_r[215] = data_r_215_sv2v_reg;
  assign data_r[214] = data_r_214_sv2v_reg;
  assign data_r[213] = data_r_213_sv2v_reg;
  assign data_r[212] = data_r_212_sv2v_reg;
  assign data_r[211] = data_r_211_sv2v_reg;
  assign data_r[210] = data_r_210_sv2v_reg;
  assign data_r[209] = data_r_209_sv2v_reg;
  assign data_r[208] = data_r_208_sv2v_reg;
  assign data_r[207] = data_r_207_sv2v_reg;
  assign data_r[206] = data_r_206_sv2v_reg;
  assign data_r[205] = data_r_205_sv2v_reg;
  assign data_r[204] = data_r_204_sv2v_reg;
  assign data_r[203] = data_r_203_sv2v_reg;
  assign data_r[202] = data_r_202_sv2v_reg;
  assign data_r[201] = data_r_201_sv2v_reg;
  assign data_r[200] = data_r_200_sv2v_reg;
  assign data_r[199] = data_r_199_sv2v_reg;
  assign data_r[198] = data_r_198_sv2v_reg;
  assign data_r[197] = data_r_197_sv2v_reg;
  assign data_r[196] = data_r_196_sv2v_reg;
  assign data_r[195] = data_r_195_sv2v_reg;
  assign data_r[194] = data_r_194_sv2v_reg;
  assign data_r[193] = data_r_193_sv2v_reg;
  assign data_r[192] = data_r_192_sv2v_reg;
  assign data_r[191] = data_r_191_sv2v_reg;
  assign data_r[190] = data_r_190_sv2v_reg;
  assign data_r[189] = data_r_189_sv2v_reg;
  assign data_r[188] = data_r_188_sv2v_reg;
  assign data_r[187] = data_r_187_sv2v_reg;
  assign data_r[186] = data_r_186_sv2v_reg;
  assign data_r[185] = data_r_185_sv2v_reg;
  assign data_r[184] = data_r_184_sv2v_reg;
  assign data_r[183] = data_r_183_sv2v_reg;
  assign data_r[182] = data_r_182_sv2v_reg;
  assign data_r[181] = data_r_181_sv2v_reg;
  assign data_r[180] = data_r_180_sv2v_reg;
  assign data_r[179] = data_r_179_sv2v_reg;
  assign data_r[178] = data_r_178_sv2v_reg;
  assign data_r[177] = data_r_177_sv2v_reg;
  assign data_r[176] = data_r_176_sv2v_reg;
  assign data_r[175] = data_r_175_sv2v_reg;
  assign data_r[174] = data_r_174_sv2v_reg;
  assign data_r[173] = data_r_173_sv2v_reg;
  assign data_r[172] = data_r_172_sv2v_reg;
  assign data_r[171] = data_r_171_sv2v_reg;
  assign data_r[170] = data_r_170_sv2v_reg;
  assign data_r[169] = data_r_169_sv2v_reg;
  assign data_r[168] = data_r_168_sv2v_reg;
  assign data_r[167] = data_r_167_sv2v_reg;
  assign data_r[166] = data_r_166_sv2v_reg;
  assign data_r[165] = data_r_165_sv2v_reg;
  assign data_r[164] = data_r_164_sv2v_reg;
  assign data_r[163] = data_r_163_sv2v_reg;
  assign data_r[162] = data_r_162_sv2v_reg;
  assign data_r[161] = data_r_161_sv2v_reg;
  assign data_r[160] = data_r_160_sv2v_reg;
  assign data_r[159] = data_r_159_sv2v_reg;
  assign data_r[158] = data_r_158_sv2v_reg;
  assign data_r[157] = data_r_157_sv2v_reg;
  assign data_r[156] = data_r_156_sv2v_reg;
  assign data_r[155] = data_r_155_sv2v_reg;
  assign data_r[154] = data_r_154_sv2v_reg;
  assign data_r[153] = data_r_153_sv2v_reg;
  assign data_r[152] = data_r_152_sv2v_reg;
  assign data_r[151] = data_r_151_sv2v_reg;
  assign data_r[150] = data_r_150_sv2v_reg;
  assign data_r[149] = data_r_149_sv2v_reg;
  assign data_r[148] = data_r_148_sv2v_reg;
  assign data_r[147] = data_r_147_sv2v_reg;
  assign data_r[146] = data_r_146_sv2v_reg;
  assign data_r[145] = data_r_145_sv2v_reg;
  assign data_r[144] = data_r_144_sv2v_reg;
  assign data_r[143] = data_r_143_sv2v_reg;
  assign data_r[142] = data_r_142_sv2v_reg;
  assign data_r[141] = data_r_141_sv2v_reg;
  assign data_r[140] = data_r_140_sv2v_reg;
  assign data_r[139] = data_r_139_sv2v_reg;
  assign data_r[138] = data_r_138_sv2v_reg;
  assign data_r[137] = data_r_137_sv2v_reg;
  assign data_r[136] = data_r_136_sv2v_reg;
  assign data_r[135] = data_r_135_sv2v_reg;
  assign data_r[134] = data_r_134_sv2v_reg;
  assign data_r[133] = data_r_133_sv2v_reg;
  assign data_r[132] = data_r_132_sv2v_reg;
  assign data_r[131] = data_r_131_sv2v_reg;
  assign data_r[130] = data_r_130_sv2v_reg;
  assign data_r[129] = data_r_129_sv2v_reg;
  assign data_r[128] = data_r_128_sv2v_reg;
  assign data_r[127] = data_r_127_sv2v_reg;
  assign data_r[126] = data_r_126_sv2v_reg;
  assign data_r[125] = data_r_125_sv2v_reg;
  assign data_r[124] = data_r_124_sv2v_reg;
  assign data_r[123] = data_r_123_sv2v_reg;
  assign data_r[122] = data_r_122_sv2v_reg;
  assign data_r[121] = data_r_121_sv2v_reg;
  assign data_r[120] = data_r_120_sv2v_reg;
  assign data_r[119] = data_r_119_sv2v_reg;
  assign data_r[118] = data_r_118_sv2v_reg;
  assign data_r[117] = data_r_117_sv2v_reg;
  assign data_r[116] = data_r_116_sv2v_reg;
  assign data_r[115] = data_r_115_sv2v_reg;
  assign data_r[114] = data_r_114_sv2v_reg;
  assign data_r[113] = data_r_113_sv2v_reg;
  assign data_r[112] = data_r_112_sv2v_reg;
  assign data_r[111] = data_r_111_sv2v_reg;
  assign data_r[110] = data_r_110_sv2v_reg;
  assign data_r[109] = data_r_109_sv2v_reg;
  assign data_r[108] = data_r_108_sv2v_reg;
  assign data_r[107] = data_r_107_sv2v_reg;
  assign data_r[106] = data_r_106_sv2v_reg;
  assign data_r[105] = data_r_105_sv2v_reg;
  assign data_r[104] = data_r_104_sv2v_reg;
  assign data_r[103] = data_r_103_sv2v_reg;
  assign data_r[102] = data_r_102_sv2v_reg;
  assign data_r[101] = data_r_101_sv2v_reg;
  assign data_r[100] = data_r_100_sv2v_reg;
  assign data_r[99] = data_r_99_sv2v_reg;
  assign data_r[98] = data_r_98_sv2v_reg;
  assign data_r[97] = data_r_97_sv2v_reg;
  assign data_r[96] = data_r_96_sv2v_reg;
  assign data_r[95] = data_r_95_sv2v_reg;
  assign data_r[94] = data_r_94_sv2v_reg;
  assign data_r[93] = data_r_93_sv2v_reg;
  assign data_r[92] = data_r_92_sv2v_reg;
  assign data_r[91] = data_r_91_sv2v_reg;
  assign data_r[90] = data_r_90_sv2v_reg;
  assign data_r[89] = data_r_89_sv2v_reg;
  assign data_r[88] = data_r_88_sv2v_reg;
  assign data_r[87] = data_r_87_sv2v_reg;
  assign data_r[86] = data_r_86_sv2v_reg;
  assign data_r[85] = data_r_85_sv2v_reg;
  assign data_r[84] = data_r_84_sv2v_reg;
  assign data_r[83] = data_r_83_sv2v_reg;
  assign data_r[82] = data_r_82_sv2v_reg;
  assign data_r[81] = data_r_81_sv2v_reg;
  assign data_r[80] = data_r_80_sv2v_reg;
  assign data_r[79] = data_r_79_sv2v_reg;
  assign data_r[78] = data_r_78_sv2v_reg;
  assign data_r[77] = data_r_77_sv2v_reg;
  assign data_r[76] = data_r_76_sv2v_reg;
  assign data_r[75] = data_r_75_sv2v_reg;
  assign data_r[74] = data_r_74_sv2v_reg;
  assign data_r[73] = data_r_73_sv2v_reg;
  assign data_r[72] = data_r_72_sv2v_reg;
  assign data_r[71] = data_r_71_sv2v_reg;
  assign data_r[70] = data_r_70_sv2v_reg;
  assign data_r[69] = data_r_69_sv2v_reg;
  assign data_r[68] = data_r_68_sv2v_reg;
  assign data_r[67] = data_r_67_sv2v_reg;
  assign data_r[66] = data_r_66_sv2v_reg;
  assign data_r[65] = data_r_65_sv2v_reg;
  assign data_r[64] = data_r_64_sv2v_reg;
  assign data_r[63] = data_r_63_sv2v_reg;
  assign data_r[62] = data_r_62_sv2v_reg;
  assign data_r[61] = data_r_61_sv2v_reg;
  assign data_r[60] = data_r_60_sv2v_reg;
  assign data_r[59] = data_r_59_sv2v_reg;
  assign data_r[58] = data_r_58_sv2v_reg;
  assign data_r[57] = data_r_57_sv2v_reg;
  assign data_r[56] = data_r_56_sv2v_reg;
  assign data_r[55] = data_r_55_sv2v_reg;
  assign data_r[54] = data_r_54_sv2v_reg;
  assign data_r[53] = data_r_53_sv2v_reg;
  assign data_r[52] = data_r_52_sv2v_reg;
  assign data_r[51] = data_r_51_sv2v_reg;
  assign data_r[50] = data_r_50_sv2v_reg;
  assign data_r[49] = data_r_49_sv2v_reg;
  assign data_r[48] = data_r_48_sv2v_reg;
  assign data_r[47] = data_r_47_sv2v_reg;
  assign data_r[46] = data_r_46_sv2v_reg;
  assign data_r[45] = data_r_45_sv2v_reg;
  assign data_r[44] = data_r_44_sv2v_reg;
  assign data_r[43] = data_r_43_sv2v_reg;
  assign data_r[42] = data_r_42_sv2v_reg;
  assign data_r[41] = data_r_41_sv2v_reg;
  assign data_r[40] = data_r_40_sv2v_reg;
  assign data_r[39] = data_r_39_sv2v_reg;
  assign data_r[38] = data_r_38_sv2v_reg;
  assign data_r[37] = data_r_37_sv2v_reg;
  assign data_r[36] = data_r_36_sv2v_reg;
  assign data_r[35] = data_r_35_sv2v_reg;
  assign data_r[34] = data_r_34_sv2v_reg;
  assign data_r[33] = data_r_33_sv2v_reg;
  assign data_r[32] = data_r_32_sv2v_reg;
  assign data_r[31] = data_r_31_sv2v_reg;
  assign data_r[30] = data_r_30_sv2v_reg;
  assign data_r[29] = data_r_29_sv2v_reg;
  assign data_r[28] = data_r_28_sv2v_reg;
  assign data_r[27] = data_r_27_sv2v_reg;
  assign data_r[26] = data_r_26_sv2v_reg;
  assign data_r[25] = data_r_25_sv2v_reg;
  assign data_r[24] = data_r_24_sv2v_reg;
  assign data_r[23] = data_r_23_sv2v_reg;
  assign data_r[22] = data_r_22_sv2v_reg;
  assign data_r[21] = data_r_21_sv2v_reg;
  assign data_r[20] = data_r_20_sv2v_reg;
  assign data_r[19] = data_r_19_sv2v_reg;
  assign data_r[18] = data_r_18_sv2v_reg;
  assign data_r[17] = data_r_17_sv2v_reg;
  assign data_r[16] = data_r_16_sv2v_reg;
  assign data_r[15] = data_r_15_sv2v_reg;
  assign data_r[14] = data_r_14_sv2v_reg;
  assign data_r[13] = data_r_13_sv2v_reg;
  assign data_r[12] = data_r_12_sv2v_reg;
  assign data_r[11] = data_r_11_sv2v_reg;
  assign data_r[10] = data_r_10_sv2v_reg;
  assign data_r[9] = data_r_9_sv2v_reg;
  assign data_r[8] = data_r_8_sv2v_reg;
  assign data_r[7] = data_r_7_sv2v_reg;
  assign data_r[6] = data_r_6_sv2v_reg;
  assign data_r[5] = data_r_5_sv2v_reg;
  assign data_r[4] = data_r_4_sv2v_reg;
  assign data_r[3] = data_r_3_sv2v_reg;
  assign data_r[2] = data_r_2_sv2v_reg;
  assign data_r[1] = data_r_1_sv2v_reg;
  assign data_r[0] = data_r_0_sv2v_reg;
  assign data_nn[31] = (N2882)? data_o[31] : 
                       (N2884)? data_o[63] : 
                       (N2886)? data_o[95] : 
                       (N2888)? data_o[127] : 
                       (N2890)? data_o[159] : 
                       (N2892)? data_o[191] : 
                       (N2894)? data_o[223] : 
                       (N2896)? data_o[255] : 
                       (N2898)? data_o[287] : 
                       (N2900)? data_o[319] : 
                       (N2902)? data_o[351] : 
                       (N2904)? data_o[383] : 
                       (N2906)? data_o[415] : 
                       (N2908)? data_o[447] : 
                       (N2910)? data_o[479] : 
                       (N2912)? data_o[511] : 
                       (N2914)? data_o[543] : 
                       (N2916)? data_o[575] : 
                       (N2918)? data_o[607] : 
                       (N2920)? data_o[639] : 
                       (N2922)? data_o[671] : 
                       (N2924)? data_o[703] : 
                       (N2926)? data_o[735] : 
                       (N2928)? data_o[767] : 
                       (N2930)? data_o[799] : 
                       (N2932)? data_o[831] : 
                       (N2934)? data_o[863] : 
                       (N2936)? data_o[895] : 
                       (N2938)? data_o[927] : 
                       (N2940)? data_o[959] : 
                       (N2942)? data_o[991] : 
                       (N2944)? data_o[1023] : 
                       (N2946)? data_o[1055] : 
                       (N2948)? data_o[1087] : 
                       (N2950)? data_o[1119] : 
                       (N2952)? data_o[1151] : 
                       (N2954)? data_o[1183] : 
                       (N2956)? data_o[1215] : 
                       (N2958)? data_o[1247] : 
                       (N2960)? data_o[1279] : 
                       (N2962)? data_o[1311] : 
                       (N2964)? data_o[1343] : 
                       (N2966)? data_o[1375] : 
                       (N2968)? data_o[1407] : 
                       (N2970)? data_o[1439] : 
                       (N2972)? data_o[1471] : 
                       (N2974)? data_o[1503] : 
                       (N2976)? data_o[1535] : 
                       (N2978)? data_o[1567] : 
                       (N2980)? data_o[1599] : 
                       (N2982)? data_o[1631] : 
                       (N2984)? data_o[1663] : 
                       (N2986)? data_o[1695] : 
                       (N2988)? data_o[1727] : 
                       (N2990)? data_o[1759] : 
                       (N2992)? data_o[1791] : 
                       (N2994)? data_o[1823] : 
                       (N2996)? data_o[1855] : 
                       (N2998)? data_o[1887] : 
                       (N3000)? data_o[1919] : 
                       (N3002)? data_o[1951] : 
                       (N3004)? data_o[1983] : 
                       (N3006)? data_o[2015] : 
                       (N3008)? data_o[2047] : 
                       (N2883)? data_n_64__31_ : 
                       (N2885)? data_n_65__31_ : 
                       (N2887)? data_n_66__31_ : 
                       (N2889)? data_n_67__31_ : 
                       (N2891)? data_n_68__31_ : 
                       (N2893)? data_n_69__31_ : 
                       (N2895)? data_n_70__31_ : 
                       (N2897)? data_n_71__31_ : 
                       (N2899)? data_n_72__31_ : 
                       (N2901)? data_n_73__31_ : 
                       (N2903)? data_n_74__31_ : 
                       (N2905)? data_n_75__31_ : 
                       (N2907)? data_n_76__31_ : 
                       (N2909)? data_n_77__31_ : 
                       (N2911)? data_n_78__31_ : 
                       (N2913)? data_n_79__31_ : 
                       (N2915)? data_n_80__31_ : 
                       (N2917)? data_n_81__31_ : 
                       (N2919)? data_n_82__31_ : 
                       (N2921)? data_n_83__31_ : 
                       (N2923)? data_n_84__31_ : 
                       (N2925)? data_n_85__31_ : 
                       (N2927)? data_n_86__31_ : 
                       (N2929)? data_n_87__31_ : 
                       (N2931)? data_n_88__31_ : 
                       (N2933)? data_n_89__31_ : 
                       (N2935)? data_n_90__31_ : 
                       (N2937)? data_n_91__31_ : 
                       (N2939)? data_n_92__31_ : 
                       (N2941)? data_n_93__31_ : 
                       (N2943)? data_n_94__31_ : 
                       (N2945)? data_n_95__31_ : 
                       (N2947)? data_n_96__31_ : 
                       (N2949)? data_n_97__31_ : 
                       (N2951)? data_n_98__31_ : 
                       (N2953)? data_n_99__31_ : 
                       (N2955)? data_n_100__31_ : 
                       (N2957)? data_n_101__31_ : 
                       (N2959)? data_n_102__31_ : 
                       (N2961)? data_n_103__31_ : 
                       (N2963)? data_n_104__31_ : 
                       (N2965)? data_n_105__31_ : 
                       (N2967)? data_n_106__31_ : 
                       (N2969)? data_n_107__31_ : 
                       (N2971)? data_n_108__31_ : 
                       (N2973)? data_n_109__31_ : 
                       (N2975)? data_n_110__31_ : 
                       (N2977)? data_n_111__31_ : 
                       (N2979)? data_n_112__31_ : 
                       (N2981)? data_n_113__31_ : 
                       (N2983)? data_n_114__31_ : 
                       (N2985)? data_n_115__31_ : 
                       (N2987)? data_n_116__31_ : 
                       (N2989)? data_n_117__31_ : 
                       (N2991)? data_n_118__31_ : 
                       (N2993)? data_n_119__31_ : 
                       (N2995)? data_n_120__31_ : 
                       (N2997)? data_n_121__31_ : 
                       (N2999)? data_n_122__31_ : 
                       (N3001)? data_n_123__31_ : 
                       (N3003)? data_n_124__31_ : 
                       (N3005)? data_n_125__31_ : 
                       (N3007)? data_n_126__31_ : 
                       (N3009)? data_n_127__31_ : 1'b0;
  assign data_nn[30] = (N2882)? data_o[30] : 
                       (N2884)? data_o[62] : 
                       (N2886)? data_o[94] : 
                       (N2888)? data_o[126] : 
                       (N2890)? data_o[158] : 
                       (N2892)? data_o[190] : 
                       (N2894)? data_o[222] : 
                       (N2896)? data_o[254] : 
                       (N2898)? data_o[286] : 
                       (N2900)? data_o[318] : 
                       (N2902)? data_o[350] : 
                       (N2904)? data_o[382] : 
                       (N2906)? data_o[414] : 
                       (N2908)? data_o[446] : 
                       (N2910)? data_o[478] : 
                       (N2912)? data_o[510] : 
                       (N2914)? data_o[542] : 
                       (N2916)? data_o[574] : 
                       (N2918)? data_o[606] : 
                       (N2920)? data_o[638] : 
                       (N2922)? data_o[670] : 
                       (N2924)? data_o[702] : 
                       (N2926)? data_o[734] : 
                       (N2928)? data_o[766] : 
                       (N2930)? data_o[798] : 
                       (N2932)? data_o[830] : 
                       (N2934)? data_o[862] : 
                       (N2936)? data_o[894] : 
                       (N2938)? data_o[926] : 
                       (N2940)? data_o[958] : 
                       (N2942)? data_o[990] : 
                       (N2944)? data_o[1022] : 
                       (N2946)? data_o[1054] : 
                       (N2948)? data_o[1086] : 
                       (N2950)? data_o[1118] : 
                       (N2952)? data_o[1150] : 
                       (N2954)? data_o[1182] : 
                       (N2956)? data_o[1214] : 
                       (N2958)? data_o[1246] : 
                       (N2960)? data_o[1278] : 
                       (N2962)? data_o[1310] : 
                       (N2964)? data_o[1342] : 
                       (N2966)? data_o[1374] : 
                       (N2968)? data_o[1406] : 
                       (N2970)? data_o[1438] : 
                       (N2972)? data_o[1470] : 
                       (N2974)? data_o[1502] : 
                       (N2976)? data_o[1534] : 
                       (N2978)? data_o[1566] : 
                       (N2980)? data_o[1598] : 
                       (N2982)? data_o[1630] : 
                       (N2984)? data_o[1662] : 
                       (N2986)? data_o[1694] : 
                       (N2988)? data_o[1726] : 
                       (N2990)? data_o[1758] : 
                       (N2992)? data_o[1790] : 
                       (N2994)? data_o[1822] : 
                       (N2996)? data_o[1854] : 
                       (N2998)? data_o[1886] : 
                       (N3000)? data_o[1918] : 
                       (N3002)? data_o[1950] : 
                       (N3004)? data_o[1982] : 
                       (N3006)? data_o[2014] : 
                       (N3008)? data_o[2046] : 
                       (N2883)? data_n_64__30_ : 
                       (N2885)? data_n_65__30_ : 
                       (N2887)? data_n_66__30_ : 
                       (N2889)? data_n_67__30_ : 
                       (N2891)? data_n_68__30_ : 
                       (N2893)? data_n_69__30_ : 
                       (N2895)? data_n_70__30_ : 
                       (N2897)? data_n_71__30_ : 
                       (N2899)? data_n_72__30_ : 
                       (N2901)? data_n_73__30_ : 
                       (N2903)? data_n_74__30_ : 
                       (N2905)? data_n_75__30_ : 
                       (N2907)? data_n_76__30_ : 
                       (N2909)? data_n_77__30_ : 
                       (N2911)? data_n_78__30_ : 
                       (N2913)? data_n_79__30_ : 
                       (N2915)? data_n_80__30_ : 
                       (N2917)? data_n_81__30_ : 
                       (N2919)? data_n_82__30_ : 
                       (N2921)? data_n_83__30_ : 
                       (N2923)? data_n_84__30_ : 
                       (N2925)? data_n_85__30_ : 
                       (N2927)? data_n_86__30_ : 
                       (N2929)? data_n_87__30_ : 
                       (N2931)? data_n_88__30_ : 
                       (N2933)? data_n_89__30_ : 
                       (N2935)? data_n_90__30_ : 
                       (N2937)? data_n_91__30_ : 
                       (N2939)? data_n_92__30_ : 
                       (N2941)? data_n_93__30_ : 
                       (N2943)? data_n_94__30_ : 
                       (N2945)? data_n_95__30_ : 
                       (N2947)? data_n_96__30_ : 
                       (N2949)? data_n_97__30_ : 
                       (N2951)? data_n_98__30_ : 
                       (N2953)? data_n_99__30_ : 
                       (N2955)? data_n_100__30_ : 
                       (N2957)? data_n_101__30_ : 
                       (N2959)? data_n_102__30_ : 
                       (N2961)? data_n_103__30_ : 
                       (N2963)? data_n_104__30_ : 
                       (N2965)? data_n_105__30_ : 
                       (N2967)? data_n_106__30_ : 
                       (N2969)? data_n_107__30_ : 
                       (N2971)? data_n_108__30_ : 
                       (N2973)? data_n_109__30_ : 
                       (N2975)? data_n_110__30_ : 
                       (N2977)? data_n_111__30_ : 
                       (N2979)? data_n_112__30_ : 
                       (N2981)? data_n_113__30_ : 
                       (N2983)? data_n_114__30_ : 
                       (N2985)? data_n_115__30_ : 
                       (N2987)? data_n_116__30_ : 
                       (N2989)? data_n_117__30_ : 
                       (N2991)? data_n_118__30_ : 
                       (N2993)? data_n_119__30_ : 
                       (N2995)? data_n_120__30_ : 
                       (N2997)? data_n_121__30_ : 
                       (N2999)? data_n_122__30_ : 
                       (N3001)? data_n_123__30_ : 
                       (N3003)? data_n_124__30_ : 
                       (N3005)? data_n_125__30_ : 
                       (N3007)? data_n_126__30_ : 
                       (N3009)? data_n_127__30_ : 1'b0;
  assign data_nn[29] = (N2882)? data_o[29] : 
                       (N2884)? data_o[61] : 
                       (N2886)? data_o[93] : 
                       (N2888)? data_o[125] : 
                       (N2890)? data_o[157] : 
                       (N2892)? data_o[189] : 
                       (N2894)? data_o[221] : 
                       (N2896)? data_o[253] : 
                       (N2898)? data_o[285] : 
                       (N2900)? data_o[317] : 
                       (N2902)? data_o[349] : 
                       (N2904)? data_o[381] : 
                       (N2906)? data_o[413] : 
                       (N2908)? data_o[445] : 
                       (N2910)? data_o[477] : 
                       (N2912)? data_o[509] : 
                       (N2914)? data_o[541] : 
                       (N2916)? data_o[573] : 
                       (N2918)? data_o[605] : 
                       (N2920)? data_o[637] : 
                       (N2922)? data_o[669] : 
                       (N2924)? data_o[701] : 
                       (N2926)? data_o[733] : 
                       (N2928)? data_o[765] : 
                       (N2930)? data_o[797] : 
                       (N2932)? data_o[829] : 
                       (N2934)? data_o[861] : 
                       (N2936)? data_o[893] : 
                       (N2938)? data_o[925] : 
                       (N2940)? data_o[957] : 
                       (N2942)? data_o[989] : 
                       (N2944)? data_o[1021] : 
                       (N2946)? data_o[1053] : 
                       (N2948)? data_o[1085] : 
                       (N2950)? data_o[1117] : 
                       (N2952)? data_o[1149] : 
                       (N2954)? data_o[1181] : 
                       (N2956)? data_o[1213] : 
                       (N2958)? data_o[1245] : 
                       (N2960)? data_o[1277] : 
                       (N2962)? data_o[1309] : 
                       (N2964)? data_o[1341] : 
                       (N2966)? data_o[1373] : 
                       (N2968)? data_o[1405] : 
                       (N2970)? data_o[1437] : 
                       (N2972)? data_o[1469] : 
                       (N2974)? data_o[1501] : 
                       (N2976)? data_o[1533] : 
                       (N2978)? data_o[1565] : 
                       (N2980)? data_o[1597] : 
                       (N2982)? data_o[1629] : 
                       (N2984)? data_o[1661] : 
                       (N2986)? data_o[1693] : 
                       (N2988)? data_o[1725] : 
                       (N2990)? data_o[1757] : 
                       (N2992)? data_o[1789] : 
                       (N2994)? data_o[1821] : 
                       (N2996)? data_o[1853] : 
                       (N2998)? data_o[1885] : 
                       (N3000)? data_o[1917] : 
                       (N3002)? data_o[1949] : 
                       (N3004)? data_o[1981] : 
                       (N3006)? data_o[2013] : 
                       (N3008)? data_o[2045] : 
                       (N2883)? data_n_64__29_ : 
                       (N2885)? data_n_65__29_ : 
                       (N2887)? data_n_66__29_ : 
                       (N2889)? data_n_67__29_ : 
                       (N2891)? data_n_68__29_ : 
                       (N2893)? data_n_69__29_ : 
                       (N2895)? data_n_70__29_ : 
                       (N2897)? data_n_71__29_ : 
                       (N2899)? data_n_72__29_ : 
                       (N2901)? data_n_73__29_ : 
                       (N2903)? data_n_74__29_ : 
                       (N2905)? data_n_75__29_ : 
                       (N2907)? data_n_76__29_ : 
                       (N2909)? data_n_77__29_ : 
                       (N2911)? data_n_78__29_ : 
                       (N2913)? data_n_79__29_ : 
                       (N2915)? data_n_80__29_ : 
                       (N2917)? data_n_81__29_ : 
                       (N2919)? data_n_82__29_ : 
                       (N2921)? data_n_83__29_ : 
                       (N2923)? data_n_84__29_ : 
                       (N2925)? data_n_85__29_ : 
                       (N2927)? data_n_86__29_ : 
                       (N2929)? data_n_87__29_ : 
                       (N2931)? data_n_88__29_ : 
                       (N2933)? data_n_89__29_ : 
                       (N2935)? data_n_90__29_ : 
                       (N2937)? data_n_91__29_ : 
                       (N2939)? data_n_92__29_ : 
                       (N2941)? data_n_93__29_ : 
                       (N2943)? data_n_94__29_ : 
                       (N2945)? data_n_95__29_ : 
                       (N2947)? data_n_96__29_ : 
                       (N2949)? data_n_97__29_ : 
                       (N2951)? data_n_98__29_ : 
                       (N2953)? data_n_99__29_ : 
                       (N2955)? data_n_100__29_ : 
                       (N2957)? data_n_101__29_ : 
                       (N2959)? data_n_102__29_ : 
                       (N2961)? data_n_103__29_ : 
                       (N2963)? data_n_104__29_ : 
                       (N2965)? data_n_105__29_ : 
                       (N2967)? data_n_106__29_ : 
                       (N2969)? data_n_107__29_ : 
                       (N2971)? data_n_108__29_ : 
                       (N2973)? data_n_109__29_ : 
                       (N2975)? data_n_110__29_ : 
                       (N2977)? data_n_111__29_ : 
                       (N2979)? data_n_112__29_ : 
                       (N2981)? data_n_113__29_ : 
                       (N2983)? data_n_114__29_ : 
                       (N2985)? data_n_115__29_ : 
                       (N2987)? data_n_116__29_ : 
                       (N2989)? data_n_117__29_ : 
                       (N2991)? data_n_118__29_ : 
                       (N2993)? data_n_119__29_ : 
                       (N2995)? data_n_120__29_ : 
                       (N2997)? data_n_121__29_ : 
                       (N2999)? data_n_122__29_ : 
                       (N3001)? data_n_123__29_ : 
                       (N3003)? data_n_124__29_ : 
                       (N3005)? data_n_125__29_ : 
                       (N3007)? data_n_126__29_ : 
                       (N3009)? data_n_127__29_ : 1'b0;
  assign data_nn[28] = (N2882)? data_o[28] : 
                       (N2884)? data_o[60] : 
                       (N2886)? data_o[92] : 
                       (N2888)? data_o[124] : 
                       (N2890)? data_o[156] : 
                       (N2892)? data_o[188] : 
                       (N2894)? data_o[220] : 
                       (N2896)? data_o[252] : 
                       (N2898)? data_o[284] : 
                       (N2900)? data_o[316] : 
                       (N2902)? data_o[348] : 
                       (N2904)? data_o[380] : 
                       (N2906)? data_o[412] : 
                       (N2908)? data_o[444] : 
                       (N2910)? data_o[476] : 
                       (N2912)? data_o[508] : 
                       (N2914)? data_o[540] : 
                       (N2916)? data_o[572] : 
                       (N2918)? data_o[604] : 
                       (N2920)? data_o[636] : 
                       (N2922)? data_o[668] : 
                       (N2924)? data_o[700] : 
                       (N2926)? data_o[732] : 
                       (N2928)? data_o[764] : 
                       (N2930)? data_o[796] : 
                       (N2932)? data_o[828] : 
                       (N2934)? data_o[860] : 
                       (N2936)? data_o[892] : 
                       (N2938)? data_o[924] : 
                       (N2940)? data_o[956] : 
                       (N2942)? data_o[988] : 
                       (N2944)? data_o[1020] : 
                       (N2946)? data_o[1052] : 
                       (N2948)? data_o[1084] : 
                       (N2950)? data_o[1116] : 
                       (N2952)? data_o[1148] : 
                       (N2954)? data_o[1180] : 
                       (N2956)? data_o[1212] : 
                       (N2958)? data_o[1244] : 
                       (N2960)? data_o[1276] : 
                       (N2962)? data_o[1308] : 
                       (N2964)? data_o[1340] : 
                       (N2966)? data_o[1372] : 
                       (N2968)? data_o[1404] : 
                       (N2970)? data_o[1436] : 
                       (N2972)? data_o[1468] : 
                       (N2974)? data_o[1500] : 
                       (N2976)? data_o[1532] : 
                       (N2978)? data_o[1564] : 
                       (N2980)? data_o[1596] : 
                       (N2982)? data_o[1628] : 
                       (N2984)? data_o[1660] : 
                       (N2986)? data_o[1692] : 
                       (N2988)? data_o[1724] : 
                       (N2990)? data_o[1756] : 
                       (N2992)? data_o[1788] : 
                       (N2994)? data_o[1820] : 
                       (N2996)? data_o[1852] : 
                       (N2998)? data_o[1884] : 
                       (N3000)? data_o[1916] : 
                       (N3002)? data_o[1948] : 
                       (N3004)? data_o[1980] : 
                       (N3006)? data_o[2012] : 
                       (N3008)? data_o[2044] : 
                       (N2883)? data_n_64__28_ : 
                       (N2885)? data_n_65__28_ : 
                       (N2887)? data_n_66__28_ : 
                       (N2889)? data_n_67__28_ : 
                       (N2891)? data_n_68__28_ : 
                       (N2893)? data_n_69__28_ : 
                       (N2895)? data_n_70__28_ : 
                       (N2897)? data_n_71__28_ : 
                       (N2899)? data_n_72__28_ : 
                       (N2901)? data_n_73__28_ : 
                       (N2903)? data_n_74__28_ : 
                       (N2905)? data_n_75__28_ : 
                       (N2907)? data_n_76__28_ : 
                       (N2909)? data_n_77__28_ : 
                       (N2911)? data_n_78__28_ : 
                       (N2913)? data_n_79__28_ : 
                       (N2915)? data_n_80__28_ : 
                       (N2917)? data_n_81__28_ : 
                       (N2919)? data_n_82__28_ : 
                       (N2921)? data_n_83__28_ : 
                       (N2923)? data_n_84__28_ : 
                       (N2925)? data_n_85__28_ : 
                       (N2927)? data_n_86__28_ : 
                       (N2929)? data_n_87__28_ : 
                       (N2931)? data_n_88__28_ : 
                       (N2933)? data_n_89__28_ : 
                       (N2935)? data_n_90__28_ : 
                       (N2937)? data_n_91__28_ : 
                       (N2939)? data_n_92__28_ : 
                       (N2941)? data_n_93__28_ : 
                       (N2943)? data_n_94__28_ : 
                       (N2945)? data_n_95__28_ : 
                       (N2947)? data_n_96__28_ : 
                       (N2949)? data_n_97__28_ : 
                       (N2951)? data_n_98__28_ : 
                       (N2953)? data_n_99__28_ : 
                       (N2955)? data_n_100__28_ : 
                       (N2957)? data_n_101__28_ : 
                       (N2959)? data_n_102__28_ : 
                       (N2961)? data_n_103__28_ : 
                       (N2963)? data_n_104__28_ : 
                       (N2965)? data_n_105__28_ : 
                       (N2967)? data_n_106__28_ : 
                       (N2969)? data_n_107__28_ : 
                       (N2971)? data_n_108__28_ : 
                       (N2973)? data_n_109__28_ : 
                       (N2975)? data_n_110__28_ : 
                       (N2977)? data_n_111__28_ : 
                       (N2979)? data_n_112__28_ : 
                       (N2981)? data_n_113__28_ : 
                       (N2983)? data_n_114__28_ : 
                       (N2985)? data_n_115__28_ : 
                       (N2987)? data_n_116__28_ : 
                       (N2989)? data_n_117__28_ : 
                       (N2991)? data_n_118__28_ : 
                       (N2993)? data_n_119__28_ : 
                       (N2995)? data_n_120__28_ : 
                       (N2997)? data_n_121__28_ : 
                       (N2999)? data_n_122__28_ : 
                       (N3001)? data_n_123__28_ : 
                       (N3003)? data_n_124__28_ : 
                       (N3005)? data_n_125__28_ : 
                       (N3007)? data_n_126__28_ : 
                       (N3009)? data_n_127__28_ : 1'b0;
  assign data_nn[27] = (N2882)? data_o[27] : 
                       (N2884)? data_o[59] : 
                       (N2886)? data_o[91] : 
                       (N2888)? data_o[123] : 
                       (N2890)? data_o[155] : 
                       (N2892)? data_o[187] : 
                       (N2894)? data_o[219] : 
                       (N2896)? data_o[251] : 
                       (N2898)? data_o[283] : 
                       (N2900)? data_o[315] : 
                       (N2902)? data_o[347] : 
                       (N2904)? data_o[379] : 
                       (N2906)? data_o[411] : 
                       (N2908)? data_o[443] : 
                       (N2910)? data_o[475] : 
                       (N2912)? data_o[507] : 
                       (N2914)? data_o[539] : 
                       (N2916)? data_o[571] : 
                       (N2918)? data_o[603] : 
                       (N2920)? data_o[635] : 
                       (N2922)? data_o[667] : 
                       (N2924)? data_o[699] : 
                       (N2926)? data_o[731] : 
                       (N2928)? data_o[763] : 
                       (N2930)? data_o[795] : 
                       (N2932)? data_o[827] : 
                       (N2934)? data_o[859] : 
                       (N2936)? data_o[891] : 
                       (N2938)? data_o[923] : 
                       (N2940)? data_o[955] : 
                       (N2942)? data_o[987] : 
                       (N2944)? data_o[1019] : 
                       (N2946)? data_o[1051] : 
                       (N2948)? data_o[1083] : 
                       (N2950)? data_o[1115] : 
                       (N2952)? data_o[1147] : 
                       (N2954)? data_o[1179] : 
                       (N2956)? data_o[1211] : 
                       (N2958)? data_o[1243] : 
                       (N2960)? data_o[1275] : 
                       (N2962)? data_o[1307] : 
                       (N2964)? data_o[1339] : 
                       (N2966)? data_o[1371] : 
                       (N2968)? data_o[1403] : 
                       (N2970)? data_o[1435] : 
                       (N2972)? data_o[1467] : 
                       (N2974)? data_o[1499] : 
                       (N2976)? data_o[1531] : 
                       (N2978)? data_o[1563] : 
                       (N2980)? data_o[1595] : 
                       (N2982)? data_o[1627] : 
                       (N2984)? data_o[1659] : 
                       (N2986)? data_o[1691] : 
                       (N2988)? data_o[1723] : 
                       (N2990)? data_o[1755] : 
                       (N2992)? data_o[1787] : 
                       (N2994)? data_o[1819] : 
                       (N2996)? data_o[1851] : 
                       (N2998)? data_o[1883] : 
                       (N3000)? data_o[1915] : 
                       (N3002)? data_o[1947] : 
                       (N3004)? data_o[1979] : 
                       (N3006)? data_o[2011] : 
                       (N3008)? data_o[2043] : 
                       (N2883)? data_n_64__27_ : 
                       (N2885)? data_n_65__27_ : 
                       (N2887)? data_n_66__27_ : 
                       (N2889)? data_n_67__27_ : 
                       (N2891)? data_n_68__27_ : 
                       (N2893)? data_n_69__27_ : 
                       (N2895)? data_n_70__27_ : 
                       (N2897)? data_n_71__27_ : 
                       (N2899)? data_n_72__27_ : 
                       (N2901)? data_n_73__27_ : 
                       (N2903)? data_n_74__27_ : 
                       (N2905)? data_n_75__27_ : 
                       (N2907)? data_n_76__27_ : 
                       (N2909)? data_n_77__27_ : 
                       (N2911)? data_n_78__27_ : 
                       (N2913)? data_n_79__27_ : 
                       (N2915)? data_n_80__27_ : 
                       (N2917)? data_n_81__27_ : 
                       (N2919)? data_n_82__27_ : 
                       (N2921)? data_n_83__27_ : 
                       (N2923)? data_n_84__27_ : 
                       (N2925)? data_n_85__27_ : 
                       (N2927)? data_n_86__27_ : 
                       (N2929)? data_n_87__27_ : 
                       (N2931)? data_n_88__27_ : 
                       (N2933)? data_n_89__27_ : 
                       (N2935)? data_n_90__27_ : 
                       (N2937)? data_n_91__27_ : 
                       (N2939)? data_n_92__27_ : 
                       (N2941)? data_n_93__27_ : 
                       (N2943)? data_n_94__27_ : 
                       (N2945)? data_n_95__27_ : 
                       (N2947)? data_n_96__27_ : 
                       (N2949)? data_n_97__27_ : 
                       (N2951)? data_n_98__27_ : 
                       (N2953)? data_n_99__27_ : 
                       (N2955)? data_n_100__27_ : 
                       (N2957)? data_n_101__27_ : 
                       (N2959)? data_n_102__27_ : 
                       (N2961)? data_n_103__27_ : 
                       (N2963)? data_n_104__27_ : 
                       (N2965)? data_n_105__27_ : 
                       (N2967)? data_n_106__27_ : 
                       (N2969)? data_n_107__27_ : 
                       (N2971)? data_n_108__27_ : 
                       (N2973)? data_n_109__27_ : 
                       (N2975)? data_n_110__27_ : 
                       (N2977)? data_n_111__27_ : 
                       (N2979)? data_n_112__27_ : 
                       (N2981)? data_n_113__27_ : 
                       (N2983)? data_n_114__27_ : 
                       (N2985)? data_n_115__27_ : 
                       (N2987)? data_n_116__27_ : 
                       (N2989)? data_n_117__27_ : 
                       (N2991)? data_n_118__27_ : 
                       (N2993)? data_n_119__27_ : 
                       (N2995)? data_n_120__27_ : 
                       (N2997)? data_n_121__27_ : 
                       (N2999)? data_n_122__27_ : 
                       (N3001)? data_n_123__27_ : 
                       (N3003)? data_n_124__27_ : 
                       (N3005)? data_n_125__27_ : 
                       (N3007)? data_n_126__27_ : 
                       (N3009)? data_n_127__27_ : 1'b0;
  assign data_nn[26] = (N2882)? data_o[26] : 
                       (N2884)? data_o[58] : 
                       (N2886)? data_o[90] : 
                       (N2888)? data_o[122] : 
                       (N2890)? data_o[154] : 
                       (N2892)? data_o[186] : 
                       (N2894)? data_o[218] : 
                       (N2896)? data_o[250] : 
                       (N2898)? data_o[282] : 
                       (N2900)? data_o[314] : 
                       (N2902)? data_o[346] : 
                       (N2904)? data_o[378] : 
                       (N2906)? data_o[410] : 
                       (N2908)? data_o[442] : 
                       (N2910)? data_o[474] : 
                       (N2912)? data_o[506] : 
                       (N2914)? data_o[538] : 
                       (N2916)? data_o[570] : 
                       (N2918)? data_o[602] : 
                       (N2920)? data_o[634] : 
                       (N2922)? data_o[666] : 
                       (N2924)? data_o[698] : 
                       (N2926)? data_o[730] : 
                       (N2928)? data_o[762] : 
                       (N2930)? data_o[794] : 
                       (N2932)? data_o[826] : 
                       (N2934)? data_o[858] : 
                       (N2936)? data_o[890] : 
                       (N2938)? data_o[922] : 
                       (N2940)? data_o[954] : 
                       (N2942)? data_o[986] : 
                       (N2944)? data_o[1018] : 
                       (N2946)? data_o[1050] : 
                       (N2948)? data_o[1082] : 
                       (N2950)? data_o[1114] : 
                       (N2952)? data_o[1146] : 
                       (N2954)? data_o[1178] : 
                       (N2956)? data_o[1210] : 
                       (N2958)? data_o[1242] : 
                       (N2960)? data_o[1274] : 
                       (N2962)? data_o[1306] : 
                       (N2964)? data_o[1338] : 
                       (N2966)? data_o[1370] : 
                       (N2968)? data_o[1402] : 
                       (N2970)? data_o[1434] : 
                       (N2972)? data_o[1466] : 
                       (N2974)? data_o[1498] : 
                       (N2976)? data_o[1530] : 
                       (N2978)? data_o[1562] : 
                       (N2980)? data_o[1594] : 
                       (N2982)? data_o[1626] : 
                       (N2984)? data_o[1658] : 
                       (N2986)? data_o[1690] : 
                       (N2988)? data_o[1722] : 
                       (N2990)? data_o[1754] : 
                       (N2992)? data_o[1786] : 
                       (N2994)? data_o[1818] : 
                       (N2996)? data_o[1850] : 
                       (N2998)? data_o[1882] : 
                       (N3000)? data_o[1914] : 
                       (N3002)? data_o[1946] : 
                       (N3004)? data_o[1978] : 
                       (N3006)? data_o[2010] : 
                       (N3008)? data_o[2042] : 
                       (N2883)? data_n_64__26_ : 
                       (N2885)? data_n_65__26_ : 
                       (N2887)? data_n_66__26_ : 
                       (N2889)? data_n_67__26_ : 
                       (N2891)? data_n_68__26_ : 
                       (N2893)? data_n_69__26_ : 
                       (N2895)? data_n_70__26_ : 
                       (N2897)? data_n_71__26_ : 
                       (N2899)? data_n_72__26_ : 
                       (N2901)? data_n_73__26_ : 
                       (N2903)? data_n_74__26_ : 
                       (N2905)? data_n_75__26_ : 
                       (N2907)? data_n_76__26_ : 
                       (N2909)? data_n_77__26_ : 
                       (N2911)? data_n_78__26_ : 
                       (N2913)? data_n_79__26_ : 
                       (N2915)? data_n_80__26_ : 
                       (N2917)? data_n_81__26_ : 
                       (N2919)? data_n_82__26_ : 
                       (N2921)? data_n_83__26_ : 
                       (N2923)? data_n_84__26_ : 
                       (N2925)? data_n_85__26_ : 
                       (N2927)? data_n_86__26_ : 
                       (N2929)? data_n_87__26_ : 
                       (N2931)? data_n_88__26_ : 
                       (N2933)? data_n_89__26_ : 
                       (N2935)? data_n_90__26_ : 
                       (N2937)? data_n_91__26_ : 
                       (N2939)? data_n_92__26_ : 
                       (N2941)? data_n_93__26_ : 
                       (N2943)? data_n_94__26_ : 
                       (N2945)? data_n_95__26_ : 
                       (N2947)? data_n_96__26_ : 
                       (N2949)? data_n_97__26_ : 
                       (N2951)? data_n_98__26_ : 
                       (N2953)? data_n_99__26_ : 
                       (N2955)? data_n_100__26_ : 
                       (N2957)? data_n_101__26_ : 
                       (N2959)? data_n_102__26_ : 
                       (N2961)? data_n_103__26_ : 
                       (N2963)? data_n_104__26_ : 
                       (N2965)? data_n_105__26_ : 
                       (N2967)? data_n_106__26_ : 
                       (N2969)? data_n_107__26_ : 
                       (N2971)? data_n_108__26_ : 
                       (N2973)? data_n_109__26_ : 
                       (N2975)? data_n_110__26_ : 
                       (N2977)? data_n_111__26_ : 
                       (N2979)? data_n_112__26_ : 
                       (N2981)? data_n_113__26_ : 
                       (N2983)? data_n_114__26_ : 
                       (N2985)? data_n_115__26_ : 
                       (N2987)? data_n_116__26_ : 
                       (N2989)? data_n_117__26_ : 
                       (N2991)? data_n_118__26_ : 
                       (N2993)? data_n_119__26_ : 
                       (N2995)? data_n_120__26_ : 
                       (N2997)? data_n_121__26_ : 
                       (N2999)? data_n_122__26_ : 
                       (N3001)? data_n_123__26_ : 
                       (N3003)? data_n_124__26_ : 
                       (N3005)? data_n_125__26_ : 
                       (N3007)? data_n_126__26_ : 
                       (N3009)? data_n_127__26_ : 1'b0;
  assign data_nn[25] = (N2882)? data_o[25] : 
                       (N2884)? data_o[57] : 
                       (N2886)? data_o[89] : 
                       (N2888)? data_o[121] : 
                       (N2890)? data_o[153] : 
                       (N2892)? data_o[185] : 
                       (N2894)? data_o[217] : 
                       (N2896)? data_o[249] : 
                       (N2898)? data_o[281] : 
                       (N2900)? data_o[313] : 
                       (N2902)? data_o[345] : 
                       (N2904)? data_o[377] : 
                       (N2906)? data_o[409] : 
                       (N2908)? data_o[441] : 
                       (N2910)? data_o[473] : 
                       (N2912)? data_o[505] : 
                       (N2914)? data_o[537] : 
                       (N2916)? data_o[569] : 
                       (N2918)? data_o[601] : 
                       (N2920)? data_o[633] : 
                       (N2922)? data_o[665] : 
                       (N2924)? data_o[697] : 
                       (N2926)? data_o[729] : 
                       (N2928)? data_o[761] : 
                       (N2930)? data_o[793] : 
                       (N2932)? data_o[825] : 
                       (N2934)? data_o[857] : 
                       (N2936)? data_o[889] : 
                       (N2938)? data_o[921] : 
                       (N2940)? data_o[953] : 
                       (N2942)? data_o[985] : 
                       (N2944)? data_o[1017] : 
                       (N2946)? data_o[1049] : 
                       (N2948)? data_o[1081] : 
                       (N2950)? data_o[1113] : 
                       (N2952)? data_o[1145] : 
                       (N2954)? data_o[1177] : 
                       (N2956)? data_o[1209] : 
                       (N2958)? data_o[1241] : 
                       (N2960)? data_o[1273] : 
                       (N2962)? data_o[1305] : 
                       (N2964)? data_o[1337] : 
                       (N2966)? data_o[1369] : 
                       (N2968)? data_o[1401] : 
                       (N2970)? data_o[1433] : 
                       (N2972)? data_o[1465] : 
                       (N2974)? data_o[1497] : 
                       (N2976)? data_o[1529] : 
                       (N2978)? data_o[1561] : 
                       (N2980)? data_o[1593] : 
                       (N2982)? data_o[1625] : 
                       (N2984)? data_o[1657] : 
                       (N2986)? data_o[1689] : 
                       (N2988)? data_o[1721] : 
                       (N2990)? data_o[1753] : 
                       (N2992)? data_o[1785] : 
                       (N2994)? data_o[1817] : 
                       (N2996)? data_o[1849] : 
                       (N2998)? data_o[1881] : 
                       (N3000)? data_o[1913] : 
                       (N3002)? data_o[1945] : 
                       (N3004)? data_o[1977] : 
                       (N3006)? data_o[2009] : 
                       (N3008)? data_o[2041] : 
                       (N2883)? data_n_64__25_ : 
                       (N2885)? data_n_65__25_ : 
                       (N2887)? data_n_66__25_ : 
                       (N2889)? data_n_67__25_ : 
                       (N2891)? data_n_68__25_ : 
                       (N2893)? data_n_69__25_ : 
                       (N2895)? data_n_70__25_ : 
                       (N2897)? data_n_71__25_ : 
                       (N2899)? data_n_72__25_ : 
                       (N2901)? data_n_73__25_ : 
                       (N2903)? data_n_74__25_ : 
                       (N2905)? data_n_75__25_ : 
                       (N2907)? data_n_76__25_ : 
                       (N2909)? data_n_77__25_ : 
                       (N2911)? data_n_78__25_ : 
                       (N2913)? data_n_79__25_ : 
                       (N2915)? data_n_80__25_ : 
                       (N2917)? data_n_81__25_ : 
                       (N2919)? data_n_82__25_ : 
                       (N2921)? data_n_83__25_ : 
                       (N2923)? data_n_84__25_ : 
                       (N2925)? data_n_85__25_ : 
                       (N2927)? data_n_86__25_ : 
                       (N2929)? data_n_87__25_ : 
                       (N2931)? data_n_88__25_ : 
                       (N2933)? data_n_89__25_ : 
                       (N2935)? data_n_90__25_ : 
                       (N2937)? data_n_91__25_ : 
                       (N2939)? data_n_92__25_ : 
                       (N2941)? data_n_93__25_ : 
                       (N2943)? data_n_94__25_ : 
                       (N2945)? data_n_95__25_ : 
                       (N2947)? data_n_96__25_ : 
                       (N2949)? data_n_97__25_ : 
                       (N2951)? data_n_98__25_ : 
                       (N2953)? data_n_99__25_ : 
                       (N2955)? data_n_100__25_ : 
                       (N2957)? data_n_101__25_ : 
                       (N2959)? data_n_102__25_ : 
                       (N2961)? data_n_103__25_ : 
                       (N2963)? data_n_104__25_ : 
                       (N2965)? data_n_105__25_ : 
                       (N2967)? data_n_106__25_ : 
                       (N2969)? data_n_107__25_ : 
                       (N2971)? data_n_108__25_ : 
                       (N2973)? data_n_109__25_ : 
                       (N2975)? data_n_110__25_ : 
                       (N2977)? data_n_111__25_ : 
                       (N2979)? data_n_112__25_ : 
                       (N2981)? data_n_113__25_ : 
                       (N2983)? data_n_114__25_ : 
                       (N2985)? data_n_115__25_ : 
                       (N2987)? data_n_116__25_ : 
                       (N2989)? data_n_117__25_ : 
                       (N2991)? data_n_118__25_ : 
                       (N2993)? data_n_119__25_ : 
                       (N2995)? data_n_120__25_ : 
                       (N2997)? data_n_121__25_ : 
                       (N2999)? data_n_122__25_ : 
                       (N3001)? data_n_123__25_ : 
                       (N3003)? data_n_124__25_ : 
                       (N3005)? data_n_125__25_ : 
                       (N3007)? data_n_126__25_ : 
                       (N3009)? data_n_127__25_ : 1'b0;
  assign data_nn[24] = (N2882)? data_o[24] : 
                       (N2884)? data_o[56] : 
                       (N2886)? data_o[88] : 
                       (N2888)? data_o[120] : 
                       (N2890)? data_o[152] : 
                       (N2892)? data_o[184] : 
                       (N2894)? data_o[216] : 
                       (N2896)? data_o[248] : 
                       (N2898)? data_o[280] : 
                       (N2900)? data_o[312] : 
                       (N2902)? data_o[344] : 
                       (N2904)? data_o[376] : 
                       (N2906)? data_o[408] : 
                       (N2908)? data_o[440] : 
                       (N2910)? data_o[472] : 
                       (N2912)? data_o[504] : 
                       (N2914)? data_o[536] : 
                       (N2916)? data_o[568] : 
                       (N2918)? data_o[600] : 
                       (N2920)? data_o[632] : 
                       (N2922)? data_o[664] : 
                       (N2924)? data_o[696] : 
                       (N2926)? data_o[728] : 
                       (N2928)? data_o[760] : 
                       (N2930)? data_o[792] : 
                       (N2932)? data_o[824] : 
                       (N2934)? data_o[856] : 
                       (N2936)? data_o[888] : 
                       (N2938)? data_o[920] : 
                       (N2940)? data_o[952] : 
                       (N2942)? data_o[984] : 
                       (N2944)? data_o[1016] : 
                       (N2946)? data_o[1048] : 
                       (N2948)? data_o[1080] : 
                       (N2950)? data_o[1112] : 
                       (N2952)? data_o[1144] : 
                       (N2954)? data_o[1176] : 
                       (N2956)? data_o[1208] : 
                       (N2958)? data_o[1240] : 
                       (N2960)? data_o[1272] : 
                       (N2962)? data_o[1304] : 
                       (N2964)? data_o[1336] : 
                       (N2966)? data_o[1368] : 
                       (N2968)? data_o[1400] : 
                       (N2970)? data_o[1432] : 
                       (N2972)? data_o[1464] : 
                       (N2974)? data_o[1496] : 
                       (N2976)? data_o[1528] : 
                       (N2978)? data_o[1560] : 
                       (N2980)? data_o[1592] : 
                       (N2982)? data_o[1624] : 
                       (N2984)? data_o[1656] : 
                       (N2986)? data_o[1688] : 
                       (N2988)? data_o[1720] : 
                       (N2990)? data_o[1752] : 
                       (N2992)? data_o[1784] : 
                       (N2994)? data_o[1816] : 
                       (N2996)? data_o[1848] : 
                       (N2998)? data_o[1880] : 
                       (N3000)? data_o[1912] : 
                       (N3002)? data_o[1944] : 
                       (N3004)? data_o[1976] : 
                       (N3006)? data_o[2008] : 
                       (N3008)? data_o[2040] : 
                       (N2883)? data_n_64__24_ : 
                       (N2885)? data_n_65__24_ : 
                       (N2887)? data_n_66__24_ : 
                       (N2889)? data_n_67__24_ : 
                       (N2891)? data_n_68__24_ : 
                       (N2893)? data_n_69__24_ : 
                       (N2895)? data_n_70__24_ : 
                       (N2897)? data_n_71__24_ : 
                       (N2899)? data_n_72__24_ : 
                       (N2901)? data_n_73__24_ : 
                       (N2903)? data_n_74__24_ : 
                       (N2905)? data_n_75__24_ : 
                       (N2907)? data_n_76__24_ : 
                       (N2909)? data_n_77__24_ : 
                       (N2911)? data_n_78__24_ : 
                       (N2913)? data_n_79__24_ : 
                       (N2915)? data_n_80__24_ : 
                       (N2917)? data_n_81__24_ : 
                       (N2919)? data_n_82__24_ : 
                       (N2921)? data_n_83__24_ : 
                       (N2923)? data_n_84__24_ : 
                       (N2925)? data_n_85__24_ : 
                       (N2927)? data_n_86__24_ : 
                       (N2929)? data_n_87__24_ : 
                       (N2931)? data_n_88__24_ : 
                       (N2933)? data_n_89__24_ : 
                       (N2935)? data_n_90__24_ : 
                       (N2937)? data_n_91__24_ : 
                       (N2939)? data_n_92__24_ : 
                       (N2941)? data_n_93__24_ : 
                       (N2943)? data_n_94__24_ : 
                       (N2945)? data_n_95__24_ : 
                       (N2947)? data_n_96__24_ : 
                       (N2949)? data_n_97__24_ : 
                       (N2951)? data_n_98__24_ : 
                       (N2953)? data_n_99__24_ : 
                       (N2955)? data_n_100__24_ : 
                       (N2957)? data_n_101__24_ : 
                       (N2959)? data_n_102__24_ : 
                       (N2961)? data_n_103__24_ : 
                       (N2963)? data_n_104__24_ : 
                       (N2965)? data_n_105__24_ : 
                       (N2967)? data_n_106__24_ : 
                       (N2969)? data_n_107__24_ : 
                       (N2971)? data_n_108__24_ : 
                       (N2973)? data_n_109__24_ : 
                       (N2975)? data_n_110__24_ : 
                       (N2977)? data_n_111__24_ : 
                       (N2979)? data_n_112__24_ : 
                       (N2981)? data_n_113__24_ : 
                       (N2983)? data_n_114__24_ : 
                       (N2985)? data_n_115__24_ : 
                       (N2987)? data_n_116__24_ : 
                       (N2989)? data_n_117__24_ : 
                       (N2991)? data_n_118__24_ : 
                       (N2993)? data_n_119__24_ : 
                       (N2995)? data_n_120__24_ : 
                       (N2997)? data_n_121__24_ : 
                       (N2999)? data_n_122__24_ : 
                       (N3001)? data_n_123__24_ : 
                       (N3003)? data_n_124__24_ : 
                       (N3005)? data_n_125__24_ : 
                       (N3007)? data_n_126__24_ : 
                       (N3009)? data_n_127__24_ : 1'b0;
  assign data_nn[23] = (N2882)? data_o[23] : 
                       (N2884)? data_o[55] : 
                       (N2886)? data_o[87] : 
                       (N2888)? data_o[119] : 
                       (N2890)? data_o[151] : 
                       (N2892)? data_o[183] : 
                       (N2894)? data_o[215] : 
                       (N2896)? data_o[247] : 
                       (N2898)? data_o[279] : 
                       (N2900)? data_o[311] : 
                       (N2902)? data_o[343] : 
                       (N2904)? data_o[375] : 
                       (N2906)? data_o[407] : 
                       (N2908)? data_o[439] : 
                       (N2910)? data_o[471] : 
                       (N2912)? data_o[503] : 
                       (N2914)? data_o[535] : 
                       (N2916)? data_o[567] : 
                       (N2918)? data_o[599] : 
                       (N2920)? data_o[631] : 
                       (N2922)? data_o[663] : 
                       (N2924)? data_o[695] : 
                       (N2926)? data_o[727] : 
                       (N2928)? data_o[759] : 
                       (N2930)? data_o[791] : 
                       (N2932)? data_o[823] : 
                       (N2934)? data_o[855] : 
                       (N2936)? data_o[887] : 
                       (N2938)? data_o[919] : 
                       (N2940)? data_o[951] : 
                       (N2942)? data_o[983] : 
                       (N2944)? data_o[1015] : 
                       (N2946)? data_o[1047] : 
                       (N2948)? data_o[1079] : 
                       (N2950)? data_o[1111] : 
                       (N2952)? data_o[1143] : 
                       (N2954)? data_o[1175] : 
                       (N2956)? data_o[1207] : 
                       (N2958)? data_o[1239] : 
                       (N2960)? data_o[1271] : 
                       (N2962)? data_o[1303] : 
                       (N2964)? data_o[1335] : 
                       (N2966)? data_o[1367] : 
                       (N2968)? data_o[1399] : 
                       (N2970)? data_o[1431] : 
                       (N2972)? data_o[1463] : 
                       (N2974)? data_o[1495] : 
                       (N2976)? data_o[1527] : 
                       (N2978)? data_o[1559] : 
                       (N2980)? data_o[1591] : 
                       (N2982)? data_o[1623] : 
                       (N2984)? data_o[1655] : 
                       (N2986)? data_o[1687] : 
                       (N2988)? data_o[1719] : 
                       (N2990)? data_o[1751] : 
                       (N2992)? data_o[1783] : 
                       (N2994)? data_o[1815] : 
                       (N2996)? data_o[1847] : 
                       (N2998)? data_o[1879] : 
                       (N3000)? data_o[1911] : 
                       (N3002)? data_o[1943] : 
                       (N3004)? data_o[1975] : 
                       (N3006)? data_o[2007] : 
                       (N3008)? data_o[2039] : 
                       (N2883)? data_n_64__23_ : 
                       (N2885)? data_n_65__23_ : 
                       (N2887)? data_n_66__23_ : 
                       (N2889)? data_n_67__23_ : 
                       (N2891)? data_n_68__23_ : 
                       (N2893)? data_n_69__23_ : 
                       (N2895)? data_n_70__23_ : 
                       (N2897)? data_n_71__23_ : 
                       (N2899)? data_n_72__23_ : 
                       (N2901)? data_n_73__23_ : 
                       (N2903)? data_n_74__23_ : 
                       (N2905)? data_n_75__23_ : 
                       (N2907)? data_n_76__23_ : 
                       (N2909)? data_n_77__23_ : 
                       (N2911)? data_n_78__23_ : 
                       (N2913)? data_n_79__23_ : 
                       (N2915)? data_n_80__23_ : 
                       (N2917)? data_n_81__23_ : 
                       (N2919)? data_n_82__23_ : 
                       (N2921)? data_n_83__23_ : 
                       (N2923)? data_n_84__23_ : 
                       (N2925)? data_n_85__23_ : 
                       (N2927)? data_n_86__23_ : 
                       (N2929)? data_n_87__23_ : 
                       (N2931)? data_n_88__23_ : 
                       (N2933)? data_n_89__23_ : 
                       (N2935)? data_n_90__23_ : 
                       (N2937)? data_n_91__23_ : 
                       (N2939)? data_n_92__23_ : 
                       (N2941)? data_n_93__23_ : 
                       (N2943)? data_n_94__23_ : 
                       (N2945)? data_n_95__23_ : 
                       (N2947)? data_n_96__23_ : 
                       (N2949)? data_n_97__23_ : 
                       (N2951)? data_n_98__23_ : 
                       (N2953)? data_n_99__23_ : 
                       (N2955)? data_n_100__23_ : 
                       (N2957)? data_n_101__23_ : 
                       (N2959)? data_n_102__23_ : 
                       (N2961)? data_n_103__23_ : 
                       (N2963)? data_n_104__23_ : 
                       (N2965)? data_n_105__23_ : 
                       (N2967)? data_n_106__23_ : 
                       (N2969)? data_n_107__23_ : 
                       (N2971)? data_n_108__23_ : 
                       (N2973)? data_n_109__23_ : 
                       (N2975)? data_n_110__23_ : 
                       (N2977)? data_n_111__23_ : 
                       (N2979)? data_n_112__23_ : 
                       (N2981)? data_n_113__23_ : 
                       (N2983)? data_n_114__23_ : 
                       (N2985)? data_n_115__23_ : 
                       (N2987)? data_n_116__23_ : 
                       (N2989)? data_n_117__23_ : 
                       (N2991)? data_n_118__23_ : 
                       (N2993)? data_n_119__23_ : 
                       (N2995)? data_n_120__23_ : 
                       (N2997)? data_n_121__23_ : 
                       (N2999)? data_n_122__23_ : 
                       (N3001)? data_n_123__23_ : 
                       (N3003)? data_n_124__23_ : 
                       (N3005)? data_n_125__23_ : 
                       (N3007)? data_n_126__23_ : 
                       (N3009)? data_n_127__23_ : 1'b0;
  assign data_nn[22] = (N2882)? data_o[22] : 
                       (N2884)? data_o[54] : 
                       (N2886)? data_o[86] : 
                       (N2888)? data_o[118] : 
                       (N2890)? data_o[150] : 
                       (N2892)? data_o[182] : 
                       (N2894)? data_o[214] : 
                       (N2896)? data_o[246] : 
                       (N2898)? data_o[278] : 
                       (N2900)? data_o[310] : 
                       (N2902)? data_o[342] : 
                       (N2904)? data_o[374] : 
                       (N2906)? data_o[406] : 
                       (N2908)? data_o[438] : 
                       (N2910)? data_o[470] : 
                       (N2912)? data_o[502] : 
                       (N2914)? data_o[534] : 
                       (N2916)? data_o[566] : 
                       (N2918)? data_o[598] : 
                       (N2920)? data_o[630] : 
                       (N2922)? data_o[662] : 
                       (N2924)? data_o[694] : 
                       (N2926)? data_o[726] : 
                       (N2928)? data_o[758] : 
                       (N2930)? data_o[790] : 
                       (N2932)? data_o[822] : 
                       (N2934)? data_o[854] : 
                       (N2936)? data_o[886] : 
                       (N2938)? data_o[918] : 
                       (N2940)? data_o[950] : 
                       (N2942)? data_o[982] : 
                       (N2944)? data_o[1014] : 
                       (N2946)? data_o[1046] : 
                       (N2948)? data_o[1078] : 
                       (N2950)? data_o[1110] : 
                       (N2952)? data_o[1142] : 
                       (N2954)? data_o[1174] : 
                       (N2956)? data_o[1206] : 
                       (N2958)? data_o[1238] : 
                       (N2960)? data_o[1270] : 
                       (N2962)? data_o[1302] : 
                       (N2964)? data_o[1334] : 
                       (N2966)? data_o[1366] : 
                       (N2968)? data_o[1398] : 
                       (N2970)? data_o[1430] : 
                       (N2972)? data_o[1462] : 
                       (N2974)? data_o[1494] : 
                       (N2976)? data_o[1526] : 
                       (N2978)? data_o[1558] : 
                       (N2980)? data_o[1590] : 
                       (N2982)? data_o[1622] : 
                       (N2984)? data_o[1654] : 
                       (N2986)? data_o[1686] : 
                       (N2988)? data_o[1718] : 
                       (N2990)? data_o[1750] : 
                       (N2992)? data_o[1782] : 
                       (N2994)? data_o[1814] : 
                       (N2996)? data_o[1846] : 
                       (N2998)? data_o[1878] : 
                       (N3000)? data_o[1910] : 
                       (N3002)? data_o[1942] : 
                       (N3004)? data_o[1974] : 
                       (N3006)? data_o[2006] : 
                       (N3008)? data_o[2038] : 
                       (N2883)? data_n_64__22_ : 
                       (N2885)? data_n_65__22_ : 
                       (N2887)? data_n_66__22_ : 
                       (N2889)? data_n_67__22_ : 
                       (N2891)? data_n_68__22_ : 
                       (N2893)? data_n_69__22_ : 
                       (N2895)? data_n_70__22_ : 
                       (N2897)? data_n_71__22_ : 
                       (N2899)? data_n_72__22_ : 
                       (N2901)? data_n_73__22_ : 
                       (N2903)? data_n_74__22_ : 
                       (N2905)? data_n_75__22_ : 
                       (N2907)? data_n_76__22_ : 
                       (N2909)? data_n_77__22_ : 
                       (N2911)? data_n_78__22_ : 
                       (N2913)? data_n_79__22_ : 
                       (N2915)? data_n_80__22_ : 
                       (N2917)? data_n_81__22_ : 
                       (N2919)? data_n_82__22_ : 
                       (N2921)? data_n_83__22_ : 
                       (N2923)? data_n_84__22_ : 
                       (N2925)? data_n_85__22_ : 
                       (N2927)? data_n_86__22_ : 
                       (N2929)? data_n_87__22_ : 
                       (N2931)? data_n_88__22_ : 
                       (N2933)? data_n_89__22_ : 
                       (N2935)? data_n_90__22_ : 
                       (N2937)? data_n_91__22_ : 
                       (N2939)? data_n_92__22_ : 
                       (N2941)? data_n_93__22_ : 
                       (N2943)? data_n_94__22_ : 
                       (N2945)? data_n_95__22_ : 
                       (N2947)? data_n_96__22_ : 
                       (N2949)? data_n_97__22_ : 
                       (N2951)? data_n_98__22_ : 
                       (N2953)? data_n_99__22_ : 
                       (N2955)? data_n_100__22_ : 
                       (N2957)? data_n_101__22_ : 
                       (N2959)? data_n_102__22_ : 
                       (N2961)? data_n_103__22_ : 
                       (N2963)? data_n_104__22_ : 
                       (N2965)? data_n_105__22_ : 
                       (N2967)? data_n_106__22_ : 
                       (N2969)? data_n_107__22_ : 
                       (N2971)? data_n_108__22_ : 
                       (N2973)? data_n_109__22_ : 
                       (N2975)? data_n_110__22_ : 
                       (N2977)? data_n_111__22_ : 
                       (N2979)? data_n_112__22_ : 
                       (N2981)? data_n_113__22_ : 
                       (N2983)? data_n_114__22_ : 
                       (N2985)? data_n_115__22_ : 
                       (N2987)? data_n_116__22_ : 
                       (N2989)? data_n_117__22_ : 
                       (N2991)? data_n_118__22_ : 
                       (N2993)? data_n_119__22_ : 
                       (N2995)? data_n_120__22_ : 
                       (N2997)? data_n_121__22_ : 
                       (N2999)? data_n_122__22_ : 
                       (N3001)? data_n_123__22_ : 
                       (N3003)? data_n_124__22_ : 
                       (N3005)? data_n_125__22_ : 
                       (N3007)? data_n_126__22_ : 
                       (N3009)? data_n_127__22_ : 1'b0;
  assign data_nn[21] = (N2882)? data_o[21] : 
                       (N2884)? data_o[53] : 
                       (N2886)? data_o[85] : 
                       (N2888)? data_o[117] : 
                       (N2890)? data_o[149] : 
                       (N2892)? data_o[181] : 
                       (N2894)? data_o[213] : 
                       (N2896)? data_o[245] : 
                       (N2898)? data_o[277] : 
                       (N2900)? data_o[309] : 
                       (N2902)? data_o[341] : 
                       (N2904)? data_o[373] : 
                       (N2906)? data_o[405] : 
                       (N2908)? data_o[437] : 
                       (N2910)? data_o[469] : 
                       (N2912)? data_o[501] : 
                       (N2914)? data_o[533] : 
                       (N2916)? data_o[565] : 
                       (N2918)? data_o[597] : 
                       (N2920)? data_o[629] : 
                       (N2922)? data_o[661] : 
                       (N2924)? data_o[693] : 
                       (N2926)? data_o[725] : 
                       (N2928)? data_o[757] : 
                       (N2930)? data_o[789] : 
                       (N2932)? data_o[821] : 
                       (N2934)? data_o[853] : 
                       (N2936)? data_o[885] : 
                       (N2938)? data_o[917] : 
                       (N2940)? data_o[949] : 
                       (N2942)? data_o[981] : 
                       (N2944)? data_o[1013] : 
                       (N2946)? data_o[1045] : 
                       (N2948)? data_o[1077] : 
                       (N2950)? data_o[1109] : 
                       (N2952)? data_o[1141] : 
                       (N2954)? data_o[1173] : 
                       (N2956)? data_o[1205] : 
                       (N2958)? data_o[1237] : 
                       (N2960)? data_o[1269] : 
                       (N2962)? data_o[1301] : 
                       (N2964)? data_o[1333] : 
                       (N2966)? data_o[1365] : 
                       (N2968)? data_o[1397] : 
                       (N2970)? data_o[1429] : 
                       (N2972)? data_o[1461] : 
                       (N2974)? data_o[1493] : 
                       (N2976)? data_o[1525] : 
                       (N2978)? data_o[1557] : 
                       (N2980)? data_o[1589] : 
                       (N2982)? data_o[1621] : 
                       (N2984)? data_o[1653] : 
                       (N2986)? data_o[1685] : 
                       (N2988)? data_o[1717] : 
                       (N2990)? data_o[1749] : 
                       (N2992)? data_o[1781] : 
                       (N2994)? data_o[1813] : 
                       (N2996)? data_o[1845] : 
                       (N2998)? data_o[1877] : 
                       (N3000)? data_o[1909] : 
                       (N3002)? data_o[1941] : 
                       (N3004)? data_o[1973] : 
                       (N3006)? data_o[2005] : 
                       (N3008)? data_o[2037] : 
                       (N2883)? data_n_64__21_ : 
                       (N2885)? data_n_65__21_ : 
                       (N2887)? data_n_66__21_ : 
                       (N2889)? data_n_67__21_ : 
                       (N2891)? data_n_68__21_ : 
                       (N2893)? data_n_69__21_ : 
                       (N2895)? data_n_70__21_ : 
                       (N2897)? data_n_71__21_ : 
                       (N2899)? data_n_72__21_ : 
                       (N2901)? data_n_73__21_ : 
                       (N2903)? data_n_74__21_ : 
                       (N2905)? data_n_75__21_ : 
                       (N2907)? data_n_76__21_ : 
                       (N2909)? data_n_77__21_ : 
                       (N2911)? data_n_78__21_ : 
                       (N2913)? data_n_79__21_ : 
                       (N2915)? data_n_80__21_ : 
                       (N2917)? data_n_81__21_ : 
                       (N2919)? data_n_82__21_ : 
                       (N2921)? data_n_83__21_ : 
                       (N2923)? data_n_84__21_ : 
                       (N2925)? data_n_85__21_ : 
                       (N2927)? data_n_86__21_ : 
                       (N2929)? data_n_87__21_ : 
                       (N2931)? data_n_88__21_ : 
                       (N2933)? data_n_89__21_ : 
                       (N2935)? data_n_90__21_ : 
                       (N2937)? data_n_91__21_ : 
                       (N2939)? data_n_92__21_ : 
                       (N2941)? data_n_93__21_ : 
                       (N2943)? data_n_94__21_ : 
                       (N2945)? data_n_95__21_ : 
                       (N2947)? data_n_96__21_ : 
                       (N2949)? data_n_97__21_ : 
                       (N2951)? data_n_98__21_ : 
                       (N2953)? data_n_99__21_ : 
                       (N2955)? data_n_100__21_ : 
                       (N2957)? data_n_101__21_ : 
                       (N2959)? data_n_102__21_ : 
                       (N2961)? data_n_103__21_ : 
                       (N2963)? data_n_104__21_ : 
                       (N2965)? data_n_105__21_ : 
                       (N2967)? data_n_106__21_ : 
                       (N2969)? data_n_107__21_ : 
                       (N2971)? data_n_108__21_ : 
                       (N2973)? data_n_109__21_ : 
                       (N2975)? data_n_110__21_ : 
                       (N2977)? data_n_111__21_ : 
                       (N2979)? data_n_112__21_ : 
                       (N2981)? data_n_113__21_ : 
                       (N2983)? data_n_114__21_ : 
                       (N2985)? data_n_115__21_ : 
                       (N2987)? data_n_116__21_ : 
                       (N2989)? data_n_117__21_ : 
                       (N2991)? data_n_118__21_ : 
                       (N2993)? data_n_119__21_ : 
                       (N2995)? data_n_120__21_ : 
                       (N2997)? data_n_121__21_ : 
                       (N2999)? data_n_122__21_ : 
                       (N3001)? data_n_123__21_ : 
                       (N3003)? data_n_124__21_ : 
                       (N3005)? data_n_125__21_ : 
                       (N3007)? data_n_126__21_ : 
                       (N3009)? data_n_127__21_ : 1'b0;
  assign data_nn[20] = (N2882)? data_o[20] : 
                       (N2884)? data_o[52] : 
                       (N2886)? data_o[84] : 
                       (N2888)? data_o[116] : 
                       (N2890)? data_o[148] : 
                       (N2892)? data_o[180] : 
                       (N2894)? data_o[212] : 
                       (N2896)? data_o[244] : 
                       (N2898)? data_o[276] : 
                       (N2900)? data_o[308] : 
                       (N2902)? data_o[340] : 
                       (N2904)? data_o[372] : 
                       (N2906)? data_o[404] : 
                       (N2908)? data_o[436] : 
                       (N2910)? data_o[468] : 
                       (N2912)? data_o[500] : 
                       (N2914)? data_o[532] : 
                       (N2916)? data_o[564] : 
                       (N2918)? data_o[596] : 
                       (N2920)? data_o[628] : 
                       (N2922)? data_o[660] : 
                       (N2924)? data_o[692] : 
                       (N2926)? data_o[724] : 
                       (N2928)? data_o[756] : 
                       (N2930)? data_o[788] : 
                       (N2932)? data_o[820] : 
                       (N2934)? data_o[852] : 
                       (N2936)? data_o[884] : 
                       (N2938)? data_o[916] : 
                       (N2940)? data_o[948] : 
                       (N2942)? data_o[980] : 
                       (N2944)? data_o[1012] : 
                       (N2946)? data_o[1044] : 
                       (N2948)? data_o[1076] : 
                       (N2950)? data_o[1108] : 
                       (N2952)? data_o[1140] : 
                       (N2954)? data_o[1172] : 
                       (N2956)? data_o[1204] : 
                       (N2958)? data_o[1236] : 
                       (N2960)? data_o[1268] : 
                       (N2962)? data_o[1300] : 
                       (N2964)? data_o[1332] : 
                       (N2966)? data_o[1364] : 
                       (N2968)? data_o[1396] : 
                       (N2970)? data_o[1428] : 
                       (N2972)? data_o[1460] : 
                       (N2974)? data_o[1492] : 
                       (N2976)? data_o[1524] : 
                       (N2978)? data_o[1556] : 
                       (N2980)? data_o[1588] : 
                       (N2982)? data_o[1620] : 
                       (N2984)? data_o[1652] : 
                       (N2986)? data_o[1684] : 
                       (N2988)? data_o[1716] : 
                       (N2990)? data_o[1748] : 
                       (N2992)? data_o[1780] : 
                       (N2994)? data_o[1812] : 
                       (N2996)? data_o[1844] : 
                       (N2998)? data_o[1876] : 
                       (N3000)? data_o[1908] : 
                       (N3002)? data_o[1940] : 
                       (N3004)? data_o[1972] : 
                       (N3006)? data_o[2004] : 
                       (N3008)? data_o[2036] : 
                       (N2883)? data_n_64__20_ : 
                       (N2885)? data_n_65__20_ : 
                       (N2887)? data_n_66__20_ : 
                       (N2889)? data_n_67__20_ : 
                       (N2891)? data_n_68__20_ : 
                       (N2893)? data_n_69__20_ : 
                       (N2895)? data_n_70__20_ : 
                       (N2897)? data_n_71__20_ : 
                       (N2899)? data_n_72__20_ : 
                       (N2901)? data_n_73__20_ : 
                       (N2903)? data_n_74__20_ : 
                       (N2905)? data_n_75__20_ : 
                       (N2907)? data_n_76__20_ : 
                       (N2909)? data_n_77__20_ : 
                       (N2911)? data_n_78__20_ : 
                       (N2913)? data_n_79__20_ : 
                       (N2915)? data_n_80__20_ : 
                       (N2917)? data_n_81__20_ : 
                       (N2919)? data_n_82__20_ : 
                       (N2921)? data_n_83__20_ : 
                       (N2923)? data_n_84__20_ : 
                       (N2925)? data_n_85__20_ : 
                       (N2927)? data_n_86__20_ : 
                       (N2929)? data_n_87__20_ : 
                       (N2931)? data_n_88__20_ : 
                       (N2933)? data_n_89__20_ : 
                       (N2935)? data_n_90__20_ : 
                       (N2937)? data_n_91__20_ : 
                       (N2939)? data_n_92__20_ : 
                       (N2941)? data_n_93__20_ : 
                       (N2943)? data_n_94__20_ : 
                       (N2945)? data_n_95__20_ : 
                       (N2947)? data_n_96__20_ : 
                       (N2949)? data_n_97__20_ : 
                       (N2951)? data_n_98__20_ : 
                       (N2953)? data_n_99__20_ : 
                       (N2955)? data_n_100__20_ : 
                       (N2957)? data_n_101__20_ : 
                       (N2959)? data_n_102__20_ : 
                       (N2961)? data_n_103__20_ : 
                       (N2963)? data_n_104__20_ : 
                       (N2965)? data_n_105__20_ : 
                       (N2967)? data_n_106__20_ : 
                       (N2969)? data_n_107__20_ : 
                       (N2971)? data_n_108__20_ : 
                       (N2973)? data_n_109__20_ : 
                       (N2975)? data_n_110__20_ : 
                       (N2977)? data_n_111__20_ : 
                       (N2979)? data_n_112__20_ : 
                       (N2981)? data_n_113__20_ : 
                       (N2983)? data_n_114__20_ : 
                       (N2985)? data_n_115__20_ : 
                       (N2987)? data_n_116__20_ : 
                       (N2989)? data_n_117__20_ : 
                       (N2991)? data_n_118__20_ : 
                       (N2993)? data_n_119__20_ : 
                       (N2995)? data_n_120__20_ : 
                       (N2997)? data_n_121__20_ : 
                       (N2999)? data_n_122__20_ : 
                       (N3001)? data_n_123__20_ : 
                       (N3003)? data_n_124__20_ : 
                       (N3005)? data_n_125__20_ : 
                       (N3007)? data_n_126__20_ : 
                       (N3009)? data_n_127__20_ : 1'b0;
  assign data_nn[19] = (N2882)? data_o[19] : 
                       (N2884)? data_o[51] : 
                       (N2886)? data_o[83] : 
                       (N2888)? data_o[115] : 
                       (N2890)? data_o[147] : 
                       (N2892)? data_o[179] : 
                       (N2894)? data_o[211] : 
                       (N2896)? data_o[243] : 
                       (N2898)? data_o[275] : 
                       (N2900)? data_o[307] : 
                       (N2902)? data_o[339] : 
                       (N2904)? data_o[371] : 
                       (N2906)? data_o[403] : 
                       (N2908)? data_o[435] : 
                       (N2910)? data_o[467] : 
                       (N2912)? data_o[499] : 
                       (N2914)? data_o[531] : 
                       (N2916)? data_o[563] : 
                       (N2918)? data_o[595] : 
                       (N2920)? data_o[627] : 
                       (N2922)? data_o[659] : 
                       (N2924)? data_o[691] : 
                       (N2926)? data_o[723] : 
                       (N2928)? data_o[755] : 
                       (N2930)? data_o[787] : 
                       (N2932)? data_o[819] : 
                       (N2934)? data_o[851] : 
                       (N2936)? data_o[883] : 
                       (N2938)? data_o[915] : 
                       (N2940)? data_o[947] : 
                       (N2942)? data_o[979] : 
                       (N2944)? data_o[1011] : 
                       (N2946)? data_o[1043] : 
                       (N2948)? data_o[1075] : 
                       (N2950)? data_o[1107] : 
                       (N2952)? data_o[1139] : 
                       (N2954)? data_o[1171] : 
                       (N2956)? data_o[1203] : 
                       (N2958)? data_o[1235] : 
                       (N2960)? data_o[1267] : 
                       (N2962)? data_o[1299] : 
                       (N2964)? data_o[1331] : 
                       (N2966)? data_o[1363] : 
                       (N2968)? data_o[1395] : 
                       (N2970)? data_o[1427] : 
                       (N2972)? data_o[1459] : 
                       (N2974)? data_o[1491] : 
                       (N2976)? data_o[1523] : 
                       (N2978)? data_o[1555] : 
                       (N2980)? data_o[1587] : 
                       (N2982)? data_o[1619] : 
                       (N2984)? data_o[1651] : 
                       (N2986)? data_o[1683] : 
                       (N2988)? data_o[1715] : 
                       (N2990)? data_o[1747] : 
                       (N2992)? data_o[1779] : 
                       (N2994)? data_o[1811] : 
                       (N2996)? data_o[1843] : 
                       (N2998)? data_o[1875] : 
                       (N3000)? data_o[1907] : 
                       (N3002)? data_o[1939] : 
                       (N3004)? data_o[1971] : 
                       (N3006)? data_o[2003] : 
                       (N3008)? data_o[2035] : 
                       (N2883)? data_n_64__19_ : 
                       (N2885)? data_n_65__19_ : 
                       (N2887)? data_n_66__19_ : 
                       (N2889)? data_n_67__19_ : 
                       (N2891)? data_n_68__19_ : 
                       (N2893)? data_n_69__19_ : 
                       (N2895)? data_n_70__19_ : 
                       (N2897)? data_n_71__19_ : 
                       (N2899)? data_n_72__19_ : 
                       (N2901)? data_n_73__19_ : 
                       (N2903)? data_n_74__19_ : 
                       (N2905)? data_n_75__19_ : 
                       (N2907)? data_n_76__19_ : 
                       (N2909)? data_n_77__19_ : 
                       (N2911)? data_n_78__19_ : 
                       (N2913)? data_n_79__19_ : 
                       (N2915)? data_n_80__19_ : 
                       (N2917)? data_n_81__19_ : 
                       (N2919)? data_n_82__19_ : 
                       (N2921)? data_n_83__19_ : 
                       (N2923)? data_n_84__19_ : 
                       (N2925)? data_n_85__19_ : 
                       (N2927)? data_n_86__19_ : 
                       (N2929)? data_n_87__19_ : 
                       (N2931)? data_n_88__19_ : 
                       (N2933)? data_n_89__19_ : 
                       (N2935)? data_n_90__19_ : 
                       (N2937)? data_n_91__19_ : 
                       (N2939)? data_n_92__19_ : 
                       (N2941)? data_n_93__19_ : 
                       (N2943)? data_n_94__19_ : 
                       (N2945)? data_n_95__19_ : 
                       (N2947)? data_n_96__19_ : 
                       (N2949)? data_n_97__19_ : 
                       (N2951)? data_n_98__19_ : 
                       (N2953)? data_n_99__19_ : 
                       (N2955)? data_n_100__19_ : 
                       (N2957)? data_n_101__19_ : 
                       (N2959)? data_n_102__19_ : 
                       (N2961)? data_n_103__19_ : 
                       (N2963)? data_n_104__19_ : 
                       (N2965)? data_n_105__19_ : 
                       (N2967)? data_n_106__19_ : 
                       (N2969)? data_n_107__19_ : 
                       (N2971)? data_n_108__19_ : 
                       (N2973)? data_n_109__19_ : 
                       (N2975)? data_n_110__19_ : 
                       (N2977)? data_n_111__19_ : 
                       (N2979)? data_n_112__19_ : 
                       (N2981)? data_n_113__19_ : 
                       (N2983)? data_n_114__19_ : 
                       (N2985)? data_n_115__19_ : 
                       (N2987)? data_n_116__19_ : 
                       (N2989)? data_n_117__19_ : 
                       (N2991)? data_n_118__19_ : 
                       (N2993)? data_n_119__19_ : 
                       (N2995)? data_n_120__19_ : 
                       (N2997)? data_n_121__19_ : 
                       (N2999)? data_n_122__19_ : 
                       (N3001)? data_n_123__19_ : 
                       (N3003)? data_n_124__19_ : 
                       (N3005)? data_n_125__19_ : 
                       (N3007)? data_n_126__19_ : 
                       (N3009)? data_n_127__19_ : 1'b0;
  assign data_nn[18] = (N2882)? data_o[18] : 
                       (N2884)? data_o[50] : 
                       (N2886)? data_o[82] : 
                       (N2888)? data_o[114] : 
                       (N2890)? data_o[146] : 
                       (N2892)? data_o[178] : 
                       (N2894)? data_o[210] : 
                       (N2896)? data_o[242] : 
                       (N2898)? data_o[274] : 
                       (N2900)? data_o[306] : 
                       (N2902)? data_o[338] : 
                       (N2904)? data_o[370] : 
                       (N2906)? data_o[402] : 
                       (N2908)? data_o[434] : 
                       (N2910)? data_o[466] : 
                       (N2912)? data_o[498] : 
                       (N2914)? data_o[530] : 
                       (N2916)? data_o[562] : 
                       (N2918)? data_o[594] : 
                       (N2920)? data_o[626] : 
                       (N2922)? data_o[658] : 
                       (N2924)? data_o[690] : 
                       (N2926)? data_o[722] : 
                       (N2928)? data_o[754] : 
                       (N2930)? data_o[786] : 
                       (N2932)? data_o[818] : 
                       (N2934)? data_o[850] : 
                       (N2936)? data_o[882] : 
                       (N2938)? data_o[914] : 
                       (N2940)? data_o[946] : 
                       (N2942)? data_o[978] : 
                       (N2944)? data_o[1010] : 
                       (N2946)? data_o[1042] : 
                       (N2948)? data_o[1074] : 
                       (N2950)? data_o[1106] : 
                       (N2952)? data_o[1138] : 
                       (N2954)? data_o[1170] : 
                       (N2956)? data_o[1202] : 
                       (N2958)? data_o[1234] : 
                       (N2960)? data_o[1266] : 
                       (N2962)? data_o[1298] : 
                       (N2964)? data_o[1330] : 
                       (N2966)? data_o[1362] : 
                       (N2968)? data_o[1394] : 
                       (N2970)? data_o[1426] : 
                       (N2972)? data_o[1458] : 
                       (N2974)? data_o[1490] : 
                       (N2976)? data_o[1522] : 
                       (N2978)? data_o[1554] : 
                       (N2980)? data_o[1586] : 
                       (N2982)? data_o[1618] : 
                       (N2984)? data_o[1650] : 
                       (N2986)? data_o[1682] : 
                       (N2988)? data_o[1714] : 
                       (N2990)? data_o[1746] : 
                       (N2992)? data_o[1778] : 
                       (N2994)? data_o[1810] : 
                       (N2996)? data_o[1842] : 
                       (N2998)? data_o[1874] : 
                       (N3000)? data_o[1906] : 
                       (N3002)? data_o[1938] : 
                       (N3004)? data_o[1970] : 
                       (N3006)? data_o[2002] : 
                       (N3008)? data_o[2034] : 
                       (N2883)? data_n_64__18_ : 
                       (N2885)? data_n_65__18_ : 
                       (N2887)? data_n_66__18_ : 
                       (N2889)? data_n_67__18_ : 
                       (N2891)? data_n_68__18_ : 
                       (N2893)? data_n_69__18_ : 
                       (N2895)? data_n_70__18_ : 
                       (N2897)? data_n_71__18_ : 
                       (N2899)? data_n_72__18_ : 
                       (N2901)? data_n_73__18_ : 
                       (N2903)? data_n_74__18_ : 
                       (N2905)? data_n_75__18_ : 
                       (N2907)? data_n_76__18_ : 
                       (N2909)? data_n_77__18_ : 
                       (N2911)? data_n_78__18_ : 
                       (N2913)? data_n_79__18_ : 
                       (N2915)? data_n_80__18_ : 
                       (N2917)? data_n_81__18_ : 
                       (N2919)? data_n_82__18_ : 
                       (N2921)? data_n_83__18_ : 
                       (N2923)? data_n_84__18_ : 
                       (N2925)? data_n_85__18_ : 
                       (N2927)? data_n_86__18_ : 
                       (N2929)? data_n_87__18_ : 
                       (N2931)? data_n_88__18_ : 
                       (N2933)? data_n_89__18_ : 
                       (N2935)? data_n_90__18_ : 
                       (N2937)? data_n_91__18_ : 
                       (N2939)? data_n_92__18_ : 
                       (N2941)? data_n_93__18_ : 
                       (N2943)? data_n_94__18_ : 
                       (N2945)? data_n_95__18_ : 
                       (N2947)? data_n_96__18_ : 
                       (N2949)? data_n_97__18_ : 
                       (N2951)? data_n_98__18_ : 
                       (N2953)? data_n_99__18_ : 
                       (N2955)? data_n_100__18_ : 
                       (N2957)? data_n_101__18_ : 
                       (N2959)? data_n_102__18_ : 
                       (N2961)? data_n_103__18_ : 
                       (N2963)? data_n_104__18_ : 
                       (N2965)? data_n_105__18_ : 
                       (N2967)? data_n_106__18_ : 
                       (N2969)? data_n_107__18_ : 
                       (N2971)? data_n_108__18_ : 
                       (N2973)? data_n_109__18_ : 
                       (N2975)? data_n_110__18_ : 
                       (N2977)? data_n_111__18_ : 
                       (N2979)? data_n_112__18_ : 
                       (N2981)? data_n_113__18_ : 
                       (N2983)? data_n_114__18_ : 
                       (N2985)? data_n_115__18_ : 
                       (N2987)? data_n_116__18_ : 
                       (N2989)? data_n_117__18_ : 
                       (N2991)? data_n_118__18_ : 
                       (N2993)? data_n_119__18_ : 
                       (N2995)? data_n_120__18_ : 
                       (N2997)? data_n_121__18_ : 
                       (N2999)? data_n_122__18_ : 
                       (N3001)? data_n_123__18_ : 
                       (N3003)? data_n_124__18_ : 
                       (N3005)? data_n_125__18_ : 
                       (N3007)? data_n_126__18_ : 
                       (N3009)? data_n_127__18_ : 1'b0;
  assign data_nn[17] = (N2882)? data_o[17] : 
                       (N2884)? data_o[49] : 
                       (N2886)? data_o[81] : 
                       (N2888)? data_o[113] : 
                       (N2890)? data_o[145] : 
                       (N2892)? data_o[177] : 
                       (N2894)? data_o[209] : 
                       (N2896)? data_o[241] : 
                       (N2898)? data_o[273] : 
                       (N2900)? data_o[305] : 
                       (N2902)? data_o[337] : 
                       (N2904)? data_o[369] : 
                       (N2906)? data_o[401] : 
                       (N2908)? data_o[433] : 
                       (N2910)? data_o[465] : 
                       (N2912)? data_o[497] : 
                       (N2914)? data_o[529] : 
                       (N2916)? data_o[561] : 
                       (N2918)? data_o[593] : 
                       (N2920)? data_o[625] : 
                       (N2922)? data_o[657] : 
                       (N2924)? data_o[689] : 
                       (N2926)? data_o[721] : 
                       (N2928)? data_o[753] : 
                       (N2930)? data_o[785] : 
                       (N2932)? data_o[817] : 
                       (N2934)? data_o[849] : 
                       (N2936)? data_o[881] : 
                       (N2938)? data_o[913] : 
                       (N2940)? data_o[945] : 
                       (N2942)? data_o[977] : 
                       (N2944)? data_o[1009] : 
                       (N2946)? data_o[1041] : 
                       (N2948)? data_o[1073] : 
                       (N2950)? data_o[1105] : 
                       (N2952)? data_o[1137] : 
                       (N2954)? data_o[1169] : 
                       (N2956)? data_o[1201] : 
                       (N2958)? data_o[1233] : 
                       (N2960)? data_o[1265] : 
                       (N2962)? data_o[1297] : 
                       (N2964)? data_o[1329] : 
                       (N2966)? data_o[1361] : 
                       (N2968)? data_o[1393] : 
                       (N2970)? data_o[1425] : 
                       (N2972)? data_o[1457] : 
                       (N2974)? data_o[1489] : 
                       (N2976)? data_o[1521] : 
                       (N2978)? data_o[1553] : 
                       (N2980)? data_o[1585] : 
                       (N2982)? data_o[1617] : 
                       (N2984)? data_o[1649] : 
                       (N2986)? data_o[1681] : 
                       (N2988)? data_o[1713] : 
                       (N2990)? data_o[1745] : 
                       (N2992)? data_o[1777] : 
                       (N2994)? data_o[1809] : 
                       (N2996)? data_o[1841] : 
                       (N2998)? data_o[1873] : 
                       (N3000)? data_o[1905] : 
                       (N3002)? data_o[1937] : 
                       (N3004)? data_o[1969] : 
                       (N3006)? data_o[2001] : 
                       (N3008)? data_o[2033] : 
                       (N2883)? data_n_64__17_ : 
                       (N2885)? data_n_65__17_ : 
                       (N2887)? data_n_66__17_ : 
                       (N2889)? data_n_67__17_ : 
                       (N2891)? data_n_68__17_ : 
                       (N2893)? data_n_69__17_ : 
                       (N2895)? data_n_70__17_ : 
                       (N2897)? data_n_71__17_ : 
                       (N2899)? data_n_72__17_ : 
                       (N2901)? data_n_73__17_ : 
                       (N2903)? data_n_74__17_ : 
                       (N2905)? data_n_75__17_ : 
                       (N2907)? data_n_76__17_ : 
                       (N2909)? data_n_77__17_ : 
                       (N2911)? data_n_78__17_ : 
                       (N2913)? data_n_79__17_ : 
                       (N2915)? data_n_80__17_ : 
                       (N2917)? data_n_81__17_ : 
                       (N2919)? data_n_82__17_ : 
                       (N2921)? data_n_83__17_ : 
                       (N2923)? data_n_84__17_ : 
                       (N2925)? data_n_85__17_ : 
                       (N2927)? data_n_86__17_ : 
                       (N2929)? data_n_87__17_ : 
                       (N2931)? data_n_88__17_ : 
                       (N2933)? data_n_89__17_ : 
                       (N2935)? data_n_90__17_ : 
                       (N2937)? data_n_91__17_ : 
                       (N2939)? data_n_92__17_ : 
                       (N2941)? data_n_93__17_ : 
                       (N2943)? data_n_94__17_ : 
                       (N2945)? data_n_95__17_ : 
                       (N2947)? data_n_96__17_ : 
                       (N2949)? data_n_97__17_ : 
                       (N2951)? data_n_98__17_ : 
                       (N2953)? data_n_99__17_ : 
                       (N2955)? data_n_100__17_ : 
                       (N2957)? data_n_101__17_ : 
                       (N2959)? data_n_102__17_ : 
                       (N2961)? data_n_103__17_ : 
                       (N2963)? data_n_104__17_ : 
                       (N2965)? data_n_105__17_ : 
                       (N2967)? data_n_106__17_ : 
                       (N2969)? data_n_107__17_ : 
                       (N2971)? data_n_108__17_ : 
                       (N2973)? data_n_109__17_ : 
                       (N2975)? data_n_110__17_ : 
                       (N2977)? data_n_111__17_ : 
                       (N2979)? data_n_112__17_ : 
                       (N2981)? data_n_113__17_ : 
                       (N2983)? data_n_114__17_ : 
                       (N2985)? data_n_115__17_ : 
                       (N2987)? data_n_116__17_ : 
                       (N2989)? data_n_117__17_ : 
                       (N2991)? data_n_118__17_ : 
                       (N2993)? data_n_119__17_ : 
                       (N2995)? data_n_120__17_ : 
                       (N2997)? data_n_121__17_ : 
                       (N2999)? data_n_122__17_ : 
                       (N3001)? data_n_123__17_ : 
                       (N3003)? data_n_124__17_ : 
                       (N3005)? data_n_125__17_ : 
                       (N3007)? data_n_126__17_ : 
                       (N3009)? data_n_127__17_ : 1'b0;
  assign data_nn[16] = (N2882)? data_o[16] : 
                       (N2884)? data_o[48] : 
                       (N2886)? data_o[80] : 
                       (N2888)? data_o[112] : 
                       (N2890)? data_o[144] : 
                       (N2892)? data_o[176] : 
                       (N2894)? data_o[208] : 
                       (N2896)? data_o[240] : 
                       (N2898)? data_o[272] : 
                       (N2900)? data_o[304] : 
                       (N2902)? data_o[336] : 
                       (N2904)? data_o[368] : 
                       (N2906)? data_o[400] : 
                       (N2908)? data_o[432] : 
                       (N2910)? data_o[464] : 
                       (N2912)? data_o[496] : 
                       (N2914)? data_o[528] : 
                       (N2916)? data_o[560] : 
                       (N2918)? data_o[592] : 
                       (N2920)? data_o[624] : 
                       (N2922)? data_o[656] : 
                       (N2924)? data_o[688] : 
                       (N2926)? data_o[720] : 
                       (N2928)? data_o[752] : 
                       (N2930)? data_o[784] : 
                       (N2932)? data_o[816] : 
                       (N2934)? data_o[848] : 
                       (N2936)? data_o[880] : 
                       (N2938)? data_o[912] : 
                       (N2940)? data_o[944] : 
                       (N2942)? data_o[976] : 
                       (N2944)? data_o[1008] : 
                       (N2946)? data_o[1040] : 
                       (N2948)? data_o[1072] : 
                       (N2950)? data_o[1104] : 
                       (N2952)? data_o[1136] : 
                       (N2954)? data_o[1168] : 
                       (N2956)? data_o[1200] : 
                       (N2958)? data_o[1232] : 
                       (N2960)? data_o[1264] : 
                       (N2962)? data_o[1296] : 
                       (N2964)? data_o[1328] : 
                       (N2966)? data_o[1360] : 
                       (N2968)? data_o[1392] : 
                       (N2970)? data_o[1424] : 
                       (N2972)? data_o[1456] : 
                       (N2974)? data_o[1488] : 
                       (N2976)? data_o[1520] : 
                       (N2978)? data_o[1552] : 
                       (N2980)? data_o[1584] : 
                       (N2982)? data_o[1616] : 
                       (N2984)? data_o[1648] : 
                       (N2986)? data_o[1680] : 
                       (N2988)? data_o[1712] : 
                       (N2990)? data_o[1744] : 
                       (N2992)? data_o[1776] : 
                       (N2994)? data_o[1808] : 
                       (N2996)? data_o[1840] : 
                       (N2998)? data_o[1872] : 
                       (N3000)? data_o[1904] : 
                       (N3002)? data_o[1936] : 
                       (N3004)? data_o[1968] : 
                       (N3006)? data_o[2000] : 
                       (N3008)? data_o[2032] : 
                       (N2883)? data_n_64__16_ : 
                       (N2885)? data_n_65__16_ : 
                       (N2887)? data_n_66__16_ : 
                       (N2889)? data_n_67__16_ : 
                       (N2891)? data_n_68__16_ : 
                       (N2893)? data_n_69__16_ : 
                       (N2895)? data_n_70__16_ : 
                       (N2897)? data_n_71__16_ : 
                       (N2899)? data_n_72__16_ : 
                       (N2901)? data_n_73__16_ : 
                       (N2903)? data_n_74__16_ : 
                       (N2905)? data_n_75__16_ : 
                       (N2907)? data_n_76__16_ : 
                       (N2909)? data_n_77__16_ : 
                       (N2911)? data_n_78__16_ : 
                       (N2913)? data_n_79__16_ : 
                       (N2915)? data_n_80__16_ : 
                       (N2917)? data_n_81__16_ : 
                       (N2919)? data_n_82__16_ : 
                       (N2921)? data_n_83__16_ : 
                       (N2923)? data_n_84__16_ : 
                       (N2925)? data_n_85__16_ : 
                       (N2927)? data_n_86__16_ : 
                       (N2929)? data_n_87__16_ : 
                       (N2931)? data_n_88__16_ : 
                       (N2933)? data_n_89__16_ : 
                       (N2935)? data_n_90__16_ : 
                       (N2937)? data_n_91__16_ : 
                       (N2939)? data_n_92__16_ : 
                       (N2941)? data_n_93__16_ : 
                       (N2943)? data_n_94__16_ : 
                       (N2945)? data_n_95__16_ : 
                       (N2947)? data_n_96__16_ : 
                       (N2949)? data_n_97__16_ : 
                       (N2951)? data_n_98__16_ : 
                       (N2953)? data_n_99__16_ : 
                       (N2955)? data_n_100__16_ : 
                       (N2957)? data_n_101__16_ : 
                       (N2959)? data_n_102__16_ : 
                       (N2961)? data_n_103__16_ : 
                       (N2963)? data_n_104__16_ : 
                       (N2965)? data_n_105__16_ : 
                       (N2967)? data_n_106__16_ : 
                       (N2969)? data_n_107__16_ : 
                       (N2971)? data_n_108__16_ : 
                       (N2973)? data_n_109__16_ : 
                       (N2975)? data_n_110__16_ : 
                       (N2977)? data_n_111__16_ : 
                       (N2979)? data_n_112__16_ : 
                       (N2981)? data_n_113__16_ : 
                       (N2983)? data_n_114__16_ : 
                       (N2985)? data_n_115__16_ : 
                       (N2987)? data_n_116__16_ : 
                       (N2989)? data_n_117__16_ : 
                       (N2991)? data_n_118__16_ : 
                       (N2993)? data_n_119__16_ : 
                       (N2995)? data_n_120__16_ : 
                       (N2997)? data_n_121__16_ : 
                       (N2999)? data_n_122__16_ : 
                       (N3001)? data_n_123__16_ : 
                       (N3003)? data_n_124__16_ : 
                       (N3005)? data_n_125__16_ : 
                       (N3007)? data_n_126__16_ : 
                       (N3009)? data_n_127__16_ : 1'b0;
  assign data_nn[15] = (N2882)? data_o[15] : 
                       (N2884)? data_o[47] : 
                       (N2886)? data_o[79] : 
                       (N2888)? data_o[111] : 
                       (N2890)? data_o[143] : 
                       (N2892)? data_o[175] : 
                       (N2894)? data_o[207] : 
                       (N2896)? data_o[239] : 
                       (N2898)? data_o[271] : 
                       (N2900)? data_o[303] : 
                       (N2902)? data_o[335] : 
                       (N2904)? data_o[367] : 
                       (N2906)? data_o[399] : 
                       (N2908)? data_o[431] : 
                       (N2910)? data_o[463] : 
                       (N2912)? data_o[495] : 
                       (N2914)? data_o[527] : 
                       (N2916)? data_o[559] : 
                       (N2918)? data_o[591] : 
                       (N2920)? data_o[623] : 
                       (N2922)? data_o[655] : 
                       (N2924)? data_o[687] : 
                       (N2926)? data_o[719] : 
                       (N2928)? data_o[751] : 
                       (N2930)? data_o[783] : 
                       (N2932)? data_o[815] : 
                       (N2934)? data_o[847] : 
                       (N2936)? data_o[879] : 
                       (N2938)? data_o[911] : 
                       (N2940)? data_o[943] : 
                       (N2942)? data_o[975] : 
                       (N2944)? data_o[1007] : 
                       (N2946)? data_o[1039] : 
                       (N2948)? data_o[1071] : 
                       (N2950)? data_o[1103] : 
                       (N2952)? data_o[1135] : 
                       (N2954)? data_o[1167] : 
                       (N2956)? data_o[1199] : 
                       (N2958)? data_o[1231] : 
                       (N2960)? data_o[1263] : 
                       (N2962)? data_o[1295] : 
                       (N2964)? data_o[1327] : 
                       (N2966)? data_o[1359] : 
                       (N2968)? data_o[1391] : 
                       (N2970)? data_o[1423] : 
                       (N2972)? data_o[1455] : 
                       (N2974)? data_o[1487] : 
                       (N2976)? data_o[1519] : 
                       (N2978)? data_o[1551] : 
                       (N2980)? data_o[1583] : 
                       (N2982)? data_o[1615] : 
                       (N2984)? data_o[1647] : 
                       (N2986)? data_o[1679] : 
                       (N2988)? data_o[1711] : 
                       (N2990)? data_o[1743] : 
                       (N2992)? data_o[1775] : 
                       (N2994)? data_o[1807] : 
                       (N2996)? data_o[1839] : 
                       (N2998)? data_o[1871] : 
                       (N3000)? data_o[1903] : 
                       (N3002)? data_o[1935] : 
                       (N3004)? data_o[1967] : 
                       (N3006)? data_o[1999] : 
                       (N3008)? data_o[2031] : 
                       (N2883)? data_n_64__15_ : 
                       (N2885)? data_n_65__15_ : 
                       (N2887)? data_n_66__15_ : 
                       (N2889)? data_n_67__15_ : 
                       (N2891)? data_n_68__15_ : 
                       (N2893)? data_n_69__15_ : 
                       (N2895)? data_n_70__15_ : 
                       (N2897)? data_n_71__15_ : 
                       (N2899)? data_n_72__15_ : 
                       (N2901)? data_n_73__15_ : 
                       (N2903)? data_n_74__15_ : 
                       (N2905)? data_n_75__15_ : 
                       (N2907)? data_n_76__15_ : 
                       (N2909)? data_n_77__15_ : 
                       (N2911)? data_n_78__15_ : 
                       (N2913)? data_n_79__15_ : 
                       (N2915)? data_n_80__15_ : 
                       (N2917)? data_n_81__15_ : 
                       (N2919)? data_n_82__15_ : 
                       (N2921)? data_n_83__15_ : 
                       (N2923)? data_n_84__15_ : 
                       (N2925)? data_n_85__15_ : 
                       (N2927)? data_n_86__15_ : 
                       (N2929)? data_n_87__15_ : 
                       (N2931)? data_n_88__15_ : 
                       (N2933)? data_n_89__15_ : 
                       (N2935)? data_n_90__15_ : 
                       (N2937)? data_n_91__15_ : 
                       (N2939)? data_n_92__15_ : 
                       (N2941)? data_n_93__15_ : 
                       (N2943)? data_n_94__15_ : 
                       (N2945)? data_n_95__15_ : 
                       (N2947)? data_n_96__15_ : 
                       (N2949)? data_n_97__15_ : 
                       (N2951)? data_n_98__15_ : 
                       (N2953)? data_n_99__15_ : 
                       (N2955)? data_n_100__15_ : 
                       (N2957)? data_n_101__15_ : 
                       (N2959)? data_n_102__15_ : 
                       (N2961)? data_n_103__15_ : 
                       (N2963)? data_n_104__15_ : 
                       (N2965)? data_n_105__15_ : 
                       (N2967)? data_n_106__15_ : 
                       (N2969)? data_n_107__15_ : 
                       (N2971)? data_n_108__15_ : 
                       (N2973)? data_n_109__15_ : 
                       (N2975)? data_n_110__15_ : 
                       (N2977)? data_n_111__15_ : 
                       (N2979)? data_n_112__15_ : 
                       (N2981)? data_n_113__15_ : 
                       (N2983)? data_n_114__15_ : 
                       (N2985)? data_n_115__15_ : 
                       (N2987)? data_n_116__15_ : 
                       (N2989)? data_n_117__15_ : 
                       (N2991)? data_n_118__15_ : 
                       (N2993)? data_n_119__15_ : 
                       (N2995)? data_n_120__15_ : 
                       (N2997)? data_n_121__15_ : 
                       (N2999)? data_n_122__15_ : 
                       (N3001)? data_n_123__15_ : 
                       (N3003)? data_n_124__15_ : 
                       (N3005)? data_n_125__15_ : 
                       (N3007)? data_n_126__15_ : 
                       (N3009)? data_n_127__15_ : 1'b0;
  assign data_nn[14] = (N2882)? data_o[14] : 
                       (N2884)? data_o[46] : 
                       (N2886)? data_o[78] : 
                       (N2888)? data_o[110] : 
                       (N2890)? data_o[142] : 
                       (N2892)? data_o[174] : 
                       (N2894)? data_o[206] : 
                       (N2896)? data_o[238] : 
                       (N2898)? data_o[270] : 
                       (N2900)? data_o[302] : 
                       (N2902)? data_o[334] : 
                       (N2904)? data_o[366] : 
                       (N2906)? data_o[398] : 
                       (N2908)? data_o[430] : 
                       (N2910)? data_o[462] : 
                       (N2912)? data_o[494] : 
                       (N2914)? data_o[526] : 
                       (N2916)? data_o[558] : 
                       (N2918)? data_o[590] : 
                       (N2920)? data_o[622] : 
                       (N2922)? data_o[654] : 
                       (N2924)? data_o[686] : 
                       (N2926)? data_o[718] : 
                       (N2928)? data_o[750] : 
                       (N2930)? data_o[782] : 
                       (N2932)? data_o[814] : 
                       (N2934)? data_o[846] : 
                       (N2936)? data_o[878] : 
                       (N2938)? data_o[910] : 
                       (N2940)? data_o[942] : 
                       (N2942)? data_o[974] : 
                       (N2944)? data_o[1006] : 
                       (N2946)? data_o[1038] : 
                       (N2948)? data_o[1070] : 
                       (N2950)? data_o[1102] : 
                       (N2952)? data_o[1134] : 
                       (N2954)? data_o[1166] : 
                       (N2956)? data_o[1198] : 
                       (N2958)? data_o[1230] : 
                       (N2960)? data_o[1262] : 
                       (N2962)? data_o[1294] : 
                       (N2964)? data_o[1326] : 
                       (N2966)? data_o[1358] : 
                       (N2968)? data_o[1390] : 
                       (N2970)? data_o[1422] : 
                       (N2972)? data_o[1454] : 
                       (N2974)? data_o[1486] : 
                       (N2976)? data_o[1518] : 
                       (N2978)? data_o[1550] : 
                       (N2980)? data_o[1582] : 
                       (N2982)? data_o[1614] : 
                       (N2984)? data_o[1646] : 
                       (N2986)? data_o[1678] : 
                       (N2988)? data_o[1710] : 
                       (N2990)? data_o[1742] : 
                       (N2992)? data_o[1774] : 
                       (N2994)? data_o[1806] : 
                       (N2996)? data_o[1838] : 
                       (N2998)? data_o[1870] : 
                       (N3000)? data_o[1902] : 
                       (N3002)? data_o[1934] : 
                       (N3004)? data_o[1966] : 
                       (N3006)? data_o[1998] : 
                       (N3008)? data_o[2030] : 
                       (N2883)? data_n_64__14_ : 
                       (N2885)? data_n_65__14_ : 
                       (N2887)? data_n_66__14_ : 
                       (N2889)? data_n_67__14_ : 
                       (N2891)? data_n_68__14_ : 
                       (N2893)? data_n_69__14_ : 
                       (N2895)? data_n_70__14_ : 
                       (N2897)? data_n_71__14_ : 
                       (N2899)? data_n_72__14_ : 
                       (N2901)? data_n_73__14_ : 
                       (N2903)? data_n_74__14_ : 
                       (N2905)? data_n_75__14_ : 
                       (N2907)? data_n_76__14_ : 
                       (N2909)? data_n_77__14_ : 
                       (N2911)? data_n_78__14_ : 
                       (N2913)? data_n_79__14_ : 
                       (N2915)? data_n_80__14_ : 
                       (N2917)? data_n_81__14_ : 
                       (N2919)? data_n_82__14_ : 
                       (N2921)? data_n_83__14_ : 
                       (N2923)? data_n_84__14_ : 
                       (N2925)? data_n_85__14_ : 
                       (N2927)? data_n_86__14_ : 
                       (N2929)? data_n_87__14_ : 
                       (N2931)? data_n_88__14_ : 
                       (N2933)? data_n_89__14_ : 
                       (N2935)? data_n_90__14_ : 
                       (N2937)? data_n_91__14_ : 
                       (N2939)? data_n_92__14_ : 
                       (N2941)? data_n_93__14_ : 
                       (N2943)? data_n_94__14_ : 
                       (N2945)? data_n_95__14_ : 
                       (N2947)? data_n_96__14_ : 
                       (N2949)? data_n_97__14_ : 
                       (N2951)? data_n_98__14_ : 
                       (N2953)? data_n_99__14_ : 
                       (N2955)? data_n_100__14_ : 
                       (N2957)? data_n_101__14_ : 
                       (N2959)? data_n_102__14_ : 
                       (N2961)? data_n_103__14_ : 
                       (N2963)? data_n_104__14_ : 
                       (N2965)? data_n_105__14_ : 
                       (N2967)? data_n_106__14_ : 
                       (N2969)? data_n_107__14_ : 
                       (N2971)? data_n_108__14_ : 
                       (N2973)? data_n_109__14_ : 
                       (N2975)? data_n_110__14_ : 
                       (N2977)? data_n_111__14_ : 
                       (N2979)? data_n_112__14_ : 
                       (N2981)? data_n_113__14_ : 
                       (N2983)? data_n_114__14_ : 
                       (N2985)? data_n_115__14_ : 
                       (N2987)? data_n_116__14_ : 
                       (N2989)? data_n_117__14_ : 
                       (N2991)? data_n_118__14_ : 
                       (N2993)? data_n_119__14_ : 
                       (N2995)? data_n_120__14_ : 
                       (N2997)? data_n_121__14_ : 
                       (N2999)? data_n_122__14_ : 
                       (N3001)? data_n_123__14_ : 
                       (N3003)? data_n_124__14_ : 
                       (N3005)? data_n_125__14_ : 
                       (N3007)? data_n_126__14_ : 
                       (N3009)? data_n_127__14_ : 1'b0;
  assign data_nn[13] = (N2882)? data_o[13] : 
                       (N2884)? data_o[45] : 
                       (N2886)? data_o[77] : 
                       (N2888)? data_o[109] : 
                       (N2890)? data_o[141] : 
                       (N2892)? data_o[173] : 
                       (N2894)? data_o[205] : 
                       (N2896)? data_o[237] : 
                       (N2898)? data_o[269] : 
                       (N2900)? data_o[301] : 
                       (N2902)? data_o[333] : 
                       (N2904)? data_o[365] : 
                       (N2906)? data_o[397] : 
                       (N2908)? data_o[429] : 
                       (N2910)? data_o[461] : 
                       (N2912)? data_o[493] : 
                       (N2914)? data_o[525] : 
                       (N2916)? data_o[557] : 
                       (N2918)? data_o[589] : 
                       (N2920)? data_o[621] : 
                       (N2922)? data_o[653] : 
                       (N2924)? data_o[685] : 
                       (N2926)? data_o[717] : 
                       (N2928)? data_o[749] : 
                       (N2930)? data_o[781] : 
                       (N2932)? data_o[813] : 
                       (N2934)? data_o[845] : 
                       (N2936)? data_o[877] : 
                       (N2938)? data_o[909] : 
                       (N2940)? data_o[941] : 
                       (N2942)? data_o[973] : 
                       (N2944)? data_o[1005] : 
                       (N2946)? data_o[1037] : 
                       (N2948)? data_o[1069] : 
                       (N2950)? data_o[1101] : 
                       (N2952)? data_o[1133] : 
                       (N2954)? data_o[1165] : 
                       (N2956)? data_o[1197] : 
                       (N2958)? data_o[1229] : 
                       (N2960)? data_o[1261] : 
                       (N2962)? data_o[1293] : 
                       (N2964)? data_o[1325] : 
                       (N2966)? data_o[1357] : 
                       (N2968)? data_o[1389] : 
                       (N2970)? data_o[1421] : 
                       (N2972)? data_o[1453] : 
                       (N2974)? data_o[1485] : 
                       (N2976)? data_o[1517] : 
                       (N2978)? data_o[1549] : 
                       (N2980)? data_o[1581] : 
                       (N2982)? data_o[1613] : 
                       (N2984)? data_o[1645] : 
                       (N2986)? data_o[1677] : 
                       (N2988)? data_o[1709] : 
                       (N2990)? data_o[1741] : 
                       (N2992)? data_o[1773] : 
                       (N2994)? data_o[1805] : 
                       (N2996)? data_o[1837] : 
                       (N2998)? data_o[1869] : 
                       (N3000)? data_o[1901] : 
                       (N3002)? data_o[1933] : 
                       (N3004)? data_o[1965] : 
                       (N3006)? data_o[1997] : 
                       (N3008)? data_o[2029] : 
                       (N2883)? data_n_64__13_ : 
                       (N2885)? data_n_65__13_ : 
                       (N2887)? data_n_66__13_ : 
                       (N2889)? data_n_67__13_ : 
                       (N2891)? data_n_68__13_ : 
                       (N2893)? data_n_69__13_ : 
                       (N2895)? data_n_70__13_ : 
                       (N2897)? data_n_71__13_ : 
                       (N2899)? data_n_72__13_ : 
                       (N2901)? data_n_73__13_ : 
                       (N2903)? data_n_74__13_ : 
                       (N2905)? data_n_75__13_ : 
                       (N2907)? data_n_76__13_ : 
                       (N2909)? data_n_77__13_ : 
                       (N2911)? data_n_78__13_ : 
                       (N2913)? data_n_79__13_ : 
                       (N2915)? data_n_80__13_ : 
                       (N2917)? data_n_81__13_ : 
                       (N2919)? data_n_82__13_ : 
                       (N2921)? data_n_83__13_ : 
                       (N2923)? data_n_84__13_ : 
                       (N2925)? data_n_85__13_ : 
                       (N2927)? data_n_86__13_ : 
                       (N2929)? data_n_87__13_ : 
                       (N2931)? data_n_88__13_ : 
                       (N2933)? data_n_89__13_ : 
                       (N2935)? data_n_90__13_ : 
                       (N2937)? data_n_91__13_ : 
                       (N2939)? data_n_92__13_ : 
                       (N2941)? data_n_93__13_ : 
                       (N2943)? data_n_94__13_ : 
                       (N2945)? data_n_95__13_ : 
                       (N2947)? data_n_96__13_ : 
                       (N2949)? data_n_97__13_ : 
                       (N2951)? data_n_98__13_ : 
                       (N2953)? data_n_99__13_ : 
                       (N2955)? data_n_100__13_ : 
                       (N2957)? data_n_101__13_ : 
                       (N2959)? data_n_102__13_ : 
                       (N2961)? data_n_103__13_ : 
                       (N2963)? data_n_104__13_ : 
                       (N2965)? data_n_105__13_ : 
                       (N2967)? data_n_106__13_ : 
                       (N2969)? data_n_107__13_ : 
                       (N2971)? data_n_108__13_ : 
                       (N2973)? data_n_109__13_ : 
                       (N2975)? data_n_110__13_ : 
                       (N2977)? data_n_111__13_ : 
                       (N2979)? data_n_112__13_ : 
                       (N2981)? data_n_113__13_ : 
                       (N2983)? data_n_114__13_ : 
                       (N2985)? data_n_115__13_ : 
                       (N2987)? data_n_116__13_ : 
                       (N2989)? data_n_117__13_ : 
                       (N2991)? data_n_118__13_ : 
                       (N2993)? data_n_119__13_ : 
                       (N2995)? data_n_120__13_ : 
                       (N2997)? data_n_121__13_ : 
                       (N2999)? data_n_122__13_ : 
                       (N3001)? data_n_123__13_ : 
                       (N3003)? data_n_124__13_ : 
                       (N3005)? data_n_125__13_ : 
                       (N3007)? data_n_126__13_ : 
                       (N3009)? data_n_127__13_ : 1'b0;
  assign data_nn[12] = (N2882)? data_o[12] : 
                       (N2884)? data_o[44] : 
                       (N2886)? data_o[76] : 
                       (N2888)? data_o[108] : 
                       (N2890)? data_o[140] : 
                       (N2892)? data_o[172] : 
                       (N2894)? data_o[204] : 
                       (N2896)? data_o[236] : 
                       (N2898)? data_o[268] : 
                       (N2900)? data_o[300] : 
                       (N2902)? data_o[332] : 
                       (N2904)? data_o[364] : 
                       (N2906)? data_o[396] : 
                       (N2908)? data_o[428] : 
                       (N2910)? data_o[460] : 
                       (N2912)? data_o[492] : 
                       (N2914)? data_o[524] : 
                       (N2916)? data_o[556] : 
                       (N2918)? data_o[588] : 
                       (N2920)? data_o[620] : 
                       (N2922)? data_o[652] : 
                       (N2924)? data_o[684] : 
                       (N2926)? data_o[716] : 
                       (N2928)? data_o[748] : 
                       (N2930)? data_o[780] : 
                       (N2932)? data_o[812] : 
                       (N2934)? data_o[844] : 
                       (N2936)? data_o[876] : 
                       (N2938)? data_o[908] : 
                       (N2940)? data_o[940] : 
                       (N2942)? data_o[972] : 
                       (N2944)? data_o[1004] : 
                       (N2946)? data_o[1036] : 
                       (N2948)? data_o[1068] : 
                       (N2950)? data_o[1100] : 
                       (N2952)? data_o[1132] : 
                       (N2954)? data_o[1164] : 
                       (N2956)? data_o[1196] : 
                       (N2958)? data_o[1228] : 
                       (N2960)? data_o[1260] : 
                       (N2962)? data_o[1292] : 
                       (N2964)? data_o[1324] : 
                       (N2966)? data_o[1356] : 
                       (N2968)? data_o[1388] : 
                       (N2970)? data_o[1420] : 
                       (N2972)? data_o[1452] : 
                       (N2974)? data_o[1484] : 
                       (N2976)? data_o[1516] : 
                       (N2978)? data_o[1548] : 
                       (N2980)? data_o[1580] : 
                       (N2982)? data_o[1612] : 
                       (N2984)? data_o[1644] : 
                       (N2986)? data_o[1676] : 
                       (N2988)? data_o[1708] : 
                       (N2990)? data_o[1740] : 
                       (N2992)? data_o[1772] : 
                       (N2994)? data_o[1804] : 
                       (N2996)? data_o[1836] : 
                       (N2998)? data_o[1868] : 
                       (N3000)? data_o[1900] : 
                       (N3002)? data_o[1932] : 
                       (N3004)? data_o[1964] : 
                       (N3006)? data_o[1996] : 
                       (N3008)? data_o[2028] : 
                       (N2883)? data_n_64__12_ : 
                       (N2885)? data_n_65__12_ : 
                       (N2887)? data_n_66__12_ : 
                       (N2889)? data_n_67__12_ : 
                       (N2891)? data_n_68__12_ : 
                       (N2893)? data_n_69__12_ : 
                       (N2895)? data_n_70__12_ : 
                       (N2897)? data_n_71__12_ : 
                       (N2899)? data_n_72__12_ : 
                       (N2901)? data_n_73__12_ : 
                       (N2903)? data_n_74__12_ : 
                       (N2905)? data_n_75__12_ : 
                       (N2907)? data_n_76__12_ : 
                       (N2909)? data_n_77__12_ : 
                       (N2911)? data_n_78__12_ : 
                       (N2913)? data_n_79__12_ : 
                       (N2915)? data_n_80__12_ : 
                       (N2917)? data_n_81__12_ : 
                       (N2919)? data_n_82__12_ : 
                       (N2921)? data_n_83__12_ : 
                       (N2923)? data_n_84__12_ : 
                       (N2925)? data_n_85__12_ : 
                       (N2927)? data_n_86__12_ : 
                       (N2929)? data_n_87__12_ : 
                       (N2931)? data_n_88__12_ : 
                       (N2933)? data_n_89__12_ : 
                       (N2935)? data_n_90__12_ : 
                       (N2937)? data_n_91__12_ : 
                       (N2939)? data_n_92__12_ : 
                       (N2941)? data_n_93__12_ : 
                       (N2943)? data_n_94__12_ : 
                       (N2945)? data_n_95__12_ : 
                       (N2947)? data_n_96__12_ : 
                       (N2949)? data_n_97__12_ : 
                       (N2951)? data_n_98__12_ : 
                       (N2953)? data_n_99__12_ : 
                       (N2955)? data_n_100__12_ : 
                       (N2957)? data_n_101__12_ : 
                       (N2959)? data_n_102__12_ : 
                       (N2961)? data_n_103__12_ : 
                       (N2963)? data_n_104__12_ : 
                       (N2965)? data_n_105__12_ : 
                       (N2967)? data_n_106__12_ : 
                       (N2969)? data_n_107__12_ : 
                       (N2971)? data_n_108__12_ : 
                       (N2973)? data_n_109__12_ : 
                       (N2975)? data_n_110__12_ : 
                       (N2977)? data_n_111__12_ : 
                       (N2979)? data_n_112__12_ : 
                       (N2981)? data_n_113__12_ : 
                       (N2983)? data_n_114__12_ : 
                       (N2985)? data_n_115__12_ : 
                       (N2987)? data_n_116__12_ : 
                       (N2989)? data_n_117__12_ : 
                       (N2991)? data_n_118__12_ : 
                       (N2993)? data_n_119__12_ : 
                       (N2995)? data_n_120__12_ : 
                       (N2997)? data_n_121__12_ : 
                       (N2999)? data_n_122__12_ : 
                       (N3001)? data_n_123__12_ : 
                       (N3003)? data_n_124__12_ : 
                       (N3005)? data_n_125__12_ : 
                       (N3007)? data_n_126__12_ : 
                       (N3009)? data_n_127__12_ : 1'b0;
  assign data_nn[11] = (N2882)? data_o[11] : 
                       (N2884)? data_o[43] : 
                       (N2886)? data_o[75] : 
                       (N2888)? data_o[107] : 
                       (N2890)? data_o[139] : 
                       (N2892)? data_o[171] : 
                       (N2894)? data_o[203] : 
                       (N2896)? data_o[235] : 
                       (N2898)? data_o[267] : 
                       (N2900)? data_o[299] : 
                       (N2902)? data_o[331] : 
                       (N2904)? data_o[363] : 
                       (N2906)? data_o[395] : 
                       (N2908)? data_o[427] : 
                       (N2910)? data_o[459] : 
                       (N2912)? data_o[491] : 
                       (N2914)? data_o[523] : 
                       (N2916)? data_o[555] : 
                       (N2918)? data_o[587] : 
                       (N2920)? data_o[619] : 
                       (N2922)? data_o[651] : 
                       (N2924)? data_o[683] : 
                       (N2926)? data_o[715] : 
                       (N2928)? data_o[747] : 
                       (N2930)? data_o[779] : 
                       (N2932)? data_o[811] : 
                       (N2934)? data_o[843] : 
                       (N2936)? data_o[875] : 
                       (N2938)? data_o[907] : 
                       (N2940)? data_o[939] : 
                       (N2942)? data_o[971] : 
                       (N2944)? data_o[1003] : 
                       (N2946)? data_o[1035] : 
                       (N2948)? data_o[1067] : 
                       (N2950)? data_o[1099] : 
                       (N2952)? data_o[1131] : 
                       (N2954)? data_o[1163] : 
                       (N2956)? data_o[1195] : 
                       (N2958)? data_o[1227] : 
                       (N2960)? data_o[1259] : 
                       (N2962)? data_o[1291] : 
                       (N2964)? data_o[1323] : 
                       (N2966)? data_o[1355] : 
                       (N2968)? data_o[1387] : 
                       (N2970)? data_o[1419] : 
                       (N2972)? data_o[1451] : 
                       (N2974)? data_o[1483] : 
                       (N2976)? data_o[1515] : 
                       (N2978)? data_o[1547] : 
                       (N2980)? data_o[1579] : 
                       (N2982)? data_o[1611] : 
                       (N2984)? data_o[1643] : 
                       (N2986)? data_o[1675] : 
                       (N2988)? data_o[1707] : 
                       (N2990)? data_o[1739] : 
                       (N2992)? data_o[1771] : 
                       (N2994)? data_o[1803] : 
                       (N2996)? data_o[1835] : 
                       (N2998)? data_o[1867] : 
                       (N3000)? data_o[1899] : 
                       (N3002)? data_o[1931] : 
                       (N3004)? data_o[1963] : 
                       (N3006)? data_o[1995] : 
                       (N3008)? data_o[2027] : 
                       (N2883)? data_n_64__11_ : 
                       (N2885)? data_n_65__11_ : 
                       (N2887)? data_n_66__11_ : 
                       (N2889)? data_n_67__11_ : 
                       (N2891)? data_n_68__11_ : 
                       (N2893)? data_n_69__11_ : 
                       (N2895)? data_n_70__11_ : 
                       (N2897)? data_n_71__11_ : 
                       (N2899)? data_n_72__11_ : 
                       (N2901)? data_n_73__11_ : 
                       (N2903)? data_n_74__11_ : 
                       (N2905)? data_n_75__11_ : 
                       (N2907)? data_n_76__11_ : 
                       (N2909)? data_n_77__11_ : 
                       (N2911)? data_n_78__11_ : 
                       (N2913)? data_n_79__11_ : 
                       (N2915)? data_n_80__11_ : 
                       (N2917)? data_n_81__11_ : 
                       (N2919)? data_n_82__11_ : 
                       (N2921)? data_n_83__11_ : 
                       (N2923)? data_n_84__11_ : 
                       (N2925)? data_n_85__11_ : 
                       (N2927)? data_n_86__11_ : 
                       (N2929)? data_n_87__11_ : 
                       (N2931)? data_n_88__11_ : 
                       (N2933)? data_n_89__11_ : 
                       (N2935)? data_n_90__11_ : 
                       (N2937)? data_n_91__11_ : 
                       (N2939)? data_n_92__11_ : 
                       (N2941)? data_n_93__11_ : 
                       (N2943)? data_n_94__11_ : 
                       (N2945)? data_n_95__11_ : 
                       (N2947)? data_n_96__11_ : 
                       (N2949)? data_n_97__11_ : 
                       (N2951)? data_n_98__11_ : 
                       (N2953)? data_n_99__11_ : 
                       (N2955)? data_n_100__11_ : 
                       (N2957)? data_n_101__11_ : 
                       (N2959)? data_n_102__11_ : 
                       (N2961)? data_n_103__11_ : 
                       (N2963)? data_n_104__11_ : 
                       (N2965)? data_n_105__11_ : 
                       (N2967)? data_n_106__11_ : 
                       (N2969)? data_n_107__11_ : 
                       (N2971)? data_n_108__11_ : 
                       (N2973)? data_n_109__11_ : 
                       (N2975)? data_n_110__11_ : 
                       (N2977)? data_n_111__11_ : 
                       (N2979)? data_n_112__11_ : 
                       (N2981)? data_n_113__11_ : 
                       (N2983)? data_n_114__11_ : 
                       (N2985)? data_n_115__11_ : 
                       (N2987)? data_n_116__11_ : 
                       (N2989)? data_n_117__11_ : 
                       (N2991)? data_n_118__11_ : 
                       (N2993)? data_n_119__11_ : 
                       (N2995)? data_n_120__11_ : 
                       (N2997)? data_n_121__11_ : 
                       (N2999)? data_n_122__11_ : 
                       (N3001)? data_n_123__11_ : 
                       (N3003)? data_n_124__11_ : 
                       (N3005)? data_n_125__11_ : 
                       (N3007)? data_n_126__11_ : 
                       (N3009)? data_n_127__11_ : 1'b0;
  assign data_nn[10] = (N2882)? data_o[10] : 
                       (N2884)? data_o[42] : 
                       (N2886)? data_o[74] : 
                       (N2888)? data_o[106] : 
                       (N2890)? data_o[138] : 
                       (N2892)? data_o[170] : 
                       (N2894)? data_o[202] : 
                       (N2896)? data_o[234] : 
                       (N2898)? data_o[266] : 
                       (N2900)? data_o[298] : 
                       (N2902)? data_o[330] : 
                       (N2904)? data_o[362] : 
                       (N2906)? data_o[394] : 
                       (N2908)? data_o[426] : 
                       (N2910)? data_o[458] : 
                       (N2912)? data_o[490] : 
                       (N2914)? data_o[522] : 
                       (N2916)? data_o[554] : 
                       (N2918)? data_o[586] : 
                       (N2920)? data_o[618] : 
                       (N2922)? data_o[650] : 
                       (N2924)? data_o[682] : 
                       (N2926)? data_o[714] : 
                       (N2928)? data_o[746] : 
                       (N2930)? data_o[778] : 
                       (N2932)? data_o[810] : 
                       (N2934)? data_o[842] : 
                       (N2936)? data_o[874] : 
                       (N2938)? data_o[906] : 
                       (N2940)? data_o[938] : 
                       (N2942)? data_o[970] : 
                       (N2944)? data_o[1002] : 
                       (N2946)? data_o[1034] : 
                       (N2948)? data_o[1066] : 
                       (N2950)? data_o[1098] : 
                       (N2952)? data_o[1130] : 
                       (N2954)? data_o[1162] : 
                       (N2956)? data_o[1194] : 
                       (N2958)? data_o[1226] : 
                       (N2960)? data_o[1258] : 
                       (N2962)? data_o[1290] : 
                       (N2964)? data_o[1322] : 
                       (N2966)? data_o[1354] : 
                       (N2968)? data_o[1386] : 
                       (N2970)? data_o[1418] : 
                       (N2972)? data_o[1450] : 
                       (N2974)? data_o[1482] : 
                       (N2976)? data_o[1514] : 
                       (N2978)? data_o[1546] : 
                       (N2980)? data_o[1578] : 
                       (N2982)? data_o[1610] : 
                       (N2984)? data_o[1642] : 
                       (N2986)? data_o[1674] : 
                       (N2988)? data_o[1706] : 
                       (N2990)? data_o[1738] : 
                       (N2992)? data_o[1770] : 
                       (N2994)? data_o[1802] : 
                       (N2996)? data_o[1834] : 
                       (N2998)? data_o[1866] : 
                       (N3000)? data_o[1898] : 
                       (N3002)? data_o[1930] : 
                       (N3004)? data_o[1962] : 
                       (N3006)? data_o[1994] : 
                       (N3008)? data_o[2026] : 
                       (N2883)? data_n_64__10_ : 
                       (N2885)? data_n_65__10_ : 
                       (N2887)? data_n_66__10_ : 
                       (N2889)? data_n_67__10_ : 
                       (N2891)? data_n_68__10_ : 
                       (N2893)? data_n_69__10_ : 
                       (N2895)? data_n_70__10_ : 
                       (N2897)? data_n_71__10_ : 
                       (N2899)? data_n_72__10_ : 
                       (N2901)? data_n_73__10_ : 
                       (N2903)? data_n_74__10_ : 
                       (N2905)? data_n_75__10_ : 
                       (N2907)? data_n_76__10_ : 
                       (N2909)? data_n_77__10_ : 
                       (N2911)? data_n_78__10_ : 
                       (N2913)? data_n_79__10_ : 
                       (N2915)? data_n_80__10_ : 
                       (N2917)? data_n_81__10_ : 
                       (N2919)? data_n_82__10_ : 
                       (N2921)? data_n_83__10_ : 
                       (N2923)? data_n_84__10_ : 
                       (N2925)? data_n_85__10_ : 
                       (N2927)? data_n_86__10_ : 
                       (N2929)? data_n_87__10_ : 
                       (N2931)? data_n_88__10_ : 
                       (N2933)? data_n_89__10_ : 
                       (N2935)? data_n_90__10_ : 
                       (N2937)? data_n_91__10_ : 
                       (N2939)? data_n_92__10_ : 
                       (N2941)? data_n_93__10_ : 
                       (N2943)? data_n_94__10_ : 
                       (N2945)? data_n_95__10_ : 
                       (N2947)? data_n_96__10_ : 
                       (N2949)? data_n_97__10_ : 
                       (N2951)? data_n_98__10_ : 
                       (N2953)? data_n_99__10_ : 
                       (N2955)? data_n_100__10_ : 
                       (N2957)? data_n_101__10_ : 
                       (N2959)? data_n_102__10_ : 
                       (N2961)? data_n_103__10_ : 
                       (N2963)? data_n_104__10_ : 
                       (N2965)? data_n_105__10_ : 
                       (N2967)? data_n_106__10_ : 
                       (N2969)? data_n_107__10_ : 
                       (N2971)? data_n_108__10_ : 
                       (N2973)? data_n_109__10_ : 
                       (N2975)? data_n_110__10_ : 
                       (N2977)? data_n_111__10_ : 
                       (N2979)? data_n_112__10_ : 
                       (N2981)? data_n_113__10_ : 
                       (N2983)? data_n_114__10_ : 
                       (N2985)? data_n_115__10_ : 
                       (N2987)? data_n_116__10_ : 
                       (N2989)? data_n_117__10_ : 
                       (N2991)? data_n_118__10_ : 
                       (N2993)? data_n_119__10_ : 
                       (N2995)? data_n_120__10_ : 
                       (N2997)? data_n_121__10_ : 
                       (N2999)? data_n_122__10_ : 
                       (N3001)? data_n_123__10_ : 
                       (N3003)? data_n_124__10_ : 
                       (N3005)? data_n_125__10_ : 
                       (N3007)? data_n_126__10_ : 
                       (N3009)? data_n_127__10_ : 1'b0;
  assign data_nn[9] = (N2882)? data_o[9] : 
                      (N2884)? data_o[41] : 
                      (N2886)? data_o[73] : 
                      (N2888)? data_o[105] : 
                      (N2890)? data_o[137] : 
                      (N2892)? data_o[169] : 
                      (N2894)? data_o[201] : 
                      (N2896)? data_o[233] : 
                      (N2898)? data_o[265] : 
                      (N2900)? data_o[297] : 
                      (N2902)? data_o[329] : 
                      (N2904)? data_o[361] : 
                      (N2906)? data_o[393] : 
                      (N2908)? data_o[425] : 
                      (N2910)? data_o[457] : 
                      (N2912)? data_o[489] : 
                      (N2914)? data_o[521] : 
                      (N2916)? data_o[553] : 
                      (N2918)? data_o[585] : 
                      (N2920)? data_o[617] : 
                      (N2922)? data_o[649] : 
                      (N2924)? data_o[681] : 
                      (N2926)? data_o[713] : 
                      (N2928)? data_o[745] : 
                      (N2930)? data_o[777] : 
                      (N2932)? data_o[809] : 
                      (N2934)? data_o[841] : 
                      (N2936)? data_o[873] : 
                      (N2938)? data_o[905] : 
                      (N2940)? data_o[937] : 
                      (N2942)? data_o[969] : 
                      (N2944)? data_o[1001] : 
                      (N2946)? data_o[1033] : 
                      (N2948)? data_o[1065] : 
                      (N2950)? data_o[1097] : 
                      (N2952)? data_o[1129] : 
                      (N2954)? data_o[1161] : 
                      (N2956)? data_o[1193] : 
                      (N2958)? data_o[1225] : 
                      (N2960)? data_o[1257] : 
                      (N2962)? data_o[1289] : 
                      (N2964)? data_o[1321] : 
                      (N2966)? data_o[1353] : 
                      (N2968)? data_o[1385] : 
                      (N2970)? data_o[1417] : 
                      (N2972)? data_o[1449] : 
                      (N2974)? data_o[1481] : 
                      (N2976)? data_o[1513] : 
                      (N2978)? data_o[1545] : 
                      (N2980)? data_o[1577] : 
                      (N2982)? data_o[1609] : 
                      (N2984)? data_o[1641] : 
                      (N2986)? data_o[1673] : 
                      (N2988)? data_o[1705] : 
                      (N2990)? data_o[1737] : 
                      (N2992)? data_o[1769] : 
                      (N2994)? data_o[1801] : 
                      (N2996)? data_o[1833] : 
                      (N2998)? data_o[1865] : 
                      (N3000)? data_o[1897] : 
                      (N3002)? data_o[1929] : 
                      (N3004)? data_o[1961] : 
                      (N3006)? data_o[1993] : 
                      (N3008)? data_o[2025] : 
                      (N2883)? data_n_64__9_ : 
                      (N2885)? data_n_65__9_ : 
                      (N2887)? data_n_66__9_ : 
                      (N2889)? data_n_67__9_ : 
                      (N2891)? data_n_68__9_ : 
                      (N2893)? data_n_69__9_ : 
                      (N2895)? data_n_70__9_ : 
                      (N2897)? data_n_71__9_ : 
                      (N2899)? data_n_72__9_ : 
                      (N2901)? data_n_73__9_ : 
                      (N2903)? data_n_74__9_ : 
                      (N2905)? data_n_75__9_ : 
                      (N2907)? data_n_76__9_ : 
                      (N2909)? data_n_77__9_ : 
                      (N2911)? data_n_78__9_ : 
                      (N2913)? data_n_79__9_ : 
                      (N2915)? data_n_80__9_ : 
                      (N2917)? data_n_81__9_ : 
                      (N2919)? data_n_82__9_ : 
                      (N2921)? data_n_83__9_ : 
                      (N2923)? data_n_84__9_ : 
                      (N2925)? data_n_85__9_ : 
                      (N2927)? data_n_86__9_ : 
                      (N2929)? data_n_87__9_ : 
                      (N2931)? data_n_88__9_ : 
                      (N2933)? data_n_89__9_ : 
                      (N2935)? data_n_90__9_ : 
                      (N2937)? data_n_91__9_ : 
                      (N2939)? data_n_92__9_ : 
                      (N2941)? data_n_93__9_ : 
                      (N2943)? data_n_94__9_ : 
                      (N2945)? data_n_95__9_ : 
                      (N2947)? data_n_96__9_ : 
                      (N2949)? data_n_97__9_ : 
                      (N2951)? data_n_98__9_ : 
                      (N2953)? data_n_99__9_ : 
                      (N2955)? data_n_100__9_ : 
                      (N2957)? data_n_101__9_ : 
                      (N2959)? data_n_102__9_ : 
                      (N2961)? data_n_103__9_ : 
                      (N2963)? data_n_104__9_ : 
                      (N2965)? data_n_105__9_ : 
                      (N2967)? data_n_106__9_ : 
                      (N2969)? data_n_107__9_ : 
                      (N2971)? data_n_108__9_ : 
                      (N2973)? data_n_109__9_ : 
                      (N2975)? data_n_110__9_ : 
                      (N2977)? data_n_111__9_ : 
                      (N2979)? data_n_112__9_ : 
                      (N2981)? data_n_113__9_ : 
                      (N2983)? data_n_114__9_ : 
                      (N2985)? data_n_115__9_ : 
                      (N2987)? data_n_116__9_ : 
                      (N2989)? data_n_117__9_ : 
                      (N2991)? data_n_118__9_ : 
                      (N2993)? data_n_119__9_ : 
                      (N2995)? data_n_120__9_ : 
                      (N2997)? data_n_121__9_ : 
                      (N2999)? data_n_122__9_ : 
                      (N3001)? data_n_123__9_ : 
                      (N3003)? data_n_124__9_ : 
                      (N3005)? data_n_125__9_ : 
                      (N3007)? data_n_126__9_ : 
                      (N3009)? data_n_127__9_ : 1'b0;
  assign data_nn[8] = (N2882)? data_o[8] : 
                      (N2884)? data_o[40] : 
                      (N2886)? data_o[72] : 
                      (N2888)? data_o[104] : 
                      (N2890)? data_o[136] : 
                      (N2892)? data_o[168] : 
                      (N2894)? data_o[200] : 
                      (N2896)? data_o[232] : 
                      (N2898)? data_o[264] : 
                      (N2900)? data_o[296] : 
                      (N2902)? data_o[328] : 
                      (N2904)? data_o[360] : 
                      (N2906)? data_o[392] : 
                      (N2908)? data_o[424] : 
                      (N2910)? data_o[456] : 
                      (N2912)? data_o[488] : 
                      (N2914)? data_o[520] : 
                      (N2916)? data_o[552] : 
                      (N2918)? data_o[584] : 
                      (N2920)? data_o[616] : 
                      (N2922)? data_o[648] : 
                      (N2924)? data_o[680] : 
                      (N2926)? data_o[712] : 
                      (N2928)? data_o[744] : 
                      (N2930)? data_o[776] : 
                      (N2932)? data_o[808] : 
                      (N2934)? data_o[840] : 
                      (N2936)? data_o[872] : 
                      (N2938)? data_o[904] : 
                      (N2940)? data_o[936] : 
                      (N2942)? data_o[968] : 
                      (N2944)? data_o[1000] : 
                      (N2946)? data_o[1032] : 
                      (N2948)? data_o[1064] : 
                      (N2950)? data_o[1096] : 
                      (N2952)? data_o[1128] : 
                      (N2954)? data_o[1160] : 
                      (N2956)? data_o[1192] : 
                      (N2958)? data_o[1224] : 
                      (N2960)? data_o[1256] : 
                      (N2962)? data_o[1288] : 
                      (N2964)? data_o[1320] : 
                      (N2966)? data_o[1352] : 
                      (N2968)? data_o[1384] : 
                      (N2970)? data_o[1416] : 
                      (N2972)? data_o[1448] : 
                      (N2974)? data_o[1480] : 
                      (N2976)? data_o[1512] : 
                      (N2978)? data_o[1544] : 
                      (N2980)? data_o[1576] : 
                      (N2982)? data_o[1608] : 
                      (N2984)? data_o[1640] : 
                      (N2986)? data_o[1672] : 
                      (N2988)? data_o[1704] : 
                      (N2990)? data_o[1736] : 
                      (N2992)? data_o[1768] : 
                      (N2994)? data_o[1800] : 
                      (N2996)? data_o[1832] : 
                      (N2998)? data_o[1864] : 
                      (N3000)? data_o[1896] : 
                      (N3002)? data_o[1928] : 
                      (N3004)? data_o[1960] : 
                      (N3006)? data_o[1992] : 
                      (N3008)? data_o[2024] : 
                      (N2883)? data_n_64__8_ : 
                      (N2885)? data_n_65__8_ : 
                      (N2887)? data_n_66__8_ : 
                      (N2889)? data_n_67__8_ : 
                      (N2891)? data_n_68__8_ : 
                      (N2893)? data_n_69__8_ : 
                      (N2895)? data_n_70__8_ : 
                      (N2897)? data_n_71__8_ : 
                      (N2899)? data_n_72__8_ : 
                      (N2901)? data_n_73__8_ : 
                      (N2903)? data_n_74__8_ : 
                      (N2905)? data_n_75__8_ : 
                      (N2907)? data_n_76__8_ : 
                      (N2909)? data_n_77__8_ : 
                      (N2911)? data_n_78__8_ : 
                      (N2913)? data_n_79__8_ : 
                      (N2915)? data_n_80__8_ : 
                      (N2917)? data_n_81__8_ : 
                      (N2919)? data_n_82__8_ : 
                      (N2921)? data_n_83__8_ : 
                      (N2923)? data_n_84__8_ : 
                      (N2925)? data_n_85__8_ : 
                      (N2927)? data_n_86__8_ : 
                      (N2929)? data_n_87__8_ : 
                      (N2931)? data_n_88__8_ : 
                      (N2933)? data_n_89__8_ : 
                      (N2935)? data_n_90__8_ : 
                      (N2937)? data_n_91__8_ : 
                      (N2939)? data_n_92__8_ : 
                      (N2941)? data_n_93__8_ : 
                      (N2943)? data_n_94__8_ : 
                      (N2945)? data_n_95__8_ : 
                      (N2947)? data_n_96__8_ : 
                      (N2949)? data_n_97__8_ : 
                      (N2951)? data_n_98__8_ : 
                      (N2953)? data_n_99__8_ : 
                      (N2955)? data_n_100__8_ : 
                      (N2957)? data_n_101__8_ : 
                      (N2959)? data_n_102__8_ : 
                      (N2961)? data_n_103__8_ : 
                      (N2963)? data_n_104__8_ : 
                      (N2965)? data_n_105__8_ : 
                      (N2967)? data_n_106__8_ : 
                      (N2969)? data_n_107__8_ : 
                      (N2971)? data_n_108__8_ : 
                      (N2973)? data_n_109__8_ : 
                      (N2975)? data_n_110__8_ : 
                      (N2977)? data_n_111__8_ : 
                      (N2979)? data_n_112__8_ : 
                      (N2981)? data_n_113__8_ : 
                      (N2983)? data_n_114__8_ : 
                      (N2985)? data_n_115__8_ : 
                      (N2987)? data_n_116__8_ : 
                      (N2989)? data_n_117__8_ : 
                      (N2991)? data_n_118__8_ : 
                      (N2993)? data_n_119__8_ : 
                      (N2995)? data_n_120__8_ : 
                      (N2997)? data_n_121__8_ : 
                      (N2999)? data_n_122__8_ : 
                      (N3001)? data_n_123__8_ : 
                      (N3003)? data_n_124__8_ : 
                      (N3005)? data_n_125__8_ : 
                      (N3007)? data_n_126__8_ : 
                      (N3009)? data_n_127__8_ : 1'b0;
  assign data_nn[7] = (N2882)? data_o[7] : 
                      (N2884)? data_o[39] : 
                      (N2886)? data_o[71] : 
                      (N2888)? data_o[103] : 
                      (N2890)? data_o[135] : 
                      (N2892)? data_o[167] : 
                      (N2894)? data_o[199] : 
                      (N2896)? data_o[231] : 
                      (N2898)? data_o[263] : 
                      (N2900)? data_o[295] : 
                      (N2902)? data_o[327] : 
                      (N2904)? data_o[359] : 
                      (N2906)? data_o[391] : 
                      (N2908)? data_o[423] : 
                      (N2910)? data_o[455] : 
                      (N2912)? data_o[487] : 
                      (N2914)? data_o[519] : 
                      (N2916)? data_o[551] : 
                      (N2918)? data_o[583] : 
                      (N2920)? data_o[615] : 
                      (N2922)? data_o[647] : 
                      (N2924)? data_o[679] : 
                      (N2926)? data_o[711] : 
                      (N2928)? data_o[743] : 
                      (N2930)? data_o[775] : 
                      (N2932)? data_o[807] : 
                      (N2934)? data_o[839] : 
                      (N2936)? data_o[871] : 
                      (N2938)? data_o[903] : 
                      (N2940)? data_o[935] : 
                      (N2942)? data_o[967] : 
                      (N2944)? data_o[999] : 
                      (N2946)? data_o[1031] : 
                      (N2948)? data_o[1063] : 
                      (N2950)? data_o[1095] : 
                      (N2952)? data_o[1127] : 
                      (N2954)? data_o[1159] : 
                      (N2956)? data_o[1191] : 
                      (N2958)? data_o[1223] : 
                      (N2960)? data_o[1255] : 
                      (N2962)? data_o[1287] : 
                      (N2964)? data_o[1319] : 
                      (N2966)? data_o[1351] : 
                      (N2968)? data_o[1383] : 
                      (N2970)? data_o[1415] : 
                      (N2972)? data_o[1447] : 
                      (N2974)? data_o[1479] : 
                      (N2976)? data_o[1511] : 
                      (N2978)? data_o[1543] : 
                      (N2980)? data_o[1575] : 
                      (N2982)? data_o[1607] : 
                      (N2984)? data_o[1639] : 
                      (N2986)? data_o[1671] : 
                      (N2988)? data_o[1703] : 
                      (N2990)? data_o[1735] : 
                      (N2992)? data_o[1767] : 
                      (N2994)? data_o[1799] : 
                      (N2996)? data_o[1831] : 
                      (N2998)? data_o[1863] : 
                      (N3000)? data_o[1895] : 
                      (N3002)? data_o[1927] : 
                      (N3004)? data_o[1959] : 
                      (N3006)? data_o[1991] : 
                      (N3008)? data_o[2023] : 
                      (N2883)? data_n_64__7_ : 
                      (N2885)? data_n_65__7_ : 
                      (N2887)? data_n_66__7_ : 
                      (N2889)? data_n_67__7_ : 
                      (N2891)? data_n_68__7_ : 
                      (N2893)? data_n_69__7_ : 
                      (N2895)? data_n_70__7_ : 
                      (N2897)? data_n_71__7_ : 
                      (N2899)? data_n_72__7_ : 
                      (N2901)? data_n_73__7_ : 
                      (N2903)? data_n_74__7_ : 
                      (N2905)? data_n_75__7_ : 
                      (N2907)? data_n_76__7_ : 
                      (N2909)? data_n_77__7_ : 
                      (N2911)? data_n_78__7_ : 
                      (N2913)? data_n_79__7_ : 
                      (N2915)? data_n_80__7_ : 
                      (N2917)? data_n_81__7_ : 
                      (N2919)? data_n_82__7_ : 
                      (N2921)? data_n_83__7_ : 
                      (N2923)? data_n_84__7_ : 
                      (N2925)? data_n_85__7_ : 
                      (N2927)? data_n_86__7_ : 
                      (N2929)? data_n_87__7_ : 
                      (N2931)? data_n_88__7_ : 
                      (N2933)? data_n_89__7_ : 
                      (N2935)? data_n_90__7_ : 
                      (N2937)? data_n_91__7_ : 
                      (N2939)? data_n_92__7_ : 
                      (N2941)? data_n_93__7_ : 
                      (N2943)? data_n_94__7_ : 
                      (N2945)? data_n_95__7_ : 
                      (N2947)? data_n_96__7_ : 
                      (N2949)? data_n_97__7_ : 
                      (N2951)? data_n_98__7_ : 
                      (N2953)? data_n_99__7_ : 
                      (N2955)? data_n_100__7_ : 
                      (N2957)? data_n_101__7_ : 
                      (N2959)? data_n_102__7_ : 
                      (N2961)? data_n_103__7_ : 
                      (N2963)? data_n_104__7_ : 
                      (N2965)? data_n_105__7_ : 
                      (N2967)? data_n_106__7_ : 
                      (N2969)? data_n_107__7_ : 
                      (N2971)? data_n_108__7_ : 
                      (N2973)? data_n_109__7_ : 
                      (N2975)? data_n_110__7_ : 
                      (N2977)? data_n_111__7_ : 
                      (N2979)? data_n_112__7_ : 
                      (N2981)? data_n_113__7_ : 
                      (N2983)? data_n_114__7_ : 
                      (N2985)? data_n_115__7_ : 
                      (N2987)? data_n_116__7_ : 
                      (N2989)? data_n_117__7_ : 
                      (N2991)? data_n_118__7_ : 
                      (N2993)? data_n_119__7_ : 
                      (N2995)? data_n_120__7_ : 
                      (N2997)? data_n_121__7_ : 
                      (N2999)? data_n_122__7_ : 
                      (N3001)? data_n_123__7_ : 
                      (N3003)? data_n_124__7_ : 
                      (N3005)? data_n_125__7_ : 
                      (N3007)? data_n_126__7_ : 
                      (N3009)? data_n_127__7_ : 1'b0;
  assign data_nn[6] = (N2882)? data_o[6] : 
                      (N2884)? data_o[38] : 
                      (N2886)? data_o[70] : 
                      (N2888)? data_o[102] : 
                      (N2890)? data_o[134] : 
                      (N2892)? data_o[166] : 
                      (N2894)? data_o[198] : 
                      (N2896)? data_o[230] : 
                      (N2898)? data_o[262] : 
                      (N2900)? data_o[294] : 
                      (N2902)? data_o[326] : 
                      (N2904)? data_o[358] : 
                      (N2906)? data_o[390] : 
                      (N2908)? data_o[422] : 
                      (N2910)? data_o[454] : 
                      (N2912)? data_o[486] : 
                      (N2914)? data_o[518] : 
                      (N2916)? data_o[550] : 
                      (N2918)? data_o[582] : 
                      (N2920)? data_o[614] : 
                      (N2922)? data_o[646] : 
                      (N2924)? data_o[678] : 
                      (N2926)? data_o[710] : 
                      (N2928)? data_o[742] : 
                      (N2930)? data_o[774] : 
                      (N2932)? data_o[806] : 
                      (N2934)? data_o[838] : 
                      (N2936)? data_o[870] : 
                      (N2938)? data_o[902] : 
                      (N2940)? data_o[934] : 
                      (N2942)? data_o[966] : 
                      (N2944)? data_o[998] : 
                      (N2946)? data_o[1030] : 
                      (N2948)? data_o[1062] : 
                      (N2950)? data_o[1094] : 
                      (N2952)? data_o[1126] : 
                      (N2954)? data_o[1158] : 
                      (N2956)? data_o[1190] : 
                      (N2958)? data_o[1222] : 
                      (N2960)? data_o[1254] : 
                      (N2962)? data_o[1286] : 
                      (N2964)? data_o[1318] : 
                      (N2966)? data_o[1350] : 
                      (N2968)? data_o[1382] : 
                      (N2970)? data_o[1414] : 
                      (N2972)? data_o[1446] : 
                      (N2974)? data_o[1478] : 
                      (N2976)? data_o[1510] : 
                      (N2978)? data_o[1542] : 
                      (N2980)? data_o[1574] : 
                      (N2982)? data_o[1606] : 
                      (N2984)? data_o[1638] : 
                      (N2986)? data_o[1670] : 
                      (N2988)? data_o[1702] : 
                      (N2990)? data_o[1734] : 
                      (N2992)? data_o[1766] : 
                      (N2994)? data_o[1798] : 
                      (N2996)? data_o[1830] : 
                      (N2998)? data_o[1862] : 
                      (N3000)? data_o[1894] : 
                      (N3002)? data_o[1926] : 
                      (N3004)? data_o[1958] : 
                      (N3006)? data_o[1990] : 
                      (N3008)? data_o[2022] : 
                      (N2883)? data_n_64__6_ : 
                      (N2885)? data_n_65__6_ : 
                      (N2887)? data_n_66__6_ : 
                      (N2889)? data_n_67__6_ : 
                      (N2891)? data_n_68__6_ : 
                      (N2893)? data_n_69__6_ : 
                      (N2895)? data_n_70__6_ : 
                      (N2897)? data_n_71__6_ : 
                      (N2899)? data_n_72__6_ : 
                      (N2901)? data_n_73__6_ : 
                      (N2903)? data_n_74__6_ : 
                      (N2905)? data_n_75__6_ : 
                      (N2907)? data_n_76__6_ : 
                      (N2909)? data_n_77__6_ : 
                      (N2911)? data_n_78__6_ : 
                      (N2913)? data_n_79__6_ : 
                      (N2915)? data_n_80__6_ : 
                      (N2917)? data_n_81__6_ : 
                      (N2919)? data_n_82__6_ : 
                      (N2921)? data_n_83__6_ : 
                      (N2923)? data_n_84__6_ : 
                      (N2925)? data_n_85__6_ : 
                      (N2927)? data_n_86__6_ : 
                      (N2929)? data_n_87__6_ : 
                      (N2931)? data_n_88__6_ : 
                      (N2933)? data_n_89__6_ : 
                      (N2935)? data_n_90__6_ : 
                      (N2937)? data_n_91__6_ : 
                      (N2939)? data_n_92__6_ : 
                      (N2941)? data_n_93__6_ : 
                      (N2943)? data_n_94__6_ : 
                      (N2945)? data_n_95__6_ : 
                      (N2947)? data_n_96__6_ : 
                      (N2949)? data_n_97__6_ : 
                      (N2951)? data_n_98__6_ : 
                      (N2953)? data_n_99__6_ : 
                      (N2955)? data_n_100__6_ : 
                      (N2957)? data_n_101__6_ : 
                      (N2959)? data_n_102__6_ : 
                      (N2961)? data_n_103__6_ : 
                      (N2963)? data_n_104__6_ : 
                      (N2965)? data_n_105__6_ : 
                      (N2967)? data_n_106__6_ : 
                      (N2969)? data_n_107__6_ : 
                      (N2971)? data_n_108__6_ : 
                      (N2973)? data_n_109__6_ : 
                      (N2975)? data_n_110__6_ : 
                      (N2977)? data_n_111__6_ : 
                      (N2979)? data_n_112__6_ : 
                      (N2981)? data_n_113__6_ : 
                      (N2983)? data_n_114__6_ : 
                      (N2985)? data_n_115__6_ : 
                      (N2987)? data_n_116__6_ : 
                      (N2989)? data_n_117__6_ : 
                      (N2991)? data_n_118__6_ : 
                      (N2993)? data_n_119__6_ : 
                      (N2995)? data_n_120__6_ : 
                      (N2997)? data_n_121__6_ : 
                      (N2999)? data_n_122__6_ : 
                      (N3001)? data_n_123__6_ : 
                      (N3003)? data_n_124__6_ : 
                      (N3005)? data_n_125__6_ : 
                      (N3007)? data_n_126__6_ : 
                      (N3009)? data_n_127__6_ : 1'b0;
  assign data_nn[5] = (N2882)? data_o[5] : 
                      (N2884)? data_o[37] : 
                      (N2886)? data_o[69] : 
                      (N2888)? data_o[101] : 
                      (N2890)? data_o[133] : 
                      (N2892)? data_o[165] : 
                      (N2894)? data_o[197] : 
                      (N2896)? data_o[229] : 
                      (N2898)? data_o[261] : 
                      (N2900)? data_o[293] : 
                      (N2902)? data_o[325] : 
                      (N2904)? data_o[357] : 
                      (N2906)? data_o[389] : 
                      (N2908)? data_o[421] : 
                      (N2910)? data_o[453] : 
                      (N2912)? data_o[485] : 
                      (N2914)? data_o[517] : 
                      (N2916)? data_o[549] : 
                      (N2918)? data_o[581] : 
                      (N2920)? data_o[613] : 
                      (N2922)? data_o[645] : 
                      (N2924)? data_o[677] : 
                      (N2926)? data_o[709] : 
                      (N2928)? data_o[741] : 
                      (N2930)? data_o[773] : 
                      (N2932)? data_o[805] : 
                      (N2934)? data_o[837] : 
                      (N2936)? data_o[869] : 
                      (N2938)? data_o[901] : 
                      (N2940)? data_o[933] : 
                      (N2942)? data_o[965] : 
                      (N2944)? data_o[997] : 
                      (N2946)? data_o[1029] : 
                      (N2948)? data_o[1061] : 
                      (N2950)? data_o[1093] : 
                      (N2952)? data_o[1125] : 
                      (N2954)? data_o[1157] : 
                      (N2956)? data_o[1189] : 
                      (N2958)? data_o[1221] : 
                      (N2960)? data_o[1253] : 
                      (N2962)? data_o[1285] : 
                      (N2964)? data_o[1317] : 
                      (N2966)? data_o[1349] : 
                      (N2968)? data_o[1381] : 
                      (N2970)? data_o[1413] : 
                      (N2972)? data_o[1445] : 
                      (N2974)? data_o[1477] : 
                      (N2976)? data_o[1509] : 
                      (N2978)? data_o[1541] : 
                      (N2980)? data_o[1573] : 
                      (N2982)? data_o[1605] : 
                      (N2984)? data_o[1637] : 
                      (N2986)? data_o[1669] : 
                      (N2988)? data_o[1701] : 
                      (N2990)? data_o[1733] : 
                      (N2992)? data_o[1765] : 
                      (N2994)? data_o[1797] : 
                      (N2996)? data_o[1829] : 
                      (N2998)? data_o[1861] : 
                      (N3000)? data_o[1893] : 
                      (N3002)? data_o[1925] : 
                      (N3004)? data_o[1957] : 
                      (N3006)? data_o[1989] : 
                      (N3008)? data_o[2021] : 
                      (N2883)? data_n_64__5_ : 
                      (N2885)? data_n_65__5_ : 
                      (N2887)? data_n_66__5_ : 
                      (N2889)? data_n_67__5_ : 
                      (N2891)? data_n_68__5_ : 
                      (N2893)? data_n_69__5_ : 
                      (N2895)? data_n_70__5_ : 
                      (N2897)? data_n_71__5_ : 
                      (N2899)? data_n_72__5_ : 
                      (N2901)? data_n_73__5_ : 
                      (N2903)? data_n_74__5_ : 
                      (N2905)? data_n_75__5_ : 
                      (N2907)? data_n_76__5_ : 
                      (N2909)? data_n_77__5_ : 
                      (N2911)? data_n_78__5_ : 
                      (N2913)? data_n_79__5_ : 
                      (N2915)? data_n_80__5_ : 
                      (N2917)? data_n_81__5_ : 
                      (N2919)? data_n_82__5_ : 
                      (N2921)? data_n_83__5_ : 
                      (N2923)? data_n_84__5_ : 
                      (N2925)? data_n_85__5_ : 
                      (N2927)? data_n_86__5_ : 
                      (N2929)? data_n_87__5_ : 
                      (N2931)? data_n_88__5_ : 
                      (N2933)? data_n_89__5_ : 
                      (N2935)? data_n_90__5_ : 
                      (N2937)? data_n_91__5_ : 
                      (N2939)? data_n_92__5_ : 
                      (N2941)? data_n_93__5_ : 
                      (N2943)? data_n_94__5_ : 
                      (N2945)? data_n_95__5_ : 
                      (N2947)? data_n_96__5_ : 
                      (N2949)? data_n_97__5_ : 
                      (N2951)? data_n_98__5_ : 
                      (N2953)? data_n_99__5_ : 
                      (N2955)? data_n_100__5_ : 
                      (N2957)? data_n_101__5_ : 
                      (N2959)? data_n_102__5_ : 
                      (N2961)? data_n_103__5_ : 
                      (N2963)? data_n_104__5_ : 
                      (N2965)? data_n_105__5_ : 
                      (N2967)? data_n_106__5_ : 
                      (N2969)? data_n_107__5_ : 
                      (N2971)? data_n_108__5_ : 
                      (N2973)? data_n_109__5_ : 
                      (N2975)? data_n_110__5_ : 
                      (N2977)? data_n_111__5_ : 
                      (N2979)? data_n_112__5_ : 
                      (N2981)? data_n_113__5_ : 
                      (N2983)? data_n_114__5_ : 
                      (N2985)? data_n_115__5_ : 
                      (N2987)? data_n_116__5_ : 
                      (N2989)? data_n_117__5_ : 
                      (N2991)? data_n_118__5_ : 
                      (N2993)? data_n_119__5_ : 
                      (N2995)? data_n_120__5_ : 
                      (N2997)? data_n_121__5_ : 
                      (N2999)? data_n_122__5_ : 
                      (N3001)? data_n_123__5_ : 
                      (N3003)? data_n_124__5_ : 
                      (N3005)? data_n_125__5_ : 
                      (N3007)? data_n_126__5_ : 
                      (N3009)? data_n_127__5_ : 1'b0;
  assign data_nn[4] = (N2882)? data_o[4] : 
                      (N2884)? data_o[36] : 
                      (N2886)? data_o[68] : 
                      (N2888)? data_o[100] : 
                      (N2890)? data_o[132] : 
                      (N2892)? data_o[164] : 
                      (N2894)? data_o[196] : 
                      (N2896)? data_o[228] : 
                      (N2898)? data_o[260] : 
                      (N2900)? data_o[292] : 
                      (N2902)? data_o[324] : 
                      (N2904)? data_o[356] : 
                      (N2906)? data_o[388] : 
                      (N2908)? data_o[420] : 
                      (N2910)? data_o[452] : 
                      (N2912)? data_o[484] : 
                      (N2914)? data_o[516] : 
                      (N2916)? data_o[548] : 
                      (N2918)? data_o[580] : 
                      (N2920)? data_o[612] : 
                      (N2922)? data_o[644] : 
                      (N2924)? data_o[676] : 
                      (N2926)? data_o[708] : 
                      (N2928)? data_o[740] : 
                      (N2930)? data_o[772] : 
                      (N2932)? data_o[804] : 
                      (N2934)? data_o[836] : 
                      (N2936)? data_o[868] : 
                      (N2938)? data_o[900] : 
                      (N2940)? data_o[932] : 
                      (N2942)? data_o[964] : 
                      (N2944)? data_o[996] : 
                      (N2946)? data_o[1028] : 
                      (N2948)? data_o[1060] : 
                      (N2950)? data_o[1092] : 
                      (N2952)? data_o[1124] : 
                      (N2954)? data_o[1156] : 
                      (N2956)? data_o[1188] : 
                      (N2958)? data_o[1220] : 
                      (N2960)? data_o[1252] : 
                      (N2962)? data_o[1284] : 
                      (N2964)? data_o[1316] : 
                      (N2966)? data_o[1348] : 
                      (N2968)? data_o[1380] : 
                      (N2970)? data_o[1412] : 
                      (N2972)? data_o[1444] : 
                      (N2974)? data_o[1476] : 
                      (N2976)? data_o[1508] : 
                      (N2978)? data_o[1540] : 
                      (N2980)? data_o[1572] : 
                      (N2982)? data_o[1604] : 
                      (N2984)? data_o[1636] : 
                      (N2986)? data_o[1668] : 
                      (N2988)? data_o[1700] : 
                      (N2990)? data_o[1732] : 
                      (N2992)? data_o[1764] : 
                      (N2994)? data_o[1796] : 
                      (N2996)? data_o[1828] : 
                      (N2998)? data_o[1860] : 
                      (N3000)? data_o[1892] : 
                      (N3002)? data_o[1924] : 
                      (N3004)? data_o[1956] : 
                      (N3006)? data_o[1988] : 
                      (N3008)? data_o[2020] : 
                      (N2883)? data_n_64__4_ : 
                      (N2885)? data_n_65__4_ : 
                      (N2887)? data_n_66__4_ : 
                      (N2889)? data_n_67__4_ : 
                      (N2891)? data_n_68__4_ : 
                      (N2893)? data_n_69__4_ : 
                      (N2895)? data_n_70__4_ : 
                      (N2897)? data_n_71__4_ : 
                      (N2899)? data_n_72__4_ : 
                      (N2901)? data_n_73__4_ : 
                      (N2903)? data_n_74__4_ : 
                      (N2905)? data_n_75__4_ : 
                      (N2907)? data_n_76__4_ : 
                      (N2909)? data_n_77__4_ : 
                      (N2911)? data_n_78__4_ : 
                      (N2913)? data_n_79__4_ : 
                      (N2915)? data_n_80__4_ : 
                      (N2917)? data_n_81__4_ : 
                      (N2919)? data_n_82__4_ : 
                      (N2921)? data_n_83__4_ : 
                      (N2923)? data_n_84__4_ : 
                      (N2925)? data_n_85__4_ : 
                      (N2927)? data_n_86__4_ : 
                      (N2929)? data_n_87__4_ : 
                      (N2931)? data_n_88__4_ : 
                      (N2933)? data_n_89__4_ : 
                      (N2935)? data_n_90__4_ : 
                      (N2937)? data_n_91__4_ : 
                      (N2939)? data_n_92__4_ : 
                      (N2941)? data_n_93__4_ : 
                      (N2943)? data_n_94__4_ : 
                      (N2945)? data_n_95__4_ : 
                      (N2947)? data_n_96__4_ : 
                      (N2949)? data_n_97__4_ : 
                      (N2951)? data_n_98__4_ : 
                      (N2953)? data_n_99__4_ : 
                      (N2955)? data_n_100__4_ : 
                      (N2957)? data_n_101__4_ : 
                      (N2959)? data_n_102__4_ : 
                      (N2961)? data_n_103__4_ : 
                      (N2963)? data_n_104__4_ : 
                      (N2965)? data_n_105__4_ : 
                      (N2967)? data_n_106__4_ : 
                      (N2969)? data_n_107__4_ : 
                      (N2971)? data_n_108__4_ : 
                      (N2973)? data_n_109__4_ : 
                      (N2975)? data_n_110__4_ : 
                      (N2977)? data_n_111__4_ : 
                      (N2979)? data_n_112__4_ : 
                      (N2981)? data_n_113__4_ : 
                      (N2983)? data_n_114__4_ : 
                      (N2985)? data_n_115__4_ : 
                      (N2987)? data_n_116__4_ : 
                      (N2989)? data_n_117__4_ : 
                      (N2991)? data_n_118__4_ : 
                      (N2993)? data_n_119__4_ : 
                      (N2995)? data_n_120__4_ : 
                      (N2997)? data_n_121__4_ : 
                      (N2999)? data_n_122__4_ : 
                      (N3001)? data_n_123__4_ : 
                      (N3003)? data_n_124__4_ : 
                      (N3005)? data_n_125__4_ : 
                      (N3007)? data_n_126__4_ : 
                      (N3009)? data_n_127__4_ : 1'b0;
  assign data_nn[3] = (N2882)? data_o[3] : 
                      (N2884)? data_o[35] : 
                      (N2886)? data_o[67] : 
                      (N2888)? data_o[99] : 
                      (N2890)? data_o[131] : 
                      (N2892)? data_o[163] : 
                      (N2894)? data_o[195] : 
                      (N2896)? data_o[227] : 
                      (N2898)? data_o[259] : 
                      (N2900)? data_o[291] : 
                      (N2902)? data_o[323] : 
                      (N2904)? data_o[355] : 
                      (N2906)? data_o[387] : 
                      (N2908)? data_o[419] : 
                      (N2910)? data_o[451] : 
                      (N2912)? data_o[483] : 
                      (N2914)? data_o[515] : 
                      (N2916)? data_o[547] : 
                      (N2918)? data_o[579] : 
                      (N2920)? data_o[611] : 
                      (N2922)? data_o[643] : 
                      (N2924)? data_o[675] : 
                      (N2926)? data_o[707] : 
                      (N2928)? data_o[739] : 
                      (N2930)? data_o[771] : 
                      (N2932)? data_o[803] : 
                      (N2934)? data_o[835] : 
                      (N2936)? data_o[867] : 
                      (N2938)? data_o[899] : 
                      (N2940)? data_o[931] : 
                      (N2942)? data_o[963] : 
                      (N2944)? data_o[995] : 
                      (N2946)? data_o[1027] : 
                      (N2948)? data_o[1059] : 
                      (N2950)? data_o[1091] : 
                      (N2952)? data_o[1123] : 
                      (N2954)? data_o[1155] : 
                      (N2956)? data_o[1187] : 
                      (N2958)? data_o[1219] : 
                      (N2960)? data_o[1251] : 
                      (N2962)? data_o[1283] : 
                      (N2964)? data_o[1315] : 
                      (N2966)? data_o[1347] : 
                      (N2968)? data_o[1379] : 
                      (N2970)? data_o[1411] : 
                      (N2972)? data_o[1443] : 
                      (N2974)? data_o[1475] : 
                      (N2976)? data_o[1507] : 
                      (N2978)? data_o[1539] : 
                      (N2980)? data_o[1571] : 
                      (N2982)? data_o[1603] : 
                      (N2984)? data_o[1635] : 
                      (N2986)? data_o[1667] : 
                      (N2988)? data_o[1699] : 
                      (N2990)? data_o[1731] : 
                      (N2992)? data_o[1763] : 
                      (N2994)? data_o[1795] : 
                      (N2996)? data_o[1827] : 
                      (N2998)? data_o[1859] : 
                      (N3000)? data_o[1891] : 
                      (N3002)? data_o[1923] : 
                      (N3004)? data_o[1955] : 
                      (N3006)? data_o[1987] : 
                      (N3008)? data_o[2019] : 
                      (N2883)? data_n_64__3_ : 
                      (N2885)? data_n_65__3_ : 
                      (N2887)? data_n_66__3_ : 
                      (N2889)? data_n_67__3_ : 
                      (N2891)? data_n_68__3_ : 
                      (N2893)? data_n_69__3_ : 
                      (N2895)? data_n_70__3_ : 
                      (N2897)? data_n_71__3_ : 
                      (N2899)? data_n_72__3_ : 
                      (N2901)? data_n_73__3_ : 
                      (N2903)? data_n_74__3_ : 
                      (N2905)? data_n_75__3_ : 
                      (N2907)? data_n_76__3_ : 
                      (N2909)? data_n_77__3_ : 
                      (N2911)? data_n_78__3_ : 
                      (N2913)? data_n_79__3_ : 
                      (N2915)? data_n_80__3_ : 
                      (N2917)? data_n_81__3_ : 
                      (N2919)? data_n_82__3_ : 
                      (N2921)? data_n_83__3_ : 
                      (N2923)? data_n_84__3_ : 
                      (N2925)? data_n_85__3_ : 
                      (N2927)? data_n_86__3_ : 
                      (N2929)? data_n_87__3_ : 
                      (N2931)? data_n_88__3_ : 
                      (N2933)? data_n_89__3_ : 
                      (N2935)? data_n_90__3_ : 
                      (N2937)? data_n_91__3_ : 
                      (N2939)? data_n_92__3_ : 
                      (N2941)? data_n_93__3_ : 
                      (N2943)? data_n_94__3_ : 
                      (N2945)? data_n_95__3_ : 
                      (N2947)? data_n_96__3_ : 
                      (N2949)? data_n_97__3_ : 
                      (N2951)? data_n_98__3_ : 
                      (N2953)? data_n_99__3_ : 
                      (N2955)? data_n_100__3_ : 
                      (N2957)? data_n_101__3_ : 
                      (N2959)? data_n_102__3_ : 
                      (N2961)? data_n_103__3_ : 
                      (N2963)? data_n_104__3_ : 
                      (N2965)? data_n_105__3_ : 
                      (N2967)? data_n_106__3_ : 
                      (N2969)? data_n_107__3_ : 
                      (N2971)? data_n_108__3_ : 
                      (N2973)? data_n_109__3_ : 
                      (N2975)? data_n_110__3_ : 
                      (N2977)? data_n_111__3_ : 
                      (N2979)? data_n_112__3_ : 
                      (N2981)? data_n_113__3_ : 
                      (N2983)? data_n_114__3_ : 
                      (N2985)? data_n_115__3_ : 
                      (N2987)? data_n_116__3_ : 
                      (N2989)? data_n_117__3_ : 
                      (N2991)? data_n_118__3_ : 
                      (N2993)? data_n_119__3_ : 
                      (N2995)? data_n_120__3_ : 
                      (N2997)? data_n_121__3_ : 
                      (N2999)? data_n_122__3_ : 
                      (N3001)? data_n_123__3_ : 
                      (N3003)? data_n_124__3_ : 
                      (N3005)? data_n_125__3_ : 
                      (N3007)? data_n_126__3_ : 
                      (N3009)? data_n_127__3_ : 1'b0;
  assign data_nn[2] = (N2882)? data_o[2] : 
                      (N2884)? data_o[34] : 
                      (N2886)? data_o[66] : 
                      (N2888)? data_o[98] : 
                      (N2890)? data_o[130] : 
                      (N2892)? data_o[162] : 
                      (N2894)? data_o[194] : 
                      (N2896)? data_o[226] : 
                      (N2898)? data_o[258] : 
                      (N2900)? data_o[290] : 
                      (N2902)? data_o[322] : 
                      (N2904)? data_o[354] : 
                      (N2906)? data_o[386] : 
                      (N2908)? data_o[418] : 
                      (N2910)? data_o[450] : 
                      (N2912)? data_o[482] : 
                      (N2914)? data_o[514] : 
                      (N2916)? data_o[546] : 
                      (N2918)? data_o[578] : 
                      (N2920)? data_o[610] : 
                      (N2922)? data_o[642] : 
                      (N2924)? data_o[674] : 
                      (N2926)? data_o[706] : 
                      (N2928)? data_o[738] : 
                      (N2930)? data_o[770] : 
                      (N2932)? data_o[802] : 
                      (N2934)? data_o[834] : 
                      (N2936)? data_o[866] : 
                      (N2938)? data_o[898] : 
                      (N2940)? data_o[930] : 
                      (N2942)? data_o[962] : 
                      (N2944)? data_o[994] : 
                      (N2946)? data_o[1026] : 
                      (N2948)? data_o[1058] : 
                      (N2950)? data_o[1090] : 
                      (N2952)? data_o[1122] : 
                      (N2954)? data_o[1154] : 
                      (N2956)? data_o[1186] : 
                      (N2958)? data_o[1218] : 
                      (N2960)? data_o[1250] : 
                      (N2962)? data_o[1282] : 
                      (N2964)? data_o[1314] : 
                      (N2966)? data_o[1346] : 
                      (N2968)? data_o[1378] : 
                      (N2970)? data_o[1410] : 
                      (N2972)? data_o[1442] : 
                      (N2974)? data_o[1474] : 
                      (N2976)? data_o[1506] : 
                      (N2978)? data_o[1538] : 
                      (N2980)? data_o[1570] : 
                      (N2982)? data_o[1602] : 
                      (N2984)? data_o[1634] : 
                      (N2986)? data_o[1666] : 
                      (N2988)? data_o[1698] : 
                      (N2990)? data_o[1730] : 
                      (N2992)? data_o[1762] : 
                      (N2994)? data_o[1794] : 
                      (N2996)? data_o[1826] : 
                      (N2998)? data_o[1858] : 
                      (N3000)? data_o[1890] : 
                      (N3002)? data_o[1922] : 
                      (N3004)? data_o[1954] : 
                      (N3006)? data_o[1986] : 
                      (N3008)? data_o[2018] : 
                      (N2883)? data_n_64__2_ : 
                      (N2885)? data_n_65__2_ : 
                      (N2887)? data_n_66__2_ : 
                      (N2889)? data_n_67__2_ : 
                      (N2891)? data_n_68__2_ : 
                      (N2893)? data_n_69__2_ : 
                      (N2895)? data_n_70__2_ : 
                      (N2897)? data_n_71__2_ : 
                      (N2899)? data_n_72__2_ : 
                      (N2901)? data_n_73__2_ : 
                      (N2903)? data_n_74__2_ : 
                      (N2905)? data_n_75__2_ : 
                      (N2907)? data_n_76__2_ : 
                      (N2909)? data_n_77__2_ : 
                      (N2911)? data_n_78__2_ : 
                      (N2913)? data_n_79__2_ : 
                      (N2915)? data_n_80__2_ : 
                      (N2917)? data_n_81__2_ : 
                      (N2919)? data_n_82__2_ : 
                      (N2921)? data_n_83__2_ : 
                      (N2923)? data_n_84__2_ : 
                      (N2925)? data_n_85__2_ : 
                      (N2927)? data_n_86__2_ : 
                      (N2929)? data_n_87__2_ : 
                      (N2931)? data_n_88__2_ : 
                      (N2933)? data_n_89__2_ : 
                      (N2935)? data_n_90__2_ : 
                      (N2937)? data_n_91__2_ : 
                      (N2939)? data_n_92__2_ : 
                      (N2941)? data_n_93__2_ : 
                      (N2943)? data_n_94__2_ : 
                      (N2945)? data_n_95__2_ : 
                      (N2947)? data_n_96__2_ : 
                      (N2949)? data_n_97__2_ : 
                      (N2951)? data_n_98__2_ : 
                      (N2953)? data_n_99__2_ : 
                      (N2955)? data_n_100__2_ : 
                      (N2957)? data_n_101__2_ : 
                      (N2959)? data_n_102__2_ : 
                      (N2961)? data_n_103__2_ : 
                      (N2963)? data_n_104__2_ : 
                      (N2965)? data_n_105__2_ : 
                      (N2967)? data_n_106__2_ : 
                      (N2969)? data_n_107__2_ : 
                      (N2971)? data_n_108__2_ : 
                      (N2973)? data_n_109__2_ : 
                      (N2975)? data_n_110__2_ : 
                      (N2977)? data_n_111__2_ : 
                      (N2979)? data_n_112__2_ : 
                      (N2981)? data_n_113__2_ : 
                      (N2983)? data_n_114__2_ : 
                      (N2985)? data_n_115__2_ : 
                      (N2987)? data_n_116__2_ : 
                      (N2989)? data_n_117__2_ : 
                      (N2991)? data_n_118__2_ : 
                      (N2993)? data_n_119__2_ : 
                      (N2995)? data_n_120__2_ : 
                      (N2997)? data_n_121__2_ : 
                      (N2999)? data_n_122__2_ : 
                      (N3001)? data_n_123__2_ : 
                      (N3003)? data_n_124__2_ : 
                      (N3005)? data_n_125__2_ : 
                      (N3007)? data_n_126__2_ : 
                      (N3009)? data_n_127__2_ : 1'b0;
  assign data_nn[1] = (N2882)? data_o[1] : 
                      (N2884)? data_o[33] : 
                      (N2886)? data_o[65] : 
                      (N2888)? data_o[97] : 
                      (N2890)? data_o[129] : 
                      (N2892)? data_o[161] : 
                      (N2894)? data_o[193] : 
                      (N2896)? data_o[225] : 
                      (N2898)? data_o[257] : 
                      (N2900)? data_o[289] : 
                      (N2902)? data_o[321] : 
                      (N2904)? data_o[353] : 
                      (N2906)? data_o[385] : 
                      (N2908)? data_o[417] : 
                      (N2910)? data_o[449] : 
                      (N2912)? data_o[481] : 
                      (N2914)? data_o[513] : 
                      (N2916)? data_o[545] : 
                      (N2918)? data_o[577] : 
                      (N2920)? data_o[609] : 
                      (N2922)? data_o[641] : 
                      (N2924)? data_o[673] : 
                      (N2926)? data_o[705] : 
                      (N2928)? data_o[737] : 
                      (N2930)? data_o[769] : 
                      (N2932)? data_o[801] : 
                      (N2934)? data_o[833] : 
                      (N2936)? data_o[865] : 
                      (N2938)? data_o[897] : 
                      (N2940)? data_o[929] : 
                      (N2942)? data_o[961] : 
                      (N2944)? data_o[993] : 
                      (N2946)? data_o[1025] : 
                      (N2948)? data_o[1057] : 
                      (N2950)? data_o[1089] : 
                      (N2952)? data_o[1121] : 
                      (N2954)? data_o[1153] : 
                      (N2956)? data_o[1185] : 
                      (N2958)? data_o[1217] : 
                      (N2960)? data_o[1249] : 
                      (N2962)? data_o[1281] : 
                      (N2964)? data_o[1313] : 
                      (N2966)? data_o[1345] : 
                      (N2968)? data_o[1377] : 
                      (N2970)? data_o[1409] : 
                      (N2972)? data_o[1441] : 
                      (N2974)? data_o[1473] : 
                      (N2976)? data_o[1505] : 
                      (N2978)? data_o[1537] : 
                      (N2980)? data_o[1569] : 
                      (N2982)? data_o[1601] : 
                      (N2984)? data_o[1633] : 
                      (N2986)? data_o[1665] : 
                      (N2988)? data_o[1697] : 
                      (N2990)? data_o[1729] : 
                      (N2992)? data_o[1761] : 
                      (N2994)? data_o[1793] : 
                      (N2996)? data_o[1825] : 
                      (N2998)? data_o[1857] : 
                      (N3000)? data_o[1889] : 
                      (N3002)? data_o[1921] : 
                      (N3004)? data_o[1953] : 
                      (N3006)? data_o[1985] : 
                      (N3008)? data_o[2017] : 
                      (N2883)? data_n_64__1_ : 
                      (N2885)? data_n_65__1_ : 
                      (N2887)? data_n_66__1_ : 
                      (N2889)? data_n_67__1_ : 
                      (N2891)? data_n_68__1_ : 
                      (N2893)? data_n_69__1_ : 
                      (N2895)? data_n_70__1_ : 
                      (N2897)? data_n_71__1_ : 
                      (N2899)? data_n_72__1_ : 
                      (N2901)? data_n_73__1_ : 
                      (N2903)? data_n_74__1_ : 
                      (N2905)? data_n_75__1_ : 
                      (N2907)? data_n_76__1_ : 
                      (N2909)? data_n_77__1_ : 
                      (N2911)? data_n_78__1_ : 
                      (N2913)? data_n_79__1_ : 
                      (N2915)? data_n_80__1_ : 
                      (N2917)? data_n_81__1_ : 
                      (N2919)? data_n_82__1_ : 
                      (N2921)? data_n_83__1_ : 
                      (N2923)? data_n_84__1_ : 
                      (N2925)? data_n_85__1_ : 
                      (N2927)? data_n_86__1_ : 
                      (N2929)? data_n_87__1_ : 
                      (N2931)? data_n_88__1_ : 
                      (N2933)? data_n_89__1_ : 
                      (N2935)? data_n_90__1_ : 
                      (N2937)? data_n_91__1_ : 
                      (N2939)? data_n_92__1_ : 
                      (N2941)? data_n_93__1_ : 
                      (N2943)? data_n_94__1_ : 
                      (N2945)? data_n_95__1_ : 
                      (N2947)? data_n_96__1_ : 
                      (N2949)? data_n_97__1_ : 
                      (N2951)? data_n_98__1_ : 
                      (N2953)? data_n_99__1_ : 
                      (N2955)? data_n_100__1_ : 
                      (N2957)? data_n_101__1_ : 
                      (N2959)? data_n_102__1_ : 
                      (N2961)? data_n_103__1_ : 
                      (N2963)? data_n_104__1_ : 
                      (N2965)? data_n_105__1_ : 
                      (N2967)? data_n_106__1_ : 
                      (N2969)? data_n_107__1_ : 
                      (N2971)? data_n_108__1_ : 
                      (N2973)? data_n_109__1_ : 
                      (N2975)? data_n_110__1_ : 
                      (N2977)? data_n_111__1_ : 
                      (N2979)? data_n_112__1_ : 
                      (N2981)? data_n_113__1_ : 
                      (N2983)? data_n_114__1_ : 
                      (N2985)? data_n_115__1_ : 
                      (N2987)? data_n_116__1_ : 
                      (N2989)? data_n_117__1_ : 
                      (N2991)? data_n_118__1_ : 
                      (N2993)? data_n_119__1_ : 
                      (N2995)? data_n_120__1_ : 
                      (N2997)? data_n_121__1_ : 
                      (N2999)? data_n_122__1_ : 
                      (N3001)? data_n_123__1_ : 
                      (N3003)? data_n_124__1_ : 
                      (N3005)? data_n_125__1_ : 
                      (N3007)? data_n_126__1_ : 
                      (N3009)? data_n_127__1_ : 1'b0;
  assign data_nn[0] = (N2882)? data_o[0] : 
                      (N2884)? data_o[32] : 
                      (N2886)? data_o[64] : 
                      (N2888)? data_o[96] : 
                      (N2890)? data_o[128] : 
                      (N2892)? data_o[160] : 
                      (N2894)? data_o[192] : 
                      (N2896)? data_o[224] : 
                      (N2898)? data_o[256] : 
                      (N2900)? data_o[288] : 
                      (N2902)? data_o[320] : 
                      (N2904)? data_o[352] : 
                      (N2906)? data_o[384] : 
                      (N2908)? data_o[416] : 
                      (N2910)? data_o[448] : 
                      (N2912)? data_o[480] : 
                      (N2914)? data_o[512] : 
                      (N2916)? data_o[544] : 
                      (N2918)? data_o[576] : 
                      (N2920)? data_o[608] : 
                      (N2922)? data_o[640] : 
                      (N2924)? data_o[672] : 
                      (N2926)? data_o[704] : 
                      (N2928)? data_o[736] : 
                      (N2930)? data_o[768] : 
                      (N2932)? data_o[800] : 
                      (N2934)? data_o[832] : 
                      (N2936)? data_o[864] : 
                      (N2938)? data_o[896] : 
                      (N2940)? data_o[928] : 
                      (N2942)? data_o[960] : 
                      (N2944)? data_o[992] : 
                      (N2946)? data_o[1024] : 
                      (N2948)? data_o[1056] : 
                      (N2950)? data_o[1088] : 
                      (N2952)? data_o[1120] : 
                      (N2954)? data_o[1152] : 
                      (N2956)? data_o[1184] : 
                      (N2958)? data_o[1216] : 
                      (N2960)? data_o[1248] : 
                      (N2962)? data_o[1280] : 
                      (N2964)? data_o[1312] : 
                      (N2966)? data_o[1344] : 
                      (N2968)? data_o[1376] : 
                      (N2970)? data_o[1408] : 
                      (N2972)? data_o[1440] : 
                      (N2974)? data_o[1472] : 
                      (N2976)? data_o[1504] : 
                      (N2978)? data_o[1536] : 
                      (N2980)? data_o[1568] : 
                      (N2982)? data_o[1600] : 
                      (N2984)? data_o[1632] : 
                      (N2986)? data_o[1664] : 
                      (N2988)? data_o[1696] : 
                      (N2990)? data_o[1728] : 
                      (N2992)? data_o[1760] : 
                      (N2994)? data_o[1792] : 
                      (N2996)? data_o[1824] : 
                      (N2998)? data_o[1856] : 
                      (N3000)? data_o[1888] : 
                      (N3002)? data_o[1920] : 
                      (N3004)? data_o[1952] : 
                      (N3006)? data_o[1984] : 
                      (N3008)? data_o[2016] : 
                      (N2883)? data_n_64__0_ : 
                      (N2885)? data_n_65__0_ : 
                      (N2887)? data_n_66__0_ : 
                      (N2889)? data_n_67__0_ : 
                      (N2891)? data_n_68__0_ : 
                      (N2893)? data_n_69__0_ : 
                      (N2895)? data_n_70__0_ : 
                      (N2897)? data_n_71__0_ : 
                      (N2899)? data_n_72__0_ : 
                      (N2901)? data_n_73__0_ : 
                      (N2903)? data_n_74__0_ : 
                      (N2905)? data_n_75__0_ : 
                      (N2907)? data_n_76__0_ : 
                      (N2909)? data_n_77__0_ : 
                      (N2911)? data_n_78__0_ : 
                      (N2913)? data_n_79__0_ : 
                      (N2915)? data_n_80__0_ : 
                      (N2917)? data_n_81__0_ : 
                      (N2919)? data_n_82__0_ : 
                      (N2921)? data_n_83__0_ : 
                      (N2923)? data_n_84__0_ : 
                      (N2925)? data_n_85__0_ : 
                      (N2927)? data_n_86__0_ : 
                      (N2929)? data_n_87__0_ : 
                      (N2931)? data_n_88__0_ : 
                      (N2933)? data_n_89__0_ : 
                      (N2935)? data_n_90__0_ : 
                      (N2937)? data_n_91__0_ : 
                      (N2939)? data_n_92__0_ : 
                      (N2941)? data_n_93__0_ : 
                      (N2943)? data_n_94__0_ : 
                      (N2945)? data_n_95__0_ : 
                      (N2947)? data_n_96__0_ : 
                      (N2949)? data_n_97__0_ : 
                      (N2951)? data_n_98__0_ : 
                      (N2953)? data_n_99__0_ : 
                      (N2955)? data_n_100__0_ : 
                      (N2957)? data_n_101__0_ : 
                      (N2959)? data_n_102__0_ : 
                      (N2961)? data_n_103__0_ : 
                      (N2963)? data_n_104__0_ : 
                      (N2965)? data_n_105__0_ : 
                      (N2967)? data_n_106__0_ : 
                      (N2969)? data_n_107__0_ : 
                      (N2971)? data_n_108__0_ : 
                      (N2973)? data_n_109__0_ : 
                      (N2975)? data_n_110__0_ : 
                      (N2977)? data_n_111__0_ : 
                      (N2979)? data_n_112__0_ : 
                      (N2981)? data_n_113__0_ : 
                      (N2983)? data_n_114__0_ : 
                      (N2985)? data_n_115__0_ : 
                      (N2987)? data_n_116__0_ : 
                      (N2989)? data_n_117__0_ : 
                      (N2991)? data_n_118__0_ : 
                      (N2993)? data_n_119__0_ : 
                      (N2995)? data_n_120__0_ : 
                      (N2997)? data_n_121__0_ : 
                      (N2999)? data_n_122__0_ : 
                      (N3001)? data_n_123__0_ : 
                      (N3003)? data_n_124__0_ : 
                      (N3005)? data_n_125__0_ : 
                      (N3007)? data_n_126__0_ : 
                      (N3009)? data_n_127__0_ : 1'b0;
  assign { N2237, N2236, N2235, N2234, N2233, N2232, N2231 } = num_els_r + N2230;
  assign num_els_n = { N2237, N2236, N2235, N2234, N2233, N2232, N2231 } - yumi_cnt_i;
  assign N5376 = ~num_els_r[6];
  assign N5377 = num_els_r[4] & num_els_r[5];
  assign N5378 = N0 & num_els_r[5];
  assign N0 = ~num_els_r[4];
  assign N5379 = num_els_r[4] & N1;
  assign N1 = ~num_els_r[5];
  assign N5380 = N2 & N3;
  assign N2 = ~num_els_r[4];
  assign N3 = ~num_els_r[5];
  assign N5381 = num_els_r[6] & N5377;
  assign N5382 = num_els_r[6] & N5378;
  assign N5383 = num_els_r[6] & N5379;
  assign N5384 = num_els_r[6] & N5380;
  assign N5385 = N5376 & N5377;
  assign N5386 = N5376 & N5378;
  assign N5387 = N5376 & N5379;
  assign N5388 = N5376 & N5380;
  assign N5389 = num_els_r[2] & num_els_r[3];
  assign N5390 = N4 & num_els_r[3];
  assign N4 = ~num_els_r[2];
  assign N5391 = num_els_r[2] & N5;
  assign N5 = ~num_els_r[3];
  assign N5392 = N6 & N7;
  assign N6 = ~num_els_r[2];
  assign N7 = ~num_els_r[3];
  assign N5393 = num_els_r[0] & num_els_r[1];
  assign N5394 = N8 & num_els_r[1];
  assign N8 = ~num_els_r[0];
  assign N5395 = num_els_r[0] & N9;
  assign N9 = ~num_els_r[1];
  assign N5396 = N10 & N11;
  assign N10 = ~num_els_r[0];
  assign N11 = ~num_els_r[1];
  assign N5397 = N5389 & N5393;
  assign N5398 = N5389 & N5394;
  assign N5399 = N5389 & N5395;
  assign N5400 = N5389 & N5396;
  assign N5401 = N5390 & N5393;
  assign N5402 = N5390 & N5394;
  assign N5403 = N5390 & N5395;
  assign N5404 = N5390 & N5396;
  assign N5405 = N5391 & N5393;
  assign N5406 = N5391 & N5394;
  assign N5407 = N5391 & N5395;
  assign N5408 = N5391 & N5396;
  assign N5409 = N5392 & N5393;
  assign N5410 = N5392 & N5394;
  assign N5411 = N5392 & N5395;
  assign N5412 = N5392 & N5396;
  assign N2365 = N5381 & N5397;
  assign N2364 = N5381 & N5398;
  assign N2363 = N5381 & N5399;
  assign N2362 = N5381 & N5400;
  assign N2361 = N5381 & N5401;
  assign N2360 = N5381 & N5402;
  assign N2359 = N5381 & N5403;
  assign N2358 = N5381 & N5404;
  assign N2357 = N5381 & N5405;
  assign N2356 = N5381 & N5406;
  assign N2355 = N5381 & N5407;
  assign N2354 = N5381 & N5408;
  assign N2353 = N5381 & N5409;
  assign N2352 = N5381 & N5410;
  assign N2351 = N5381 & N5411;
  assign N2350 = N5381 & N5412;
  assign N2349 = N5382 & N5397;
  assign N2348 = N5382 & N5398;
  assign N2347 = N5382 & N5399;
  assign N2346 = N5382 & N5400;
  assign N2345 = N5382 & N5401;
  assign N2344 = N5382 & N5402;
  assign N2343 = N5382 & N5403;
  assign N2342 = N5382 & N5404;
  assign N2341 = N5382 & N5405;
  assign N2340 = N5382 & N5406;
  assign N2339 = N5382 & N5407;
  assign N2338 = N5382 & N5408;
  assign N2337 = N5382 & N5409;
  assign N2336 = N5382 & N5410;
  assign N2335 = N5382 & N5411;
  assign N2334 = N5382 & N5412;
  assign N2333 = N5383 & N5397;
  assign N2332 = N5383 & N5398;
  assign N2331 = N5383 & N5399;
  assign N2330 = N5383 & N5400;
  assign N2329 = N5383 & N5401;
  assign N2328 = N5383 & N5402;
  assign N2327 = N5383 & N5403;
  assign N2326 = N5383 & N5404;
  assign N2325 = N5383 & N5405;
  assign N2324 = N5383 & N5406;
  assign N2323 = N5383 & N5407;
  assign N2322 = N5383 & N5408;
  assign N2321 = N5383 & N5409;
  assign N2320 = N5383 & N5410;
  assign N2319 = N5383 & N5411;
  assign N2318 = N5383 & N5412;
  assign N2317 = N5384 & N5397;
  assign N2316 = N5384 & N5398;
  assign N2315 = N5384 & N5399;
  assign N2314 = N5384 & N5400;
  assign N2313 = N5384 & N5401;
  assign N2312 = N5384 & N5402;
  assign N2311 = N5384 & N5403;
  assign N2310 = N5384 & N5404;
  assign N2309 = N5384 & N5405;
  assign N2308 = N5384 & N5406;
  assign N2307 = N5384 & N5407;
  assign N2306 = N5384 & N5408;
  assign N2305 = N5384 & N5409;
  assign N2304 = N5384 & N5410;
  assign N2303 = N5384 & N5411;
  assign N2302 = N5384 & N5412;
  assign N2301 = N5385 & N5397;
  assign N2300 = N5385 & N5398;
  assign N2299 = N5385 & N5399;
  assign N2298 = N5385 & N5400;
  assign N2297 = N5385 & N5401;
  assign N2296 = N5385 & N5402;
  assign N2295 = N5385 & N5403;
  assign N2294 = N5385 & N5404;
  assign N2293 = N5385 & N5405;
  assign N2292 = N5385 & N5406;
  assign N2291 = N5385 & N5407;
  assign N2290 = N5385 & N5408;
  assign N2289 = N5385 & N5409;
  assign N2288 = N5385 & N5410;
  assign N2287 = N5385 & N5411;
  assign N2286 = N5385 & N5412;
  assign N2285 = N5386 & N5397;
  assign N2284 = N5386 & N5398;
  assign N2283 = N5386 & N5399;
  assign N2282 = N5386 & N5400;
  assign N2281 = N5386 & N5401;
  assign N2280 = N5386 & N5402;
  assign N2279 = N5386 & N5403;
  assign N2278 = N5386 & N5404;
  assign N2277 = N5386 & N5405;
  assign N2276 = N5386 & N5406;
  assign N2275 = N5386 & N5407;
  assign N2274 = N5386 & N5408;
  assign N2273 = N5386 & N5409;
  assign N2272 = N5386 & N5410;
  assign N2271 = N5386 & N5411;
  assign N2270 = N5386 & N5412;
  assign N2269 = N5387 & N5397;
  assign N2268 = N5387 & N5398;
  assign N2267 = N5387 & N5399;
  assign N2266 = N5387 & N5400;
  assign N2265 = N5387 & N5401;
  assign N2264 = N5387 & N5402;
  assign N2263 = N5387 & N5403;
  assign N2262 = N5387 & N5404;
  assign N2261 = N5387 & N5405;
  assign N2260 = N5387 & N5406;
  assign N2259 = N5387 & N5407;
  assign N2258 = N5387 & N5408;
  assign N2257 = N5387 & N5409;
  assign N2256 = N5387 & N5410;
  assign N2255 = N5387 & N5411;
  assign N2254 = N5387 & N5412;
  assign N2253 = N5388 & N5397;
  assign N2252 = N5388 & N5398;
  assign N2251 = N5388 & N5399;
  assign N2250 = N5388 & N5400;
  assign N2249 = N5388 & N5401;
  assign N2248 = N5388 & N5402;
  assign N2247 = N5388 & N5403;
  assign N2246 = N5388 & N5404;
  assign N2245 = N5388 & N5405;
  assign N2244 = N5388 & N5406;
  assign N2243 = N5388 & N5407;
  assign N2242 = N5388 & N5408;
  assign N2241 = N5388 & N5409;
  assign N2240 = N5388 & N5410;
  assign N2239 = N5388 & N5411;
  assign N2238 = N5388 & N5412;
  assign N5413 = num_els_r[4] & num_els_r[5];
  assign N5414 = N12 & num_els_r[5];
  assign N12 = ~num_els_r[4];
  assign N5415 = num_els_r[4] & N13;
  assign N13 = ~num_els_r[5];
  assign N5416 = N14 & N15;
  assign N14 = ~num_els_r[4];
  assign N15 = ~num_els_r[5];
  assign N5417 = num_els_r[6] & N5413;
  assign N5418 = num_els_r[6] & N5414;
  assign N5419 = num_els_r[6] & N5415;
  assign N5420 = num_els_r[6] & N5416;
  assign N5421 = N5376 & N5413;
  assign N5422 = N5376 & N5414;
  assign N5423 = N5376 & N5415;
  assign N5424 = N5376 & N5416;
  assign N5425 = num_els_r[2] & num_els_r[3];
  assign N5426 = N16 & num_els_r[3];
  assign N16 = ~num_els_r[2];
  assign N5427 = num_els_r[2] & N17;
  assign N17 = ~num_els_r[3];
  assign N5428 = N18 & N19;
  assign N18 = ~num_els_r[2];
  assign N19 = ~num_els_r[3];
  assign N5429 = num_els_r[0] & num_els_r[1];
  assign N5430 = N20 & num_els_r[1];
  assign N20 = ~num_els_r[0];
  assign N5431 = num_els_r[0] & N21;
  assign N21 = ~num_els_r[1];
  assign N5432 = N22 & N23;
  assign N22 = ~num_els_r[0];
  assign N23 = ~num_els_r[1];
  assign N5433 = N5425 & N5429;
  assign N5434 = N5425 & N5430;
  assign N5435 = N5425 & N5431;
  assign N5436 = N5425 & N5432;
  assign N5437 = N5426 & N5429;
  assign N5438 = N5426 & N5430;
  assign N5439 = N5426 & N5431;
  assign N5440 = N5426 & N5432;
  assign N5441 = N5427 & N5429;
  assign N5442 = N5427 & N5430;
  assign N5443 = N5427 & N5431;
  assign N5444 = N5427 & N5432;
  assign N5445 = N5428 & N5429;
  assign N5446 = N5428 & N5430;
  assign N5447 = N5428 & N5431;
  assign N5448 = N5428 & N5432;
  assign N2621 = N5417 & N5433;
  assign N2620 = N5417 & N5434;
  assign N2619 = N5417 & N5435;
  assign N2618 = N5417 & N5436;
  assign N2617 = N5417 & N5437;
  assign N2616 = N5417 & N5438;
  assign N2615 = N5417 & N5439;
  assign N2614 = N5417 & N5440;
  assign N2613 = N5417 & N5441;
  assign N2612 = N5417 & N5442;
  assign N2611 = N5417 & N5443;
  assign N2610 = N5417 & N5444;
  assign N2609 = N5417 & N5445;
  assign N2608 = N5417 & N5446;
  assign N2607 = N5417 & N5447;
  assign N2606 = N5417 & N5448;
  assign N2605 = N5418 & N5433;
  assign N2604 = N5418 & N5434;
  assign N2603 = N5418 & N5435;
  assign N2602 = N5418 & N5436;
  assign N2601 = N5418 & N5437;
  assign N2600 = N5418 & N5438;
  assign N2599 = N5418 & N5439;
  assign N2598 = N5418 & N5440;
  assign N2597 = N5418 & N5441;
  assign N2596 = N5418 & N5442;
  assign N2595 = N5418 & N5443;
  assign N2594 = N5418 & N5444;
  assign N2593 = N5418 & N5445;
  assign N2592 = N5418 & N5446;
  assign N2591 = N5418 & N5447;
  assign N2590 = N5418 & N5448;
  assign N2589 = N5419 & N5433;
  assign N2588 = N5419 & N5434;
  assign N2587 = N5419 & N5435;
  assign N2586 = N5419 & N5436;
  assign N2585 = N5419 & N5437;
  assign N2584 = N5419 & N5438;
  assign N2583 = N5419 & N5439;
  assign N2582 = N5419 & N5440;
  assign N2581 = N5419 & N5441;
  assign N2580 = N5419 & N5442;
  assign N2579 = N5419 & N5443;
  assign N2578 = N5419 & N5444;
  assign N2577 = N5419 & N5445;
  assign N2576 = N5419 & N5446;
  assign N2575 = N5419 & N5447;
  assign N2574 = N5419 & N5448;
  assign N2573 = N5420 & N5433;
  assign N2572 = N5420 & N5434;
  assign N2571 = N5420 & N5435;
  assign N2570 = N5420 & N5436;
  assign N2569 = N5420 & N5437;
  assign N2568 = N5420 & N5438;
  assign N2567 = N5420 & N5439;
  assign N2566 = N5420 & N5440;
  assign N2565 = N5420 & N5441;
  assign N2564 = N5420 & N5442;
  assign N2563 = N5420 & N5443;
  assign N2562 = N5420 & N5444;
  assign N2561 = N5420 & N5445;
  assign N2560 = N5420 & N5446;
  assign N2559 = N5420 & N5447;
  assign N2558 = N5420 & N5448;
  assign N2557 = N5421 & N5433;
  assign N2556 = N5421 & N5434;
  assign N2555 = N5421 & N5435;
  assign N2554 = N5421 & N5436;
  assign N2553 = N5421 & N5437;
  assign N2552 = N5421 & N5438;
  assign N2551 = N5421 & N5439;
  assign N2550 = N5421 & N5440;
  assign N2549 = N5421 & N5441;
  assign N2548 = N5421 & N5442;
  assign N2547 = N5421 & N5443;
  assign N2546 = N5421 & N5444;
  assign N2545 = N5421 & N5445;
  assign N2544 = N5421 & N5446;
  assign N2543 = N5421 & N5447;
  assign N2542 = N5421 & N5448;
  assign N2541 = N5422 & N5433;
  assign N2540 = N5422 & N5434;
  assign N2539 = N5422 & N5435;
  assign N2538 = N5422 & N5436;
  assign N2537 = N5422 & N5437;
  assign N2536 = N5422 & N5438;
  assign N2535 = N5422 & N5439;
  assign N2534 = N5422 & N5440;
  assign N2533 = N5422 & N5441;
  assign N2532 = N5422 & N5442;
  assign N2531 = N5422 & N5443;
  assign N2530 = N5422 & N5444;
  assign N2529 = N5422 & N5445;
  assign N2528 = N5422 & N5446;
  assign N2527 = N5422 & N5447;
  assign N2526 = N5422 & N5448;
  assign N2525 = N5423 & N5433;
  assign N2524 = N5423 & N5434;
  assign N2523 = N5423 & N5435;
  assign N2522 = N5423 & N5436;
  assign N2521 = N5423 & N5437;
  assign N2520 = N5423 & N5438;
  assign N2519 = N5423 & N5439;
  assign N2518 = N5423 & N5440;
  assign N2517 = N5423 & N5441;
  assign N2516 = N5423 & N5442;
  assign N2515 = N5423 & N5443;
  assign N2514 = N5423 & N5444;
  assign N2513 = N5423 & N5445;
  assign N2512 = N5423 & N5446;
  assign N2511 = N5423 & N5447;
  assign N2510 = N5423 & N5448;
  assign N2509 = N5424 & N5433;
  assign N2508 = N5424 & N5434;
  assign N2507 = N5424 & N5435;
  assign N2506 = N5424 & N5436;
  assign N2505 = N5424 & N5437;
  assign N2504 = N5424 & N5438;
  assign N2503 = N5424 & N5439;
  assign N2502 = N5424 & N5440;
  assign N2501 = N5424 & N5441;
  assign N2500 = N5424 & N5442;
  assign N2499 = N5424 & N5443;
  assign N2498 = N5424 & N5444;
  assign N2497 = N5424 & N5445;
  assign N2496 = N5424 & N5446;
  assign N2495 = N5424 & N5447;
  assign N2494 = N5424 & N5448;
  assign N5449 = N5461 & N5512;
  assign N5450 = N5461 & N5513;
  assign N5451 = N5461 & N5514;
  assign N5452 = N5461 & N5515;
  assign N3127 = N5461 & N5516;
  assign N3126 = N5461 & N5517;
  assign N3125 = N5461 & N5518;
  assign N3124 = N5461 & N5519;
  assign N3123 = N5461 & N5520;
  assign N3122 = N5461 & N5521;
  assign N3121 = N5462 & N5506;
  assign N3120 = N5462 & N5507;
  assign N3119 = N5462 & N5508;
  assign N3118 = N5462 & N5509;
  assign N3117 = N5462 & N5510;
  assign N3116 = N5462 & N5511;
  assign N3115 = N5462 & N5512;
  assign N3114 = N5462 & N5513;
  assign N3113 = N5462 & N5514;
  assign N3112 = N5462 & N5515;
  assign N3111 = N5462 & N5516;
  assign N3110 = N5462 & N5517;
  assign N3109 = N5462 & N5518;
  assign N3108 = N5462 & N5519;
  assign N3107 = N5462 & N5520;
  assign N3106 = N5462 & N5521;
  assign N3105 = N5463 & N5506;
  assign N3104 = N5463 & N5507;
  assign N3103 = N5463 & N5508;
  assign N3102 = N5463 & N5509;
  assign N3101 = N5463 & N5510;
  assign N3100 = N5463 & N5511;
  assign N3099 = N5463 & N5512;
  assign N3098 = N5463 & N5513;
  assign N3097 = N5463 & N5514;
  assign N3096 = N5463 & N5515;
  assign N3095 = N5463 & N5516;
  assign N3094 = N5463 & N5517;
  assign N3093 = N5463 & N5518;
  assign N3092 = N5463 & N5519;
  assign N3091 = N5463 & N5520;
  assign N3090 = N5463 & N5521;
  assign N3089 = N5464 & N5506;
  assign N3088 = N5464 & N5507;
  assign N3087 = N5464 & N5508;
  assign N3086 = N5464 & N5509;
  assign N3085 = N5464 & N5510;
  assign N3084 = N5464 & N5511;
  assign N3083 = N5464 & N5512;
  assign N3082 = N5464 & N5513;
  assign N3081 = N5464 & N5514;
  assign N3080 = N5464 & N5515;
  assign N3079 = N5464 & N5516;
  assign N3078 = N5464 & N5517;
  assign N3077 = N5464 & N5518;
  assign N3076 = N5464 & N5519;
  assign N3075 = N5464 & N5520;
  assign N3074 = N5464 & N5521;
  assign N3073 = N5465 & N5506;
  assign N3072 = N5465 & N5507;
  assign N3071 = N5465 & N5508;
  assign N3070 = N5465 & N5509;
  assign N3069 = N5465 & N5510;
  assign N3068 = N5465 & N5511;
  assign N3067 = N5465 & N5512;
  assign N3066 = N5465 & N5513;
  assign N3065 = N5465 & N5514;
  assign N3064 = N5465 & N5515;
  assign N3063 = N5465 & N5516;
  assign N3062 = N5465 & N5517;
  assign N3061 = N5465 & N5518;
  assign N3060 = N5465 & N5519;
  assign N3059 = N5465 & N5520;
  assign N3058 = N5465 & N5521;
  assign N3057 = N5466 & N5506;
  assign N3056 = N5466 & N5507;
  assign N3055 = N5466 & N5508;
  assign N3054 = N5466 & N5509;
  assign N3053 = N5466 & N5510;
  assign N3052 = N5466 & N5511;
  assign N3051 = N5466 & N5512;
  assign N3050 = N5466 & N5513;
  assign N3049 = N5466 & N5514;
  assign N3048 = N5466 & N5515;
  assign N3047 = N5466 & N5516;
  assign N3046 = N5466 & N5517;
  assign N3045 = N5466 & N5518;
  assign N3044 = N5466 & N5519;
  assign N3043 = N5466 & N5520;
  assign N3042 = N5466 & N5521;
  assign N3041 = N5467 & N5506;
  assign N3040 = N5467 & N5507;
  assign N3039 = N5467 & N5508;
  assign N3038 = N5467 & N5509;
  assign N3037 = N5467 & N5510;
  assign N3036 = N5467 & N5511;
  assign N3035 = N5467 & N5512;
  assign N3034 = N5467 & N5513;
  assign N3033 = N5467 & N5514;
  assign N3032 = N5467 & N5515;
  assign N3031 = N5467 & N5516;
  assign N3030 = N5467 & N5517;
  assign N3029 = N5467 & N5518;
  assign N3028 = N5467 & N5519;
  assign N3027 = N5467 & N5520;
  assign N3026 = N5467 & N5521;
  assign N3025 = N5468 & N5506;
  assign N3024 = N5468 & N5507;
  assign N3023 = N5468 & N5508;
  assign N3022 = N5468 & N5509;
  assign N3021 = N5468 & N5510;
  assign N3020 = N5468 & N5511;
  assign N3019 = N5468 & N5512;
  assign N3018 = N5468 & N5513;
  assign N3017 = N5468 & N5514;
  assign N3016 = N5468 & N5515;
  assign N3015 = N5468 & N5516;
  assign N3014 = N5468 & N5517;
  assign N3013 = N5468 & N5518;
  assign N3012 = N5468 & N5519;
  assign N3011 = N5468 & N5520;
  assign N3010 = N5468 & N5521;
  assign N5453 = yumi_cnt_i[6] & N5486;
  assign N5454 = yumi_cnt_i[6] & N5487;
  assign N5455 = yumi_cnt_i[6] & N5488;
  assign N5456 = yumi_cnt_i[6] & N5489;
  assign N5457 = N5485 & N5486;
  assign N5458 = N5485 & N5487;
  assign N5459 = N5485 & N5488;
  assign N5460 = N5485 & N5489;
  assign N3244 = N5453 & N5517;
  assign N3243 = N5453 & N5518;
  assign N3242 = N5453 & N5519;
  assign N3241 = N5453 & N5520;
  assign N3240 = N5453 & N5521;
  assign N3239 = N5454 & N5506;
  assign N3238 = N5454 & N5507;
  assign N3237 = N5454 & N5508;
  assign N3236 = N5454 & N5509;
  assign N3235 = N5454 & N5510;
  assign N3234 = N5454 & N5511;
  assign N3233 = N5454 & N5512;
  assign N3232 = N5454 & N5513;
  assign N3231 = N5454 & N5514;
  assign N3230 = N5454 & N5515;
  assign N3229 = N5454 & N5516;
  assign N3228 = N5454 & N5517;
  assign N3227 = N5454 & N5518;
  assign N3226 = N5454 & N5519;
  assign N3225 = N5454 & N5520;
  assign N3224 = N5454 & N5521;
  assign N3223 = N5455 & N5506;
  assign N3222 = N5455 & N5507;
  assign N3221 = N5455 & N5508;
  assign N3220 = N5455 & N5509;
  assign N3219 = N5455 & N5510;
  assign N3218 = N5455 & N5511;
  assign N3217 = N5455 & N5512;
  assign N3216 = N5455 & N5513;
  assign N3215 = N5455 & N5514;
  assign N3214 = N5455 & N5515;
  assign N3213 = N5455 & N5516;
  assign N3212 = N5455 & N5517;
  assign N3211 = N5455 & N5518;
  assign N3210 = N5455 & N5519;
  assign N3209 = N5455 & N5520;
  assign N3208 = N5455 & N5521;
  assign N3207 = N5456 & N5506;
  assign N3206 = N5456 & N5507;
  assign N3205 = N5456 & N5508;
  assign N3204 = N5456 & N5509;
  assign N3203 = N5456 & N5510;
  assign N3202 = N5456 & N5511;
  assign N3201 = N5456 & N5512;
  assign N3200 = N5456 & N5513;
  assign N3199 = N5456 & N5514;
  assign N3198 = N5456 & N5515;
  assign N3197 = N5456 & N5516;
  assign N3196 = N5456 & N5517;
  assign N3195 = N5456 & N5518;
  assign N3194 = N5456 & N5519;
  assign N3193 = N5456 & N5520;
  assign N3192 = N5456 & N5521;
  assign N3191 = N5457 & N5506;
  assign N3190 = N5457 & N5507;
  assign N3189 = N5457 & N5508;
  assign N3188 = N5457 & N5509;
  assign N3187 = N5457 & N5510;
  assign N3186 = N5457 & N5511;
  assign N3185 = N5457 & N5512;
  assign N3184 = N5457 & N5513;
  assign N3183 = N5457 & N5514;
  assign N3182 = N5457 & N5515;
  assign N3181 = N5457 & N5516;
  assign N3180 = N5457 & N5517;
  assign N3179 = N5457 & N5518;
  assign N3178 = N5457 & N5519;
  assign N3177 = N5457 & N5520;
  assign N3176 = N5457 & N5521;
  assign N3175 = N5458 & N5506;
  assign N3174 = N5458 & N5507;
  assign N3173 = N5458 & N5508;
  assign N3172 = N5458 & N5509;
  assign N3171 = N5458 & N5510;
  assign N3170 = N5458 & N5511;
  assign N3169 = N5458 & N5512;
  assign N3168 = N5458 & N5513;
  assign N3167 = N5458 & N5514;
  assign N3166 = N5458 & N5515;
  assign N3165 = N5458 & N5516;
  assign N3164 = N5458 & N5517;
  assign N3163 = N5458 & N5518;
  assign N3162 = N5458 & N5519;
  assign N3161 = N5458 & N5520;
  assign N3160 = N5458 & N5521;
  assign N3159 = N5459 & N5506;
  assign N3158 = N5459 & N5507;
  assign N3157 = N5459 & N5508;
  assign N3156 = N5459 & N5509;
  assign N3155 = N5459 & N5510;
  assign N3154 = N5459 & N5511;
  assign N3153 = N5459 & N5512;
  assign N3152 = N5459 & N5513;
  assign N3151 = N5459 & N5514;
  assign N3150 = N5459 & N5515;
  assign N3149 = N5459 & N5516;
  assign N3148 = N5459 & N5517;
  assign N3147 = N5459 & N5518;
  assign N3146 = N5459 & N5519;
  assign N3145 = N5459 & N5520;
  assign N3144 = N5459 & N5521;
  assign N3143 = N5460 & N5506;
  assign N3142 = N5460 & N5507;
  assign N3141 = N5460 & N5508;
  assign N3140 = N5460 & N5509;
  assign N3139 = N5460 & N5510;
  assign N3138 = N5460 & N5511;
  assign N3137 = N5460 & N5512;
  assign N3136 = N5460 & N5513;
  assign N3135 = N5460 & N5514;
  assign N3134 = N5460 & N5515;
  assign N3133 = N5460 & N5516;
  assign N3132 = N5460 & N5517;
  assign N3131 = N5460 & N5518;
  assign N3130 = N5460 & N5519;
  assign N3129 = N5460 & N5520;
  assign N3128 = N5460 & N5521;
  assign N5461 = yumi_cnt_i[6] & N5486;
  assign N5462 = yumi_cnt_i[6] & N5487;
  assign N5463 = yumi_cnt_i[6] & N5488;
  assign N5464 = yumi_cnt_i[6] & N5489;
  assign N5465 = N5485 & N5486;
  assign N5466 = N5485 & N5487;
  assign N5467 = N5485 & N5488;
  assign N5468 = N5485 & N5489;
  assign N5469 = N5498 & N5502;
  assign N5470 = N5498 & N5503;
  assign N5471 = N5498 & N5504;
  assign N5472 = N5498 & N5505;
  assign N5473 = N5499 & N5502;
  assign N5474 = N5499 & N5503;
  assign N5475 = N5499 & N5504;
  assign N5476 = N5499 & N5505;
  assign N5477 = N5500 & N5502;
  assign N5478 = N5500 & N5503;
  assign N5479 = N5500 & N5504;
  assign N5480 = N5500 & N5505;
  assign N5481 = N5501 & N5502;
  assign N5482 = N5501 & N5503;
  assign N5483 = N5501 & N5504;
  assign N5484 = N5501 & N5505;
  assign N3360 = N5461 & N5481;
  assign N3359 = N5461 & N5482;
  assign N3358 = N5461 & N5483;
  assign N3357 = N5461 & N5484;
  assign N3356 = N5462 & N5469;
  assign N3355 = N5462 & N5470;
  assign N3354 = N5462 & N5471;
  assign N3353 = N5462 & N5472;
  assign N3352 = N5462 & N5473;
  assign N3351 = N5462 & N5474;
  assign N3350 = N5462 & N5475;
  assign N3349 = N5462 & N5476;
  assign N3348 = N5462 & N5477;
  assign N3347 = N5462 & N5478;
  assign N3346 = N5462 & N5479;
  assign N3345 = N5462 & N5480;
  assign N3344 = N5462 & N5481;
  assign N3343 = N5462 & N5482;
  assign N3342 = N5462 & N5483;
  assign N3341 = N5462 & N5484;
  assign N3340 = N5463 & N5469;
  assign N3339 = N5463 & N5470;
  assign N3338 = N5463 & N5471;
  assign N3337 = N5463 & N5472;
  assign N3336 = N5463 & N5473;
  assign N3335 = N5463 & N5474;
  assign N3334 = N5463 & N5475;
  assign N3333 = N5463 & N5476;
  assign N3332 = N5463 & N5477;
  assign N3331 = N5463 & N5478;
  assign N3330 = N5463 & N5479;
  assign N3329 = N5463 & N5480;
  assign N3328 = N5463 & N5481;
  assign N3327 = N5463 & N5482;
  assign N3326 = N5463 & N5483;
  assign N3325 = N5463 & N5484;
  assign N3324 = N5464 & N5469;
  assign N3323 = N5464 & N5470;
  assign N3322 = N5464 & N5471;
  assign N3321 = N5464 & N5472;
  assign N3320 = N5464 & N5473;
  assign N3319 = N5464 & N5474;
  assign N3318 = N5464 & N5475;
  assign N3317 = N5464 & N5476;
  assign N3316 = N5464 & N5477;
  assign N3315 = N5464 & N5478;
  assign N3314 = N5464 & N5479;
  assign N3313 = N5464 & N5480;
  assign N3312 = N5464 & N5481;
  assign N3311 = N5464 & N5482;
  assign N3310 = N5464 & N5483;
  assign N3309 = N5464 & N5484;
  assign N3308 = N5465 & N5469;
  assign N3307 = N5465 & N5470;
  assign N3306 = N5465 & N5471;
  assign N3305 = N5465 & N5472;
  assign N3304 = N5465 & N5473;
  assign N3303 = N5465 & N5474;
  assign N3302 = N5465 & N5475;
  assign N3301 = N5465 & N5476;
  assign N3300 = N5465 & N5477;
  assign N3299 = N5465 & N5478;
  assign N3298 = N5465 & N5479;
  assign N3297 = N5465 & N5480;
  assign N3296 = N5465 & N5481;
  assign N3295 = N5465 & N5482;
  assign N3294 = N5465 & N5483;
  assign N3293 = N5465 & N5484;
  assign N3292 = N5466 & N5469;
  assign N3291 = N5466 & N5470;
  assign N3290 = N5466 & N5471;
  assign N3289 = N5466 & N5472;
  assign N3288 = N5466 & N5473;
  assign N3287 = N5466 & N5474;
  assign N3286 = N5466 & N5475;
  assign N3285 = N5466 & N5476;
  assign N3284 = N5466 & N5477;
  assign N3283 = N5466 & N5478;
  assign N3282 = N5466 & N5479;
  assign N3281 = N5466 & N5480;
  assign N3280 = N5466 & N5481;
  assign N3279 = N5466 & N5482;
  assign N3278 = N5466 & N5483;
  assign N3277 = N5466 & N5484;
  assign N3276 = N5467 & N5469;
  assign N3275 = N5467 & N5470;
  assign N3274 = N5467 & N5471;
  assign N3273 = N5467 & N5472;
  assign N3272 = N5467 & N5473;
  assign N3271 = N5467 & N5474;
  assign N3270 = N5467 & N5475;
  assign N3269 = N5467 & N5476;
  assign N3268 = N5467 & N5477;
  assign N3267 = N5467 & N5478;
  assign N3266 = N5467 & N5479;
  assign N3265 = N5467 & N5480;
  assign N3264 = N5467 & N5481;
  assign N3263 = N5467 & N5482;
  assign N3262 = N5467 & N5483;
  assign N3261 = N5467 & N5484;
  assign N3260 = N5468 & N5469;
  assign N3259 = N5468 & N5470;
  assign N3258 = N5468 & N5471;
  assign N3257 = N5468 & N5472;
  assign N3256 = N5468 & N5473;
  assign N3255 = N5468 & N5474;
  assign N3254 = N5468 & N5475;
  assign N3253 = N5468 & N5476;
  assign N3252 = N5468 & N5477;
  assign N3251 = N5468 & N5478;
  assign N3250 = N5468 & N5479;
  assign N3249 = N5468 & N5480;
  assign N3248 = N5468 & N5481;
  assign N3247 = N5468 & N5482;
  assign N3246 = N5468 & N5483;
  assign N3245 = N5468 & N5484;
  assign N5485 = ~yumi_cnt_i[6];
  assign N5486 = yumi_cnt_i[4] & yumi_cnt_i[5];
  assign N5487 = N24 & yumi_cnt_i[5];
  assign N24 = ~yumi_cnt_i[4];
  assign N5488 = yumi_cnt_i[4] & N25;
  assign N25 = ~yumi_cnt_i[5];
  assign N5489 = N26 & N27;
  assign N26 = ~yumi_cnt_i[4];
  assign N27 = ~yumi_cnt_i[5];
  assign N5490 = yumi_cnt_i[6] & N5486;
  assign N5491 = yumi_cnt_i[6] & N5487;
  assign N5492 = yumi_cnt_i[6] & N5488;
  assign N5493 = yumi_cnt_i[6] & N5489;
  assign N5494 = N5485 & N5486;
  assign N5495 = N5485 & N5487;
  assign N5496 = N5485 & N5488;
  assign N5497 = N5485 & N5489;
  assign N5498 = yumi_cnt_i[2] & yumi_cnt_i[3];
  assign N5499 = N28 & yumi_cnt_i[3];
  assign N28 = ~yumi_cnt_i[2];
  assign N5500 = yumi_cnt_i[2] & N29;
  assign N29 = ~yumi_cnt_i[3];
  assign N5501 = N30 & N31;
  assign N30 = ~yumi_cnt_i[2];
  assign N31 = ~yumi_cnt_i[3];
  assign N5502 = yumi_cnt_i[0] & yumi_cnt_i[1];
  assign N5503 = N32 & yumi_cnt_i[1];
  assign N32 = ~yumi_cnt_i[0];
  assign N5504 = yumi_cnt_i[0] & N33;
  assign N33 = ~yumi_cnt_i[1];
  assign N5505 = N34 & N35;
  assign N34 = ~yumi_cnt_i[0];
  assign N35 = ~yumi_cnt_i[1];
  assign N5506 = N5498 & N5502;
  assign N5507 = N5498 & N5503;
  assign N5508 = N5498 & N5504;
  assign N5509 = N5498 & N5505;
  assign N5510 = N5499 & N5502;
  assign N5511 = N5499 & N5503;
  assign N5512 = N5499 & N5504;
  assign N5513 = N5499 & N5505;
  assign N5514 = N5500 & N5502;
  assign N5515 = N5500 & N5503;
  assign N5516 = N5500 & N5504;
  assign N5517 = N5500 & N5505;
  assign N5518 = N5501 & N5502;
  assign N5519 = N5501 & N5503;
  assign N5520 = N5501 & N5504;
  assign N5521 = N5501 & N5505;
  assign N5522 = N5490 & N5507;
  assign N5523 = N5490 & N5508;
  assign N5524 = N5490 & N5509;
  assign N5525 = N5490 & N5510;
  assign N5526 = N5490 & N5511;
  assign N5527 = N5490 & N5512;
  assign N5528 = N5490 & N5513;
  assign N5529 = N5490 & N5514;
  assign N5530 = N5490 & N5515;
  assign N5531 = N5490 & N5516;
  assign N5532 = N5490 & N5517;
  assign N5533 = N5490 & N5518;
  assign N3475 = N5490 & N5519;
  assign N3474 = N5490 & N5520;
  assign N3473 = N5490 & N5521;
  assign N3472 = N5491 & N5506;
  assign N3471 = N5491 & N5507;
  assign N3470 = N5491 & N5508;
  assign N3469 = N5491 & N5509;
  assign N3468 = N5491 & N5510;
  assign N3467 = N5491 & N5511;
  assign N3466 = N5491 & N5512;
  assign N3465 = N5491 & N5513;
  assign N3464 = N5491 & N5514;
  assign N3463 = N5491 & N5515;
  assign N3462 = N5491 & N5516;
  assign N3461 = N5491 & N5517;
  assign N3460 = N5491 & N5518;
  assign N3459 = N5491 & N5519;
  assign N3458 = N5491 & N5520;
  assign N3457 = N5491 & N5521;
  assign N3456 = N5492 & N5506;
  assign N3455 = N5492 & N5507;
  assign N3454 = N5492 & N5508;
  assign N3453 = N5492 & N5509;
  assign N3452 = N5492 & N5510;
  assign N3451 = N5492 & N5511;
  assign N3450 = N5492 & N5512;
  assign N3449 = N5492 & N5513;
  assign N3448 = N5492 & N5514;
  assign N3447 = N5492 & N5515;
  assign N3446 = N5492 & N5516;
  assign N3445 = N5492 & N5517;
  assign N3444 = N5492 & N5518;
  assign N3443 = N5492 & N5519;
  assign N3442 = N5492 & N5520;
  assign N3441 = N5492 & N5521;
  assign N3440 = N5493 & N5506;
  assign N3439 = N5493 & N5507;
  assign N3438 = N5493 & N5508;
  assign N3437 = N5493 & N5509;
  assign N3436 = N5493 & N5510;
  assign N3435 = N5493 & N5511;
  assign N3434 = N5493 & N5512;
  assign N3433 = N5493 & N5513;
  assign N3432 = N5493 & N5514;
  assign N3431 = N5493 & N5515;
  assign N3430 = N5493 & N5516;
  assign N3429 = N5493 & N5517;
  assign N3428 = N5493 & N5518;
  assign N3427 = N5493 & N5519;
  assign N3426 = N5493 & N5520;
  assign N3425 = N5493 & N5521;
  assign N3424 = N5494 & N5506;
  assign N3423 = N5494 & N5507;
  assign N3422 = N5494 & N5508;
  assign N3421 = N5494 & N5509;
  assign N3420 = N5494 & N5510;
  assign N3419 = N5494 & N5511;
  assign N3418 = N5494 & N5512;
  assign N3417 = N5494 & N5513;
  assign N3416 = N5494 & N5514;
  assign N3415 = N5494 & N5515;
  assign N3414 = N5494 & N5516;
  assign N3413 = N5494 & N5517;
  assign N3412 = N5494 & N5518;
  assign N3411 = N5494 & N5519;
  assign N3410 = N5494 & N5520;
  assign N3409 = N5494 & N5521;
  assign N3408 = N5495 & N5506;
  assign N3407 = N5495 & N5507;
  assign N3406 = N5495 & N5508;
  assign N3405 = N5495 & N5509;
  assign N3404 = N5495 & N5510;
  assign N3403 = N5495 & N5511;
  assign N3402 = N5495 & N5512;
  assign N3401 = N5495 & N5513;
  assign N3400 = N5495 & N5514;
  assign N3399 = N5495 & N5515;
  assign N3398 = N5495 & N5516;
  assign N3397 = N5495 & N5517;
  assign N3396 = N5495 & N5518;
  assign N3395 = N5495 & N5519;
  assign N3394 = N5495 & N5520;
  assign N3393 = N5495 & N5521;
  assign N3392 = N5496 & N5506;
  assign N3391 = N5496 & N5507;
  assign N3390 = N5496 & N5508;
  assign N3389 = N5496 & N5509;
  assign N3388 = N5496 & N5510;
  assign N3387 = N5496 & N5511;
  assign N3386 = N5496 & N5512;
  assign N3385 = N5496 & N5513;
  assign N3384 = N5496 & N5514;
  assign N3383 = N5496 & N5515;
  assign N3382 = N5496 & N5516;
  assign N3381 = N5496 & N5517;
  assign N3380 = N5496 & N5518;
  assign N3379 = N5496 & N5519;
  assign N3378 = N5496 & N5520;
  assign N3377 = N5496 & N5521;
  assign N3376 = N5497 & N5506;
  assign N3375 = N5497 & N5507;
  assign N3374 = N5497 & N5508;
  assign N3373 = N5497 & N5509;
  assign N3372 = N5497 & N5510;
  assign N3371 = N5497 & N5511;
  assign N3370 = N5497 & N5512;
  assign N3369 = N5497 & N5513;
  assign N3368 = N5497 & N5514;
  assign N3367 = N5497 & N5515;
  assign N3366 = N5497 & N5516;
  assign N3365 = N5497 & N5517;
  assign N3364 = N5497 & N5518;
  assign N3363 = N5497 & N5519;
  assign N3362 = N5497 & N5520;
  assign N3361 = N5497 & N5521;
  assign N5534 = N5712 & N5626;
  assign N5535 = N5712 & N5627;
  assign N5536 = N5713 & N5612;
  assign N5537 = N5713 & N5613;
  assign N3521 = N5713 & N5614;
  assign N3520 = N5713 & N5615;
  assign N3519 = N5713 & N5616;
  assign N3518 = N5713 & N5617;
  assign N3517 = N5713 & N5618;
  assign N3516 = N5713 & N5619;
  assign N3515 = N5713 & N5620;
  assign N3514 = N5713 & N5621;
  assign N3513 = N5713 & N5622;
  assign N3512 = N5713 & N5623;
  assign N3511 = N5713 & N5624;
  assign N3510 = N5713 & N5625;
  assign N3509 = N5713 & N5626;
  assign N3508 = N5713 & N5627;
  assign N3507 = N5714 & N5612;
  assign N3506 = N5714 & N5613;
  assign N3505 = N5714 & N5614;
  assign N3504 = N5714 & N5615;
  assign N3503 = N5714 & N5616;
  assign N3502 = N5714 & N5617;
  assign N3501 = N5714 & N5618;
  assign N3500 = N5714 & N5619;
  assign N3499 = N5714 & N5620;
  assign N3498 = N5714 & N5621;
  assign N3497 = N5714 & N5622;
  assign N3496 = N5714 & N5623;
  assign N3495 = N5714 & N5624;
  assign N3494 = N5714 & N5625;
  assign N3493 = N5714 & N5626;
  assign N3492 = N5714 & N5627;
  assign N3491 = N5715 & N5612;
  assign N3490 = N5715 & N5613;
  assign N3489 = N5715 & N5614;
  assign N3488 = N5715 & N5615;
  assign N3487 = N5715 & N5616;
  assign N3486 = N5715 & N5617;
  assign N3485 = N5715 & N5618;
  assign N3484 = N5715 & N5619;
  assign N3483 = N5715 & N5620;
  assign N3482 = N5715 & N5621;
  assign N3481 = N5715 & N5622;
  assign N3480 = N5715 & N5623;
  assign N3479 = N5715 & N5624;
  assign N3478 = N5715 & N5625;
  assign N3477 = N5715 & N5626;
  assign N3476 = N5715 & N5627;
  assign N5538 = N5685 & N5615;
  assign N5539 = N5685 & N5616;
  assign N5540 = N5685 & N5617;
  assign N5541 = N5685 & N5618;
  assign N3626 = N5685 & N5619;
  assign N3625 = N5685 & N5620;
  assign N3624 = N5685 & N5621;
  assign N3623 = N5685 & N5622;
  assign N3622 = N5685 & N5623;
  assign N3621 = N5685 & N5624;
  assign N3620 = N5685 & N5625;
  assign N3619 = N5685 & N5626;
  assign N3618 = N5685 & N5627;
  assign N3617 = N5686 & N5612;
  assign N3616 = N5686 & N5613;
  assign N3615 = N5686 & N5614;
  assign N3614 = N5686 & N5615;
  assign N3613 = N5686 & N5616;
  assign N3612 = N5686 & N5617;
  assign N3611 = N5686 & N5618;
  assign N3610 = N5686 & N5619;
  assign N3609 = N5686 & N5620;
  assign N3608 = N5686 & N5621;
  assign N3607 = N5686 & N5622;
  assign N3606 = N5686 & N5623;
  assign N3605 = N5686 & N5624;
  assign N3604 = N5686 & N5625;
  assign N3603 = N5686 & N5626;
  assign N3602 = N5686 & N5627;
  assign N3601 = N5687 & N5612;
  assign N3600 = N5687 & N5613;
  assign N3599 = N5687 & N5614;
  assign N3598 = N5687 & N5615;
  assign N3597 = N5687 & N5616;
  assign N3596 = N5687 & N5617;
  assign N3595 = N5687 & N5618;
  assign N3594 = N5687 & N5619;
  assign N3593 = N5687 & N5620;
  assign N3592 = N5687 & N5621;
  assign N3591 = N5687 & N5622;
  assign N3590 = N5687 & N5623;
  assign N3589 = N5687 & N5624;
  assign N3588 = N5687 & N5625;
  assign N3587 = N5687 & N5626;
  assign N3586 = N5687 & N5627;
  assign N3585 = N5577 & N5612;
  assign N3584 = N5577 & N5613;
  assign N3583 = N5577 & N5614;
  assign N3582 = N5577 & N5615;
  assign N3581 = N5577 & N5616;
  assign N3580 = N5577 & N5617;
  assign N3579 = N5577 & N5618;
  assign N3578 = N5577 & N5619;
  assign N3577 = N5577 & N5620;
  assign N3576 = N5577 & N5621;
  assign N3575 = N5577 & N5622;
  assign N3574 = N5577 & N5623;
  assign N3573 = N5577 & N5624;
  assign N3572 = N5577 & N5625;
  assign N3571 = N5577 & N5626;
  assign N3570 = N5577 & N5627;
  assign N3569 = N5578 & N5612;
  assign N3568 = N5578 & N5613;
  assign N3567 = N5578 & N5614;
  assign N3566 = N5578 & N5615;
  assign N3565 = N5578 & N5616;
  assign N3564 = N5578 & N5617;
  assign N3563 = N5578 & N5618;
  assign N3562 = N5578 & N5619;
  assign N3561 = N5578 & N5620;
  assign N3560 = N5578 & N5621;
  assign N3559 = N5578 & N5622;
  assign N3558 = N5578 & N5623;
  assign N3557 = N5578 & N5624;
  assign N3556 = N5578 & N5625;
  assign N3555 = N5578 & N5626;
  assign N3554 = N5578 & N5627;
  assign N3553 = N5579 & N5612;
  assign N3552 = N5579 & N5613;
  assign N3551 = N5579 & N5614;
  assign N3550 = N5579 & N5615;
  assign N3549 = N5579 & N5616;
  assign N3548 = N5579 & N5617;
  assign N3547 = N5579 & N5618;
  assign N3546 = N5579 & N5619;
  assign N3545 = N5579 & N5620;
  assign N3544 = N5579 & N5621;
  assign N3543 = N5579 & N5622;
  assign N3542 = N5579 & N5623;
  assign N3541 = N5579 & N5624;
  assign N3540 = N5579 & N5625;
  assign N3539 = N5579 & N5626;
  assign N3538 = N5579 & N5627;
  assign N3537 = N5580 & N5612;
  assign N3536 = N5580 & N5613;
  assign N3535 = N5580 & N5614;
  assign N3534 = N5580 & N5615;
  assign N3533 = N5580 & N5616;
  assign N3532 = N5580 & N5617;
  assign N3531 = N5580 & N5618;
  assign N3530 = N5580 & N5619;
  assign N3529 = N5580 & N5620;
  assign N3528 = N5580 & N5621;
  assign N3527 = N5580 & N5622;
  assign N3526 = N5580 & N5623;
  assign N3525 = N5580 & N5624;
  assign N3524 = N5580 & N5625;
  assign N3523 = N5580 & N5626;
  assign N3522 = N5580 & N5627;
  assign N3730 = N5662 & N5620;
  assign N3729 = N5662 & N5621;
  assign N3728 = N5662 & N5622;
  assign N3727 = N5662 & N5623;
  assign N3726 = N5662 & N5624;
  assign N3725 = N5662 & N5625;
  assign N3724 = N5662 & N5626;
  assign N3723 = N5662 & N5627;
  assign N3722 = N5663 & N5612;
  assign N3721 = N5663 & N5613;
  assign N3720 = N5663 & N5614;
  assign N3719 = N5663 & N5615;
  assign N3718 = N5663 & N5616;
  assign N3717 = N5663 & N5617;
  assign N3716 = N5663 & N5618;
  assign N3715 = N5663 & N5619;
  assign N3714 = N5663 & N5620;
  assign N3713 = N5663 & N5621;
  assign N3712 = N5663 & N5622;
  assign N3711 = N5663 & N5623;
  assign N3710 = N5663 & N5624;
  assign N3709 = N5663 & N5625;
  assign N3708 = N5663 & N5626;
  assign N3707 = N5663 & N5627;
  assign N3706 = N5664 & N5612;
  assign N3705 = N5664 & N5613;
  assign N3704 = N5664 & N5614;
  assign N3703 = N5664 & N5615;
  assign N3702 = N5664 & N5616;
  assign N3701 = N5664 & N5617;
  assign N3700 = N5664 & N5618;
  assign N3699 = N5664 & N5619;
  assign N3698 = N5664 & N5620;
  assign N3697 = N5664 & N5621;
  assign N3696 = N5664 & N5622;
  assign N3695 = N5664 & N5623;
  assign N3694 = N5664 & N5624;
  assign N3693 = N5664 & N5625;
  assign N3692 = N5664 & N5626;
  assign N3691 = N5664 & N5627;
  assign N3690 = N5557 & N5612;
  assign N3689 = N5557 & N5613;
  assign N3688 = N5557 & N5614;
  assign N3687 = N5557 & N5615;
  assign N3686 = N5557 & N5616;
  assign N3685 = N5557 & N5617;
  assign N3684 = N5557 & N5618;
  assign N3683 = N5557 & N5619;
  assign N3682 = N5557 & N5620;
  assign N3681 = N5557 & N5621;
  assign N3680 = N5557 & N5622;
  assign N3679 = N5557 & N5623;
  assign N3678 = N5557 & N5624;
  assign N3677 = N5557 & N5625;
  assign N3676 = N5557 & N5626;
  assign N3675 = N5557 & N5627;
  assign N3674 = N5558 & N5612;
  assign N3673 = N5558 & N5613;
  assign N3672 = N5558 & N5614;
  assign N3671 = N5558 & N5615;
  assign N3670 = N5558 & N5616;
  assign N3669 = N5558 & N5617;
  assign N3668 = N5558 & N5618;
  assign N3667 = N5558 & N5619;
  assign N3666 = N5558 & N5620;
  assign N3665 = N5558 & N5621;
  assign N3664 = N5558 & N5622;
  assign N3663 = N5558 & N5623;
  assign N3662 = N5558 & N5624;
  assign N3661 = N5558 & N5625;
  assign N3660 = N5558 & N5626;
  assign N3659 = N5558 & N5627;
  assign N3658 = N5559 & N5612;
  assign N3657 = N5559 & N5613;
  assign N3656 = N5559 & N5614;
  assign N3655 = N5559 & N5615;
  assign N3654 = N5559 & N5616;
  assign N3653 = N5559 & N5617;
  assign N3652 = N5559 & N5618;
  assign N3651 = N5559 & N5619;
  assign N3650 = N5559 & N5620;
  assign N3649 = N5559 & N5621;
  assign N3648 = N5559 & N5622;
  assign N3647 = N5559 & N5623;
  assign N3646 = N5559 & N5624;
  assign N3645 = N5559 & N5625;
  assign N3644 = N5559 & N5626;
  assign N3643 = N5559 & N5627;
  assign N3642 = N5560 & N5612;
  assign N3641 = N5560 & N5613;
  assign N3640 = N5560 & N5614;
  assign N3639 = N5560 & N5615;
  assign N3638 = N5560 & N5616;
  assign N3637 = N5560 & N5617;
  assign N3636 = N5560 & N5618;
  assign N3635 = N5560 & N5619;
  assign N3634 = N5560 & N5620;
  assign N3633 = N5560 & N5621;
  assign N3632 = N5560 & N5622;
  assign N3631 = N5560 & N5623;
  assign N3630 = N5560 & N5624;
  assign N3629 = N5560 & N5625;
  assign N3628 = N5560 & N5626;
  assign N3627 = N5560 & N5627;
  assign N5542 = N5662 & N5590;
  assign N5543 = N5662 & N5591;
  assign N5544 = N5662 & N5592;
  assign N3830 = N5662 & N5593;
  assign N3829 = N5662 & N5594;
  assign N3828 = N5662 & N5595;
  assign N3827 = N5662 & N5596;
  assign N3826 = N5663 & N5581;
  assign N3825 = N5663 & N5582;
  assign N3824 = N5663 & N5583;
  assign N3823 = N5663 & N5584;
  assign N3822 = N5663 & N5585;
  assign N3821 = N5663 & N5586;
  assign N3820 = N5663 & N5587;
  assign N3819 = N5663 & N5588;
  assign N3818 = N5663 & N5589;
  assign N3817 = N5663 & N5590;
  assign N3816 = N5663 & N5591;
  assign N3815 = N5663 & N5592;
  assign N3814 = N5663 & N5593;
  assign N3813 = N5663 & N5594;
  assign N3812 = N5663 & N5595;
  assign N3811 = N5663 & N5596;
  assign N3810 = N5664 & N5581;
  assign N3809 = N5664 & N5582;
  assign N3808 = N5664 & N5583;
  assign N3807 = N5664 & N5584;
  assign N3806 = N5664 & N5585;
  assign N3805 = N5664 & N5586;
  assign N3804 = N5664 & N5587;
  assign N3803 = N5664 & N5588;
  assign N3802 = N5664 & N5589;
  assign N3801 = N5664 & N5590;
  assign N3800 = N5664 & N5591;
  assign N3799 = N5664 & N5592;
  assign N3798 = N5664 & N5593;
  assign N3797 = N5664 & N5594;
  assign N3796 = N5664 & N5595;
  assign N3795 = N5664 & N5596;
  assign N3794 = N5557 & N5581;
  assign N3793 = N5557 & N5582;
  assign N3792 = N5557 & N5583;
  assign N3791 = N5557 & N5584;
  assign N3790 = N5557 & N5585;
  assign N3789 = N5557 & N5586;
  assign N3788 = N5557 & N5587;
  assign N3787 = N5557 & N5588;
  assign N3786 = N5557 & N5589;
  assign N3785 = N5557 & N5590;
  assign N3784 = N5557 & N5591;
  assign N3783 = N5557 & N5592;
  assign N3782 = N5557 & N5593;
  assign N3781 = N5557 & N5594;
  assign N3780 = N5557 & N5595;
  assign N3779 = N5557 & N5596;
  assign N3778 = N5558 & N5581;
  assign N3777 = N5558 & N5582;
  assign N3776 = N5558 & N5583;
  assign N3775 = N5558 & N5584;
  assign N3774 = N5558 & N5585;
  assign N3773 = N5558 & N5586;
  assign N3772 = N5558 & N5587;
  assign N3771 = N5558 & N5588;
  assign N3770 = N5558 & N5589;
  assign N3769 = N5558 & N5590;
  assign N3768 = N5558 & N5591;
  assign N3767 = N5558 & N5592;
  assign N3766 = N5558 & N5593;
  assign N3765 = N5558 & N5594;
  assign N3764 = N5558 & N5595;
  assign N3763 = N5558 & N5596;
  assign N3762 = N5559 & N5581;
  assign N3761 = N5559 & N5582;
  assign N3760 = N5559 & N5583;
  assign N3759 = N5559 & N5584;
  assign N3758 = N5559 & N5585;
  assign N3757 = N5559 & N5586;
  assign N3756 = N5559 & N5587;
  assign N3755 = N5559 & N5588;
  assign N3754 = N5559 & N5589;
  assign N3753 = N5559 & N5590;
  assign N3752 = N5559 & N5591;
  assign N3751 = N5559 & N5592;
  assign N3750 = N5559 & N5593;
  assign N3749 = N5559 & N5594;
  assign N3748 = N5559 & N5595;
  assign N3747 = N5559 & N5596;
  assign N3746 = N5560 & N5581;
  assign N3745 = N5560 & N5582;
  assign N3744 = N5560 & N5583;
  assign N3743 = N5560 & N5584;
  assign N3742 = N5560 & N5585;
  assign N3741 = N5560 & N5586;
  assign N3740 = N5560 & N5587;
  assign N3739 = N5560 & N5588;
  assign N3738 = N5560 & N5589;
  assign N3737 = N5560 & N5590;
  assign N3736 = N5560 & N5591;
  assign N3735 = N5560 & N5592;
  assign N3734 = N5560 & N5593;
  assign N3733 = N5560 & N5594;
  assign N3732 = N5560 & N5595;
  assign N3731 = N5560 & N5596;
  assign N5545 = N5655 & N5594;
  assign N5546 = N5655 & N5595;
  assign N5547 = N5655 & N5596;
  assign N5548 = N5656 & N5581;
  assign N3861 = N5656 & N5582;
  assign N3860 = N5656 & N5583;
  assign N3859 = N5656 & N5584;
  assign N3858 = N5656 & N5585;
  assign N3857 = N5656 & N5586;
  assign N3856 = N5656 & N5587;
  assign N3855 = N5656 & N5588;
  assign N3854 = N5656 & N5589;
  assign N3853 = N5656 & N5590;
  assign N3852 = N5656 & N5591;
  assign N3851 = N5656 & N5592;
  assign N3850 = N5656 & N5593;
  assign N3849 = N5656 & N5594;
  assign N3848 = N5656 & N5595;
  assign N3847 = N5656 & N5596;
  assign N3846 = N5657 & N5581;
  assign N3845 = N5657 & N5582;
  assign N3844 = N5657 & N5583;
  assign N3843 = N5657 & N5584;
  assign N3842 = N5657 & N5585;
  assign N3841 = N5657 & N5586;
  assign N3840 = N5657 & N5587;
  assign N3839 = N5657 & N5588;
  assign N3838 = N5657 & N5589;
  assign N3837 = N5657 & N5590;
  assign N3836 = N5657 & N5591;
  assign N3835 = N5657 & N5592;
  assign N3834 = N5657 & N5593;
  assign N3833 = N5657 & N5594;
  assign N3832 = N5657 & N5595;
  assign N3831 = N5657 & N5596;
  assign N5549 = N5485 & N5708;
  assign N5550 = N5485 & N5709;
  assign N5551 = N5485 & N5710;
  assign N5552 = N5485 & N5711;
  assign N3925 = N5549 & N5581;
  assign N3924 = N5549 & N5582;
  assign N3923 = N5549 & N5583;
  assign N3922 = N5549 & N5584;
  assign N3921 = N5549 & N5585;
  assign N3920 = N5549 & N5586;
  assign N3919 = N5549 & N5587;
  assign N3918 = N5549 & N5588;
  assign N3917 = N5549 & N5589;
  assign N3916 = N5549 & N5590;
  assign N3915 = N5549 & N5591;
  assign N3914 = N5549 & N5592;
  assign N3913 = N5549 & N5593;
  assign N3912 = N5549 & N5594;
  assign N3911 = N5549 & N5595;
  assign N3910 = N5549 & N5596;
  assign N3909 = N5550 & N5581;
  assign N3908 = N5550 & N5582;
  assign N3907 = N5550 & N5583;
  assign N3906 = N5550 & N5584;
  assign N3905 = N5550 & N5585;
  assign N3904 = N5550 & N5586;
  assign N3903 = N5550 & N5587;
  assign N3902 = N5550 & N5588;
  assign N3901 = N5550 & N5589;
  assign N3900 = N5550 & N5590;
  assign N3899 = N5550 & N5591;
  assign N3898 = N5550 & N5592;
  assign N3897 = N5550 & N5593;
  assign N3896 = N5550 & N5594;
  assign N3895 = N5550 & N5595;
  assign N3894 = N5550 & N5596;
  assign N3893 = N5551 & N5581;
  assign N3892 = N5551 & N5582;
  assign N3891 = N5551 & N5583;
  assign N3890 = N5551 & N5584;
  assign N3889 = N5551 & N5585;
  assign N3888 = N5551 & N5586;
  assign N3887 = N5551 & N5587;
  assign N3886 = N5551 & N5588;
  assign N3885 = N5551 & N5589;
  assign N3884 = N5551 & N5590;
  assign N3883 = N5551 & N5591;
  assign N3882 = N5551 & N5592;
  assign N3881 = N5551 & N5593;
  assign N3880 = N5551 & N5594;
  assign N3879 = N5551 & N5595;
  assign N3878 = N5551 & N5596;
  assign N3877 = N5552 & N5581;
  assign N3876 = N5552 & N5582;
  assign N3875 = N5552 & N5583;
  assign N3874 = N5552 & N5584;
  assign N3873 = N5552 & N5585;
  assign N3872 = N5552 & N5586;
  assign N3871 = N5552 & N5587;
  assign N3870 = N5552 & N5588;
  assign N3869 = N5552 & N5589;
  assign N3868 = N5552 & N5590;
  assign N3867 = N5552 & N5591;
  assign N3866 = N5552 & N5592;
  assign N3865 = N5552 & N5593;
  assign N3864 = N5552 & N5594;
  assign N3863 = N5552 & N5595;
  assign N3862 = N5552 & N5596;
  assign N5553 = N5485 & N5708;
  assign N5554 = N5485 & N5709;
  assign N5555 = N5485 & N5710;
  assign N5556 = N5485 & N5711;
  assign N3989 = N5553 & N5581;
  assign N3988 = N5553 & N5582;
  assign N3987 = N5553 & N5583;
  assign N3986 = N5553 & N5584;
  assign N3985 = N5553 & N5585;
  assign N3984 = N5553 & N5586;
  assign N3983 = N5553 & N5587;
  assign N3982 = N5553 & N5588;
  assign N3981 = N5553 & N5589;
  assign N3980 = N5553 & N5590;
  assign N3979 = N5553 & N5591;
  assign N3978 = N5553 & N5592;
  assign N3977 = N5553 & N5593;
  assign N3976 = N5553 & N5594;
  assign N3975 = N5553 & N5595;
  assign N3974 = N5553 & N5596;
  assign N3973 = N5554 & N5581;
  assign N3972 = N5554 & N5582;
  assign N3971 = N5554 & N5583;
  assign N3970 = N5554 & N5584;
  assign N3969 = N5554 & N5585;
  assign N3968 = N5554 & N5586;
  assign N3967 = N5554 & N5587;
  assign N3966 = N5554 & N5588;
  assign N3965 = N5554 & N5589;
  assign N3964 = N5554 & N5590;
  assign N3963 = N5554 & N5591;
  assign N3962 = N5554 & N5592;
  assign N3961 = N5554 & N5593;
  assign N3960 = N5554 & N5594;
  assign N3959 = N5554 & N5595;
  assign N3958 = N5554 & N5596;
  assign N3957 = N5555 & N5581;
  assign N3956 = N5555 & N5582;
  assign N3955 = N5555 & N5583;
  assign N3954 = N5555 & N5584;
  assign N3953 = N5555 & N5585;
  assign N3952 = N5555 & N5586;
  assign N3951 = N5555 & N5587;
  assign N3950 = N5555 & N5588;
  assign N3949 = N5555 & N5589;
  assign N3948 = N5555 & N5590;
  assign N3947 = N5555 & N5591;
  assign N3946 = N5555 & N5592;
  assign N3945 = N5555 & N5593;
  assign N3944 = N5555 & N5594;
  assign N3943 = N5555 & N5595;
  assign N3942 = N5555 & N5596;
  assign N3941 = N5556 & N5581;
  assign N3940 = N5556 & N5582;
  assign N3939 = N5556 & N5583;
  assign N3938 = N5556 & N5584;
  assign N3937 = N5556 & N5585;
  assign N3936 = N5556 & N5586;
  assign N3935 = N5556 & N5587;
  assign N3934 = N5556 & N5588;
  assign N3933 = N5556 & N5589;
  assign N3932 = N5556 & N5590;
  assign N3931 = N5556 & N5591;
  assign N3930 = N5556 & N5592;
  assign N3929 = N5556 & N5593;
  assign N3928 = N5556 & N5594;
  assign N3927 = N5556 & N5595;
  assign N3926 = N5556 & N5596;
  assign N5557 = N5485 & N5708;
  assign N5558 = N5485 & N5709;
  assign N5559 = N5485 & N5710;
  assign N5560 = N5485 & N5711;
  assign N5561 = N5604 & N5608;
  assign N5562 = N5604 & N5609;
  assign N5563 = N5604 & N5610;
  assign N5564 = N5604 & N5611;
  assign N5565 = N5605 & N5608;
  assign N5566 = N5605 & N5609;
  assign N5567 = N5605 & N5610;
  assign N5568 = N5605 & N5611;
  assign N5569 = N5606 & N5608;
  assign N5570 = N5606 & N5609;
  assign N5571 = N5606 & N5610;
  assign N5572 = N5606 & N5611;
  assign N5573 = N5607 & N5608;
  assign N5574 = N5607 & N5609;
  assign N5575 = N5607 & N5610;
  assign N5576 = N5607 & N5611;
  assign N4081 = N5649 & N5565;
  assign N4080 = N5649 & N5566;
  assign N4079 = N5649 & N5567;
  assign N4078 = N5649 & N5568;
  assign N4077 = N5649 & N5569;
  assign N4076 = N5649 & N5570;
  assign N4075 = N5649 & N5571;
  assign N4074 = N5649 & N5572;
  assign N4073 = N5649 & N5573;
  assign N4072 = N5649 & N5574;
  assign N4071 = N5649 & N5575;
  assign N4070 = N5649 & N5576;
  assign N4069 = N5650 & N5561;
  assign N4068 = N5650 & N5562;
  assign N4067 = N5650 & N5563;
  assign N4066 = N5650 & N5564;
  assign N4065 = N5650 & N5565;
  assign N4064 = N5650 & N5566;
  assign N4063 = N5650 & N5567;
  assign N4062 = N5650 & N5568;
  assign N4061 = N5650 & N5569;
  assign N4060 = N5650 & N5570;
  assign N4059 = N5650 & N5571;
  assign N4058 = N5650 & N5572;
  assign N4057 = N5650 & N5573;
  assign N4056 = N5650 & N5574;
  assign N4055 = N5650 & N5575;
  assign N4054 = N5650 & N5576;
  assign N4053 = N5557 & N5561;
  assign N4052 = N5557 & N5562;
  assign N4051 = N5557 & N5563;
  assign N4050 = N5557 & N5564;
  assign N4049 = N5557 & N5565;
  assign N4048 = N5557 & N5566;
  assign N4047 = N5557 & N5567;
  assign N4046 = N5557 & N5568;
  assign N4045 = N5557 & N5569;
  assign N4044 = N5557 & N5570;
  assign N4043 = N5557 & N5571;
  assign N4042 = N5557 & N5572;
  assign N4041 = N5557 & N5573;
  assign N4040 = N5557 & N5574;
  assign N4039 = N5557 & N5575;
  assign N4038 = N5557 & N5576;
  assign N4037 = N5558 & N5561;
  assign N4036 = N5558 & N5562;
  assign N4035 = N5558 & N5563;
  assign N4034 = N5558 & N5564;
  assign N4033 = N5558 & N5565;
  assign N4032 = N5558 & N5566;
  assign N4031 = N5558 & N5567;
  assign N4030 = N5558 & N5568;
  assign N4029 = N5558 & N5569;
  assign N4028 = N5558 & N5570;
  assign N4027 = N5558 & N5571;
  assign N4026 = N5558 & N5572;
  assign N4025 = N5558 & N5573;
  assign N4024 = N5558 & N5574;
  assign N4023 = N5558 & N5575;
  assign N4022 = N5558 & N5576;
  assign N4021 = N5559 & N5561;
  assign N4020 = N5559 & N5562;
  assign N4019 = N5559 & N5563;
  assign N4018 = N5559 & N5564;
  assign N4017 = N5559 & N5565;
  assign N4016 = N5559 & N5566;
  assign N4015 = N5559 & N5567;
  assign N4014 = N5559 & N5568;
  assign N4013 = N5559 & N5569;
  assign N4012 = N5559 & N5570;
  assign N4011 = N5559 & N5571;
  assign N4010 = N5559 & N5572;
  assign N4009 = N5559 & N5573;
  assign N4008 = N5559 & N5574;
  assign N4007 = N5559 & N5575;
  assign N4006 = N5559 & N5576;
  assign N4005 = N5560 & N5561;
  assign N4004 = N5560 & N5562;
  assign N4003 = N5560 & N5563;
  assign N4002 = N5560 & N5564;
  assign N4001 = N5560 & N5565;
  assign N4000 = N5560 & N5566;
  assign N3999 = N5560 & N5567;
  assign N3998 = N5560 & N5568;
  assign N3997 = N5560 & N5569;
  assign N3996 = N5560 & N5570;
  assign N3995 = N5560 & N5571;
  assign N3994 = N5560 & N5572;
  assign N3993 = N5560 & N5573;
  assign N3992 = N5560 & N5574;
  assign N3991 = N5560 & N5575;
  assign N3990 = N5560 & N5576;
  assign N5577 = N5485 & N5708;
  assign N5578 = N5485 & N5709;
  assign N5579 = N5485 & N5710;
  assign N5580 = N5485 & N5711;
  assign N5581 = N5604 & N5608;
  assign N5582 = N5604 & N5609;
  assign N5583 = N5604 & N5610;
  assign N5584 = N5604 & N5611;
  assign N5585 = N5605 & N5608;
  assign N5586 = N5605 & N5609;
  assign N5587 = N5605 & N5610;
  assign N5588 = N5605 & N5611;
  assign N5589 = N5606 & N5608;
  assign N5590 = N5606 & N5609;
  assign N5591 = N5606 & N5610;
  assign N5592 = N5606 & N5611;
  assign N5593 = N5607 & N5608;
  assign N5594 = N5607 & N5609;
  assign N5595 = N5607 & N5610;
  assign N5596 = N5607 & N5611;
  assign N5597 = N5649 & N5583;
  assign N5598 = N5649 & N5584;
  assign N5599 = N5649 & N5585;
  assign N4172 = N5649 & N5586;
  assign N4171 = N5649 & N5587;
  assign N4170 = N5649 & N5588;
  assign N4169 = N5649 & N5589;
  assign N4168 = N5649 & N5590;
  assign N4167 = N5649 & N5591;
  assign N4166 = N5649 & N5592;
  assign N4165 = N5649 & N5593;
  assign N4164 = N5649 & N5594;
  assign N4163 = N5649 & N5595;
  assign N4162 = N5649 & N5596;
  assign N4161 = N5650 & N5581;
  assign N4160 = N5650 & N5582;
  assign N4159 = N5650 & N5583;
  assign N4158 = N5650 & N5584;
  assign N4157 = N5650 & N5585;
  assign N4156 = N5650 & N5586;
  assign N4155 = N5650 & N5587;
  assign N4154 = N5650 & N5588;
  assign N4153 = N5650 & N5589;
  assign N4152 = N5650 & N5590;
  assign N4151 = N5650 & N5591;
  assign N4150 = N5650 & N5592;
  assign N4149 = N5650 & N5593;
  assign N4148 = N5650 & N5594;
  assign N4147 = N5650 & N5595;
  assign N4146 = N5650 & N5596;
  assign N4145 = N5577 & N5581;
  assign N4144 = N5577 & N5582;
  assign N4143 = N5577 & N5583;
  assign N4142 = N5577 & N5584;
  assign N4141 = N5577 & N5585;
  assign N4140 = N5577 & N5586;
  assign N4139 = N5577 & N5587;
  assign N4138 = N5577 & N5588;
  assign N4137 = N5577 & N5589;
  assign N4136 = N5577 & N5590;
  assign N4135 = N5577 & N5591;
  assign N4134 = N5577 & N5592;
  assign N4133 = N5577 & N5593;
  assign N4132 = N5577 & N5594;
  assign N4131 = N5577 & N5595;
  assign N4130 = N5577 & N5596;
  assign N4129 = N5578 & N5581;
  assign N4128 = N5578 & N5582;
  assign N4127 = N5578 & N5583;
  assign N4126 = N5578 & N5584;
  assign N4125 = N5578 & N5585;
  assign N4124 = N5578 & N5586;
  assign N4123 = N5578 & N5587;
  assign N4122 = N5578 & N5588;
  assign N4121 = N5578 & N5589;
  assign N4120 = N5578 & N5590;
  assign N4119 = N5578 & N5591;
  assign N4118 = N5578 & N5592;
  assign N4117 = N5578 & N5593;
  assign N4116 = N5578 & N5594;
  assign N4115 = N5578 & N5595;
  assign N4114 = N5578 & N5596;
  assign N4113 = N5579 & N5581;
  assign N4112 = N5579 & N5582;
  assign N4111 = N5579 & N5583;
  assign N4110 = N5579 & N5584;
  assign N4109 = N5579 & N5585;
  assign N4108 = N5579 & N5586;
  assign N4107 = N5579 & N5587;
  assign N4106 = N5579 & N5588;
  assign N4105 = N5579 & N5589;
  assign N4104 = N5579 & N5590;
  assign N4103 = N5579 & N5591;
  assign N4102 = N5579 & N5592;
  assign N4101 = N5579 & N5593;
  assign N4100 = N5579 & N5594;
  assign N4099 = N5579 & N5595;
  assign N4098 = N5579 & N5596;
  assign N4097 = N5580 & N5581;
  assign N4096 = N5580 & N5582;
  assign N4095 = N5580 & N5583;
  assign N4094 = N5580 & N5584;
  assign N4093 = N5580 & N5585;
  assign N4092 = N5580 & N5586;
  assign N4091 = N5580 & N5587;
  assign N4090 = N5580 & N5588;
  assign N4089 = N5580 & N5589;
  assign N4088 = N5580 & N5590;
  assign N4087 = N5580 & N5591;
  assign N4086 = N5580 & N5592;
  assign N4085 = N5580 & N5593;
  assign N4084 = N5580 & N5594;
  assign N4083 = N5580 & N5595;
  assign N4082 = N5580 & N5596;
  assign N5600 = N5485 & N5708;
  assign N5601 = N5485 & N5709;
  assign N5602 = N5485 & N5710;
  assign N5603 = N5485 & N5711;
  assign N5604 = yumi_cnt_i[2] & yumi_cnt_i[3];
  assign N5605 = N36 & yumi_cnt_i[3];
  assign N36 = ~yumi_cnt_i[2];
  assign N5606 = yumi_cnt_i[2] & N37;
  assign N37 = ~yumi_cnt_i[3];
  assign N5607 = N38 & N39;
  assign N38 = ~yumi_cnt_i[2];
  assign N39 = ~yumi_cnt_i[3];
  assign N5608 = yumi_cnt_i[0] & yumi_cnt_i[1];
  assign N5609 = N40 & yumi_cnt_i[1];
  assign N40 = ~yumi_cnt_i[0];
  assign N5610 = yumi_cnt_i[0] & N41;
  assign N41 = ~yumi_cnt_i[1];
  assign N5611 = N42 & N43;
  assign N42 = ~yumi_cnt_i[0];
  assign N43 = ~yumi_cnt_i[1];
  assign N5612 = N5604 & N5608;
  assign N5613 = N5604 & N5609;
  assign N5614 = N5604 & N5610;
  assign N5615 = N5604 & N5611;
  assign N5616 = N5605 & N5608;
  assign N5617 = N5605 & N5609;
  assign N5618 = N5605 & N5610;
  assign N5619 = N5605 & N5611;
  assign N5620 = N5606 & N5608;
  assign N5621 = N5606 & N5609;
  assign N5622 = N5606 & N5610;
  assign N5623 = N5606 & N5611;
  assign N5624 = N5607 & N5608;
  assign N5625 = N5607 & N5609;
  assign N5626 = N5607 & N5610;
  assign N5627 = N5607 & N5611;
  assign N4262 = N5649 & N5618;
  assign N4261 = N5649 & N5619;
  assign N4260 = N5649 & N5620;
  assign N4259 = N5649 & N5621;
  assign N4258 = N5649 & N5622;
  assign N4257 = N5649 & N5623;
  assign N4256 = N5649 & N5624;
  assign N4255 = N5649 & N5625;
  assign N4254 = N5649 & N5626;
  assign N4253 = N5649 & N5627;
  assign N4252 = N5650 & N5612;
  assign N4251 = N5650 & N5613;
  assign N4250 = N5650 & N5614;
  assign N4249 = N5650 & N5615;
  assign N4248 = N5650 & N5616;
  assign N4247 = N5650 & N5617;
  assign N4246 = N5650 & N5618;
  assign N4245 = N5650 & N5619;
  assign N4244 = N5650 & N5620;
  assign N4243 = N5650 & N5621;
  assign N4242 = N5650 & N5622;
  assign N4241 = N5650 & N5623;
  assign N4240 = N5650 & N5624;
  assign N4239 = N5650 & N5625;
  assign N4238 = N5650 & N5626;
  assign N4237 = N5650 & N5627;
  assign N4236 = N5600 & N5612;
  assign N4235 = N5600 & N5613;
  assign N4234 = N5600 & N5614;
  assign N4233 = N5600 & N5615;
  assign N4232 = N5600 & N5616;
  assign N4231 = N5600 & N5617;
  assign N4230 = N5600 & N5618;
  assign N4229 = N5600 & N5619;
  assign N4228 = N5600 & N5620;
  assign N4227 = N5600 & N5621;
  assign N4226 = N5600 & N5622;
  assign N4225 = N5600 & N5623;
  assign N4224 = N5600 & N5624;
  assign N4223 = N5600 & N5625;
  assign N4222 = N5600 & N5626;
  assign N4221 = N5600 & N5627;
  assign N4220 = N5601 & N5612;
  assign N4219 = N5601 & N5613;
  assign N4218 = N5601 & N5614;
  assign N4217 = N5601 & N5615;
  assign N4216 = N5601 & N5616;
  assign N4215 = N5601 & N5617;
  assign N4214 = N5601 & N5618;
  assign N4213 = N5601 & N5619;
  assign N4212 = N5601 & N5620;
  assign N4211 = N5601 & N5621;
  assign N4210 = N5601 & N5622;
  assign N4209 = N5601 & N5623;
  assign N4208 = N5601 & N5624;
  assign N4207 = N5601 & N5625;
  assign N4206 = N5601 & N5626;
  assign N4205 = N5601 & N5627;
  assign N4204 = N5602 & N5612;
  assign N4203 = N5602 & N5613;
  assign N4202 = N5602 & N5614;
  assign N4201 = N5602 & N5615;
  assign N4200 = N5602 & N5616;
  assign N4199 = N5602 & N5617;
  assign N4198 = N5602 & N5618;
  assign N4197 = N5602 & N5619;
  assign N4196 = N5602 & N5620;
  assign N4195 = N5602 & N5621;
  assign N4194 = N5602 & N5622;
  assign N4193 = N5602 & N5623;
  assign N4192 = N5602 & N5624;
  assign N4191 = N5602 & N5625;
  assign N4190 = N5602 & N5626;
  assign N4189 = N5602 & N5627;
  assign N4188 = N5603 & N5612;
  assign N4187 = N5603 & N5613;
  assign N4186 = N5603 & N5614;
  assign N4185 = N5603 & N5615;
  assign N4184 = N5603 & N5616;
  assign N4183 = N5603 & N5617;
  assign N4182 = N5603 & N5618;
  assign N4181 = N5603 & N5619;
  assign N4180 = N5603 & N5620;
  assign N4179 = N5603 & N5621;
  assign N4178 = N5603 & N5622;
  assign N4177 = N5603 & N5623;
  assign N4176 = N5603 & N5624;
  assign N4175 = N5603 & N5625;
  assign N4174 = N5603 & N5626;
  assign N4173 = N5603 & N5627;
  assign N5628 = N5647 & N5735;
  assign N5629 = N5647 & N5736;
  assign N5630 = N5647 & N5737;
  assign N5631 = N5647 & N5738;
  assign N4283 = N5647 & N5739;
  assign N4282 = N5647 & N5740;
  assign N4281 = N5647 & N5741;
  assign N4280 = N5647 & N5742;
  assign N4279 = N5647 & N5743;
  assign N4278 = N5648 & N5728;
  assign N4277 = N5648 & N5729;
  assign N4276 = N5648 & N5730;
  assign N4275 = N5648 & N5731;
  assign N4274 = N5648 & N5732;
  assign N4273 = N5648 & N5733;
  assign N4272 = N5648 & N5734;
  assign N4271 = N5648 & N5735;
  assign N4270 = N5648 & N5736;
  assign N4269 = N5648 & N5737;
  assign N4268 = N5648 & N5738;
  assign N4267 = N5648 & N5739;
  assign N4266 = N5648 & N5740;
  assign N4265 = N5648 & N5741;
  assign N4264 = N5648 & N5742;
  assign N4263 = N5648 & N5743;
  assign N5632 = N5645 & N5740;
  assign N5633 = N5645 & N5741;
  assign N5634 = N5645 & N5742;
  assign N5635 = N5645 & N5743;
  assign N4363 = N5646 & N5728;
  assign N4362 = N5646 & N5729;
  assign N4361 = N5646 & N5730;
  assign N4360 = N5646 & N5731;
  assign N4359 = N5646 & N5732;
  assign N4358 = N5646 & N5733;
  assign N4357 = N5646 & N5734;
  assign N4356 = N5646 & N5735;
  assign N4355 = N5646 & N5736;
  assign N4354 = N5646 & N5737;
  assign N4353 = N5646 & N5738;
  assign N4352 = N5646 & N5739;
  assign N4351 = N5646 & N5740;
  assign N4350 = N5646 & N5741;
  assign N4349 = N5646 & N5742;
  assign N4348 = N5646 & N5743;
  assign N4347 = N5688 & N5728;
  assign N4346 = N5688 & N5729;
  assign N4345 = N5688 & N5730;
  assign N4344 = N5688 & N5731;
  assign N4343 = N5688 & N5732;
  assign N4342 = N5688 & N5733;
  assign N4341 = N5688 & N5734;
  assign N4340 = N5688 & N5735;
  assign N4339 = N5688 & N5736;
  assign N4338 = N5688 & N5737;
  assign N4337 = N5688 & N5738;
  assign N4336 = N5688 & N5739;
  assign N4335 = N5688 & N5740;
  assign N4334 = N5688 & N5741;
  assign N4333 = N5688 & N5742;
  assign N4332 = N5688 & N5743;
  assign N4331 = N5689 & N5728;
  assign N4330 = N5689 & N5729;
  assign N4329 = N5689 & N5730;
  assign N4328 = N5689 & N5731;
  assign N4327 = N5689 & N5732;
  assign N4326 = N5689 & N5733;
  assign N4325 = N5689 & N5734;
  assign N4324 = N5689 & N5735;
  assign N4323 = N5689 & N5736;
  assign N4322 = N5689 & N5737;
  assign N4321 = N5689 & N5738;
  assign N4320 = N5689 & N5739;
  assign N4319 = N5689 & N5740;
  assign N4318 = N5689 & N5741;
  assign N4317 = N5689 & N5742;
  assign N4316 = N5689 & N5743;
  assign N4315 = N5690 & N5728;
  assign N4314 = N5690 & N5729;
  assign N4313 = N5690 & N5730;
  assign N4312 = N5690 & N5731;
  assign N4311 = N5690 & N5732;
  assign N4310 = N5690 & N5733;
  assign N4309 = N5690 & N5734;
  assign N4308 = N5690 & N5735;
  assign N4307 = N5690 & N5736;
  assign N4306 = N5690 & N5737;
  assign N4305 = N5690 & N5738;
  assign N4304 = N5690 & N5739;
  assign N4303 = N5690 & N5740;
  assign N4302 = N5690 & N5741;
  assign N4301 = N5690 & N5742;
  assign N4300 = N5690 & N5743;
  assign N4299 = N5691 & N5728;
  assign N4298 = N5691 & N5729;
  assign N4297 = N5691 & N5730;
  assign N4296 = N5691 & N5731;
  assign N4295 = N5691 & N5732;
  assign N4294 = N5691 & N5733;
  assign N4293 = N5691 & N5734;
  assign N4292 = N5691 & N5735;
  assign N4291 = N5691 & N5736;
  assign N4290 = N5691 & N5737;
  assign N4289 = N5691 & N5738;
  assign N4288 = N5691 & N5739;
  assign N4287 = N5691 & N5740;
  assign N4286 = N5691 & N5741;
  assign N4285 = N5691 & N5742;
  assign N4284 = N5691 & N5743;
  assign N4442 = N5638 & N5729;
  assign N4441 = N5638 & N5730;
  assign N4440 = N5638 & N5731;
  assign N4439 = N5638 & N5732;
  assign N4438 = N5638 & N5733;
  assign N4437 = N5638 & N5734;
  assign N4436 = N5638 & N5735;
  assign N4435 = N5638 & N5736;
  assign N4434 = N5638 & N5737;
  assign N4433 = N5638 & N5738;
  assign N4432 = N5638 & N5739;
  assign N4431 = N5638 & N5740;
  assign N4430 = N5638 & N5741;
  assign N4429 = N5638 & N5742;
  assign N4428 = N5638 & N5743;
  assign N4427 = N5665 & N5728;
  assign N4426 = N5665 & N5729;
  assign N4425 = N5665 & N5730;
  assign N4424 = N5665 & N5731;
  assign N4423 = N5665 & N5732;
  assign N4422 = N5665 & N5733;
  assign N4421 = N5665 & N5734;
  assign N4420 = N5665 & N5735;
  assign N4419 = N5665 & N5736;
  assign N4418 = N5665 & N5737;
  assign N4417 = N5665 & N5738;
  assign N4416 = N5665 & N5739;
  assign N4415 = N5665 & N5740;
  assign N4414 = N5665 & N5741;
  assign N4413 = N5665 & N5742;
  assign N4412 = N5665 & N5743;
  assign N4411 = N5666 & N5728;
  assign N4410 = N5666 & N5729;
  assign N4409 = N5666 & N5730;
  assign N4408 = N5666 & N5731;
  assign N4407 = N5666 & N5732;
  assign N4406 = N5666 & N5733;
  assign N4405 = N5666 & N5734;
  assign N4404 = N5666 & N5735;
  assign N4403 = N5666 & N5736;
  assign N4402 = N5666 & N5737;
  assign N4401 = N5666 & N5738;
  assign N4400 = N5666 & N5739;
  assign N4399 = N5666 & N5740;
  assign N4398 = N5666 & N5741;
  assign N4397 = N5666 & N5742;
  assign N4396 = N5666 & N5743;
  assign N4395 = N5667 & N5728;
  assign N4394 = N5667 & N5729;
  assign N4393 = N5667 & N5730;
  assign N4392 = N5667 & N5731;
  assign N4391 = N5667 & N5732;
  assign N4390 = N5667 & N5733;
  assign N4389 = N5667 & N5734;
  assign N4388 = N5667 & N5735;
  assign N4387 = N5667 & N5736;
  assign N4386 = N5667 & N5737;
  assign N4385 = N5667 & N5738;
  assign N4384 = N5667 & N5739;
  assign N4383 = N5667 & N5740;
  assign N4382 = N5667 & N5741;
  assign N4381 = N5667 & N5742;
  assign N4380 = N5667 & N5743;
  assign N4379 = N5668 & N5728;
  assign N4378 = N5668 & N5729;
  assign N4377 = N5668 & N5730;
  assign N4376 = N5668 & N5731;
  assign N4375 = N5668 & N5732;
  assign N4374 = N5668 & N5733;
  assign N4373 = N5668 & N5734;
  assign N4372 = N5668 & N5735;
  assign N4371 = N5668 & N5736;
  assign N4370 = N5668 & N5737;
  assign N4369 = N5668 & N5738;
  assign N4368 = N5668 & N5739;
  assign N4367 = N5668 & N5740;
  assign N4366 = N5668 & N5741;
  assign N4365 = N5668 & N5742;
  assign N4364 = N5668 & N5743;
  assign N4506 = N5665 & N5692;
  assign N4505 = N5665 & N5693;
  assign N4504 = N5665 & N5694;
  assign N4503 = N5665 & N5695;
  assign N4502 = N5665 & N5696;
  assign N4501 = N5665 & N5697;
  assign N4500 = N5665 & N5698;
  assign N4499 = N5665 & N5699;
  assign N4498 = N5665 & N5700;
  assign N4497 = N5665 & N5701;
  assign N4496 = N5665 & N5702;
  assign N4495 = N5665 & N5703;
  assign N4494 = N5665 & N5704;
  assign N4493 = N5665 & N5705;
  assign N4492 = N5665 & N5706;
  assign N4491 = N5665 & N5707;
  assign N4490 = N5666 & N5692;
  assign N4489 = N5666 & N5693;
  assign N4488 = N5666 & N5694;
  assign N4487 = N5666 & N5695;
  assign N4486 = N5666 & N5696;
  assign N4485 = N5666 & N5697;
  assign N4484 = N5666 & N5698;
  assign N4483 = N5666 & N5699;
  assign N4482 = N5666 & N5700;
  assign N4481 = N5666 & N5701;
  assign N4480 = N5666 & N5702;
  assign N4479 = N5666 & N5703;
  assign N4478 = N5666 & N5704;
  assign N4477 = N5666 & N5705;
  assign N4476 = N5666 & N5706;
  assign N4475 = N5666 & N5707;
  assign N4474 = N5667 & N5692;
  assign N4473 = N5667 & N5693;
  assign N4472 = N5667 & N5694;
  assign N4471 = N5667 & N5695;
  assign N4470 = N5667 & N5696;
  assign N4469 = N5667 & N5697;
  assign N4468 = N5667 & N5698;
  assign N4467 = N5667 & N5699;
  assign N4466 = N5667 & N5700;
  assign N4465 = N5667 & N5701;
  assign N4464 = N5667 & N5702;
  assign N4463 = N5667 & N5703;
  assign N4462 = N5667 & N5704;
  assign N4461 = N5667 & N5705;
  assign N4460 = N5667 & N5706;
  assign N4459 = N5667 & N5707;
  assign N4458 = N5668 & N5692;
  assign N4457 = N5668 & N5693;
  assign N4456 = N5668 & N5694;
  assign N4455 = N5668 & N5695;
  assign N4454 = N5668 & N5696;
  assign N4453 = N5668 & N5697;
  assign N4452 = N5668 & N5698;
  assign N4451 = N5668 & N5699;
  assign N4450 = N5668 & N5700;
  assign N4449 = N5668 & N5701;
  assign N4448 = N5668 & N5702;
  assign N4447 = N5668 & N5703;
  assign N4446 = N5668 & N5704;
  assign N4445 = N5668 & N5705;
  assign N4444 = N5668 & N5706;
  assign N4443 = N5668 & N5707;
  assign N5636 = yumi_cnt_i[6] & N5711;
  assign N5637 = N5636 & N5698;
  assign N4515 = N5636 & N5699;
  assign N4514 = N5636 & N5700;
  assign N4513 = N5636 & N5701;
  assign N4512 = N5636 & N5702;
  assign N4511 = N5636 & N5703;
  assign N4510 = N5636 & N5704;
  assign N4509 = N5636 & N5705;
  assign N4508 = N5636 & N5706;
  assign N4507 = N5636 & N5707;
  assign N5638 = yumi_cnt_i[6] & N5711;
  assign N5639 = N5638 & N5694;
  assign N5640 = N5638 & N5695;
  assign N5641 = N5638 & N5696;
  assign N5642 = N5638 & N5697;
  assign N5643 = N5638 & N5698;
  assign N5644 = N5638 & N5699;
  assign N4523 = N5638 & N5700;
  assign N4522 = N5638 & N5701;
  assign N4521 = N5638 & N5702;
  assign N4520 = N5638 & N5703;
  assign N4519 = N5638 & N5704;
  assign N4518 = N5638 & N5705;
  assign N4517 = N5638 & N5706;
  assign N4516 = N5638 & N5707;
  assign N5645 = yumi_cnt_i[6] & N5710;
  assign N5646 = yumi_cnt_i[6] & N5711;
  assign N4530 = N5646 & N5701;
  assign N4529 = N5646 & N5702;
  assign N4528 = N5646 & N5703;
  assign N4527 = N5646 & N5704;
  assign N4526 = N5646 & N5705;
  assign N4525 = N5646 & N5706;
  assign N4524 = N5646 & N5707;
  assign N5647 = yumi_cnt_i[6] & N5710;
  assign N5648 = yumi_cnt_i[6] & N5711;
  assign N4536 = N5648 & N5702;
  assign N4535 = N5648 & N5703;
  assign N4534 = N5648 & N5704;
  assign N4533 = N5648 & N5705;
  assign N4532 = N5648 & N5706;
  assign N4531 = N5648 & N5707;
  assign N5649 = yumi_cnt_i[6] & N5710;
  assign N5650 = yumi_cnt_i[6] & N5711;
  assign N5651 = N5485 & N5708;
  assign N5652 = N5485 & N5709;
  assign N5653 = N5485 & N5710;
  assign N5654 = N5485 & N5711;
  assign N4605 = N5650 & N5703;
  assign N4604 = N5650 & N5704;
  assign N4603 = N5650 & N5705;
  assign N4602 = N5650 & N5706;
  assign N4601 = N5650 & N5707;
  assign N4600 = N5651 & N5692;
  assign N4599 = N5651 & N5693;
  assign N4598 = N5651 & N5694;
  assign N4597 = N5651 & N5695;
  assign N4596 = N5651 & N5696;
  assign N4595 = N5651 & N5697;
  assign N4594 = N5651 & N5698;
  assign N4593 = N5651 & N5699;
  assign N4592 = N5651 & N5700;
  assign N4591 = N5651 & N5701;
  assign N4590 = N5651 & N5702;
  assign N4589 = N5651 & N5703;
  assign N4588 = N5651 & N5704;
  assign N4587 = N5651 & N5705;
  assign N4586 = N5651 & N5706;
  assign N4585 = N5651 & N5707;
  assign N4584 = N5652 & N5692;
  assign N4583 = N5652 & N5693;
  assign N4582 = N5652 & N5694;
  assign N4581 = N5652 & N5695;
  assign N4580 = N5652 & N5696;
  assign N4579 = N5652 & N5697;
  assign N4578 = N5652 & N5698;
  assign N4577 = N5652 & N5699;
  assign N4576 = N5652 & N5700;
  assign N4575 = N5652 & N5701;
  assign N4574 = N5652 & N5702;
  assign N4573 = N5652 & N5703;
  assign N4572 = N5652 & N5704;
  assign N4571 = N5652 & N5705;
  assign N4570 = N5652 & N5706;
  assign N4569 = N5652 & N5707;
  assign N4568 = N5653 & N5692;
  assign N4567 = N5653 & N5693;
  assign N4566 = N5653 & N5694;
  assign N4565 = N5653 & N5695;
  assign N4564 = N5653 & N5696;
  assign N4563 = N5653 & N5697;
  assign N4562 = N5653 & N5698;
  assign N4561 = N5653 & N5699;
  assign N4560 = N5653 & N5700;
  assign N4559 = N5653 & N5701;
  assign N4558 = N5653 & N5702;
  assign N4557 = N5653 & N5703;
  assign N4556 = N5653 & N5704;
  assign N4555 = N5653 & N5705;
  assign N4554 = N5653 & N5706;
  assign N4553 = N5653 & N5707;
  assign N4552 = N5654 & N5692;
  assign N4551 = N5654 & N5693;
  assign N4550 = N5654 & N5694;
  assign N4549 = N5654 & N5695;
  assign N4548 = N5654 & N5696;
  assign N4547 = N5654 & N5697;
  assign N4546 = N5654 & N5698;
  assign N4545 = N5654 & N5699;
  assign N4544 = N5654 & N5700;
  assign N4543 = N5654 & N5701;
  assign N4542 = N5654 & N5702;
  assign N4541 = N5654 & N5703;
  assign N4540 = N5654 & N5704;
  assign N4539 = N5654 & N5705;
  assign N4538 = N5654 & N5706;
  assign N4537 = N5654 & N5707;
  assign N5655 = yumi_cnt_i[6] & N5709;
  assign N5656 = yumi_cnt_i[6] & N5710;
  assign N5657 = yumi_cnt_i[6] & N5711;
  assign N5658 = N5485 & N5708;
  assign N5659 = N5485 & N5709;
  assign N5660 = N5485 & N5710;
  assign N5661 = N5485 & N5711;
  assign N4673 = N5657 & N5704;
  assign N4672 = N5657 & N5705;
  assign N4671 = N5657 & N5706;
  assign N4670 = N5657 & N5707;
  assign N4669 = N5658 & N5692;
  assign N4668 = N5658 & N5693;
  assign N4667 = N5658 & N5694;
  assign N4666 = N5658 & N5695;
  assign N4665 = N5658 & N5696;
  assign N4664 = N5658 & N5697;
  assign N4663 = N5658 & N5698;
  assign N4662 = N5658 & N5699;
  assign N4661 = N5658 & N5700;
  assign N4660 = N5658 & N5701;
  assign N4659 = N5658 & N5702;
  assign N4658 = N5658 & N5703;
  assign N4657 = N5658 & N5704;
  assign N4656 = N5658 & N5705;
  assign N4655 = N5658 & N5706;
  assign N4654 = N5658 & N5707;
  assign N4653 = N5659 & N5692;
  assign N4652 = N5659 & N5693;
  assign N4651 = N5659 & N5694;
  assign N4650 = N5659 & N5695;
  assign N4649 = N5659 & N5696;
  assign N4648 = N5659 & N5697;
  assign N4647 = N5659 & N5698;
  assign N4646 = N5659 & N5699;
  assign N4645 = N5659 & N5700;
  assign N4644 = N5659 & N5701;
  assign N4643 = N5659 & N5702;
  assign N4642 = N5659 & N5703;
  assign N4641 = N5659 & N5704;
  assign N4640 = N5659 & N5705;
  assign N4639 = N5659 & N5706;
  assign N4638 = N5659 & N5707;
  assign N4637 = N5660 & N5692;
  assign N4636 = N5660 & N5693;
  assign N4635 = N5660 & N5694;
  assign N4634 = N5660 & N5695;
  assign N4633 = N5660 & N5696;
  assign N4632 = N5660 & N5697;
  assign N4631 = N5660 & N5698;
  assign N4630 = N5660 & N5699;
  assign N4629 = N5660 & N5700;
  assign N4628 = N5660 & N5701;
  assign N4627 = N5660 & N5702;
  assign N4626 = N5660 & N5703;
  assign N4625 = N5660 & N5704;
  assign N4624 = N5660 & N5705;
  assign N4623 = N5660 & N5706;
  assign N4622 = N5660 & N5707;
  assign N4621 = N5661 & N5692;
  assign N4620 = N5661 & N5693;
  assign N4619 = N5661 & N5694;
  assign N4618 = N5661 & N5695;
  assign N4617 = N5661 & N5696;
  assign N4616 = N5661 & N5697;
  assign N4615 = N5661 & N5698;
  assign N4614 = N5661 & N5699;
  assign N4613 = N5661 & N5700;
  assign N4612 = N5661 & N5701;
  assign N4611 = N5661 & N5702;
  assign N4610 = N5661 & N5703;
  assign N4609 = N5661 & N5704;
  assign N4608 = N5661 & N5705;
  assign N4607 = N5661 & N5706;
  assign N4606 = N5661 & N5707;
  assign N5662 = yumi_cnt_i[6] & N5709;
  assign N5663 = yumi_cnt_i[6] & N5710;
  assign N5664 = yumi_cnt_i[6] & N5711;
  assign N5665 = N5485 & N5708;
  assign N5666 = N5485 & N5709;
  assign N5667 = N5485 & N5710;
  assign N5668 = N5485 & N5711;
  assign N5669 = N5720 & N5724;
  assign N5670 = N5720 & N5725;
  assign N5671 = N5720 & N5726;
  assign N5672 = N5720 & N5727;
  assign N5673 = N5721 & N5724;
  assign N5674 = N5721 & N5725;
  assign N5675 = N5721 & N5726;
  assign N5676 = N5721 & N5727;
  assign N5677 = N5722 & N5724;
  assign N5678 = N5722 & N5725;
  assign N5679 = N5722 & N5726;
  assign N5680 = N5722 & N5727;
  assign N5681 = N5723 & N5724;
  assign N5682 = N5723 & N5725;
  assign N5683 = N5723 & N5726;
  assign N5684 = N5723 & N5727;
  assign N4740 = N5664 & N5682;
  assign N4739 = N5664 & N5683;
  assign N4738 = N5664 & N5684;
  assign N4737 = N5665 & N5669;
  assign N4736 = N5665 & N5670;
  assign N4735 = N5665 & N5671;
  assign N4734 = N5665 & N5672;
  assign N4733 = N5665 & N5673;
  assign N4732 = N5665 & N5674;
  assign N4731 = N5665 & N5675;
  assign N4730 = N5665 & N5676;
  assign N4729 = N5665 & N5677;
  assign N4728 = N5665 & N5678;
  assign N4727 = N5665 & N5679;
  assign N4726 = N5665 & N5680;
  assign N4725 = N5665 & N5681;
  assign N4724 = N5665 & N5682;
  assign N4723 = N5665 & N5683;
  assign N4722 = N5665 & N5684;
  assign N4721 = N5666 & N5669;
  assign N4720 = N5666 & N5670;
  assign N4719 = N5666 & N5671;
  assign N4718 = N5666 & N5672;
  assign N4717 = N5666 & N5673;
  assign N4716 = N5666 & N5674;
  assign N4715 = N5666 & N5675;
  assign N4714 = N5666 & N5676;
  assign N4713 = N5666 & N5677;
  assign N4712 = N5666 & N5678;
  assign N4711 = N5666 & N5679;
  assign N4710 = N5666 & N5680;
  assign N4709 = N5666 & N5681;
  assign N4708 = N5666 & N5682;
  assign N4707 = N5666 & N5683;
  assign N4706 = N5666 & N5684;
  assign N4705 = N5667 & N5669;
  assign N4704 = N5667 & N5670;
  assign N4703 = N5667 & N5671;
  assign N4702 = N5667 & N5672;
  assign N4701 = N5667 & N5673;
  assign N4700 = N5667 & N5674;
  assign N4699 = N5667 & N5675;
  assign N4698 = N5667 & N5676;
  assign N4697 = N5667 & N5677;
  assign N4696 = N5667 & N5678;
  assign N4695 = N5667 & N5679;
  assign N4694 = N5667 & N5680;
  assign N4693 = N5667 & N5681;
  assign N4692 = N5667 & N5682;
  assign N4691 = N5667 & N5683;
  assign N4690 = N5667 & N5684;
  assign N4689 = N5668 & N5669;
  assign N4688 = N5668 & N5670;
  assign N4687 = N5668 & N5671;
  assign N4686 = N5668 & N5672;
  assign N4685 = N5668 & N5673;
  assign N4684 = N5668 & N5674;
  assign N4683 = N5668 & N5675;
  assign N4682 = N5668 & N5676;
  assign N4681 = N5668 & N5677;
  assign N4680 = N5668 & N5678;
  assign N4679 = N5668 & N5679;
  assign N4678 = N5668 & N5680;
  assign N4677 = N5668 & N5681;
  assign N4676 = N5668 & N5682;
  assign N4675 = N5668 & N5683;
  assign N4674 = N5668 & N5684;
  assign N5685 = yumi_cnt_i[6] & N5709;
  assign N5686 = yumi_cnt_i[6] & N5710;
  assign N5687 = yumi_cnt_i[6] & N5711;
  assign N5688 = N5485 & N5708;
  assign N5689 = N5485 & N5709;
  assign N5690 = N5485 & N5710;
  assign N5691 = N5485 & N5711;
  assign N5692 = N5720 & N5724;
  assign N5693 = N5720 & N5725;
  assign N5694 = N5720 & N5726;
  assign N5695 = N5720 & N5727;
  assign N5696 = N5721 & N5724;
  assign N5697 = N5721 & N5725;
  assign N5698 = N5721 & N5726;
  assign N5699 = N5721 & N5727;
  assign N5700 = N5722 & N5724;
  assign N5701 = N5722 & N5725;
  assign N5702 = N5722 & N5726;
  assign N5703 = N5722 & N5727;
  assign N5704 = N5723 & N5724;
  assign N5705 = N5723 & N5725;
  assign N5706 = N5723 & N5726;
  assign N5707 = N5723 & N5727;
  assign N4806 = N5687 & N5706;
  assign N4805 = N5687 & N5707;
  assign N4804 = N5688 & N5692;
  assign N4803 = N5688 & N5693;
  assign N4802 = N5688 & N5694;
  assign N4801 = N5688 & N5695;
  assign N4800 = N5688 & N5696;
  assign N4799 = N5688 & N5697;
  assign N4798 = N5688 & N5698;
  assign N4797 = N5688 & N5699;
  assign N4796 = N5688 & N5700;
  assign N4795 = N5688 & N5701;
  assign N4794 = N5688 & N5702;
  assign N4793 = N5688 & N5703;
  assign N4792 = N5688 & N5704;
  assign N4791 = N5688 & N5705;
  assign N4790 = N5688 & N5706;
  assign N4789 = N5688 & N5707;
  assign N4788 = N5689 & N5692;
  assign N4787 = N5689 & N5693;
  assign N4786 = N5689 & N5694;
  assign N4785 = N5689 & N5695;
  assign N4784 = N5689 & N5696;
  assign N4783 = N5689 & N5697;
  assign N4782 = N5689 & N5698;
  assign N4781 = N5689 & N5699;
  assign N4780 = N5689 & N5700;
  assign N4779 = N5689 & N5701;
  assign N4778 = N5689 & N5702;
  assign N4777 = N5689 & N5703;
  assign N4776 = N5689 & N5704;
  assign N4775 = N5689 & N5705;
  assign N4774 = N5689 & N5706;
  assign N4773 = N5689 & N5707;
  assign N4772 = N5690 & N5692;
  assign N4771 = N5690 & N5693;
  assign N4770 = N5690 & N5694;
  assign N4769 = N5690 & N5695;
  assign N4768 = N5690 & N5696;
  assign N4767 = N5690 & N5697;
  assign N4766 = N5690 & N5698;
  assign N4765 = N5690 & N5699;
  assign N4764 = N5690 & N5700;
  assign N4763 = N5690 & N5701;
  assign N4762 = N5690 & N5702;
  assign N4761 = N5690 & N5703;
  assign N4760 = N5690 & N5704;
  assign N4759 = N5690 & N5705;
  assign N4758 = N5690 & N5706;
  assign N4757 = N5690 & N5707;
  assign N4756 = N5691 & N5692;
  assign N4755 = N5691 & N5693;
  assign N4754 = N5691 & N5694;
  assign N4753 = N5691 & N5695;
  assign N4752 = N5691 & N5696;
  assign N4751 = N5691 & N5697;
  assign N4750 = N5691 & N5698;
  assign N4749 = N5691 & N5699;
  assign N4748 = N5691 & N5700;
  assign N4747 = N5691 & N5701;
  assign N4746 = N5691 & N5702;
  assign N4745 = N5691 & N5703;
  assign N4744 = N5691 & N5704;
  assign N4743 = N5691 & N5705;
  assign N4742 = N5691 & N5706;
  assign N4741 = N5691 & N5707;
  assign N5708 = yumi_cnt_i[4] & yumi_cnt_i[5];
  assign N5709 = N44 & yumi_cnt_i[5];
  assign N44 = ~yumi_cnt_i[4];
  assign N5710 = yumi_cnt_i[4] & N45;
  assign N45 = ~yumi_cnt_i[5];
  assign N5711 = N46 & N47;
  assign N46 = ~yumi_cnt_i[4];
  assign N47 = ~yumi_cnt_i[5];
  assign N5712 = yumi_cnt_i[6] & N5708;
  assign N5713 = yumi_cnt_i[6] & N5709;
  assign N5714 = yumi_cnt_i[6] & N5710;
  assign N5715 = yumi_cnt_i[6] & N5711;
  assign N5716 = N5485 & N5708;
  assign N5717 = N5485 & N5709;
  assign N5718 = N5485 & N5710;
  assign N5719 = N5485 & N5711;
  assign N5720 = yumi_cnt_i[2] & yumi_cnt_i[3];
  assign N5721 = N48 & yumi_cnt_i[3];
  assign N48 = ~yumi_cnt_i[2];
  assign N5722 = yumi_cnt_i[2] & N49;
  assign N49 = ~yumi_cnt_i[3];
  assign N5723 = N50 & N51;
  assign N50 = ~yumi_cnt_i[2];
  assign N51 = ~yumi_cnt_i[3];
  assign N5724 = yumi_cnt_i[0] & yumi_cnt_i[1];
  assign N5725 = N52 & yumi_cnt_i[1];
  assign N52 = ~yumi_cnt_i[0];
  assign N5726 = yumi_cnt_i[0] & N53;
  assign N53 = ~yumi_cnt_i[1];
  assign N5727 = N54 & N55;
  assign N54 = ~yumi_cnt_i[0];
  assign N55 = ~yumi_cnt_i[1];
  assign N5728 = N5720 & N5724;
  assign N5729 = N5720 & N5725;
  assign N5730 = N5720 & N5726;
  assign N5731 = N5720 & N5727;
  assign N5732 = N5721 & N5724;
  assign N5733 = N5721 & N5725;
  assign N5734 = N5721 & N5726;
  assign N5735 = N5721 & N5727;
  assign N5736 = N5722 & N5724;
  assign N5737 = N5722 & N5725;
  assign N5738 = N5722 & N5726;
  assign N5739 = N5722 & N5727;
  assign N5740 = N5723 & N5724;
  assign N5741 = N5723 & N5725;
  assign N5742 = N5723 & N5726;
  assign N5743 = N5723 & N5727;
  assign N4871 = N5715 & N5743;
  assign N4870 = N5716 & N5728;
  assign N4869 = N5716 & N5729;
  assign N4868 = N5716 & N5730;
  assign N4867 = N5716 & N5731;
  assign N4866 = N5716 & N5732;
  assign N4865 = N5716 & N5733;
  assign N4864 = N5716 & N5734;
  assign N4863 = N5716 & N5735;
  assign N4862 = N5716 & N5736;
  assign N4861 = N5716 & N5737;
  assign N4860 = N5716 & N5738;
  assign N4859 = N5716 & N5739;
  assign N4858 = N5716 & N5740;
  assign N4857 = N5716 & N5741;
  assign N4856 = N5716 & N5742;
  assign N4855 = N5716 & N5743;
  assign N4854 = N5717 & N5728;
  assign N4853 = N5717 & N5729;
  assign N4852 = N5717 & N5730;
  assign N4851 = N5717 & N5731;
  assign N4850 = N5717 & N5732;
  assign N4849 = N5717 & N5733;
  assign N4848 = N5717 & N5734;
  assign N4847 = N5717 & N5735;
  assign N4846 = N5717 & N5736;
  assign N4845 = N5717 & N5737;
  assign N4844 = N5717 & N5738;
  assign N4843 = N5717 & N5739;
  assign N4842 = N5717 & N5740;
  assign N4841 = N5717 & N5741;
  assign N4840 = N5717 & N5742;
  assign N4839 = N5717 & N5743;
  assign N4838 = N5718 & N5728;
  assign N4837 = N5718 & N5729;
  assign N4836 = N5718 & N5730;
  assign N4835 = N5718 & N5731;
  assign N4834 = N5718 & N5732;
  assign N4833 = N5718 & N5733;
  assign N4832 = N5718 & N5734;
  assign N4831 = N5718 & N5735;
  assign N4830 = N5718 & N5736;
  assign N4829 = N5718 & N5737;
  assign N4828 = N5718 & N5738;
  assign N4827 = N5718 & N5739;
  assign N4826 = N5718 & N5740;
  assign N4825 = N5718 & N5741;
  assign N4824 = N5718 & N5742;
  assign N4823 = N5718 & N5743;
  assign N4822 = N5719 & N5728;
  assign N4821 = N5719 & N5729;
  assign N4820 = N5719 & N5730;
  assign N4819 = N5719 & N5731;
  assign N4818 = N5719 & N5732;
  assign N4817 = N5719 & N5733;
  assign N4816 = N5719 & N5734;
  assign N4815 = N5719 & N5735;
  assign N4814 = N5719 & N5736;
  assign N4813 = N5719 & N5737;
  assign N4812 = N5719 & N5738;
  assign N4811 = N5719 & N5739;
  assign N4810 = N5719 & N5740;
  assign N4809 = N5719 & N5741;
  assign N4808 = N5719 & N5742;
  assign N4807 = N5719 & N5743;
  assign { data_o[0:0], data_o[1:1], data_o[2:2], data_o[3:3], data_o[4:4], data_o[5:5], data_o[6:6], data_o[7:7], data_o[8:8], data_o[9:9], data_o[10:10], data_o[11:11], data_o[12:12], data_o[13:13], data_o[14:14], data_o[15:15], data_o[16:16], data_o[17:17], data_o[18:18], data_o[19:19], data_o[20:20], data_o[21:21], data_o[22:22], data_o[23:23], data_o[24:24], data_o[25:25], data_o[26:26], data_o[27:27], data_o[28:28], data_o[29:29], data_o[30:30], data_o[31:31] } = (N56)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N2366)? { data_r[0:0], data_r[1:1], data_r[2:2], data_r[3:3], data_r[4:4], data_r[5:5], data_r[6:6], data_r[7:7], data_r[8:8], data_r[9:9], data_r[10:10], data_r[11:11], data_r[12:12], data_r[13:13], data_r[14:14], data_r[15:15], data_r[16:16], data_r[17:17], data_r[18:18], data_r[19:19], data_r[20:20], data_r[21:21], data_r[22:22], data_r[23:23], data_r[24:24], data_r[25:25], data_r[26:26], data_r[27:27], data_r[28:28], data_r[29:29], data_r[30:30], data_r[31:31] } : 1'b0;
  assign N56 = N2238;
  assign { data_o[32:32], data_o[33:33], data_o[34:34], data_o[35:35], data_o[36:36], data_o[37:37], data_o[38:38], data_o[39:39], data_o[40:40], data_o[41:41], data_o[42:42], data_o[43:43], data_o[44:44], data_o[45:45], data_o[46:46], data_o[47:47], data_o[48:48], data_o[49:49], data_o[50:50], data_o[51:51], data_o[52:52], data_o[53:53], data_o[54:54], data_o[55:55], data_o[56:56], data_o[57:57], data_o[58:58], data_o[59:59], data_o[60:60], data_o[61:61], data_o[62:62], data_o[63:63] } = (N57)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2367)? { data_r[32:32], data_r[33:33], data_r[34:34], data_r[35:35], data_r[36:36], data_r[37:37], data_r[38:38], data_r[39:39], data_r[40:40], data_r[41:41], data_r[42:42], data_r[43:43], data_r[44:44], data_r[45:45], data_r[46:46], data_r[47:47], data_r[48:48], data_r[49:49], data_r[50:50], data_r[51:51], data_r[52:52], data_r[53:53], data_r[54:54], data_r[55:55], data_r[56:56], data_r[57:57], data_r[58:58], data_r[59:59], data_r[60:60], data_r[61:61], data_r[62:62], data_r[63:63] } : 1'b0;
  assign N57 = N2239;
  assign { data_o[64:64], data_o[65:65], data_o[66:66], data_o[67:67], data_o[68:68], data_o[69:69], data_o[70:70], data_o[71:71], data_o[72:72], data_o[73:73], data_o[74:74], data_o[75:75], data_o[76:76], data_o[77:77], data_o[78:78], data_o[79:79], data_o[80:80], data_o[81:81], data_o[82:82], data_o[83:83], data_o[84:84], data_o[85:85], data_o[86:86], data_o[87:87], data_o[88:88], data_o[89:89], data_o[90:90], data_o[91:91], data_o[92:92], data_o[93:93], data_o[94:94], data_o[95:95] } = (N58)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2368)? { data_r[64:64], data_r[65:65], data_r[66:66], data_r[67:67], data_r[68:68], data_r[69:69], data_r[70:70], data_r[71:71], data_r[72:72], data_r[73:73], data_r[74:74], data_r[75:75], data_r[76:76], data_r[77:77], data_r[78:78], data_r[79:79], data_r[80:80], data_r[81:81], data_r[82:82], data_r[83:83], data_r[84:84], data_r[85:85], data_r[86:86], data_r[87:87], data_r[88:88], data_r[89:89], data_r[90:90], data_r[91:91], data_r[92:92], data_r[93:93], data_r[94:94], data_r[95:95] } : 1'b0;
  assign N58 = N2240;
  assign { data_o[96:96], data_o[97:97], data_o[98:98], data_o[99:99], data_o[100:100], data_o[101:101], data_o[102:102], data_o[103:103], data_o[104:104], data_o[105:105], data_o[106:106], data_o[107:107], data_o[108:108], data_o[109:109], data_o[110:110], data_o[111:111], data_o[112:112], data_o[113:113], data_o[114:114], data_o[115:115], data_o[116:116], data_o[117:117], data_o[118:118], data_o[119:119], data_o[120:120], data_o[121:121], data_o[122:122], data_o[123:123], data_o[124:124], data_o[125:125], data_o[126:126], data_o[127:127] } = (N59)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N2369)? { data_r[96:96], data_r[97:97], data_r[98:98], data_r[99:99], data_r[100:100], data_r[101:101], data_r[102:102], data_r[103:103], data_r[104:104], data_r[105:105], data_r[106:106], data_r[107:107], data_r[108:108], data_r[109:109], data_r[110:110], data_r[111:111], data_r[112:112], data_r[113:113], data_r[114:114], data_r[115:115], data_r[116:116], data_r[117:117], data_r[118:118], data_r[119:119], data_r[120:120], data_r[121:121], data_r[122:122], data_r[123:123], data_r[124:124], data_r[125:125], data_r[126:126], data_r[127:127] } : 1'b0;
  assign N59 = N2241;
  assign { data_o[128:128], data_o[129:129], data_o[130:130], data_o[131:131], data_o[132:132], data_o[133:133], data_o[134:134], data_o[135:135], data_o[136:136], data_o[137:137], data_o[138:138], data_o[139:139], data_o[140:140], data_o[141:141], data_o[142:142], data_o[143:143], data_o[144:144], data_o[145:145], data_o[146:146], data_o[147:147], data_o[148:148], data_o[149:149], data_o[150:150], data_o[151:151], data_o[152:152], data_o[153:153], data_o[154:154], data_o[155:155], data_o[156:156], data_o[157:157], data_o[158:158], data_o[159:159] } = (N60)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2370)? { data_r[128:128], data_r[129:129], data_r[130:130], data_r[131:131], data_r[132:132], data_r[133:133], data_r[134:134], data_r[135:135], data_r[136:136], data_r[137:137], data_r[138:138], data_r[139:139], data_r[140:140], data_r[141:141], data_r[142:142], data_r[143:143], data_r[144:144], data_r[145:145], data_r[146:146], data_r[147:147], data_r[148:148], data_r[149:149], data_r[150:150], data_r[151:151], data_r[152:152], data_r[153:153], data_r[154:154], data_r[155:155], data_r[156:156], data_r[157:157], data_r[158:158], data_r[159:159] } : 1'b0;
  assign N60 = N2242;
  assign { data_o[160:160], data_o[161:161], data_o[162:162], data_o[163:163], data_o[164:164], data_o[165:165], data_o[166:166], data_o[167:167], data_o[168:168], data_o[169:169], data_o[170:170], data_o[171:171], data_o[172:172], data_o[173:173], data_o[174:174], data_o[175:175], data_o[176:176], data_o[177:177], data_o[178:178], data_o[179:179], data_o[180:180], data_o[181:181], data_o[182:182], data_o[183:183], data_o[184:184], data_o[185:185], data_o[186:186], data_o[187:187], data_o[188:188], data_o[189:189], data_o[190:190], data_o[191:191] } = (N61)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2371)? { data_r[160:160], data_r[161:161], data_r[162:162], data_r[163:163], data_r[164:164], data_r[165:165], data_r[166:166], data_r[167:167], data_r[168:168], data_r[169:169], data_r[170:170], data_r[171:171], data_r[172:172], data_r[173:173], data_r[174:174], data_r[175:175], data_r[176:176], data_r[177:177], data_r[178:178], data_r[179:179], data_r[180:180], data_r[181:181], data_r[182:182], data_r[183:183], data_r[184:184], data_r[185:185], data_r[186:186], data_r[187:187], data_r[188:188], data_r[189:189], data_r[190:190], data_r[191:191] } : 1'b0;
  assign N61 = N2243;
  assign { data_o[192:192], data_o[193:193], data_o[194:194], data_o[195:195], data_o[196:196], data_o[197:197], data_o[198:198], data_o[199:199], data_o[200:200], data_o[201:201], data_o[202:202], data_o[203:203], data_o[204:204], data_o[205:205], data_o[206:206], data_o[207:207], data_o[208:208], data_o[209:209], data_o[210:210], data_o[211:211], data_o[212:212], data_o[213:213], data_o[214:214], data_o[215:215], data_o[216:216], data_o[217:217], data_o[218:218], data_o[219:219], data_o[220:220], data_o[221:221], data_o[222:222], data_o[223:223] } = (N62)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2372)? { data_r[192:192], data_r[193:193], data_r[194:194], data_r[195:195], data_r[196:196], data_r[197:197], data_r[198:198], data_r[199:199], data_r[200:200], data_r[201:201], data_r[202:202], data_r[203:203], data_r[204:204], data_r[205:205], data_r[206:206], data_r[207:207], data_r[208:208], data_r[209:209], data_r[210:210], data_r[211:211], data_r[212:212], data_r[213:213], data_r[214:214], data_r[215:215], data_r[216:216], data_r[217:217], data_r[218:218], data_r[219:219], data_r[220:220], data_r[221:221], data_r[222:222], data_r[223:223] } : 1'b0;
  assign N62 = N2244;
  assign { data_o[224:224], data_o[225:225], data_o[226:226], data_o[227:227], data_o[228:228], data_o[229:229], data_o[230:230], data_o[231:231], data_o[232:232], data_o[233:233], data_o[234:234], data_o[235:235], data_o[236:236], data_o[237:237], data_o[238:238], data_o[239:239], data_o[240:240], data_o[241:241], data_o[242:242], data_o[243:243], data_o[244:244], data_o[245:245], data_o[246:246], data_o[247:247], data_o[248:248], data_o[249:249], data_o[250:250], data_o[251:251], data_o[252:252], data_o[253:253], data_o[254:254], data_o[255:255] } = (N63)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2373)? { data_r[224:224], data_r[225:225], data_r[226:226], data_r[227:227], data_r[228:228], data_r[229:229], data_r[230:230], data_r[231:231], data_r[232:232], data_r[233:233], data_r[234:234], data_r[235:235], data_r[236:236], data_r[237:237], data_r[238:238], data_r[239:239], data_r[240:240], data_r[241:241], data_r[242:242], data_r[243:243], data_r[244:244], data_r[245:245], data_r[246:246], data_r[247:247], data_r[248:248], data_r[249:249], data_r[250:250], data_r[251:251], data_r[252:252], data_r[253:253], data_r[254:254], data_r[255:255] } : 1'b0;
  assign N63 = N2245;
  assign { data_o[256:256], data_o[257:257], data_o[258:258], data_o[259:259], data_o[260:260], data_o[261:261], data_o[262:262], data_o[263:263], data_o[264:264], data_o[265:265], data_o[266:266], data_o[267:267], data_o[268:268], data_o[269:269], data_o[270:270], data_o[271:271], data_o[272:272], data_o[273:273], data_o[274:274], data_o[275:275], data_o[276:276], data_o[277:277], data_o[278:278], data_o[279:279], data_o[280:280], data_o[281:281], data_o[282:282], data_o[283:283], data_o[284:284], data_o[285:285], data_o[286:286], data_o[287:287] } = (N64)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2374)? { data_r[256:256], data_r[257:257], data_r[258:258], data_r[259:259], data_r[260:260], data_r[261:261], data_r[262:262], data_r[263:263], data_r[264:264], data_r[265:265], data_r[266:266], data_r[267:267], data_r[268:268], data_r[269:269], data_r[270:270], data_r[271:271], data_r[272:272], data_r[273:273], data_r[274:274], data_r[275:275], data_r[276:276], data_r[277:277], data_r[278:278], data_r[279:279], data_r[280:280], data_r[281:281], data_r[282:282], data_r[283:283], data_r[284:284], data_r[285:285], data_r[286:286], data_r[287:287] } : 1'b0;
  assign N64 = N2246;
  assign { data_o[288:288], data_o[289:289], data_o[290:290], data_o[291:291], data_o[292:292], data_o[293:293], data_o[294:294], data_o[295:295], data_o[296:296], data_o[297:297], data_o[298:298], data_o[299:299], data_o[300:300], data_o[301:301], data_o[302:302], data_o[303:303], data_o[304:304], data_o[305:305], data_o[306:306], data_o[307:307], data_o[308:308], data_o[309:309], data_o[310:310], data_o[311:311], data_o[312:312], data_o[313:313], data_o[314:314], data_o[315:315], data_o[316:316], data_o[317:317], data_o[318:318], data_o[319:319] } = (N65)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2375)? { data_r[288:288], data_r[289:289], data_r[290:290], data_r[291:291], data_r[292:292], data_r[293:293], data_r[294:294], data_r[295:295], data_r[296:296], data_r[297:297], data_r[298:298], data_r[299:299], data_r[300:300], data_r[301:301], data_r[302:302], data_r[303:303], data_r[304:304], data_r[305:305], data_r[306:306], data_r[307:307], data_r[308:308], data_r[309:309], data_r[310:310], data_r[311:311], data_r[312:312], data_r[313:313], data_r[314:314], data_r[315:315], data_r[316:316], data_r[317:317], data_r[318:318], data_r[319:319] } : 1'b0;
  assign N65 = N2247;
  assign { data_o[320:320], data_o[321:321], data_o[322:322], data_o[323:323], data_o[324:324], data_o[325:325], data_o[326:326], data_o[327:327], data_o[328:328], data_o[329:329], data_o[330:330], data_o[331:331], data_o[332:332], data_o[333:333], data_o[334:334], data_o[335:335], data_o[336:336], data_o[337:337], data_o[338:338], data_o[339:339], data_o[340:340], data_o[341:341], data_o[342:342], data_o[343:343], data_o[344:344], data_o[345:345], data_o[346:346], data_o[347:347], data_o[348:348], data_o[349:349], data_o[350:350], data_o[351:351] } = (N66)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2376)? { data_r[320:320], data_r[321:321], data_r[322:322], data_r[323:323], data_r[324:324], data_r[325:325], data_r[326:326], data_r[327:327], data_r[328:328], data_r[329:329], data_r[330:330], data_r[331:331], data_r[332:332], data_r[333:333], data_r[334:334], data_r[335:335], data_r[336:336], data_r[337:337], data_r[338:338], data_r[339:339], data_r[340:340], data_r[341:341], data_r[342:342], data_r[343:343], data_r[344:344], data_r[345:345], data_r[346:346], data_r[347:347], data_r[348:348], data_r[349:349], data_r[350:350], data_r[351:351] } : 1'b0;
  assign N66 = N2248;
  assign { data_o[352:352], data_o[353:353], data_o[354:354], data_o[355:355], data_o[356:356], data_o[357:357], data_o[358:358], data_o[359:359], data_o[360:360], data_o[361:361], data_o[362:362], data_o[363:363], data_o[364:364], data_o[365:365], data_o[366:366], data_o[367:367], data_o[368:368], data_o[369:369], data_o[370:370], data_o[371:371], data_o[372:372], data_o[373:373], data_o[374:374], data_o[375:375], data_o[376:376], data_o[377:377], data_o[378:378], data_o[379:379], data_o[380:380], data_o[381:381], data_o[382:382], data_o[383:383] } = (N67)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2377)? { data_r[352:352], data_r[353:353], data_r[354:354], data_r[355:355], data_r[356:356], data_r[357:357], data_r[358:358], data_r[359:359], data_r[360:360], data_r[361:361], data_r[362:362], data_r[363:363], data_r[364:364], data_r[365:365], data_r[366:366], data_r[367:367], data_r[368:368], data_r[369:369], data_r[370:370], data_r[371:371], data_r[372:372], data_r[373:373], data_r[374:374], data_r[375:375], data_r[376:376], data_r[377:377], data_r[378:378], data_r[379:379], data_r[380:380], data_r[381:381], data_r[382:382], data_r[383:383] } : 1'b0;
  assign N67 = N2249;
  assign { data_o[384:384], data_o[385:385], data_o[386:386], data_o[387:387], data_o[388:388], data_o[389:389], data_o[390:390], data_o[391:391], data_o[392:392], data_o[393:393], data_o[394:394], data_o[395:395], data_o[396:396], data_o[397:397], data_o[398:398], data_o[399:399], data_o[400:400], data_o[401:401], data_o[402:402], data_o[403:403], data_o[404:404], data_o[405:405], data_o[406:406], data_o[407:407], data_o[408:408], data_o[409:409], data_o[410:410], data_o[411:411], data_o[412:412], data_o[413:413], data_o[414:414], data_o[415:415] } = (N68)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2378)? { data_r[384:384], data_r[385:385], data_r[386:386], data_r[387:387], data_r[388:388], data_r[389:389], data_r[390:390], data_r[391:391], data_r[392:392], data_r[393:393], data_r[394:394], data_r[395:395], data_r[396:396], data_r[397:397], data_r[398:398], data_r[399:399], data_r[400:400], data_r[401:401], data_r[402:402], data_r[403:403], data_r[404:404], data_r[405:405], data_r[406:406], data_r[407:407], data_r[408:408], data_r[409:409], data_r[410:410], data_r[411:411], data_r[412:412], data_r[413:413], data_r[414:414], data_r[415:415] } : 1'b0;
  assign N68 = N2250;
  assign { data_o[416:416], data_o[417:417], data_o[418:418], data_o[419:419], data_o[420:420], data_o[421:421], data_o[422:422], data_o[423:423], data_o[424:424], data_o[425:425], data_o[426:426], data_o[427:427], data_o[428:428], data_o[429:429], data_o[430:430], data_o[431:431], data_o[432:432], data_o[433:433], data_o[434:434], data_o[435:435], data_o[436:436], data_o[437:437], data_o[438:438], data_o[439:439], data_o[440:440], data_o[441:441], data_o[442:442], data_o[443:443], data_o[444:444], data_o[445:445], data_o[446:446], data_o[447:447] } = (N69)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2379)? { data_r[416:416], data_r[417:417], data_r[418:418], data_r[419:419], data_r[420:420], data_r[421:421], data_r[422:422], data_r[423:423], data_r[424:424], data_r[425:425], data_r[426:426], data_r[427:427], data_r[428:428], data_r[429:429], data_r[430:430], data_r[431:431], data_r[432:432], data_r[433:433], data_r[434:434], data_r[435:435], data_r[436:436], data_r[437:437], data_r[438:438], data_r[439:439], data_r[440:440], data_r[441:441], data_r[442:442], data_r[443:443], data_r[444:444], data_r[445:445], data_r[446:446], data_r[447:447] } : 1'b0;
  assign N69 = N2251;
  assign { data_o[448:448], data_o[449:449], data_o[450:450], data_o[451:451], data_o[452:452], data_o[453:453], data_o[454:454], data_o[455:455], data_o[456:456], data_o[457:457], data_o[458:458], data_o[459:459], data_o[460:460], data_o[461:461], data_o[462:462], data_o[463:463], data_o[464:464], data_o[465:465], data_o[466:466], data_o[467:467], data_o[468:468], data_o[469:469], data_o[470:470], data_o[471:471], data_o[472:472], data_o[473:473], data_o[474:474], data_o[475:475], data_o[476:476], data_o[477:477], data_o[478:478], data_o[479:479] } = (N70)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2380)? { data_r[448:448], data_r[449:449], data_r[450:450], data_r[451:451], data_r[452:452], data_r[453:453], data_r[454:454], data_r[455:455], data_r[456:456], data_r[457:457], data_r[458:458], data_r[459:459], data_r[460:460], data_r[461:461], data_r[462:462], data_r[463:463], data_r[464:464], data_r[465:465], data_r[466:466], data_r[467:467], data_r[468:468], data_r[469:469], data_r[470:470], data_r[471:471], data_r[472:472], data_r[473:473], data_r[474:474], data_r[475:475], data_r[476:476], data_r[477:477], data_r[478:478], data_r[479:479] } : 1'b0;
  assign N70 = N2252;
  assign { data_o[480:480], data_o[481:481], data_o[482:482], data_o[483:483], data_o[484:484], data_o[485:485], data_o[486:486], data_o[487:487], data_o[488:488], data_o[489:489], data_o[490:490], data_o[491:491], data_o[492:492], data_o[493:493], data_o[494:494], data_o[495:495], data_o[496:496], data_o[497:497], data_o[498:498], data_o[499:499], data_o[500:500], data_o[501:501], data_o[502:502], data_o[503:503], data_o[504:504], data_o[505:505], data_o[506:506], data_o[507:507], data_o[508:508], data_o[509:509], data_o[510:510], data_o[511:511] } = (N71)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2381)? { data_r[480:480], data_r[481:481], data_r[482:482], data_r[483:483], data_r[484:484], data_r[485:485], data_r[486:486], data_r[487:487], data_r[488:488], data_r[489:489], data_r[490:490], data_r[491:491], data_r[492:492], data_r[493:493], data_r[494:494], data_r[495:495], data_r[496:496], data_r[497:497], data_r[498:498], data_r[499:499], data_r[500:500], data_r[501:501], data_r[502:502], data_r[503:503], data_r[504:504], data_r[505:505], data_r[506:506], data_r[507:507], data_r[508:508], data_r[509:509], data_r[510:510], data_r[511:511] } : 1'b0;
  assign N71 = N2253;
  assign { data_o[512:512], data_o[513:513], data_o[514:514], data_o[515:515], data_o[516:516], data_o[517:517], data_o[518:518], data_o[519:519], data_o[520:520], data_o[521:521], data_o[522:522], data_o[523:523], data_o[524:524], data_o[525:525], data_o[526:526], data_o[527:527], data_o[528:528], data_o[529:529], data_o[530:530], data_o[531:531], data_o[532:532], data_o[533:533], data_o[534:534], data_o[535:535], data_o[536:536], data_o[537:537], data_o[538:538], data_o[539:539], data_o[540:540], data_o[541:541], data_o[542:542], data_o[543:543] } = (N72)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2382)? { data_r[512:512], data_r[513:513], data_r[514:514], data_r[515:515], data_r[516:516], data_r[517:517], data_r[518:518], data_r[519:519], data_r[520:520], data_r[521:521], data_r[522:522], data_r[523:523], data_r[524:524], data_r[525:525], data_r[526:526], data_r[527:527], data_r[528:528], data_r[529:529], data_r[530:530], data_r[531:531], data_r[532:532], data_r[533:533], data_r[534:534], data_r[535:535], data_r[536:536], data_r[537:537], data_r[538:538], data_r[539:539], data_r[540:540], data_r[541:541], data_r[542:542], data_r[543:543] } : 1'b0;
  assign N72 = N2254;
  assign { data_o[544:544], data_o[545:545], data_o[546:546], data_o[547:547], data_o[548:548], data_o[549:549], data_o[550:550], data_o[551:551], data_o[552:552], data_o[553:553], data_o[554:554], data_o[555:555], data_o[556:556], data_o[557:557], data_o[558:558], data_o[559:559], data_o[560:560], data_o[561:561], data_o[562:562], data_o[563:563], data_o[564:564], data_o[565:565], data_o[566:566], data_o[567:567], data_o[568:568], data_o[569:569], data_o[570:570], data_o[571:571], data_o[572:572], data_o[573:573], data_o[574:574], data_o[575:575] } = (N73)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2383)? { data_r[544:544], data_r[545:545], data_r[546:546], data_r[547:547], data_r[548:548], data_r[549:549], data_r[550:550], data_r[551:551], data_r[552:552], data_r[553:553], data_r[554:554], data_r[555:555], data_r[556:556], data_r[557:557], data_r[558:558], data_r[559:559], data_r[560:560], data_r[561:561], data_r[562:562], data_r[563:563], data_r[564:564], data_r[565:565], data_r[566:566], data_r[567:567], data_r[568:568], data_r[569:569], data_r[570:570], data_r[571:571], data_r[572:572], data_r[573:573], data_r[574:574], data_r[575:575] } : 1'b0;
  assign N73 = N2255;
  assign { data_o[576:576], data_o[577:577], data_o[578:578], data_o[579:579], data_o[580:580], data_o[581:581], data_o[582:582], data_o[583:583], data_o[584:584], data_o[585:585], data_o[586:586], data_o[587:587], data_o[588:588], data_o[589:589], data_o[590:590], data_o[591:591], data_o[592:592], data_o[593:593], data_o[594:594], data_o[595:595], data_o[596:596], data_o[597:597], data_o[598:598], data_o[599:599], data_o[600:600], data_o[601:601], data_o[602:602], data_o[603:603], data_o[604:604], data_o[605:605], data_o[606:606], data_o[607:607] } = (N74)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2384)? { data_r[576:576], data_r[577:577], data_r[578:578], data_r[579:579], data_r[580:580], data_r[581:581], data_r[582:582], data_r[583:583], data_r[584:584], data_r[585:585], data_r[586:586], data_r[587:587], data_r[588:588], data_r[589:589], data_r[590:590], data_r[591:591], data_r[592:592], data_r[593:593], data_r[594:594], data_r[595:595], data_r[596:596], data_r[597:597], data_r[598:598], data_r[599:599], data_r[600:600], data_r[601:601], data_r[602:602], data_r[603:603], data_r[604:604], data_r[605:605], data_r[606:606], data_r[607:607] } : 1'b0;
  assign N74 = N2256;
  assign { data_o[608:608], data_o[609:609], data_o[610:610], data_o[611:611], data_o[612:612], data_o[613:613], data_o[614:614], data_o[615:615], data_o[616:616], data_o[617:617], data_o[618:618], data_o[619:619], data_o[620:620], data_o[621:621], data_o[622:622], data_o[623:623], data_o[624:624], data_o[625:625], data_o[626:626], data_o[627:627], data_o[628:628], data_o[629:629], data_o[630:630], data_o[631:631], data_o[632:632], data_o[633:633], data_o[634:634], data_o[635:635], data_o[636:636], data_o[637:637], data_o[638:638], data_o[639:639] } = (N75)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2385)? { data_r[608:608], data_r[609:609], data_r[610:610], data_r[611:611], data_r[612:612], data_r[613:613], data_r[614:614], data_r[615:615], data_r[616:616], data_r[617:617], data_r[618:618], data_r[619:619], data_r[620:620], data_r[621:621], data_r[622:622], data_r[623:623], data_r[624:624], data_r[625:625], data_r[626:626], data_r[627:627], data_r[628:628], data_r[629:629], data_r[630:630], data_r[631:631], data_r[632:632], data_r[633:633], data_r[634:634], data_r[635:635], data_r[636:636], data_r[637:637], data_r[638:638], data_r[639:639] } : 1'b0;
  assign N75 = N2257;
  assign { data_o[640:640], data_o[641:641], data_o[642:642], data_o[643:643], data_o[644:644], data_o[645:645], data_o[646:646], data_o[647:647], data_o[648:648], data_o[649:649], data_o[650:650], data_o[651:651], data_o[652:652], data_o[653:653], data_o[654:654], data_o[655:655], data_o[656:656], data_o[657:657], data_o[658:658], data_o[659:659], data_o[660:660], data_o[661:661], data_o[662:662], data_o[663:663], data_o[664:664], data_o[665:665], data_o[666:666], data_o[667:667], data_o[668:668], data_o[669:669], data_o[670:670], data_o[671:671] } = (N76)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2386)? { data_r[640:640], data_r[641:641], data_r[642:642], data_r[643:643], data_r[644:644], data_r[645:645], data_r[646:646], data_r[647:647], data_r[648:648], data_r[649:649], data_r[650:650], data_r[651:651], data_r[652:652], data_r[653:653], data_r[654:654], data_r[655:655], data_r[656:656], data_r[657:657], data_r[658:658], data_r[659:659], data_r[660:660], data_r[661:661], data_r[662:662], data_r[663:663], data_r[664:664], data_r[665:665], data_r[666:666], data_r[667:667], data_r[668:668], data_r[669:669], data_r[670:670], data_r[671:671] } : 1'b0;
  assign N76 = N2258;
  assign { data_o[672:672], data_o[673:673], data_o[674:674], data_o[675:675], data_o[676:676], data_o[677:677], data_o[678:678], data_o[679:679], data_o[680:680], data_o[681:681], data_o[682:682], data_o[683:683], data_o[684:684], data_o[685:685], data_o[686:686], data_o[687:687], data_o[688:688], data_o[689:689], data_o[690:690], data_o[691:691], data_o[692:692], data_o[693:693], data_o[694:694], data_o[695:695], data_o[696:696], data_o[697:697], data_o[698:698], data_o[699:699], data_o[700:700], data_o[701:701], data_o[702:702], data_o[703:703] } = (N77)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2387)? { data_r[672:672], data_r[673:673], data_r[674:674], data_r[675:675], data_r[676:676], data_r[677:677], data_r[678:678], data_r[679:679], data_r[680:680], data_r[681:681], data_r[682:682], data_r[683:683], data_r[684:684], data_r[685:685], data_r[686:686], data_r[687:687], data_r[688:688], data_r[689:689], data_r[690:690], data_r[691:691], data_r[692:692], data_r[693:693], data_r[694:694], data_r[695:695], data_r[696:696], data_r[697:697], data_r[698:698], data_r[699:699], data_r[700:700], data_r[701:701], data_r[702:702], data_r[703:703] } : 1'b0;
  assign N77 = N2259;
  assign { data_o[704:704], data_o[705:705], data_o[706:706], data_o[707:707], data_o[708:708], data_o[709:709], data_o[710:710], data_o[711:711], data_o[712:712], data_o[713:713], data_o[714:714], data_o[715:715], data_o[716:716], data_o[717:717], data_o[718:718], data_o[719:719], data_o[720:720], data_o[721:721], data_o[722:722], data_o[723:723], data_o[724:724], data_o[725:725], data_o[726:726], data_o[727:727], data_o[728:728], data_o[729:729], data_o[730:730], data_o[731:731], data_o[732:732], data_o[733:733], data_o[734:734], data_o[735:735] } = (N78)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2388)? { data_r[704:704], data_r[705:705], data_r[706:706], data_r[707:707], data_r[708:708], data_r[709:709], data_r[710:710], data_r[711:711], data_r[712:712], data_r[713:713], data_r[714:714], data_r[715:715], data_r[716:716], data_r[717:717], data_r[718:718], data_r[719:719], data_r[720:720], data_r[721:721], data_r[722:722], data_r[723:723], data_r[724:724], data_r[725:725], data_r[726:726], data_r[727:727], data_r[728:728], data_r[729:729], data_r[730:730], data_r[731:731], data_r[732:732], data_r[733:733], data_r[734:734], data_r[735:735] } : 1'b0;
  assign N78 = N2260;
  assign { data_o[736:736], data_o[737:737], data_o[738:738], data_o[739:739], data_o[740:740], data_o[741:741], data_o[742:742], data_o[743:743], data_o[744:744], data_o[745:745], data_o[746:746], data_o[747:747], data_o[748:748], data_o[749:749], data_o[750:750], data_o[751:751], data_o[752:752], data_o[753:753], data_o[754:754], data_o[755:755], data_o[756:756], data_o[757:757], data_o[758:758], data_o[759:759], data_o[760:760], data_o[761:761], data_o[762:762], data_o[763:763], data_o[764:764], data_o[765:765], data_o[766:766], data_o[767:767] } = (N79)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2389)? { data_r[736:736], data_r[737:737], data_r[738:738], data_r[739:739], data_r[740:740], data_r[741:741], data_r[742:742], data_r[743:743], data_r[744:744], data_r[745:745], data_r[746:746], data_r[747:747], data_r[748:748], data_r[749:749], data_r[750:750], data_r[751:751], data_r[752:752], data_r[753:753], data_r[754:754], data_r[755:755], data_r[756:756], data_r[757:757], data_r[758:758], data_r[759:759], data_r[760:760], data_r[761:761], data_r[762:762], data_r[763:763], data_r[764:764], data_r[765:765], data_r[766:766], data_r[767:767] } : 1'b0;
  assign N79 = N2261;
  assign { data_o[768:768], data_o[769:769], data_o[770:770], data_o[771:771], data_o[772:772], data_o[773:773], data_o[774:774], data_o[775:775], data_o[776:776], data_o[777:777], data_o[778:778], data_o[779:779], data_o[780:780], data_o[781:781], data_o[782:782], data_o[783:783], data_o[784:784], data_o[785:785], data_o[786:786], data_o[787:787], data_o[788:788], data_o[789:789], data_o[790:790], data_o[791:791], data_o[792:792], data_o[793:793], data_o[794:794], data_o[795:795], data_o[796:796], data_o[797:797], data_o[798:798], data_o[799:799] } = (N80)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2390)? { data_r[768:768], data_r[769:769], data_r[770:770], data_r[771:771], data_r[772:772], data_r[773:773], data_r[774:774], data_r[775:775], data_r[776:776], data_r[777:777], data_r[778:778], data_r[779:779], data_r[780:780], data_r[781:781], data_r[782:782], data_r[783:783], data_r[784:784], data_r[785:785], data_r[786:786], data_r[787:787], data_r[788:788], data_r[789:789], data_r[790:790], data_r[791:791], data_r[792:792], data_r[793:793], data_r[794:794], data_r[795:795], data_r[796:796], data_r[797:797], data_r[798:798], data_r[799:799] } : 1'b0;
  assign N80 = N2262;
  assign { data_o[800:800], data_o[801:801], data_o[802:802], data_o[803:803], data_o[804:804], data_o[805:805], data_o[806:806], data_o[807:807], data_o[808:808], data_o[809:809], data_o[810:810], data_o[811:811], data_o[812:812], data_o[813:813], data_o[814:814], data_o[815:815], data_o[816:816], data_o[817:817], data_o[818:818], data_o[819:819], data_o[820:820], data_o[821:821], data_o[822:822], data_o[823:823], data_o[824:824], data_o[825:825], data_o[826:826], data_o[827:827], data_o[828:828], data_o[829:829], data_o[830:830], data_o[831:831] } = (N81)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2391)? { data_r[800:800], data_r[801:801], data_r[802:802], data_r[803:803], data_r[804:804], data_r[805:805], data_r[806:806], data_r[807:807], data_r[808:808], data_r[809:809], data_r[810:810], data_r[811:811], data_r[812:812], data_r[813:813], data_r[814:814], data_r[815:815], data_r[816:816], data_r[817:817], data_r[818:818], data_r[819:819], data_r[820:820], data_r[821:821], data_r[822:822], data_r[823:823], data_r[824:824], data_r[825:825], data_r[826:826], data_r[827:827], data_r[828:828], data_r[829:829], data_r[830:830], data_r[831:831] } : 1'b0;
  assign N81 = N2263;
  assign { data_o[832:832], data_o[833:833], data_o[834:834], data_o[835:835], data_o[836:836], data_o[837:837], data_o[838:838], data_o[839:839], data_o[840:840], data_o[841:841], data_o[842:842], data_o[843:843], data_o[844:844], data_o[845:845], data_o[846:846], data_o[847:847], data_o[848:848], data_o[849:849], data_o[850:850], data_o[851:851], data_o[852:852], data_o[853:853], data_o[854:854], data_o[855:855], data_o[856:856], data_o[857:857], data_o[858:858], data_o[859:859], data_o[860:860], data_o[861:861], data_o[862:862], data_o[863:863] } = (N82)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2392)? { data_r[832:832], data_r[833:833], data_r[834:834], data_r[835:835], data_r[836:836], data_r[837:837], data_r[838:838], data_r[839:839], data_r[840:840], data_r[841:841], data_r[842:842], data_r[843:843], data_r[844:844], data_r[845:845], data_r[846:846], data_r[847:847], data_r[848:848], data_r[849:849], data_r[850:850], data_r[851:851], data_r[852:852], data_r[853:853], data_r[854:854], data_r[855:855], data_r[856:856], data_r[857:857], data_r[858:858], data_r[859:859], data_r[860:860], data_r[861:861], data_r[862:862], data_r[863:863] } : 1'b0;
  assign N82 = N2264;
  assign { data_o[864:864], data_o[865:865], data_o[866:866], data_o[867:867], data_o[868:868], data_o[869:869], data_o[870:870], data_o[871:871], data_o[872:872], data_o[873:873], data_o[874:874], data_o[875:875], data_o[876:876], data_o[877:877], data_o[878:878], data_o[879:879], data_o[880:880], data_o[881:881], data_o[882:882], data_o[883:883], data_o[884:884], data_o[885:885], data_o[886:886], data_o[887:887], data_o[888:888], data_o[889:889], data_o[890:890], data_o[891:891], data_o[892:892], data_o[893:893], data_o[894:894], data_o[895:895] } = (N83)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2393)? { data_r[864:864], data_r[865:865], data_r[866:866], data_r[867:867], data_r[868:868], data_r[869:869], data_r[870:870], data_r[871:871], data_r[872:872], data_r[873:873], data_r[874:874], data_r[875:875], data_r[876:876], data_r[877:877], data_r[878:878], data_r[879:879], data_r[880:880], data_r[881:881], data_r[882:882], data_r[883:883], data_r[884:884], data_r[885:885], data_r[886:886], data_r[887:887], data_r[888:888], data_r[889:889], data_r[890:890], data_r[891:891], data_r[892:892], data_r[893:893], data_r[894:894], data_r[895:895] } : 1'b0;
  assign N83 = N2265;
  assign { data_o[896:896], data_o[897:897], data_o[898:898], data_o[899:899], data_o[900:900], data_o[901:901], data_o[902:902], data_o[903:903], data_o[904:904], data_o[905:905], data_o[906:906], data_o[907:907], data_o[908:908], data_o[909:909], data_o[910:910], data_o[911:911], data_o[912:912], data_o[913:913], data_o[914:914], data_o[915:915], data_o[916:916], data_o[917:917], data_o[918:918], data_o[919:919], data_o[920:920], data_o[921:921], data_o[922:922], data_o[923:923], data_o[924:924], data_o[925:925], data_o[926:926], data_o[927:927] } = (N84)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2394)? { data_r[896:896], data_r[897:897], data_r[898:898], data_r[899:899], data_r[900:900], data_r[901:901], data_r[902:902], data_r[903:903], data_r[904:904], data_r[905:905], data_r[906:906], data_r[907:907], data_r[908:908], data_r[909:909], data_r[910:910], data_r[911:911], data_r[912:912], data_r[913:913], data_r[914:914], data_r[915:915], data_r[916:916], data_r[917:917], data_r[918:918], data_r[919:919], data_r[920:920], data_r[921:921], data_r[922:922], data_r[923:923], data_r[924:924], data_r[925:925], data_r[926:926], data_r[927:927] } : 1'b0;
  assign N84 = N2266;
  assign { data_o[928:928], data_o[929:929], data_o[930:930], data_o[931:931], data_o[932:932], data_o[933:933], data_o[934:934], data_o[935:935], data_o[936:936], data_o[937:937], data_o[938:938], data_o[939:939], data_o[940:940], data_o[941:941], data_o[942:942], data_o[943:943], data_o[944:944], data_o[945:945], data_o[946:946], data_o[947:947], data_o[948:948], data_o[949:949], data_o[950:950], data_o[951:951], data_o[952:952], data_o[953:953], data_o[954:954], data_o[955:955], data_o[956:956], data_o[957:957], data_o[958:958], data_o[959:959] } = (N85)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2395)? { data_r[928:928], data_r[929:929], data_r[930:930], data_r[931:931], data_r[932:932], data_r[933:933], data_r[934:934], data_r[935:935], data_r[936:936], data_r[937:937], data_r[938:938], data_r[939:939], data_r[940:940], data_r[941:941], data_r[942:942], data_r[943:943], data_r[944:944], data_r[945:945], data_r[946:946], data_r[947:947], data_r[948:948], data_r[949:949], data_r[950:950], data_r[951:951], data_r[952:952], data_r[953:953], data_r[954:954], data_r[955:955], data_r[956:956], data_r[957:957], data_r[958:958], data_r[959:959] } : 1'b0;
  assign N85 = N2267;
  assign { data_o[960:960], data_o[961:961], data_o[962:962], data_o[963:963], data_o[964:964], data_o[965:965], data_o[966:966], data_o[967:967], data_o[968:968], data_o[969:969], data_o[970:970], data_o[971:971], data_o[972:972], data_o[973:973], data_o[974:974], data_o[975:975], data_o[976:976], data_o[977:977], data_o[978:978], data_o[979:979], data_o[980:980], data_o[981:981], data_o[982:982], data_o[983:983], data_o[984:984], data_o[985:985], data_o[986:986], data_o[987:987], data_o[988:988], data_o[989:989], data_o[990:990], data_o[991:991] } = (N86)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2396)? { data_r[960:960], data_r[961:961], data_r[962:962], data_r[963:963], data_r[964:964], data_r[965:965], data_r[966:966], data_r[967:967], data_r[968:968], data_r[969:969], data_r[970:970], data_r[971:971], data_r[972:972], data_r[973:973], data_r[974:974], data_r[975:975], data_r[976:976], data_r[977:977], data_r[978:978], data_r[979:979], data_r[980:980], data_r[981:981], data_r[982:982], data_r[983:983], data_r[984:984], data_r[985:985], data_r[986:986], data_r[987:987], data_r[988:988], data_r[989:989], data_r[990:990], data_r[991:991] } : 1'b0;
  assign N86 = N2268;
  assign { data_o[992:992], data_o[993:993], data_o[994:994], data_o[995:995], data_o[996:996], data_o[997:997], data_o[998:998], data_o[999:999], data_o[1000:1000], data_o[1001:1001], data_o[1002:1002], data_o[1003:1003], data_o[1004:1004], data_o[1005:1005], data_o[1006:1006], data_o[1007:1007], data_o[1008:1008], data_o[1009:1009], data_o[1010:1010], data_o[1011:1011], data_o[1012:1012], data_o[1013:1013], data_o[1014:1014], data_o[1015:1015], data_o[1016:1016], data_o[1017:1017], data_o[1018:1018], data_o[1019:1019], data_o[1020:1020], data_o[1021:1021], data_o[1022:1022], data_o[1023:1023] } = (N87)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2397)? { data_r[992:992], data_r[993:993], data_r[994:994], data_r[995:995], data_r[996:996], data_r[997:997], data_r[998:998], data_r[999:999], data_r[1000:1000], data_r[1001:1001], data_r[1002:1002], data_r[1003:1003], data_r[1004:1004], data_r[1005:1005], data_r[1006:1006], data_r[1007:1007], data_r[1008:1008], data_r[1009:1009], data_r[1010:1010], data_r[1011:1011], data_r[1012:1012], data_r[1013:1013], data_r[1014:1014], data_r[1015:1015], data_r[1016:1016], data_r[1017:1017], data_r[1018:1018], data_r[1019:1019], data_r[1020:1020], data_r[1021:1021], data_r[1022:1022], data_r[1023:1023] } : 1'b0;
  assign N87 = N2269;
  assign { data_o[1024:1024], data_o[1025:1025], data_o[1026:1026], data_o[1027:1027], data_o[1028:1028], data_o[1029:1029], data_o[1030:1030], data_o[1031:1031], data_o[1032:1032], data_o[1033:1033], data_o[1034:1034], data_o[1035:1035], data_o[1036:1036], data_o[1037:1037], data_o[1038:1038], data_o[1039:1039], data_o[1040:1040], data_o[1041:1041], data_o[1042:1042], data_o[1043:1043], data_o[1044:1044], data_o[1045:1045], data_o[1046:1046], data_o[1047:1047], data_o[1048:1048], data_o[1049:1049], data_o[1050:1050], data_o[1051:1051], data_o[1052:1052], data_o[1053:1053], data_o[1054:1054], data_o[1055:1055] } = (N88)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2398)? { data_r[1024:1024], data_r[1025:1025], data_r[1026:1026], data_r[1027:1027], data_r[1028:1028], data_r[1029:1029], data_r[1030:1030], data_r[1031:1031], data_r[1032:1032], data_r[1033:1033], data_r[1034:1034], data_r[1035:1035], data_r[1036:1036], data_r[1037:1037], data_r[1038:1038], data_r[1039:1039], data_r[1040:1040], data_r[1041:1041], data_r[1042:1042], data_r[1043:1043], data_r[1044:1044], data_r[1045:1045], data_r[1046:1046], data_r[1047:1047], data_r[1048:1048], data_r[1049:1049], data_r[1050:1050], data_r[1051:1051], data_r[1052:1052], data_r[1053:1053], data_r[1054:1054], data_r[1055:1055] } : 1'b0;
  assign N88 = N2270;
  assign { data_o[1056:1056], data_o[1057:1057], data_o[1058:1058], data_o[1059:1059], data_o[1060:1060], data_o[1061:1061], data_o[1062:1062], data_o[1063:1063], data_o[1064:1064], data_o[1065:1065], data_o[1066:1066], data_o[1067:1067], data_o[1068:1068], data_o[1069:1069], data_o[1070:1070], data_o[1071:1071], data_o[1072:1072], data_o[1073:1073], data_o[1074:1074], data_o[1075:1075], data_o[1076:1076], data_o[1077:1077], data_o[1078:1078], data_o[1079:1079], data_o[1080:1080], data_o[1081:1081], data_o[1082:1082], data_o[1083:1083], data_o[1084:1084], data_o[1085:1085], data_o[1086:1086], data_o[1087:1087] } = (N89)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2399)? { data_r[1056:1056], data_r[1057:1057], data_r[1058:1058], data_r[1059:1059], data_r[1060:1060], data_r[1061:1061], data_r[1062:1062], data_r[1063:1063], data_r[1064:1064], data_r[1065:1065], data_r[1066:1066], data_r[1067:1067], data_r[1068:1068], data_r[1069:1069], data_r[1070:1070], data_r[1071:1071], data_r[1072:1072], data_r[1073:1073], data_r[1074:1074], data_r[1075:1075], data_r[1076:1076], data_r[1077:1077], data_r[1078:1078], data_r[1079:1079], data_r[1080:1080], data_r[1081:1081], data_r[1082:1082], data_r[1083:1083], data_r[1084:1084], data_r[1085:1085], data_r[1086:1086], data_r[1087:1087] } : 1'b0;
  assign N89 = N2271;
  assign { data_o[1088:1088], data_o[1089:1089], data_o[1090:1090], data_o[1091:1091], data_o[1092:1092], data_o[1093:1093], data_o[1094:1094], data_o[1095:1095], data_o[1096:1096], data_o[1097:1097], data_o[1098:1098], data_o[1099:1099], data_o[1100:1100], data_o[1101:1101], data_o[1102:1102], data_o[1103:1103], data_o[1104:1104], data_o[1105:1105], data_o[1106:1106], data_o[1107:1107], data_o[1108:1108], data_o[1109:1109], data_o[1110:1110], data_o[1111:1111], data_o[1112:1112], data_o[1113:1113], data_o[1114:1114], data_o[1115:1115], data_o[1116:1116], data_o[1117:1117], data_o[1118:1118], data_o[1119:1119] } = (N90)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2400)? { data_r[1088:1088], data_r[1089:1089], data_r[1090:1090], data_r[1091:1091], data_r[1092:1092], data_r[1093:1093], data_r[1094:1094], data_r[1095:1095], data_r[1096:1096], data_r[1097:1097], data_r[1098:1098], data_r[1099:1099], data_r[1100:1100], data_r[1101:1101], data_r[1102:1102], data_r[1103:1103], data_r[1104:1104], data_r[1105:1105], data_r[1106:1106], data_r[1107:1107], data_r[1108:1108], data_r[1109:1109], data_r[1110:1110], data_r[1111:1111], data_r[1112:1112], data_r[1113:1113], data_r[1114:1114], data_r[1115:1115], data_r[1116:1116], data_r[1117:1117], data_r[1118:1118], data_r[1119:1119] } : 1'b0;
  assign N90 = N2272;
  assign { data_o[1120:1120], data_o[1121:1121], data_o[1122:1122], data_o[1123:1123], data_o[1124:1124], data_o[1125:1125], data_o[1126:1126], data_o[1127:1127], data_o[1128:1128], data_o[1129:1129], data_o[1130:1130], data_o[1131:1131], data_o[1132:1132], data_o[1133:1133], data_o[1134:1134], data_o[1135:1135], data_o[1136:1136], data_o[1137:1137], data_o[1138:1138], data_o[1139:1139], data_o[1140:1140], data_o[1141:1141], data_o[1142:1142], data_o[1143:1143], data_o[1144:1144], data_o[1145:1145], data_o[1146:1146], data_o[1147:1147], data_o[1148:1148], data_o[1149:1149], data_o[1150:1150], data_o[1151:1151] } = (N91)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2401)? { data_r[1120:1120], data_r[1121:1121], data_r[1122:1122], data_r[1123:1123], data_r[1124:1124], data_r[1125:1125], data_r[1126:1126], data_r[1127:1127], data_r[1128:1128], data_r[1129:1129], data_r[1130:1130], data_r[1131:1131], data_r[1132:1132], data_r[1133:1133], data_r[1134:1134], data_r[1135:1135], data_r[1136:1136], data_r[1137:1137], data_r[1138:1138], data_r[1139:1139], data_r[1140:1140], data_r[1141:1141], data_r[1142:1142], data_r[1143:1143], data_r[1144:1144], data_r[1145:1145], data_r[1146:1146], data_r[1147:1147], data_r[1148:1148], data_r[1149:1149], data_r[1150:1150], data_r[1151:1151] } : 1'b0;
  assign N91 = N2273;
  assign { data_o[1152:1152], data_o[1153:1153], data_o[1154:1154], data_o[1155:1155], data_o[1156:1156], data_o[1157:1157], data_o[1158:1158], data_o[1159:1159], data_o[1160:1160], data_o[1161:1161], data_o[1162:1162], data_o[1163:1163], data_o[1164:1164], data_o[1165:1165], data_o[1166:1166], data_o[1167:1167], data_o[1168:1168], data_o[1169:1169], data_o[1170:1170], data_o[1171:1171], data_o[1172:1172], data_o[1173:1173], data_o[1174:1174], data_o[1175:1175], data_o[1176:1176], data_o[1177:1177], data_o[1178:1178], data_o[1179:1179], data_o[1180:1180], data_o[1181:1181], data_o[1182:1182], data_o[1183:1183] } = (N92)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2402)? { data_r[1152:1152], data_r[1153:1153], data_r[1154:1154], data_r[1155:1155], data_r[1156:1156], data_r[1157:1157], data_r[1158:1158], data_r[1159:1159], data_r[1160:1160], data_r[1161:1161], data_r[1162:1162], data_r[1163:1163], data_r[1164:1164], data_r[1165:1165], data_r[1166:1166], data_r[1167:1167], data_r[1168:1168], data_r[1169:1169], data_r[1170:1170], data_r[1171:1171], data_r[1172:1172], data_r[1173:1173], data_r[1174:1174], data_r[1175:1175], data_r[1176:1176], data_r[1177:1177], data_r[1178:1178], data_r[1179:1179], data_r[1180:1180], data_r[1181:1181], data_r[1182:1182], data_r[1183:1183] } : 1'b0;
  assign N92 = N2274;
  assign { data_o[1184:1184], data_o[1185:1185], data_o[1186:1186], data_o[1187:1187], data_o[1188:1188], data_o[1189:1189], data_o[1190:1190], data_o[1191:1191], data_o[1192:1192], data_o[1193:1193], data_o[1194:1194], data_o[1195:1195], data_o[1196:1196], data_o[1197:1197], data_o[1198:1198], data_o[1199:1199], data_o[1200:1200], data_o[1201:1201], data_o[1202:1202], data_o[1203:1203], data_o[1204:1204], data_o[1205:1205], data_o[1206:1206], data_o[1207:1207], data_o[1208:1208], data_o[1209:1209], data_o[1210:1210], data_o[1211:1211], data_o[1212:1212], data_o[1213:1213], data_o[1214:1214], data_o[1215:1215] } = (N93)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2403)? { data_r[1184:1184], data_r[1185:1185], data_r[1186:1186], data_r[1187:1187], data_r[1188:1188], data_r[1189:1189], data_r[1190:1190], data_r[1191:1191], data_r[1192:1192], data_r[1193:1193], data_r[1194:1194], data_r[1195:1195], data_r[1196:1196], data_r[1197:1197], data_r[1198:1198], data_r[1199:1199], data_r[1200:1200], data_r[1201:1201], data_r[1202:1202], data_r[1203:1203], data_r[1204:1204], data_r[1205:1205], data_r[1206:1206], data_r[1207:1207], data_r[1208:1208], data_r[1209:1209], data_r[1210:1210], data_r[1211:1211], data_r[1212:1212], data_r[1213:1213], data_r[1214:1214], data_r[1215:1215] } : 1'b0;
  assign N93 = N2275;
  assign { data_o[1216:1216], data_o[1217:1217], data_o[1218:1218], data_o[1219:1219], data_o[1220:1220], data_o[1221:1221], data_o[1222:1222], data_o[1223:1223], data_o[1224:1224], data_o[1225:1225], data_o[1226:1226], data_o[1227:1227], data_o[1228:1228], data_o[1229:1229], data_o[1230:1230], data_o[1231:1231], data_o[1232:1232], data_o[1233:1233], data_o[1234:1234], data_o[1235:1235], data_o[1236:1236], data_o[1237:1237], data_o[1238:1238], data_o[1239:1239], data_o[1240:1240], data_o[1241:1241], data_o[1242:1242], data_o[1243:1243], data_o[1244:1244], data_o[1245:1245], data_o[1246:1246], data_o[1247:1247] } = (N94)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2404)? { data_r[1216:1216], data_r[1217:1217], data_r[1218:1218], data_r[1219:1219], data_r[1220:1220], data_r[1221:1221], data_r[1222:1222], data_r[1223:1223], data_r[1224:1224], data_r[1225:1225], data_r[1226:1226], data_r[1227:1227], data_r[1228:1228], data_r[1229:1229], data_r[1230:1230], data_r[1231:1231], data_r[1232:1232], data_r[1233:1233], data_r[1234:1234], data_r[1235:1235], data_r[1236:1236], data_r[1237:1237], data_r[1238:1238], data_r[1239:1239], data_r[1240:1240], data_r[1241:1241], data_r[1242:1242], data_r[1243:1243], data_r[1244:1244], data_r[1245:1245], data_r[1246:1246], data_r[1247:1247] } : 1'b0;
  assign N94 = N2276;
  assign { data_o[1248:1248], data_o[1249:1249], data_o[1250:1250], data_o[1251:1251], data_o[1252:1252], data_o[1253:1253], data_o[1254:1254], data_o[1255:1255], data_o[1256:1256], data_o[1257:1257], data_o[1258:1258], data_o[1259:1259], data_o[1260:1260], data_o[1261:1261], data_o[1262:1262], data_o[1263:1263], data_o[1264:1264], data_o[1265:1265], data_o[1266:1266], data_o[1267:1267], data_o[1268:1268], data_o[1269:1269], data_o[1270:1270], data_o[1271:1271], data_o[1272:1272], data_o[1273:1273], data_o[1274:1274], data_o[1275:1275], data_o[1276:1276], data_o[1277:1277], data_o[1278:1278], data_o[1279:1279] } = (N95)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2405)? { data_r[1248:1248], data_r[1249:1249], data_r[1250:1250], data_r[1251:1251], data_r[1252:1252], data_r[1253:1253], data_r[1254:1254], data_r[1255:1255], data_r[1256:1256], data_r[1257:1257], data_r[1258:1258], data_r[1259:1259], data_r[1260:1260], data_r[1261:1261], data_r[1262:1262], data_r[1263:1263], data_r[1264:1264], data_r[1265:1265], data_r[1266:1266], data_r[1267:1267], data_r[1268:1268], data_r[1269:1269], data_r[1270:1270], data_r[1271:1271], data_r[1272:1272], data_r[1273:1273], data_r[1274:1274], data_r[1275:1275], data_r[1276:1276], data_r[1277:1277], data_r[1278:1278], data_r[1279:1279] } : 1'b0;
  assign N95 = N2277;
  assign { data_o[1280:1280], data_o[1281:1281], data_o[1282:1282], data_o[1283:1283], data_o[1284:1284], data_o[1285:1285], data_o[1286:1286], data_o[1287:1287], data_o[1288:1288], data_o[1289:1289], data_o[1290:1290], data_o[1291:1291], data_o[1292:1292], data_o[1293:1293], data_o[1294:1294], data_o[1295:1295], data_o[1296:1296], data_o[1297:1297], data_o[1298:1298], data_o[1299:1299], data_o[1300:1300], data_o[1301:1301], data_o[1302:1302], data_o[1303:1303], data_o[1304:1304], data_o[1305:1305], data_o[1306:1306], data_o[1307:1307], data_o[1308:1308], data_o[1309:1309], data_o[1310:1310], data_o[1311:1311] } = (N96)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2406)? { data_r[1280:1280], data_r[1281:1281], data_r[1282:1282], data_r[1283:1283], data_r[1284:1284], data_r[1285:1285], data_r[1286:1286], data_r[1287:1287], data_r[1288:1288], data_r[1289:1289], data_r[1290:1290], data_r[1291:1291], data_r[1292:1292], data_r[1293:1293], data_r[1294:1294], data_r[1295:1295], data_r[1296:1296], data_r[1297:1297], data_r[1298:1298], data_r[1299:1299], data_r[1300:1300], data_r[1301:1301], data_r[1302:1302], data_r[1303:1303], data_r[1304:1304], data_r[1305:1305], data_r[1306:1306], data_r[1307:1307], data_r[1308:1308], data_r[1309:1309], data_r[1310:1310], data_r[1311:1311] } : 1'b0;
  assign N96 = N2278;
  assign { data_o[1312:1312], data_o[1313:1313], data_o[1314:1314], data_o[1315:1315], data_o[1316:1316], data_o[1317:1317], data_o[1318:1318], data_o[1319:1319], data_o[1320:1320], data_o[1321:1321], data_o[1322:1322], data_o[1323:1323], data_o[1324:1324], data_o[1325:1325], data_o[1326:1326], data_o[1327:1327], data_o[1328:1328], data_o[1329:1329], data_o[1330:1330], data_o[1331:1331], data_o[1332:1332], data_o[1333:1333], data_o[1334:1334], data_o[1335:1335], data_o[1336:1336], data_o[1337:1337], data_o[1338:1338], data_o[1339:1339], data_o[1340:1340], data_o[1341:1341], data_o[1342:1342], data_o[1343:1343] } = (N97)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2407)? { data_r[1312:1312], data_r[1313:1313], data_r[1314:1314], data_r[1315:1315], data_r[1316:1316], data_r[1317:1317], data_r[1318:1318], data_r[1319:1319], data_r[1320:1320], data_r[1321:1321], data_r[1322:1322], data_r[1323:1323], data_r[1324:1324], data_r[1325:1325], data_r[1326:1326], data_r[1327:1327], data_r[1328:1328], data_r[1329:1329], data_r[1330:1330], data_r[1331:1331], data_r[1332:1332], data_r[1333:1333], data_r[1334:1334], data_r[1335:1335], data_r[1336:1336], data_r[1337:1337], data_r[1338:1338], data_r[1339:1339], data_r[1340:1340], data_r[1341:1341], data_r[1342:1342], data_r[1343:1343] } : 1'b0;
  assign N97 = N2279;
  assign { data_o[1344:1344], data_o[1345:1345], data_o[1346:1346], data_o[1347:1347], data_o[1348:1348], data_o[1349:1349], data_o[1350:1350], data_o[1351:1351], data_o[1352:1352], data_o[1353:1353], data_o[1354:1354], data_o[1355:1355], data_o[1356:1356], data_o[1357:1357], data_o[1358:1358], data_o[1359:1359], data_o[1360:1360], data_o[1361:1361], data_o[1362:1362], data_o[1363:1363], data_o[1364:1364], data_o[1365:1365], data_o[1366:1366], data_o[1367:1367], data_o[1368:1368], data_o[1369:1369], data_o[1370:1370], data_o[1371:1371], data_o[1372:1372], data_o[1373:1373], data_o[1374:1374], data_o[1375:1375] } = (N98)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2408)? { data_r[1344:1344], data_r[1345:1345], data_r[1346:1346], data_r[1347:1347], data_r[1348:1348], data_r[1349:1349], data_r[1350:1350], data_r[1351:1351], data_r[1352:1352], data_r[1353:1353], data_r[1354:1354], data_r[1355:1355], data_r[1356:1356], data_r[1357:1357], data_r[1358:1358], data_r[1359:1359], data_r[1360:1360], data_r[1361:1361], data_r[1362:1362], data_r[1363:1363], data_r[1364:1364], data_r[1365:1365], data_r[1366:1366], data_r[1367:1367], data_r[1368:1368], data_r[1369:1369], data_r[1370:1370], data_r[1371:1371], data_r[1372:1372], data_r[1373:1373], data_r[1374:1374], data_r[1375:1375] } : 1'b0;
  assign N98 = N2280;
  assign { data_o[1376:1376], data_o[1377:1377], data_o[1378:1378], data_o[1379:1379], data_o[1380:1380], data_o[1381:1381], data_o[1382:1382], data_o[1383:1383], data_o[1384:1384], data_o[1385:1385], data_o[1386:1386], data_o[1387:1387], data_o[1388:1388], data_o[1389:1389], data_o[1390:1390], data_o[1391:1391], data_o[1392:1392], data_o[1393:1393], data_o[1394:1394], data_o[1395:1395], data_o[1396:1396], data_o[1397:1397], data_o[1398:1398], data_o[1399:1399], data_o[1400:1400], data_o[1401:1401], data_o[1402:1402], data_o[1403:1403], data_o[1404:1404], data_o[1405:1405], data_o[1406:1406], data_o[1407:1407] } = (N99)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2409)? { data_r[1376:1376], data_r[1377:1377], data_r[1378:1378], data_r[1379:1379], data_r[1380:1380], data_r[1381:1381], data_r[1382:1382], data_r[1383:1383], data_r[1384:1384], data_r[1385:1385], data_r[1386:1386], data_r[1387:1387], data_r[1388:1388], data_r[1389:1389], data_r[1390:1390], data_r[1391:1391], data_r[1392:1392], data_r[1393:1393], data_r[1394:1394], data_r[1395:1395], data_r[1396:1396], data_r[1397:1397], data_r[1398:1398], data_r[1399:1399], data_r[1400:1400], data_r[1401:1401], data_r[1402:1402], data_r[1403:1403], data_r[1404:1404], data_r[1405:1405], data_r[1406:1406], data_r[1407:1407] } : 1'b0;
  assign N99 = N2281;
  assign { data_o[1408:1408], data_o[1409:1409], data_o[1410:1410], data_o[1411:1411], data_o[1412:1412], data_o[1413:1413], data_o[1414:1414], data_o[1415:1415], data_o[1416:1416], data_o[1417:1417], data_o[1418:1418], data_o[1419:1419], data_o[1420:1420], data_o[1421:1421], data_o[1422:1422], data_o[1423:1423], data_o[1424:1424], data_o[1425:1425], data_o[1426:1426], data_o[1427:1427], data_o[1428:1428], data_o[1429:1429], data_o[1430:1430], data_o[1431:1431], data_o[1432:1432], data_o[1433:1433], data_o[1434:1434], data_o[1435:1435], data_o[1436:1436], data_o[1437:1437], data_o[1438:1438], data_o[1439:1439] } = (N100)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2410)? { data_r[1408:1408], data_r[1409:1409], data_r[1410:1410], data_r[1411:1411], data_r[1412:1412], data_r[1413:1413], data_r[1414:1414], data_r[1415:1415], data_r[1416:1416], data_r[1417:1417], data_r[1418:1418], data_r[1419:1419], data_r[1420:1420], data_r[1421:1421], data_r[1422:1422], data_r[1423:1423], data_r[1424:1424], data_r[1425:1425], data_r[1426:1426], data_r[1427:1427], data_r[1428:1428], data_r[1429:1429], data_r[1430:1430], data_r[1431:1431], data_r[1432:1432], data_r[1433:1433], data_r[1434:1434], data_r[1435:1435], data_r[1436:1436], data_r[1437:1437], data_r[1438:1438], data_r[1439:1439] } : 1'b0;
  assign N100 = N2282;
  assign { data_o[1440:1440], data_o[1441:1441], data_o[1442:1442], data_o[1443:1443], data_o[1444:1444], data_o[1445:1445], data_o[1446:1446], data_o[1447:1447], data_o[1448:1448], data_o[1449:1449], data_o[1450:1450], data_o[1451:1451], data_o[1452:1452], data_o[1453:1453], data_o[1454:1454], data_o[1455:1455], data_o[1456:1456], data_o[1457:1457], data_o[1458:1458], data_o[1459:1459], data_o[1460:1460], data_o[1461:1461], data_o[1462:1462], data_o[1463:1463], data_o[1464:1464], data_o[1465:1465], data_o[1466:1466], data_o[1467:1467], data_o[1468:1468], data_o[1469:1469], data_o[1470:1470], data_o[1471:1471] } = (N101)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2411)? { data_r[1440:1440], data_r[1441:1441], data_r[1442:1442], data_r[1443:1443], data_r[1444:1444], data_r[1445:1445], data_r[1446:1446], data_r[1447:1447], data_r[1448:1448], data_r[1449:1449], data_r[1450:1450], data_r[1451:1451], data_r[1452:1452], data_r[1453:1453], data_r[1454:1454], data_r[1455:1455], data_r[1456:1456], data_r[1457:1457], data_r[1458:1458], data_r[1459:1459], data_r[1460:1460], data_r[1461:1461], data_r[1462:1462], data_r[1463:1463], data_r[1464:1464], data_r[1465:1465], data_r[1466:1466], data_r[1467:1467], data_r[1468:1468], data_r[1469:1469], data_r[1470:1470], data_r[1471:1471] } : 1'b0;
  assign N101 = N2283;
  assign { data_o[1472:1472], data_o[1473:1473], data_o[1474:1474], data_o[1475:1475], data_o[1476:1476], data_o[1477:1477], data_o[1478:1478], data_o[1479:1479], data_o[1480:1480], data_o[1481:1481], data_o[1482:1482], data_o[1483:1483], data_o[1484:1484], data_o[1485:1485], data_o[1486:1486], data_o[1487:1487], data_o[1488:1488], data_o[1489:1489], data_o[1490:1490], data_o[1491:1491], data_o[1492:1492], data_o[1493:1493], data_o[1494:1494], data_o[1495:1495], data_o[1496:1496], data_o[1497:1497], data_o[1498:1498], data_o[1499:1499], data_o[1500:1500], data_o[1501:1501], data_o[1502:1502], data_o[1503:1503] } = (N102)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2412)? { data_r[1472:1472], data_r[1473:1473], data_r[1474:1474], data_r[1475:1475], data_r[1476:1476], data_r[1477:1477], data_r[1478:1478], data_r[1479:1479], data_r[1480:1480], data_r[1481:1481], data_r[1482:1482], data_r[1483:1483], data_r[1484:1484], data_r[1485:1485], data_r[1486:1486], data_r[1487:1487], data_r[1488:1488], data_r[1489:1489], data_r[1490:1490], data_r[1491:1491], data_r[1492:1492], data_r[1493:1493], data_r[1494:1494], data_r[1495:1495], data_r[1496:1496], data_r[1497:1497], data_r[1498:1498], data_r[1499:1499], data_r[1500:1500], data_r[1501:1501], data_r[1502:1502], data_r[1503:1503] } : 1'b0;
  assign N102 = N2284;
  assign { data_o[1504:1504], data_o[1505:1505], data_o[1506:1506], data_o[1507:1507], data_o[1508:1508], data_o[1509:1509], data_o[1510:1510], data_o[1511:1511], data_o[1512:1512], data_o[1513:1513], data_o[1514:1514], data_o[1515:1515], data_o[1516:1516], data_o[1517:1517], data_o[1518:1518], data_o[1519:1519], data_o[1520:1520], data_o[1521:1521], data_o[1522:1522], data_o[1523:1523], data_o[1524:1524], data_o[1525:1525], data_o[1526:1526], data_o[1527:1527], data_o[1528:1528], data_o[1529:1529], data_o[1530:1530], data_o[1531:1531], data_o[1532:1532], data_o[1533:1533], data_o[1534:1534], data_o[1535:1535] } = (N103)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2413)? { data_r[1504:1504], data_r[1505:1505], data_r[1506:1506], data_r[1507:1507], data_r[1508:1508], data_r[1509:1509], data_r[1510:1510], data_r[1511:1511], data_r[1512:1512], data_r[1513:1513], data_r[1514:1514], data_r[1515:1515], data_r[1516:1516], data_r[1517:1517], data_r[1518:1518], data_r[1519:1519], data_r[1520:1520], data_r[1521:1521], data_r[1522:1522], data_r[1523:1523], data_r[1524:1524], data_r[1525:1525], data_r[1526:1526], data_r[1527:1527], data_r[1528:1528], data_r[1529:1529], data_r[1530:1530], data_r[1531:1531], data_r[1532:1532], data_r[1533:1533], data_r[1534:1534], data_r[1535:1535] } : 1'b0;
  assign N103 = N2285;
  assign { data_o[1536:1536], data_o[1537:1537], data_o[1538:1538], data_o[1539:1539], data_o[1540:1540], data_o[1541:1541], data_o[1542:1542], data_o[1543:1543], data_o[1544:1544], data_o[1545:1545], data_o[1546:1546], data_o[1547:1547], data_o[1548:1548], data_o[1549:1549], data_o[1550:1550], data_o[1551:1551], data_o[1552:1552], data_o[1553:1553], data_o[1554:1554], data_o[1555:1555], data_o[1556:1556], data_o[1557:1557], data_o[1558:1558], data_o[1559:1559], data_o[1560:1560], data_o[1561:1561], data_o[1562:1562], data_o[1563:1563], data_o[1564:1564], data_o[1565:1565], data_o[1566:1566], data_o[1567:1567] } = (N104)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2414)? { data_r[1536:1536], data_r[1537:1537], data_r[1538:1538], data_r[1539:1539], data_r[1540:1540], data_r[1541:1541], data_r[1542:1542], data_r[1543:1543], data_r[1544:1544], data_r[1545:1545], data_r[1546:1546], data_r[1547:1547], data_r[1548:1548], data_r[1549:1549], data_r[1550:1550], data_r[1551:1551], data_r[1552:1552], data_r[1553:1553], data_r[1554:1554], data_r[1555:1555], data_r[1556:1556], data_r[1557:1557], data_r[1558:1558], data_r[1559:1559], data_r[1560:1560], data_r[1561:1561], data_r[1562:1562], data_r[1563:1563], data_r[1564:1564], data_r[1565:1565], data_r[1566:1566], data_r[1567:1567] } : 1'b0;
  assign N104 = N2286;
  assign { data_o[1568:1568], data_o[1569:1569], data_o[1570:1570], data_o[1571:1571], data_o[1572:1572], data_o[1573:1573], data_o[1574:1574], data_o[1575:1575], data_o[1576:1576], data_o[1577:1577], data_o[1578:1578], data_o[1579:1579], data_o[1580:1580], data_o[1581:1581], data_o[1582:1582], data_o[1583:1583], data_o[1584:1584], data_o[1585:1585], data_o[1586:1586], data_o[1587:1587], data_o[1588:1588], data_o[1589:1589], data_o[1590:1590], data_o[1591:1591], data_o[1592:1592], data_o[1593:1593], data_o[1594:1594], data_o[1595:1595], data_o[1596:1596], data_o[1597:1597], data_o[1598:1598], data_o[1599:1599] } = (N105)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2415)? { data_r[1568:1568], data_r[1569:1569], data_r[1570:1570], data_r[1571:1571], data_r[1572:1572], data_r[1573:1573], data_r[1574:1574], data_r[1575:1575], data_r[1576:1576], data_r[1577:1577], data_r[1578:1578], data_r[1579:1579], data_r[1580:1580], data_r[1581:1581], data_r[1582:1582], data_r[1583:1583], data_r[1584:1584], data_r[1585:1585], data_r[1586:1586], data_r[1587:1587], data_r[1588:1588], data_r[1589:1589], data_r[1590:1590], data_r[1591:1591], data_r[1592:1592], data_r[1593:1593], data_r[1594:1594], data_r[1595:1595], data_r[1596:1596], data_r[1597:1597], data_r[1598:1598], data_r[1599:1599] } : 1'b0;
  assign N105 = N2287;
  assign { data_o[1600:1600], data_o[1601:1601], data_o[1602:1602], data_o[1603:1603], data_o[1604:1604], data_o[1605:1605], data_o[1606:1606], data_o[1607:1607], data_o[1608:1608], data_o[1609:1609], data_o[1610:1610], data_o[1611:1611], data_o[1612:1612], data_o[1613:1613], data_o[1614:1614], data_o[1615:1615], data_o[1616:1616], data_o[1617:1617], data_o[1618:1618], data_o[1619:1619], data_o[1620:1620], data_o[1621:1621], data_o[1622:1622], data_o[1623:1623], data_o[1624:1624], data_o[1625:1625], data_o[1626:1626], data_o[1627:1627], data_o[1628:1628], data_o[1629:1629], data_o[1630:1630], data_o[1631:1631] } = (N106)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2416)? { data_r[1600:1600], data_r[1601:1601], data_r[1602:1602], data_r[1603:1603], data_r[1604:1604], data_r[1605:1605], data_r[1606:1606], data_r[1607:1607], data_r[1608:1608], data_r[1609:1609], data_r[1610:1610], data_r[1611:1611], data_r[1612:1612], data_r[1613:1613], data_r[1614:1614], data_r[1615:1615], data_r[1616:1616], data_r[1617:1617], data_r[1618:1618], data_r[1619:1619], data_r[1620:1620], data_r[1621:1621], data_r[1622:1622], data_r[1623:1623], data_r[1624:1624], data_r[1625:1625], data_r[1626:1626], data_r[1627:1627], data_r[1628:1628], data_r[1629:1629], data_r[1630:1630], data_r[1631:1631] } : 1'b0;
  assign N106 = N2288;
  assign { data_o[1632:1632], data_o[1633:1633], data_o[1634:1634], data_o[1635:1635], data_o[1636:1636], data_o[1637:1637], data_o[1638:1638], data_o[1639:1639], data_o[1640:1640], data_o[1641:1641], data_o[1642:1642], data_o[1643:1643], data_o[1644:1644], data_o[1645:1645], data_o[1646:1646], data_o[1647:1647], data_o[1648:1648], data_o[1649:1649], data_o[1650:1650], data_o[1651:1651], data_o[1652:1652], data_o[1653:1653], data_o[1654:1654], data_o[1655:1655], data_o[1656:1656], data_o[1657:1657], data_o[1658:1658], data_o[1659:1659], data_o[1660:1660], data_o[1661:1661], data_o[1662:1662], data_o[1663:1663] } = (N107)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2417)? { data_r[1632:1632], data_r[1633:1633], data_r[1634:1634], data_r[1635:1635], data_r[1636:1636], data_r[1637:1637], data_r[1638:1638], data_r[1639:1639], data_r[1640:1640], data_r[1641:1641], data_r[1642:1642], data_r[1643:1643], data_r[1644:1644], data_r[1645:1645], data_r[1646:1646], data_r[1647:1647], data_r[1648:1648], data_r[1649:1649], data_r[1650:1650], data_r[1651:1651], data_r[1652:1652], data_r[1653:1653], data_r[1654:1654], data_r[1655:1655], data_r[1656:1656], data_r[1657:1657], data_r[1658:1658], data_r[1659:1659], data_r[1660:1660], data_r[1661:1661], data_r[1662:1662], data_r[1663:1663] } : 1'b0;
  assign N107 = N2289;
  assign { data_o[1664:1664], data_o[1665:1665], data_o[1666:1666], data_o[1667:1667], data_o[1668:1668], data_o[1669:1669], data_o[1670:1670], data_o[1671:1671], data_o[1672:1672], data_o[1673:1673], data_o[1674:1674], data_o[1675:1675], data_o[1676:1676], data_o[1677:1677], data_o[1678:1678], data_o[1679:1679], data_o[1680:1680], data_o[1681:1681], data_o[1682:1682], data_o[1683:1683], data_o[1684:1684], data_o[1685:1685], data_o[1686:1686], data_o[1687:1687], data_o[1688:1688], data_o[1689:1689], data_o[1690:1690], data_o[1691:1691], data_o[1692:1692], data_o[1693:1693], data_o[1694:1694], data_o[1695:1695] } = (N108)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2418)? { data_r[1664:1664], data_r[1665:1665], data_r[1666:1666], data_r[1667:1667], data_r[1668:1668], data_r[1669:1669], data_r[1670:1670], data_r[1671:1671], data_r[1672:1672], data_r[1673:1673], data_r[1674:1674], data_r[1675:1675], data_r[1676:1676], data_r[1677:1677], data_r[1678:1678], data_r[1679:1679], data_r[1680:1680], data_r[1681:1681], data_r[1682:1682], data_r[1683:1683], data_r[1684:1684], data_r[1685:1685], data_r[1686:1686], data_r[1687:1687], data_r[1688:1688], data_r[1689:1689], data_r[1690:1690], data_r[1691:1691], data_r[1692:1692], data_r[1693:1693], data_r[1694:1694], data_r[1695:1695] } : 1'b0;
  assign N108 = N2290;
  assign { data_o[1696:1696], data_o[1697:1697], data_o[1698:1698], data_o[1699:1699], data_o[1700:1700], data_o[1701:1701], data_o[1702:1702], data_o[1703:1703], data_o[1704:1704], data_o[1705:1705], data_o[1706:1706], data_o[1707:1707], data_o[1708:1708], data_o[1709:1709], data_o[1710:1710], data_o[1711:1711], data_o[1712:1712], data_o[1713:1713], data_o[1714:1714], data_o[1715:1715], data_o[1716:1716], data_o[1717:1717], data_o[1718:1718], data_o[1719:1719], data_o[1720:1720], data_o[1721:1721], data_o[1722:1722], data_o[1723:1723], data_o[1724:1724], data_o[1725:1725], data_o[1726:1726], data_o[1727:1727] } = (N109)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2419)? { data_r[1696:1696], data_r[1697:1697], data_r[1698:1698], data_r[1699:1699], data_r[1700:1700], data_r[1701:1701], data_r[1702:1702], data_r[1703:1703], data_r[1704:1704], data_r[1705:1705], data_r[1706:1706], data_r[1707:1707], data_r[1708:1708], data_r[1709:1709], data_r[1710:1710], data_r[1711:1711], data_r[1712:1712], data_r[1713:1713], data_r[1714:1714], data_r[1715:1715], data_r[1716:1716], data_r[1717:1717], data_r[1718:1718], data_r[1719:1719], data_r[1720:1720], data_r[1721:1721], data_r[1722:1722], data_r[1723:1723], data_r[1724:1724], data_r[1725:1725], data_r[1726:1726], data_r[1727:1727] } : 1'b0;
  assign N109 = N2291;
  assign { data_o[1728:1728], data_o[1729:1729], data_o[1730:1730], data_o[1731:1731], data_o[1732:1732], data_o[1733:1733], data_o[1734:1734], data_o[1735:1735], data_o[1736:1736], data_o[1737:1737], data_o[1738:1738], data_o[1739:1739], data_o[1740:1740], data_o[1741:1741], data_o[1742:1742], data_o[1743:1743], data_o[1744:1744], data_o[1745:1745], data_o[1746:1746], data_o[1747:1747], data_o[1748:1748], data_o[1749:1749], data_o[1750:1750], data_o[1751:1751], data_o[1752:1752], data_o[1753:1753], data_o[1754:1754], data_o[1755:1755], data_o[1756:1756], data_o[1757:1757], data_o[1758:1758], data_o[1759:1759] } = (N110)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2420)? { data_r[1728:1728], data_r[1729:1729], data_r[1730:1730], data_r[1731:1731], data_r[1732:1732], data_r[1733:1733], data_r[1734:1734], data_r[1735:1735], data_r[1736:1736], data_r[1737:1737], data_r[1738:1738], data_r[1739:1739], data_r[1740:1740], data_r[1741:1741], data_r[1742:1742], data_r[1743:1743], data_r[1744:1744], data_r[1745:1745], data_r[1746:1746], data_r[1747:1747], data_r[1748:1748], data_r[1749:1749], data_r[1750:1750], data_r[1751:1751], data_r[1752:1752], data_r[1753:1753], data_r[1754:1754], data_r[1755:1755], data_r[1756:1756], data_r[1757:1757], data_r[1758:1758], data_r[1759:1759] } : 1'b0;
  assign N110 = N2292;
  assign { data_o[1760:1760], data_o[1761:1761], data_o[1762:1762], data_o[1763:1763], data_o[1764:1764], data_o[1765:1765], data_o[1766:1766], data_o[1767:1767], data_o[1768:1768], data_o[1769:1769], data_o[1770:1770], data_o[1771:1771], data_o[1772:1772], data_o[1773:1773], data_o[1774:1774], data_o[1775:1775], data_o[1776:1776], data_o[1777:1777], data_o[1778:1778], data_o[1779:1779], data_o[1780:1780], data_o[1781:1781], data_o[1782:1782], data_o[1783:1783], data_o[1784:1784], data_o[1785:1785], data_o[1786:1786], data_o[1787:1787], data_o[1788:1788], data_o[1789:1789], data_o[1790:1790], data_o[1791:1791] } = (N111)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2421)? { data_r[1760:1760], data_r[1761:1761], data_r[1762:1762], data_r[1763:1763], data_r[1764:1764], data_r[1765:1765], data_r[1766:1766], data_r[1767:1767], data_r[1768:1768], data_r[1769:1769], data_r[1770:1770], data_r[1771:1771], data_r[1772:1772], data_r[1773:1773], data_r[1774:1774], data_r[1775:1775], data_r[1776:1776], data_r[1777:1777], data_r[1778:1778], data_r[1779:1779], data_r[1780:1780], data_r[1781:1781], data_r[1782:1782], data_r[1783:1783], data_r[1784:1784], data_r[1785:1785], data_r[1786:1786], data_r[1787:1787], data_r[1788:1788], data_r[1789:1789], data_r[1790:1790], data_r[1791:1791] } : 1'b0;
  assign N111 = N2293;
  assign { data_o[1792:1792], data_o[1793:1793], data_o[1794:1794], data_o[1795:1795], data_o[1796:1796], data_o[1797:1797], data_o[1798:1798], data_o[1799:1799], data_o[1800:1800], data_o[1801:1801], data_o[1802:1802], data_o[1803:1803], data_o[1804:1804], data_o[1805:1805], data_o[1806:1806], data_o[1807:1807], data_o[1808:1808], data_o[1809:1809], data_o[1810:1810], data_o[1811:1811], data_o[1812:1812], data_o[1813:1813], data_o[1814:1814], data_o[1815:1815], data_o[1816:1816], data_o[1817:1817], data_o[1818:1818], data_o[1819:1819], data_o[1820:1820], data_o[1821:1821], data_o[1822:1822], data_o[1823:1823] } = (N112)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2422)? { data_r[1792:1792], data_r[1793:1793], data_r[1794:1794], data_r[1795:1795], data_r[1796:1796], data_r[1797:1797], data_r[1798:1798], data_r[1799:1799], data_r[1800:1800], data_r[1801:1801], data_r[1802:1802], data_r[1803:1803], data_r[1804:1804], data_r[1805:1805], data_r[1806:1806], data_r[1807:1807], data_r[1808:1808], data_r[1809:1809], data_r[1810:1810], data_r[1811:1811], data_r[1812:1812], data_r[1813:1813], data_r[1814:1814], data_r[1815:1815], data_r[1816:1816], data_r[1817:1817], data_r[1818:1818], data_r[1819:1819], data_r[1820:1820], data_r[1821:1821], data_r[1822:1822], data_r[1823:1823] } : 1'b0;
  assign N112 = N2294;
  assign { data_o[1824:1824], data_o[1825:1825], data_o[1826:1826], data_o[1827:1827], data_o[1828:1828], data_o[1829:1829], data_o[1830:1830], data_o[1831:1831], data_o[1832:1832], data_o[1833:1833], data_o[1834:1834], data_o[1835:1835], data_o[1836:1836], data_o[1837:1837], data_o[1838:1838], data_o[1839:1839], data_o[1840:1840], data_o[1841:1841], data_o[1842:1842], data_o[1843:1843], data_o[1844:1844], data_o[1845:1845], data_o[1846:1846], data_o[1847:1847], data_o[1848:1848], data_o[1849:1849], data_o[1850:1850], data_o[1851:1851], data_o[1852:1852], data_o[1853:1853], data_o[1854:1854], data_o[1855:1855] } = (N113)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2423)? { data_r[1824:1824], data_r[1825:1825], data_r[1826:1826], data_r[1827:1827], data_r[1828:1828], data_r[1829:1829], data_r[1830:1830], data_r[1831:1831], data_r[1832:1832], data_r[1833:1833], data_r[1834:1834], data_r[1835:1835], data_r[1836:1836], data_r[1837:1837], data_r[1838:1838], data_r[1839:1839], data_r[1840:1840], data_r[1841:1841], data_r[1842:1842], data_r[1843:1843], data_r[1844:1844], data_r[1845:1845], data_r[1846:1846], data_r[1847:1847], data_r[1848:1848], data_r[1849:1849], data_r[1850:1850], data_r[1851:1851], data_r[1852:1852], data_r[1853:1853], data_r[1854:1854], data_r[1855:1855] } : 1'b0;
  assign N113 = N2295;
  assign { data_o[1856:1856], data_o[1857:1857], data_o[1858:1858], data_o[1859:1859], data_o[1860:1860], data_o[1861:1861], data_o[1862:1862], data_o[1863:1863], data_o[1864:1864], data_o[1865:1865], data_o[1866:1866], data_o[1867:1867], data_o[1868:1868], data_o[1869:1869], data_o[1870:1870], data_o[1871:1871], data_o[1872:1872], data_o[1873:1873], data_o[1874:1874], data_o[1875:1875], data_o[1876:1876], data_o[1877:1877], data_o[1878:1878], data_o[1879:1879], data_o[1880:1880], data_o[1881:1881], data_o[1882:1882], data_o[1883:1883], data_o[1884:1884], data_o[1885:1885], data_o[1886:1886], data_o[1887:1887] } = (N114)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2424)? { data_r[1856:1856], data_r[1857:1857], data_r[1858:1858], data_r[1859:1859], data_r[1860:1860], data_r[1861:1861], data_r[1862:1862], data_r[1863:1863], data_r[1864:1864], data_r[1865:1865], data_r[1866:1866], data_r[1867:1867], data_r[1868:1868], data_r[1869:1869], data_r[1870:1870], data_r[1871:1871], data_r[1872:1872], data_r[1873:1873], data_r[1874:1874], data_r[1875:1875], data_r[1876:1876], data_r[1877:1877], data_r[1878:1878], data_r[1879:1879], data_r[1880:1880], data_r[1881:1881], data_r[1882:1882], data_r[1883:1883], data_r[1884:1884], data_r[1885:1885], data_r[1886:1886], data_r[1887:1887] } : 1'b0;
  assign N114 = N2296;
  assign { data_o[1888:1888], data_o[1889:1889], data_o[1890:1890], data_o[1891:1891], data_o[1892:1892], data_o[1893:1893], data_o[1894:1894], data_o[1895:1895], data_o[1896:1896], data_o[1897:1897], data_o[1898:1898], data_o[1899:1899], data_o[1900:1900], data_o[1901:1901], data_o[1902:1902], data_o[1903:1903], data_o[1904:1904], data_o[1905:1905], data_o[1906:1906], data_o[1907:1907], data_o[1908:1908], data_o[1909:1909], data_o[1910:1910], data_o[1911:1911], data_o[1912:1912], data_o[1913:1913], data_o[1914:1914], data_o[1915:1915], data_o[1916:1916], data_o[1917:1917], data_o[1918:1918], data_o[1919:1919] } = (N115)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2425)? { data_r[1888:1888], data_r[1889:1889], data_r[1890:1890], data_r[1891:1891], data_r[1892:1892], data_r[1893:1893], data_r[1894:1894], data_r[1895:1895], data_r[1896:1896], data_r[1897:1897], data_r[1898:1898], data_r[1899:1899], data_r[1900:1900], data_r[1901:1901], data_r[1902:1902], data_r[1903:1903], data_r[1904:1904], data_r[1905:1905], data_r[1906:1906], data_r[1907:1907], data_r[1908:1908], data_r[1909:1909], data_r[1910:1910], data_r[1911:1911], data_r[1912:1912], data_r[1913:1913], data_r[1914:1914], data_r[1915:1915], data_r[1916:1916], data_r[1917:1917], data_r[1918:1918], data_r[1919:1919] } : 1'b0;
  assign N115 = N2297;
  assign { data_o[1920:1920], data_o[1921:1921], data_o[1922:1922], data_o[1923:1923], data_o[1924:1924], data_o[1925:1925], data_o[1926:1926], data_o[1927:1927], data_o[1928:1928], data_o[1929:1929], data_o[1930:1930], data_o[1931:1931], data_o[1932:1932], data_o[1933:1933], data_o[1934:1934], data_o[1935:1935], data_o[1936:1936], data_o[1937:1937], data_o[1938:1938], data_o[1939:1939], data_o[1940:1940], data_o[1941:1941], data_o[1942:1942], data_o[1943:1943], data_o[1944:1944], data_o[1945:1945], data_o[1946:1946], data_o[1947:1947], data_o[1948:1948], data_o[1949:1949], data_o[1950:1950], data_o[1951:1951] } = (N116)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2426)? { data_r[1920:1920], data_r[1921:1921], data_r[1922:1922], data_r[1923:1923], data_r[1924:1924], data_r[1925:1925], data_r[1926:1926], data_r[1927:1927], data_r[1928:1928], data_r[1929:1929], data_r[1930:1930], data_r[1931:1931], data_r[1932:1932], data_r[1933:1933], data_r[1934:1934], data_r[1935:1935], data_r[1936:1936], data_r[1937:1937], data_r[1938:1938], data_r[1939:1939], data_r[1940:1940], data_r[1941:1941], data_r[1942:1942], data_r[1943:1943], data_r[1944:1944], data_r[1945:1945], data_r[1946:1946], data_r[1947:1947], data_r[1948:1948], data_r[1949:1949], data_r[1950:1950], data_r[1951:1951] } : 1'b0;
  assign N116 = N2298;
  assign { data_o[1952:1952], data_o[1953:1953], data_o[1954:1954], data_o[1955:1955], data_o[1956:1956], data_o[1957:1957], data_o[1958:1958], data_o[1959:1959], data_o[1960:1960], data_o[1961:1961], data_o[1962:1962], data_o[1963:1963], data_o[1964:1964], data_o[1965:1965], data_o[1966:1966], data_o[1967:1967], data_o[1968:1968], data_o[1969:1969], data_o[1970:1970], data_o[1971:1971], data_o[1972:1972], data_o[1973:1973], data_o[1974:1974], data_o[1975:1975], data_o[1976:1976], data_o[1977:1977], data_o[1978:1978], data_o[1979:1979], data_o[1980:1980], data_o[1981:1981], data_o[1982:1982], data_o[1983:1983] } = (N117)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2427)? { data_r[1952:1952], data_r[1953:1953], data_r[1954:1954], data_r[1955:1955], data_r[1956:1956], data_r[1957:1957], data_r[1958:1958], data_r[1959:1959], data_r[1960:1960], data_r[1961:1961], data_r[1962:1962], data_r[1963:1963], data_r[1964:1964], data_r[1965:1965], data_r[1966:1966], data_r[1967:1967], data_r[1968:1968], data_r[1969:1969], data_r[1970:1970], data_r[1971:1971], data_r[1972:1972], data_r[1973:1973], data_r[1974:1974], data_r[1975:1975], data_r[1976:1976], data_r[1977:1977], data_r[1978:1978], data_r[1979:1979], data_r[1980:1980], data_r[1981:1981], data_r[1982:1982], data_r[1983:1983] } : 1'b0;
  assign N117 = N2299;
  assign { data_o[1984:1984], data_o[1985:1985], data_o[1986:1986], data_o[1987:1987], data_o[1988:1988], data_o[1989:1989], data_o[1990:1990], data_o[1991:1991], data_o[1992:1992], data_o[1993:1993], data_o[1994:1994], data_o[1995:1995], data_o[1996:1996], data_o[1997:1997], data_o[1998:1998], data_o[1999:1999], data_o[2000:2000], data_o[2001:2001], data_o[2002:2002], data_o[2003:2003], data_o[2004:2004], data_o[2005:2005], data_o[2006:2006], data_o[2007:2007], data_o[2008:2008], data_o[2009:2009], data_o[2010:2010], data_o[2011:2011], data_o[2012:2012], data_o[2013:2013], data_o[2014:2014], data_o[2015:2015] } = (N118)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2428)? { data_r[1984:1984], data_r[1985:1985], data_r[1986:1986], data_r[1987:1987], data_r[1988:1988], data_r[1989:1989], data_r[1990:1990], data_r[1991:1991], data_r[1992:1992], data_r[1993:1993], data_r[1994:1994], data_r[1995:1995], data_r[1996:1996], data_r[1997:1997], data_r[1998:1998], data_r[1999:1999], data_r[2000:2000], data_r[2001:2001], data_r[2002:2002], data_r[2003:2003], data_r[2004:2004], data_r[2005:2005], data_r[2006:2006], data_r[2007:2007], data_r[2008:2008], data_r[2009:2009], data_r[2010:2010], data_r[2011:2011], data_r[2012:2012], data_r[2013:2013], data_r[2014:2014], data_r[2015:2015] } : 1'b0;
  assign N118 = N2300;
  assign { data_o[2016:2016], data_o[2017:2017], data_o[2018:2018], data_o[2019:2019], data_o[2020:2020], data_o[2021:2021], data_o[2022:2022], data_o[2023:2023], data_o[2024:2024], data_o[2025:2025], data_o[2026:2026], data_o[2027:2027], data_o[2028:2028], data_o[2029:2029], data_o[2030:2030], data_o[2031:2031], data_o[2032:2032], data_o[2033:2033], data_o[2034:2034], data_o[2035:2035], data_o[2036:2036], data_o[2037:2037], data_o[2038:2038], data_o[2039:2039], data_o[2040:2040], data_o[2041:2041], data_o[2042:2042], data_o[2043:2043], data_o[2044:2044], data_o[2045:2045], data_o[2046:2046], data_o[2047:2047] } = (N119)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2429)? { data_r[2016:2016], data_r[2017:2017], data_r[2018:2018], data_r[2019:2019], data_r[2020:2020], data_r[2021:2021], data_r[2022:2022], data_r[2023:2023], data_r[2024:2024], data_r[2025:2025], data_r[2026:2026], data_r[2027:2027], data_r[2028:2028], data_r[2029:2029], data_r[2030:2030], data_r[2031:2031], data_r[2032:2032], data_r[2033:2033], data_r[2034:2034], data_r[2035:2035], data_r[2036:2036], data_r[2037:2037], data_r[2038:2038], data_r[2039:2039], data_r[2040:2040], data_r[2041:2041], data_r[2042:2042], data_r[2043:2043], data_r[2044:2044], data_r[2045:2045], data_r[2046:2046], data_r[2047:2047] } : 1'b0;
  assign N119 = N2301;
  assign { data_n_64__0_, data_n_64__1_, data_n_64__2_, data_n_64__3_, data_n_64__4_, data_n_64__5_, data_n_64__6_, data_n_64__7_, data_n_64__8_, data_n_64__9_, data_n_64__10_, data_n_64__11_, data_n_64__12_, data_n_64__13_, data_n_64__14_, data_n_64__15_, data_n_64__16_, data_n_64__17_, data_n_64__18_, data_n_64__19_, data_n_64__20_, data_n_64__21_, data_n_64__22_, data_n_64__23_, data_n_64__24_, data_n_64__25_, data_n_64__26_, data_n_64__27_, data_n_64__28_, data_n_64__29_, data_n_64__30_, data_n_64__31_ } = (N120)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2430)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N120 = N2302;
  assign { data_n_65__0_, data_n_65__1_, data_n_65__2_, data_n_65__3_, data_n_65__4_, data_n_65__5_, data_n_65__6_, data_n_65__7_, data_n_65__8_, data_n_65__9_, data_n_65__10_, data_n_65__11_, data_n_65__12_, data_n_65__13_, data_n_65__14_, data_n_65__15_, data_n_65__16_, data_n_65__17_, data_n_65__18_, data_n_65__19_, data_n_65__20_, data_n_65__21_, data_n_65__22_, data_n_65__23_, data_n_65__24_, data_n_65__25_, data_n_65__26_, data_n_65__27_, data_n_65__28_, data_n_65__29_, data_n_65__30_, data_n_65__31_ } = (N121)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2431)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N121 = N2303;
  assign { data_n_66__0_, data_n_66__1_, data_n_66__2_, data_n_66__3_, data_n_66__4_, data_n_66__5_, data_n_66__6_, data_n_66__7_, data_n_66__8_, data_n_66__9_, data_n_66__10_, data_n_66__11_, data_n_66__12_, data_n_66__13_, data_n_66__14_, data_n_66__15_, data_n_66__16_, data_n_66__17_, data_n_66__18_, data_n_66__19_, data_n_66__20_, data_n_66__21_, data_n_66__22_, data_n_66__23_, data_n_66__24_, data_n_66__25_, data_n_66__26_, data_n_66__27_, data_n_66__28_, data_n_66__29_, data_n_66__30_, data_n_66__31_ } = (N122)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2432)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N122 = N2304;
  assign { data_n_67__0_, data_n_67__1_, data_n_67__2_, data_n_67__3_, data_n_67__4_, data_n_67__5_, data_n_67__6_, data_n_67__7_, data_n_67__8_, data_n_67__9_, data_n_67__10_, data_n_67__11_, data_n_67__12_, data_n_67__13_, data_n_67__14_, data_n_67__15_, data_n_67__16_, data_n_67__17_, data_n_67__18_, data_n_67__19_, data_n_67__20_, data_n_67__21_, data_n_67__22_, data_n_67__23_, data_n_67__24_, data_n_67__25_, data_n_67__26_, data_n_67__27_, data_n_67__28_, data_n_67__29_, data_n_67__30_, data_n_67__31_ } = (N123)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2433)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N123 = N2305;
  assign { data_n_68__0_, data_n_68__1_, data_n_68__2_, data_n_68__3_, data_n_68__4_, data_n_68__5_, data_n_68__6_, data_n_68__7_, data_n_68__8_, data_n_68__9_, data_n_68__10_, data_n_68__11_, data_n_68__12_, data_n_68__13_, data_n_68__14_, data_n_68__15_, data_n_68__16_, data_n_68__17_, data_n_68__18_, data_n_68__19_, data_n_68__20_, data_n_68__21_, data_n_68__22_, data_n_68__23_, data_n_68__24_, data_n_68__25_, data_n_68__26_, data_n_68__27_, data_n_68__28_, data_n_68__29_, data_n_68__30_, data_n_68__31_ } = (N124)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2434)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N124 = N2306;
  assign { data_n_69__0_, data_n_69__1_, data_n_69__2_, data_n_69__3_, data_n_69__4_, data_n_69__5_, data_n_69__6_, data_n_69__7_, data_n_69__8_, data_n_69__9_, data_n_69__10_, data_n_69__11_, data_n_69__12_, data_n_69__13_, data_n_69__14_, data_n_69__15_, data_n_69__16_, data_n_69__17_, data_n_69__18_, data_n_69__19_, data_n_69__20_, data_n_69__21_, data_n_69__22_, data_n_69__23_, data_n_69__24_, data_n_69__25_, data_n_69__26_, data_n_69__27_, data_n_69__28_, data_n_69__29_, data_n_69__30_, data_n_69__31_ } = (N125)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2435)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N125 = N2307;
  assign { data_n_70__0_, data_n_70__1_, data_n_70__2_, data_n_70__3_, data_n_70__4_, data_n_70__5_, data_n_70__6_, data_n_70__7_, data_n_70__8_, data_n_70__9_, data_n_70__10_, data_n_70__11_, data_n_70__12_, data_n_70__13_, data_n_70__14_, data_n_70__15_, data_n_70__16_, data_n_70__17_, data_n_70__18_, data_n_70__19_, data_n_70__20_, data_n_70__21_, data_n_70__22_, data_n_70__23_, data_n_70__24_, data_n_70__25_, data_n_70__26_, data_n_70__27_, data_n_70__28_, data_n_70__29_, data_n_70__30_, data_n_70__31_ } = (N126)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2436)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N126 = N2308;
  assign { data_n_71__0_, data_n_71__1_, data_n_71__2_, data_n_71__3_, data_n_71__4_, data_n_71__5_, data_n_71__6_, data_n_71__7_, data_n_71__8_, data_n_71__9_, data_n_71__10_, data_n_71__11_, data_n_71__12_, data_n_71__13_, data_n_71__14_, data_n_71__15_, data_n_71__16_, data_n_71__17_, data_n_71__18_, data_n_71__19_, data_n_71__20_, data_n_71__21_, data_n_71__22_, data_n_71__23_, data_n_71__24_, data_n_71__25_, data_n_71__26_, data_n_71__27_, data_n_71__28_, data_n_71__29_, data_n_71__30_, data_n_71__31_ } = (N127)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2437)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N127 = N2309;
  assign { data_n_72__0_, data_n_72__1_, data_n_72__2_, data_n_72__3_, data_n_72__4_, data_n_72__5_, data_n_72__6_, data_n_72__7_, data_n_72__8_, data_n_72__9_, data_n_72__10_, data_n_72__11_, data_n_72__12_, data_n_72__13_, data_n_72__14_, data_n_72__15_, data_n_72__16_, data_n_72__17_, data_n_72__18_, data_n_72__19_, data_n_72__20_, data_n_72__21_, data_n_72__22_, data_n_72__23_, data_n_72__24_, data_n_72__25_, data_n_72__26_, data_n_72__27_, data_n_72__28_, data_n_72__29_, data_n_72__30_, data_n_72__31_ } = (N128)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2438)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N128 = N2310;
  assign { data_n_73__0_, data_n_73__1_, data_n_73__2_, data_n_73__3_, data_n_73__4_, data_n_73__5_, data_n_73__6_, data_n_73__7_, data_n_73__8_, data_n_73__9_, data_n_73__10_, data_n_73__11_, data_n_73__12_, data_n_73__13_, data_n_73__14_, data_n_73__15_, data_n_73__16_, data_n_73__17_, data_n_73__18_, data_n_73__19_, data_n_73__20_, data_n_73__21_, data_n_73__22_, data_n_73__23_, data_n_73__24_, data_n_73__25_, data_n_73__26_, data_n_73__27_, data_n_73__28_, data_n_73__29_, data_n_73__30_, data_n_73__31_ } = (N129)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2439)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N129 = N2311;
  assign { data_n_74__0_, data_n_74__1_, data_n_74__2_, data_n_74__3_, data_n_74__4_, data_n_74__5_, data_n_74__6_, data_n_74__7_, data_n_74__8_, data_n_74__9_, data_n_74__10_, data_n_74__11_, data_n_74__12_, data_n_74__13_, data_n_74__14_, data_n_74__15_, data_n_74__16_, data_n_74__17_, data_n_74__18_, data_n_74__19_, data_n_74__20_, data_n_74__21_, data_n_74__22_, data_n_74__23_, data_n_74__24_, data_n_74__25_, data_n_74__26_, data_n_74__27_, data_n_74__28_, data_n_74__29_, data_n_74__30_, data_n_74__31_ } = (N130)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2440)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N130 = N2312;
  assign { data_n_75__0_, data_n_75__1_, data_n_75__2_, data_n_75__3_, data_n_75__4_, data_n_75__5_, data_n_75__6_, data_n_75__7_, data_n_75__8_, data_n_75__9_, data_n_75__10_, data_n_75__11_, data_n_75__12_, data_n_75__13_, data_n_75__14_, data_n_75__15_, data_n_75__16_, data_n_75__17_, data_n_75__18_, data_n_75__19_, data_n_75__20_, data_n_75__21_, data_n_75__22_, data_n_75__23_, data_n_75__24_, data_n_75__25_, data_n_75__26_, data_n_75__27_, data_n_75__28_, data_n_75__29_, data_n_75__30_, data_n_75__31_ } = (N131)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2441)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N131 = N2313;
  assign { data_n_76__0_, data_n_76__1_, data_n_76__2_, data_n_76__3_, data_n_76__4_, data_n_76__5_, data_n_76__6_, data_n_76__7_, data_n_76__8_, data_n_76__9_, data_n_76__10_, data_n_76__11_, data_n_76__12_, data_n_76__13_, data_n_76__14_, data_n_76__15_, data_n_76__16_, data_n_76__17_, data_n_76__18_, data_n_76__19_, data_n_76__20_, data_n_76__21_, data_n_76__22_, data_n_76__23_, data_n_76__24_, data_n_76__25_, data_n_76__26_, data_n_76__27_, data_n_76__28_, data_n_76__29_, data_n_76__30_, data_n_76__31_ } = (N132)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2442)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N132 = N2314;
  assign { data_n_77__0_, data_n_77__1_, data_n_77__2_, data_n_77__3_, data_n_77__4_, data_n_77__5_, data_n_77__6_, data_n_77__7_, data_n_77__8_, data_n_77__9_, data_n_77__10_, data_n_77__11_, data_n_77__12_, data_n_77__13_, data_n_77__14_, data_n_77__15_, data_n_77__16_, data_n_77__17_, data_n_77__18_, data_n_77__19_, data_n_77__20_, data_n_77__21_, data_n_77__22_, data_n_77__23_, data_n_77__24_, data_n_77__25_, data_n_77__26_, data_n_77__27_, data_n_77__28_, data_n_77__29_, data_n_77__30_, data_n_77__31_ } = (N133)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2443)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N133 = N2315;
  assign { data_n_78__0_, data_n_78__1_, data_n_78__2_, data_n_78__3_, data_n_78__4_, data_n_78__5_, data_n_78__6_, data_n_78__7_, data_n_78__8_, data_n_78__9_, data_n_78__10_, data_n_78__11_, data_n_78__12_, data_n_78__13_, data_n_78__14_, data_n_78__15_, data_n_78__16_, data_n_78__17_, data_n_78__18_, data_n_78__19_, data_n_78__20_, data_n_78__21_, data_n_78__22_, data_n_78__23_, data_n_78__24_, data_n_78__25_, data_n_78__26_, data_n_78__27_, data_n_78__28_, data_n_78__29_, data_n_78__30_, data_n_78__31_ } = (N134)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2444)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N134 = N2316;
  assign { data_n_79__0_, data_n_79__1_, data_n_79__2_, data_n_79__3_, data_n_79__4_, data_n_79__5_, data_n_79__6_, data_n_79__7_, data_n_79__8_, data_n_79__9_, data_n_79__10_, data_n_79__11_, data_n_79__12_, data_n_79__13_, data_n_79__14_, data_n_79__15_, data_n_79__16_, data_n_79__17_, data_n_79__18_, data_n_79__19_, data_n_79__20_, data_n_79__21_, data_n_79__22_, data_n_79__23_, data_n_79__24_, data_n_79__25_, data_n_79__26_, data_n_79__27_, data_n_79__28_, data_n_79__29_, data_n_79__30_, data_n_79__31_ } = (N135)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2445)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N135 = N2317;
  assign { data_n_80__0_, data_n_80__1_, data_n_80__2_, data_n_80__3_, data_n_80__4_, data_n_80__5_, data_n_80__6_, data_n_80__7_, data_n_80__8_, data_n_80__9_, data_n_80__10_, data_n_80__11_, data_n_80__12_, data_n_80__13_, data_n_80__14_, data_n_80__15_, data_n_80__16_, data_n_80__17_, data_n_80__18_, data_n_80__19_, data_n_80__20_, data_n_80__21_, data_n_80__22_, data_n_80__23_, data_n_80__24_, data_n_80__25_, data_n_80__26_, data_n_80__27_, data_n_80__28_, data_n_80__29_, data_n_80__30_, data_n_80__31_ } = (N136)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2446)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N136 = N2318;
  assign { data_n_81__0_, data_n_81__1_, data_n_81__2_, data_n_81__3_, data_n_81__4_, data_n_81__5_, data_n_81__6_, data_n_81__7_, data_n_81__8_, data_n_81__9_, data_n_81__10_, data_n_81__11_, data_n_81__12_, data_n_81__13_, data_n_81__14_, data_n_81__15_, data_n_81__16_, data_n_81__17_, data_n_81__18_, data_n_81__19_, data_n_81__20_, data_n_81__21_, data_n_81__22_, data_n_81__23_, data_n_81__24_, data_n_81__25_, data_n_81__26_, data_n_81__27_, data_n_81__28_, data_n_81__29_, data_n_81__30_, data_n_81__31_ } = (N137)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2447)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N137 = N2319;
  assign { data_n_82__0_, data_n_82__1_, data_n_82__2_, data_n_82__3_, data_n_82__4_, data_n_82__5_, data_n_82__6_, data_n_82__7_, data_n_82__8_, data_n_82__9_, data_n_82__10_, data_n_82__11_, data_n_82__12_, data_n_82__13_, data_n_82__14_, data_n_82__15_, data_n_82__16_, data_n_82__17_, data_n_82__18_, data_n_82__19_, data_n_82__20_, data_n_82__21_, data_n_82__22_, data_n_82__23_, data_n_82__24_, data_n_82__25_, data_n_82__26_, data_n_82__27_, data_n_82__28_, data_n_82__29_, data_n_82__30_, data_n_82__31_ } = (N138)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2448)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N138 = N2320;
  assign { data_n_83__0_, data_n_83__1_, data_n_83__2_, data_n_83__3_, data_n_83__4_, data_n_83__5_, data_n_83__6_, data_n_83__7_, data_n_83__8_, data_n_83__9_, data_n_83__10_, data_n_83__11_, data_n_83__12_, data_n_83__13_, data_n_83__14_, data_n_83__15_, data_n_83__16_, data_n_83__17_, data_n_83__18_, data_n_83__19_, data_n_83__20_, data_n_83__21_, data_n_83__22_, data_n_83__23_, data_n_83__24_, data_n_83__25_, data_n_83__26_, data_n_83__27_, data_n_83__28_, data_n_83__29_, data_n_83__30_, data_n_83__31_ } = (N139)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2449)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N139 = N2321;
  assign { data_n_84__0_, data_n_84__1_, data_n_84__2_, data_n_84__3_, data_n_84__4_, data_n_84__5_, data_n_84__6_, data_n_84__7_, data_n_84__8_, data_n_84__9_, data_n_84__10_, data_n_84__11_, data_n_84__12_, data_n_84__13_, data_n_84__14_, data_n_84__15_, data_n_84__16_, data_n_84__17_, data_n_84__18_, data_n_84__19_, data_n_84__20_, data_n_84__21_, data_n_84__22_, data_n_84__23_, data_n_84__24_, data_n_84__25_, data_n_84__26_, data_n_84__27_, data_n_84__28_, data_n_84__29_, data_n_84__30_, data_n_84__31_ } = (N140)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2450)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N140 = N2322;
  assign { data_n_85__0_, data_n_85__1_, data_n_85__2_, data_n_85__3_, data_n_85__4_, data_n_85__5_, data_n_85__6_, data_n_85__7_, data_n_85__8_, data_n_85__9_, data_n_85__10_, data_n_85__11_, data_n_85__12_, data_n_85__13_, data_n_85__14_, data_n_85__15_, data_n_85__16_, data_n_85__17_, data_n_85__18_, data_n_85__19_, data_n_85__20_, data_n_85__21_, data_n_85__22_, data_n_85__23_, data_n_85__24_, data_n_85__25_, data_n_85__26_, data_n_85__27_, data_n_85__28_, data_n_85__29_, data_n_85__30_, data_n_85__31_ } = (N141)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2451)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N141 = N2323;
  assign { data_n_86__0_, data_n_86__1_, data_n_86__2_, data_n_86__3_, data_n_86__4_, data_n_86__5_, data_n_86__6_, data_n_86__7_, data_n_86__8_, data_n_86__9_, data_n_86__10_, data_n_86__11_, data_n_86__12_, data_n_86__13_, data_n_86__14_, data_n_86__15_, data_n_86__16_, data_n_86__17_, data_n_86__18_, data_n_86__19_, data_n_86__20_, data_n_86__21_, data_n_86__22_, data_n_86__23_, data_n_86__24_, data_n_86__25_, data_n_86__26_, data_n_86__27_, data_n_86__28_, data_n_86__29_, data_n_86__30_, data_n_86__31_ } = (N142)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2452)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N142 = N2324;
  assign { data_n_87__0_, data_n_87__1_, data_n_87__2_, data_n_87__3_, data_n_87__4_, data_n_87__5_, data_n_87__6_, data_n_87__7_, data_n_87__8_, data_n_87__9_, data_n_87__10_, data_n_87__11_, data_n_87__12_, data_n_87__13_, data_n_87__14_, data_n_87__15_, data_n_87__16_, data_n_87__17_, data_n_87__18_, data_n_87__19_, data_n_87__20_, data_n_87__21_, data_n_87__22_, data_n_87__23_, data_n_87__24_, data_n_87__25_, data_n_87__26_, data_n_87__27_, data_n_87__28_, data_n_87__29_, data_n_87__30_, data_n_87__31_ } = (N143)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2453)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N143 = N2325;
  assign { data_n_88__0_, data_n_88__1_, data_n_88__2_, data_n_88__3_, data_n_88__4_, data_n_88__5_, data_n_88__6_, data_n_88__7_, data_n_88__8_, data_n_88__9_, data_n_88__10_, data_n_88__11_, data_n_88__12_, data_n_88__13_, data_n_88__14_, data_n_88__15_, data_n_88__16_, data_n_88__17_, data_n_88__18_, data_n_88__19_, data_n_88__20_, data_n_88__21_, data_n_88__22_, data_n_88__23_, data_n_88__24_, data_n_88__25_, data_n_88__26_, data_n_88__27_, data_n_88__28_, data_n_88__29_, data_n_88__30_, data_n_88__31_ } = (N144)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2454)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N144 = N2326;
  assign { data_n_89__0_, data_n_89__1_, data_n_89__2_, data_n_89__3_, data_n_89__4_, data_n_89__5_, data_n_89__6_, data_n_89__7_, data_n_89__8_, data_n_89__9_, data_n_89__10_, data_n_89__11_, data_n_89__12_, data_n_89__13_, data_n_89__14_, data_n_89__15_, data_n_89__16_, data_n_89__17_, data_n_89__18_, data_n_89__19_, data_n_89__20_, data_n_89__21_, data_n_89__22_, data_n_89__23_, data_n_89__24_, data_n_89__25_, data_n_89__26_, data_n_89__27_, data_n_89__28_, data_n_89__29_, data_n_89__30_, data_n_89__31_ } = (N145)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2455)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N145 = N2327;
  assign { data_n_90__0_, data_n_90__1_, data_n_90__2_, data_n_90__3_, data_n_90__4_, data_n_90__5_, data_n_90__6_, data_n_90__7_, data_n_90__8_, data_n_90__9_, data_n_90__10_, data_n_90__11_, data_n_90__12_, data_n_90__13_, data_n_90__14_, data_n_90__15_, data_n_90__16_, data_n_90__17_, data_n_90__18_, data_n_90__19_, data_n_90__20_, data_n_90__21_, data_n_90__22_, data_n_90__23_, data_n_90__24_, data_n_90__25_, data_n_90__26_, data_n_90__27_, data_n_90__28_, data_n_90__29_, data_n_90__30_, data_n_90__31_ } = (N146)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2456)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N146 = N2328;
  assign { data_n_91__0_, data_n_91__1_, data_n_91__2_, data_n_91__3_, data_n_91__4_, data_n_91__5_, data_n_91__6_, data_n_91__7_, data_n_91__8_, data_n_91__9_, data_n_91__10_, data_n_91__11_, data_n_91__12_, data_n_91__13_, data_n_91__14_, data_n_91__15_, data_n_91__16_, data_n_91__17_, data_n_91__18_, data_n_91__19_, data_n_91__20_, data_n_91__21_, data_n_91__22_, data_n_91__23_, data_n_91__24_, data_n_91__25_, data_n_91__26_, data_n_91__27_, data_n_91__28_, data_n_91__29_, data_n_91__30_, data_n_91__31_ } = (N147)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2457)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N147 = N2329;
  assign { data_n_92__0_, data_n_92__1_, data_n_92__2_, data_n_92__3_, data_n_92__4_, data_n_92__5_, data_n_92__6_, data_n_92__7_, data_n_92__8_, data_n_92__9_, data_n_92__10_, data_n_92__11_, data_n_92__12_, data_n_92__13_, data_n_92__14_, data_n_92__15_, data_n_92__16_, data_n_92__17_, data_n_92__18_, data_n_92__19_, data_n_92__20_, data_n_92__21_, data_n_92__22_, data_n_92__23_, data_n_92__24_, data_n_92__25_, data_n_92__26_, data_n_92__27_, data_n_92__28_, data_n_92__29_, data_n_92__30_, data_n_92__31_ } = (N148)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2458)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N148 = N2330;
  assign { data_n_93__0_, data_n_93__1_, data_n_93__2_, data_n_93__3_, data_n_93__4_, data_n_93__5_, data_n_93__6_, data_n_93__7_, data_n_93__8_, data_n_93__9_, data_n_93__10_, data_n_93__11_, data_n_93__12_, data_n_93__13_, data_n_93__14_, data_n_93__15_, data_n_93__16_, data_n_93__17_, data_n_93__18_, data_n_93__19_, data_n_93__20_, data_n_93__21_, data_n_93__22_, data_n_93__23_, data_n_93__24_, data_n_93__25_, data_n_93__26_, data_n_93__27_, data_n_93__28_, data_n_93__29_, data_n_93__30_, data_n_93__31_ } = (N149)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2459)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N149 = N2331;
  assign { data_n_94__0_, data_n_94__1_, data_n_94__2_, data_n_94__3_, data_n_94__4_, data_n_94__5_, data_n_94__6_, data_n_94__7_, data_n_94__8_, data_n_94__9_, data_n_94__10_, data_n_94__11_, data_n_94__12_, data_n_94__13_, data_n_94__14_, data_n_94__15_, data_n_94__16_, data_n_94__17_, data_n_94__18_, data_n_94__19_, data_n_94__20_, data_n_94__21_, data_n_94__22_, data_n_94__23_, data_n_94__24_, data_n_94__25_, data_n_94__26_, data_n_94__27_, data_n_94__28_, data_n_94__29_, data_n_94__30_, data_n_94__31_ } = (N150)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2460)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N150 = N2332;
  assign { data_n_95__0_, data_n_95__1_, data_n_95__2_, data_n_95__3_, data_n_95__4_, data_n_95__5_, data_n_95__6_, data_n_95__7_, data_n_95__8_, data_n_95__9_, data_n_95__10_, data_n_95__11_, data_n_95__12_, data_n_95__13_, data_n_95__14_, data_n_95__15_, data_n_95__16_, data_n_95__17_, data_n_95__18_, data_n_95__19_, data_n_95__20_, data_n_95__21_, data_n_95__22_, data_n_95__23_, data_n_95__24_, data_n_95__25_, data_n_95__26_, data_n_95__27_, data_n_95__28_, data_n_95__29_, data_n_95__30_, data_n_95__31_ } = (N151)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2461)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N151 = N2333;
  assign { data_n_96__0_, data_n_96__1_, data_n_96__2_, data_n_96__3_, data_n_96__4_, data_n_96__5_, data_n_96__6_, data_n_96__7_, data_n_96__8_, data_n_96__9_, data_n_96__10_, data_n_96__11_, data_n_96__12_, data_n_96__13_, data_n_96__14_, data_n_96__15_, data_n_96__16_, data_n_96__17_, data_n_96__18_, data_n_96__19_, data_n_96__20_, data_n_96__21_, data_n_96__22_, data_n_96__23_, data_n_96__24_, data_n_96__25_, data_n_96__26_, data_n_96__27_, data_n_96__28_, data_n_96__29_, data_n_96__30_, data_n_96__31_ } = (N152)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2462)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N152 = N2334;
  assign { data_n_97__0_, data_n_97__1_, data_n_97__2_, data_n_97__3_, data_n_97__4_, data_n_97__5_, data_n_97__6_, data_n_97__7_, data_n_97__8_, data_n_97__9_, data_n_97__10_, data_n_97__11_, data_n_97__12_, data_n_97__13_, data_n_97__14_, data_n_97__15_, data_n_97__16_, data_n_97__17_, data_n_97__18_, data_n_97__19_, data_n_97__20_, data_n_97__21_, data_n_97__22_, data_n_97__23_, data_n_97__24_, data_n_97__25_, data_n_97__26_, data_n_97__27_, data_n_97__28_, data_n_97__29_, data_n_97__30_, data_n_97__31_ } = (N153)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2463)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N153 = N2335;
  assign { data_n_98__0_, data_n_98__1_, data_n_98__2_, data_n_98__3_, data_n_98__4_, data_n_98__5_, data_n_98__6_, data_n_98__7_, data_n_98__8_, data_n_98__9_, data_n_98__10_, data_n_98__11_, data_n_98__12_, data_n_98__13_, data_n_98__14_, data_n_98__15_, data_n_98__16_, data_n_98__17_, data_n_98__18_, data_n_98__19_, data_n_98__20_, data_n_98__21_, data_n_98__22_, data_n_98__23_, data_n_98__24_, data_n_98__25_, data_n_98__26_, data_n_98__27_, data_n_98__28_, data_n_98__29_, data_n_98__30_, data_n_98__31_ } = (N154)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2464)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N154 = N2336;
  assign { data_n_99__0_, data_n_99__1_, data_n_99__2_, data_n_99__3_, data_n_99__4_, data_n_99__5_, data_n_99__6_, data_n_99__7_, data_n_99__8_, data_n_99__9_, data_n_99__10_, data_n_99__11_, data_n_99__12_, data_n_99__13_, data_n_99__14_, data_n_99__15_, data_n_99__16_, data_n_99__17_, data_n_99__18_, data_n_99__19_, data_n_99__20_, data_n_99__21_, data_n_99__22_, data_n_99__23_, data_n_99__24_, data_n_99__25_, data_n_99__26_, data_n_99__27_, data_n_99__28_, data_n_99__29_, data_n_99__30_, data_n_99__31_ } = (N155)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2465)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N155 = N2337;
  assign { data_n_100__0_, data_n_100__1_, data_n_100__2_, data_n_100__3_, data_n_100__4_, data_n_100__5_, data_n_100__6_, data_n_100__7_, data_n_100__8_, data_n_100__9_, data_n_100__10_, data_n_100__11_, data_n_100__12_, data_n_100__13_, data_n_100__14_, data_n_100__15_, data_n_100__16_, data_n_100__17_, data_n_100__18_, data_n_100__19_, data_n_100__20_, data_n_100__21_, data_n_100__22_, data_n_100__23_, data_n_100__24_, data_n_100__25_, data_n_100__26_, data_n_100__27_, data_n_100__28_, data_n_100__29_, data_n_100__30_, data_n_100__31_ } = (N156)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2466)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N156 = N2338;
  assign { data_n_101__0_, data_n_101__1_, data_n_101__2_, data_n_101__3_, data_n_101__4_, data_n_101__5_, data_n_101__6_, data_n_101__7_, data_n_101__8_, data_n_101__9_, data_n_101__10_, data_n_101__11_, data_n_101__12_, data_n_101__13_, data_n_101__14_, data_n_101__15_, data_n_101__16_, data_n_101__17_, data_n_101__18_, data_n_101__19_, data_n_101__20_, data_n_101__21_, data_n_101__22_, data_n_101__23_, data_n_101__24_, data_n_101__25_, data_n_101__26_, data_n_101__27_, data_n_101__28_, data_n_101__29_, data_n_101__30_, data_n_101__31_ } = (N157)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2467)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N157 = N2339;
  assign { data_n_102__0_, data_n_102__1_, data_n_102__2_, data_n_102__3_, data_n_102__4_, data_n_102__5_, data_n_102__6_, data_n_102__7_, data_n_102__8_, data_n_102__9_, data_n_102__10_, data_n_102__11_, data_n_102__12_, data_n_102__13_, data_n_102__14_, data_n_102__15_, data_n_102__16_, data_n_102__17_, data_n_102__18_, data_n_102__19_, data_n_102__20_, data_n_102__21_, data_n_102__22_, data_n_102__23_, data_n_102__24_, data_n_102__25_, data_n_102__26_, data_n_102__27_, data_n_102__28_, data_n_102__29_, data_n_102__30_, data_n_102__31_ } = (N158)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2468)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N158 = N2340;
  assign { data_n_103__0_, data_n_103__1_, data_n_103__2_, data_n_103__3_, data_n_103__4_, data_n_103__5_, data_n_103__6_, data_n_103__7_, data_n_103__8_, data_n_103__9_, data_n_103__10_, data_n_103__11_, data_n_103__12_, data_n_103__13_, data_n_103__14_, data_n_103__15_, data_n_103__16_, data_n_103__17_, data_n_103__18_, data_n_103__19_, data_n_103__20_, data_n_103__21_, data_n_103__22_, data_n_103__23_, data_n_103__24_, data_n_103__25_, data_n_103__26_, data_n_103__27_, data_n_103__28_, data_n_103__29_, data_n_103__30_, data_n_103__31_ } = (N159)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2469)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N159 = N2341;
  assign { data_n_104__0_, data_n_104__1_, data_n_104__2_, data_n_104__3_, data_n_104__4_, data_n_104__5_, data_n_104__6_, data_n_104__7_, data_n_104__8_, data_n_104__9_, data_n_104__10_, data_n_104__11_, data_n_104__12_, data_n_104__13_, data_n_104__14_, data_n_104__15_, data_n_104__16_, data_n_104__17_, data_n_104__18_, data_n_104__19_, data_n_104__20_, data_n_104__21_, data_n_104__22_, data_n_104__23_, data_n_104__24_, data_n_104__25_, data_n_104__26_, data_n_104__27_, data_n_104__28_, data_n_104__29_, data_n_104__30_, data_n_104__31_ } = (N160)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2470)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N160 = N2342;
  assign { data_n_105__0_, data_n_105__1_, data_n_105__2_, data_n_105__3_, data_n_105__4_, data_n_105__5_, data_n_105__6_, data_n_105__7_, data_n_105__8_, data_n_105__9_, data_n_105__10_, data_n_105__11_, data_n_105__12_, data_n_105__13_, data_n_105__14_, data_n_105__15_, data_n_105__16_, data_n_105__17_, data_n_105__18_, data_n_105__19_, data_n_105__20_, data_n_105__21_, data_n_105__22_, data_n_105__23_, data_n_105__24_, data_n_105__25_, data_n_105__26_, data_n_105__27_, data_n_105__28_, data_n_105__29_, data_n_105__30_, data_n_105__31_ } = (N161)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2471)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N161 = N2343;
  assign { data_n_106__0_, data_n_106__1_, data_n_106__2_, data_n_106__3_, data_n_106__4_, data_n_106__5_, data_n_106__6_, data_n_106__7_, data_n_106__8_, data_n_106__9_, data_n_106__10_, data_n_106__11_, data_n_106__12_, data_n_106__13_, data_n_106__14_, data_n_106__15_, data_n_106__16_, data_n_106__17_, data_n_106__18_, data_n_106__19_, data_n_106__20_, data_n_106__21_, data_n_106__22_, data_n_106__23_, data_n_106__24_, data_n_106__25_, data_n_106__26_, data_n_106__27_, data_n_106__28_, data_n_106__29_, data_n_106__30_, data_n_106__31_ } = (N162)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2472)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N162 = N2344;
  assign { data_n_107__0_, data_n_107__1_, data_n_107__2_, data_n_107__3_, data_n_107__4_, data_n_107__5_, data_n_107__6_, data_n_107__7_, data_n_107__8_, data_n_107__9_, data_n_107__10_, data_n_107__11_, data_n_107__12_, data_n_107__13_, data_n_107__14_, data_n_107__15_, data_n_107__16_, data_n_107__17_, data_n_107__18_, data_n_107__19_, data_n_107__20_, data_n_107__21_, data_n_107__22_, data_n_107__23_, data_n_107__24_, data_n_107__25_, data_n_107__26_, data_n_107__27_, data_n_107__28_, data_n_107__29_, data_n_107__30_, data_n_107__31_ } = (N163)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2473)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N163 = N2345;
  assign { data_n_108__0_, data_n_108__1_, data_n_108__2_, data_n_108__3_, data_n_108__4_, data_n_108__5_, data_n_108__6_, data_n_108__7_, data_n_108__8_, data_n_108__9_, data_n_108__10_, data_n_108__11_, data_n_108__12_, data_n_108__13_, data_n_108__14_, data_n_108__15_, data_n_108__16_, data_n_108__17_, data_n_108__18_, data_n_108__19_, data_n_108__20_, data_n_108__21_, data_n_108__22_, data_n_108__23_, data_n_108__24_, data_n_108__25_, data_n_108__26_, data_n_108__27_, data_n_108__28_, data_n_108__29_, data_n_108__30_, data_n_108__31_ } = (N164)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2474)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N164 = N2346;
  assign { data_n_109__0_, data_n_109__1_, data_n_109__2_, data_n_109__3_, data_n_109__4_, data_n_109__5_, data_n_109__6_, data_n_109__7_, data_n_109__8_, data_n_109__9_, data_n_109__10_, data_n_109__11_, data_n_109__12_, data_n_109__13_, data_n_109__14_, data_n_109__15_, data_n_109__16_, data_n_109__17_, data_n_109__18_, data_n_109__19_, data_n_109__20_, data_n_109__21_, data_n_109__22_, data_n_109__23_, data_n_109__24_, data_n_109__25_, data_n_109__26_, data_n_109__27_, data_n_109__28_, data_n_109__29_, data_n_109__30_, data_n_109__31_ } = (N165)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2475)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N165 = N2347;
  assign { data_n_110__0_, data_n_110__1_, data_n_110__2_, data_n_110__3_, data_n_110__4_, data_n_110__5_, data_n_110__6_, data_n_110__7_, data_n_110__8_, data_n_110__9_, data_n_110__10_, data_n_110__11_, data_n_110__12_, data_n_110__13_, data_n_110__14_, data_n_110__15_, data_n_110__16_, data_n_110__17_, data_n_110__18_, data_n_110__19_, data_n_110__20_, data_n_110__21_, data_n_110__22_, data_n_110__23_, data_n_110__24_, data_n_110__25_, data_n_110__26_, data_n_110__27_, data_n_110__28_, data_n_110__29_, data_n_110__30_, data_n_110__31_ } = (N166)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2476)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N166 = N2348;
  assign { data_n_111__0_, data_n_111__1_, data_n_111__2_, data_n_111__3_, data_n_111__4_, data_n_111__5_, data_n_111__6_, data_n_111__7_, data_n_111__8_, data_n_111__9_, data_n_111__10_, data_n_111__11_, data_n_111__12_, data_n_111__13_, data_n_111__14_, data_n_111__15_, data_n_111__16_, data_n_111__17_, data_n_111__18_, data_n_111__19_, data_n_111__20_, data_n_111__21_, data_n_111__22_, data_n_111__23_, data_n_111__24_, data_n_111__25_, data_n_111__26_, data_n_111__27_, data_n_111__28_, data_n_111__29_, data_n_111__30_, data_n_111__31_ } = (N167)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2477)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N167 = N2349;
  assign { data_n_112__0_, data_n_112__1_, data_n_112__2_, data_n_112__3_, data_n_112__4_, data_n_112__5_, data_n_112__6_, data_n_112__7_, data_n_112__8_, data_n_112__9_, data_n_112__10_, data_n_112__11_, data_n_112__12_, data_n_112__13_, data_n_112__14_, data_n_112__15_, data_n_112__16_, data_n_112__17_, data_n_112__18_, data_n_112__19_, data_n_112__20_, data_n_112__21_, data_n_112__22_, data_n_112__23_, data_n_112__24_, data_n_112__25_, data_n_112__26_, data_n_112__27_, data_n_112__28_, data_n_112__29_, data_n_112__30_, data_n_112__31_ } = (N168)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2478)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N168 = N2350;
  assign { data_n_113__0_, data_n_113__1_, data_n_113__2_, data_n_113__3_, data_n_113__4_, data_n_113__5_, data_n_113__6_, data_n_113__7_, data_n_113__8_, data_n_113__9_, data_n_113__10_, data_n_113__11_, data_n_113__12_, data_n_113__13_, data_n_113__14_, data_n_113__15_, data_n_113__16_, data_n_113__17_, data_n_113__18_, data_n_113__19_, data_n_113__20_, data_n_113__21_, data_n_113__22_, data_n_113__23_, data_n_113__24_, data_n_113__25_, data_n_113__26_, data_n_113__27_, data_n_113__28_, data_n_113__29_, data_n_113__30_, data_n_113__31_ } = (N169)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2479)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N169 = N2351;
  assign { data_n_114__0_, data_n_114__1_, data_n_114__2_, data_n_114__3_, data_n_114__4_, data_n_114__5_, data_n_114__6_, data_n_114__7_, data_n_114__8_, data_n_114__9_, data_n_114__10_, data_n_114__11_, data_n_114__12_, data_n_114__13_, data_n_114__14_, data_n_114__15_, data_n_114__16_, data_n_114__17_, data_n_114__18_, data_n_114__19_, data_n_114__20_, data_n_114__21_, data_n_114__22_, data_n_114__23_, data_n_114__24_, data_n_114__25_, data_n_114__26_, data_n_114__27_, data_n_114__28_, data_n_114__29_, data_n_114__30_, data_n_114__31_ } = (N170)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2480)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N170 = N2352;
  assign { data_n_115__0_, data_n_115__1_, data_n_115__2_, data_n_115__3_, data_n_115__4_, data_n_115__5_, data_n_115__6_, data_n_115__7_, data_n_115__8_, data_n_115__9_, data_n_115__10_, data_n_115__11_, data_n_115__12_, data_n_115__13_, data_n_115__14_, data_n_115__15_, data_n_115__16_, data_n_115__17_, data_n_115__18_, data_n_115__19_, data_n_115__20_, data_n_115__21_, data_n_115__22_, data_n_115__23_, data_n_115__24_, data_n_115__25_, data_n_115__26_, data_n_115__27_, data_n_115__28_, data_n_115__29_, data_n_115__30_, data_n_115__31_ } = (N171)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2481)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N171 = N2353;
  assign { data_n_116__0_, data_n_116__1_, data_n_116__2_, data_n_116__3_, data_n_116__4_, data_n_116__5_, data_n_116__6_, data_n_116__7_, data_n_116__8_, data_n_116__9_, data_n_116__10_, data_n_116__11_, data_n_116__12_, data_n_116__13_, data_n_116__14_, data_n_116__15_, data_n_116__16_, data_n_116__17_, data_n_116__18_, data_n_116__19_, data_n_116__20_, data_n_116__21_, data_n_116__22_, data_n_116__23_, data_n_116__24_, data_n_116__25_, data_n_116__26_, data_n_116__27_, data_n_116__28_, data_n_116__29_, data_n_116__30_, data_n_116__31_ } = (N172)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2482)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N172 = N2354;
  assign { data_n_117__0_, data_n_117__1_, data_n_117__2_, data_n_117__3_, data_n_117__4_, data_n_117__5_, data_n_117__6_, data_n_117__7_, data_n_117__8_, data_n_117__9_, data_n_117__10_, data_n_117__11_, data_n_117__12_, data_n_117__13_, data_n_117__14_, data_n_117__15_, data_n_117__16_, data_n_117__17_, data_n_117__18_, data_n_117__19_, data_n_117__20_, data_n_117__21_, data_n_117__22_, data_n_117__23_, data_n_117__24_, data_n_117__25_, data_n_117__26_, data_n_117__27_, data_n_117__28_, data_n_117__29_, data_n_117__30_, data_n_117__31_ } = (N173)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2483)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N173 = N2355;
  assign { data_n_118__0_, data_n_118__1_, data_n_118__2_, data_n_118__3_, data_n_118__4_, data_n_118__5_, data_n_118__6_, data_n_118__7_, data_n_118__8_, data_n_118__9_, data_n_118__10_, data_n_118__11_, data_n_118__12_, data_n_118__13_, data_n_118__14_, data_n_118__15_, data_n_118__16_, data_n_118__17_, data_n_118__18_, data_n_118__19_, data_n_118__20_, data_n_118__21_, data_n_118__22_, data_n_118__23_, data_n_118__24_, data_n_118__25_, data_n_118__26_, data_n_118__27_, data_n_118__28_, data_n_118__29_, data_n_118__30_, data_n_118__31_ } = (N174)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2484)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N174 = N2356;
  assign { data_n_119__0_, data_n_119__1_, data_n_119__2_, data_n_119__3_, data_n_119__4_, data_n_119__5_, data_n_119__6_, data_n_119__7_, data_n_119__8_, data_n_119__9_, data_n_119__10_, data_n_119__11_, data_n_119__12_, data_n_119__13_, data_n_119__14_, data_n_119__15_, data_n_119__16_, data_n_119__17_, data_n_119__18_, data_n_119__19_, data_n_119__20_, data_n_119__21_, data_n_119__22_, data_n_119__23_, data_n_119__24_, data_n_119__25_, data_n_119__26_, data_n_119__27_, data_n_119__28_, data_n_119__29_, data_n_119__30_, data_n_119__31_ } = (N175)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2485)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N175 = N2357;
  assign { data_n_120__0_, data_n_120__1_, data_n_120__2_, data_n_120__3_, data_n_120__4_, data_n_120__5_, data_n_120__6_, data_n_120__7_, data_n_120__8_, data_n_120__9_, data_n_120__10_, data_n_120__11_, data_n_120__12_, data_n_120__13_, data_n_120__14_, data_n_120__15_, data_n_120__16_, data_n_120__17_, data_n_120__18_, data_n_120__19_, data_n_120__20_, data_n_120__21_, data_n_120__22_, data_n_120__23_, data_n_120__24_, data_n_120__25_, data_n_120__26_, data_n_120__27_, data_n_120__28_, data_n_120__29_, data_n_120__30_, data_n_120__31_ } = (N176)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2486)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N176 = N2358;
  assign { data_n_121__0_, data_n_121__1_, data_n_121__2_, data_n_121__3_, data_n_121__4_, data_n_121__5_, data_n_121__6_, data_n_121__7_, data_n_121__8_, data_n_121__9_, data_n_121__10_, data_n_121__11_, data_n_121__12_, data_n_121__13_, data_n_121__14_, data_n_121__15_, data_n_121__16_, data_n_121__17_, data_n_121__18_, data_n_121__19_, data_n_121__20_, data_n_121__21_, data_n_121__22_, data_n_121__23_, data_n_121__24_, data_n_121__25_, data_n_121__26_, data_n_121__27_, data_n_121__28_, data_n_121__29_, data_n_121__30_, data_n_121__31_ } = (N177)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2487)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N177 = N2359;
  assign { data_n_122__0_, data_n_122__1_, data_n_122__2_, data_n_122__3_, data_n_122__4_, data_n_122__5_, data_n_122__6_, data_n_122__7_, data_n_122__8_, data_n_122__9_, data_n_122__10_, data_n_122__11_, data_n_122__12_, data_n_122__13_, data_n_122__14_, data_n_122__15_, data_n_122__16_, data_n_122__17_, data_n_122__18_, data_n_122__19_, data_n_122__20_, data_n_122__21_, data_n_122__22_, data_n_122__23_, data_n_122__24_, data_n_122__25_, data_n_122__26_, data_n_122__27_, data_n_122__28_, data_n_122__29_, data_n_122__30_, data_n_122__31_ } = (N178)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2488)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N178 = N2360;
  assign { data_n_123__0_, data_n_123__1_, data_n_123__2_, data_n_123__3_, data_n_123__4_, data_n_123__5_, data_n_123__6_, data_n_123__7_, data_n_123__8_, data_n_123__9_, data_n_123__10_, data_n_123__11_, data_n_123__12_, data_n_123__13_, data_n_123__14_, data_n_123__15_, data_n_123__16_, data_n_123__17_, data_n_123__18_, data_n_123__19_, data_n_123__20_, data_n_123__21_, data_n_123__22_, data_n_123__23_, data_n_123__24_, data_n_123__25_, data_n_123__26_, data_n_123__27_, data_n_123__28_, data_n_123__29_, data_n_123__30_, data_n_123__31_ } = (N179)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2489)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N179 = N2361;
  assign { data_n_124__0_, data_n_124__1_, data_n_124__2_, data_n_124__3_, data_n_124__4_, data_n_124__5_, data_n_124__6_, data_n_124__7_, data_n_124__8_, data_n_124__9_, data_n_124__10_, data_n_124__11_, data_n_124__12_, data_n_124__13_, data_n_124__14_, data_n_124__15_, data_n_124__16_, data_n_124__17_, data_n_124__18_, data_n_124__19_, data_n_124__20_, data_n_124__21_, data_n_124__22_, data_n_124__23_, data_n_124__24_, data_n_124__25_, data_n_124__26_, data_n_124__27_, data_n_124__28_, data_n_124__29_, data_n_124__30_, data_n_124__31_ } = (N180)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2490)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N180 = N2362;
  assign { data_n_125__0_, data_n_125__1_, data_n_125__2_, data_n_125__3_, data_n_125__4_, data_n_125__5_, data_n_125__6_, data_n_125__7_, data_n_125__8_, data_n_125__9_, data_n_125__10_, data_n_125__11_, data_n_125__12_, data_n_125__13_, data_n_125__14_, data_n_125__15_, data_n_125__16_, data_n_125__17_, data_n_125__18_, data_n_125__19_, data_n_125__20_, data_n_125__21_, data_n_125__22_, data_n_125__23_, data_n_125__24_, data_n_125__25_, data_n_125__26_, data_n_125__27_, data_n_125__28_, data_n_125__29_, data_n_125__30_, data_n_125__31_ } = (N181)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2491)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N181 = N2363;
  assign { data_n_126__0_, data_n_126__1_, data_n_126__2_, data_n_126__3_, data_n_126__4_, data_n_126__5_, data_n_126__6_, data_n_126__7_, data_n_126__8_, data_n_126__9_, data_n_126__10_, data_n_126__11_, data_n_126__12_, data_n_126__13_, data_n_126__14_, data_n_126__15_, data_n_126__16_, data_n_126__17_, data_n_126__18_, data_n_126__19_, data_n_126__20_, data_n_126__21_, data_n_126__22_, data_n_126__23_, data_n_126__24_, data_n_126__25_, data_n_126__26_, data_n_126__27_, data_n_126__28_, data_n_126__29_, data_n_126__30_, data_n_126__31_ } = (N182)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2492)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N182 = N2364;
  assign { data_n_127__0_, data_n_127__1_, data_n_127__2_, data_n_127__3_, data_n_127__4_, data_n_127__5_, data_n_127__6_, data_n_127__7_, data_n_127__8_, data_n_127__9_, data_n_127__10_, data_n_127__11_, data_n_127__12_, data_n_127__13_, data_n_127__14_, data_n_127__15_, data_n_127__16_, data_n_127__17_, data_n_127__18_, data_n_127__19_, data_n_127__20_, data_n_127__21_, data_n_127__22_, data_n_127__23_, data_n_127__24_, data_n_127__25_, data_n_127__26_, data_n_127__27_, data_n_127__28_, data_n_127__29_, data_n_127__30_, data_n_127__31_ } = (N183)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2493)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N183 = N2365;
  assign valid_o[0] = (N184)? N2622 : 
                      (N2623)? valid_r[0] : 1'b0;
  assign N184 = N2494;
  assign valid_o[1] = (N185)? N2622 : 
                      (N2624)? valid_r[1] : 1'b0;
  assign N185 = N2495;
  assign valid_o[2] = (N186)? N2622 : 
                      (N2625)? valid_r[2] : 1'b0;
  assign N186 = N2496;
  assign valid_o[3] = (N187)? N2622 : 
                      (N2626)? valid_r[3] : 1'b0;
  assign N187 = N2497;
  assign valid_o[4] = (N188)? N2622 : 
                      (N2627)? valid_r[4] : 1'b0;
  assign N188 = N2498;
  assign valid_o[5] = (N189)? N2622 : 
                      (N2628)? valid_r[5] : 1'b0;
  assign N189 = N2499;
  assign valid_o[6] = (N190)? N2622 : 
                      (N2629)? valid_r[6] : 1'b0;
  assign N190 = N2500;
  assign valid_o[7] = (N191)? N2622 : 
                      (N2630)? valid_r[7] : 1'b0;
  assign N191 = N2501;
  assign valid_o[8] = (N192)? N2622 : 
                      (N2631)? valid_r[8] : 1'b0;
  assign N192 = N2502;
  assign valid_o[9] = (N193)? N2622 : 
                      (N2632)? valid_r[9] : 1'b0;
  assign N193 = N2503;
  assign valid_o[10] = (N194)? N2622 : 
                       (N2633)? valid_r[10] : 1'b0;
  assign N194 = N2504;
  assign valid_o[11] = (N195)? N2622 : 
                       (N2634)? valid_r[11] : 1'b0;
  assign N195 = N2505;
  assign valid_o[12] = (N196)? N2622 : 
                       (N2635)? valid_r[12] : 1'b0;
  assign N196 = N2506;
  assign valid_o[13] = (N197)? N2622 : 
                       (N2636)? valid_r[13] : 1'b0;
  assign N197 = N2507;
  assign valid_o[14] = (N198)? N2622 : 
                       (N2637)? valid_r[14] : 1'b0;
  assign N198 = N2508;
  assign valid_o[15] = (N199)? N2622 : 
                       (N2638)? valid_r[15] : 1'b0;
  assign N199 = N2509;
  assign valid_o[16] = (N200)? N2622 : 
                       (N2639)? valid_r[16] : 1'b0;
  assign N200 = N2510;
  assign valid_o[17] = (N201)? N2622 : 
                       (N2640)? valid_r[17] : 1'b0;
  assign N201 = N2511;
  assign valid_o[18] = (N202)? N2622 : 
                       (N2641)? valid_r[18] : 1'b0;
  assign N202 = N2512;
  assign valid_o[19] = (N203)? N2622 : 
                       (N2642)? valid_r[19] : 1'b0;
  assign N203 = N2513;
  assign valid_o[20] = (N204)? N2622 : 
                       (N2643)? valid_r[20] : 1'b0;
  assign N204 = N2514;
  assign valid_o[21] = (N205)? N2622 : 
                       (N2644)? valid_r[21] : 1'b0;
  assign N205 = N2515;
  assign valid_o[22] = (N206)? N2622 : 
                       (N2645)? valid_r[22] : 1'b0;
  assign N206 = N2516;
  assign valid_o[23] = (N207)? N2622 : 
                       (N2646)? valid_r[23] : 1'b0;
  assign N207 = N2517;
  assign valid_o[24] = (N208)? N2622 : 
                       (N2647)? valid_r[24] : 1'b0;
  assign N208 = N2518;
  assign valid_o[25] = (N209)? N2622 : 
                       (N2648)? valid_r[25] : 1'b0;
  assign N209 = N2519;
  assign valid_o[26] = (N210)? N2622 : 
                       (N2649)? valid_r[26] : 1'b0;
  assign N210 = N2520;
  assign valid_o[27] = (N211)? N2622 : 
                       (N2650)? valid_r[27] : 1'b0;
  assign N211 = N2521;
  assign valid_o[28] = (N212)? N2622 : 
                       (N2651)? valid_r[28] : 1'b0;
  assign N212 = N2522;
  assign valid_o[29] = (N213)? N2622 : 
                       (N2652)? valid_r[29] : 1'b0;
  assign N213 = N2523;
  assign valid_o[30] = (N214)? N2622 : 
                       (N2653)? valid_r[30] : 1'b0;
  assign N214 = N2524;
  assign valid_o[31] = (N215)? N2622 : 
                       (N2654)? valid_r[31] : 1'b0;
  assign N215 = N2525;
  assign valid_o[32] = (N216)? N2622 : 
                       (N2655)? valid_r[32] : 1'b0;
  assign N216 = N2526;
  assign valid_o[33] = (N217)? N2622 : 
                       (N2656)? valid_r[33] : 1'b0;
  assign N217 = N2527;
  assign valid_o[34] = (N218)? N2622 : 
                       (N2657)? valid_r[34] : 1'b0;
  assign N218 = N2528;
  assign valid_o[35] = (N219)? N2622 : 
                       (N2658)? valid_r[35] : 1'b0;
  assign N219 = N2529;
  assign valid_o[36] = (N220)? N2622 : 
                       (N2659)? valid_r[36] : 1'b0;
  assign N220 = N2530;
  assign valid_o[37] = (N221)? N2622 : 
                       (N2660)? valid_r[37] : 1'b0;
  assign N221 = N2531;
  assign valid_o[38] = (N222)? N2622 : 
                       (N2661)? valid_r[38] : 1'b0;
  assign N222 = N2532;
  assign valid_o[39] = (N223)? N2622 : 
                       (N2662)? valid_r[39] : 1'b0;
  assign N223 = N2533;
  assign valid_o[40] = (N224)? N2622 : 
                       (N2663)? valid_r[40] : 1'b0;
  assign N224 = N2534;
  assign valid_o[41] = (N225)? N2622 : 
                       (N2664)? valid_r[41] : 1'b0;
  assign N225 = N2535;
  assign valid_o[42] = (N226)? N2622 : 
                       (N2665)? valid_r[42] : 1'b0;
  assign N226 = N2536;
  assign valid_o[43] = (N227)? N2622 : 
                       (N2666)? valid_r[43] : 1'b0;
  assign N227 = N2537;
  assign valid_o[44] = (N228)? N2622 : 
                       (N2667)? valid_r[44] : 1'b0;
  assign N228 = N2538;
  assign valid_o[45] = (N229)? N2622 : 
                       (N2668)? valid_r[45] : 1'b0;
  assign N229 = N2539;
  assign valid_o[46] = (N230)? N2622 : 
                       (N2669)? valid_r[46] : 1'b0;
  assign N230 = N2540;
  assign valid_o[47] = (N231)? N2622 : 
                       (N2670)? valid_r[47] : 1'b0;
  assign N231 = N2541;
  assign valid_o[48] = (N232)? N2622 : 
                       (N2671)? valid_r[48] : 1'b0;
  assign N232 = N2542;
  assign valid_o[49] = (N233)? N2622 : 
                       (N2672)? valid_r[49] : 1'b0;
  assign N233 = N2543;
  assign valid_o[50] = (N234)? N2622 : 
                       (N2673)? valid_r[50] : 1'b0;
  assign N234 = N2544;
  assign valid_o[51] = (N235)? N2622 : 
                       (N2674)? valid_r[51] : 1'b0;
  assign N235 = N2545;
  assign valid_o[52] = (N236)? N2622 : 
                       (N2675)? valid_r[52] : 1'b0;
  assign N236 = N2546;
  assign valid_o[53] = (N237)? N2622 : 
                       (N2676)? valid_r[53] : 1'b0;
  assign N237 = N2547;
  assign valid_o[54] = (N238)? N2622 : 
                       (N2677)? valid_r[54] : 1'b0;
  assign N238 = N2548;
  assign valid_o[55] = (N239)? N2622 : 
                       (N2678)? valid_r[55] : 1'b0;
  assign N239 = N2549;
  assign valid_o[56] = (N240)? N2622 : 
                       (N2679)? valid_r[56] : 1'b0;
  assign N240 = N2550;
  assign valid_o[57] = (N241)? N2622 : 
                       (N2680)? valid_r[57] : 1'b0;
  assign N241 = N2551;
  assign valid_o[58] = (N242)? N2622 : 
                       (N2681)? valid_r[58] : 1'b0;
  assign N242 = N2552;
  assign valid_o[59] = (N243)? N2622 : 
                       (N2682)? valid_r[59] : 1'b0;
  assign N243 = N2553;
  assign valid_o[60] = (N244)? N2622 : 
                       (N2683)? valid_r[60] : 1'b0;
  assign N244 = N2554;
  assign valid_o[61] = (N245)? N2622 : 
                       (N2684)? valid_r[61] : 1'b0;
  assign N245 = N2555;
  assign valid_o[62] = (N246)? N2622 : 
                       (N2685)? valid_r[62] : 1'b0;
  assign N246 = N2556;
  assign valid_o[63] = (N247)? N2622 : 
                       (N2686)? valid_r[63] : 1'b0;
  assign N247 = N2557;
  assign valid_n[64] = (N248)? N2622 : 
                       (N2687)? 1'b0 : 1'b0;
  assign N248 = N2558;
  assign valid_n[65] = (N249)? N2622 : 
                       (N2688)? 1'b0 : 1'b0;
  assign N249 = N2559;
  assign valid_n[66] = (N250)? N2622 : 
                       (N2689)? 1'b0 : 1'b0;
  assign N250 = N2560;
  assign valid_n[67] = (N251)? N2622 : 
                       (N2690)? 1'b0 : 1'b0;
  assign N251 = N2561;
  assign valid_n[68] = (N252)? N2622 : 
                       (N2691)? 1'b0 : 1'b0;
  assign N252 = N2562;
  assign valid_n[69] = (N253)? N2622 : 
                       (N2692)? 1'b0 : 1'b0;
  assign N253 = N2563;
  assign valid_n[70] = (N254)? N2622 : 
                       (N2693)? 1'b0 : 1'b0;
  assign N254 = N2564;
  assign valid_n[71] = (N255)? N2622 : 
                       (N2694)? 1'b0 : 1'b0;
  assign N255 = N2565;
  assign valid_n[72] = (N256)? N2622 : 
                       (N2695)? 1'b0 : 1'b0;
  assign N256 = N2566;
  assign valid_n[73] = (N257)? N2622 : 
                       (N2696)? 1'b0 : 1'b0;
  assign N257 = N2567;
  assign valid_n[74] = (N258)? N2622 : 
                       (N2697)? 1'b0 : 1'b0;
  assign N258 = N2568;
  assign valid_n[75] = (N259)? N2622 : 
                       (N2698)? 1'b0 : 1'b0;
  assign N259 = N2569;
  assign valid_n[76] = (N260)? N2622 : 
                       (N2699)? 1'b0 : 1'b0;
  assign N260 = N2570;
  assign valid_n[77] = (N261)? N2622 : 
                       (N2700)? 1'b0 : 1'b0;
  assign N261 = N2571;
  assign valid_n[78] = (N262)? N2622 : 
                       (N2701)? 1'b0 : 1'b0;
  assign N262 = N2572;
  assign valid_n[79] = (N263)? N2622 : 
                       (N2702)? 1'b0 : 1'b0;
  assign N263 = N2573;
  assign valid_n[80] = (N264)? N2622 : 
                       (N2703)? 1'b0 : 1'b0;
  assign N264 = N2574;
  assign valid_n[81] = (N265)? N2622 : 
                       (N2704)? 1'b0 : 1'b0;
  assign N265 = N2575;
  assign valid_n[82] = (N266)? N2622 : 
                       (N2705)? 1'b0 : 1'b0;
  assign N266 = N2576;
  assign valid_n[83] = (N267)? N2622 : 
                       (N2706)? 1'b0 : 1'b0;
  assign N267 = N2577;
  assign valid_n[84] = (N268)? N2622 : 
                       (N2707)? 1'b0 : 1'b0;
  assign N268 = N2578;
  assign valid_n[85] = (N269)? N2622 : 
                       (N2708)? 1'b0 : 1'b0;
  assign N269 = N2579;
  assign valid_n[86] = (N270)? N2622 : 
                       (N2709)? 1'b0 : 1'b0;
  assign N270 = N2580;
  assign valid_n[87] = (N271)? N2622 : 
                       (N2710)? 1'b0 : 1'b0;
  assign N271 = N2581;
  assign valid_n[88] = (N272)? N2622 : 
                       (N2711)? 1'b0 : 1'b0;
  assign N272 = N2582;
  assign valid_n[89] = (N273)? N2622 : 
                       (N2712)? 1'b0 : 1'b0;
  assign N273 = N2583;
  assign valid_n[90] = (N274)? N2622 : 
                       (N2713)? 1'b0 : 1'b0;
  assign N274 = N2584;
  assign valid_n[91] = (N275)? N2622 : 
                       (N2714)? 1'b0 : 1'b0;
  assign N275 = N2585;
  assign valid_n[92] = (N276)? N2622 : 
                       (N2715)? 1'b0 : 1'b0;
  assign N276 = N2586;
  assign valid_n[93] = (N277)? N2622 : 
                       (N2716)? 1'b0 : 1'b0;
  assign N277 = N2587;
  assign valid_n[94] = (N278)? N2622 : 
                       (N2717)? 1'b0 : 1'b0;
  assign N278 = N2588;
  assign valid_n[95] = (N279)? N2622 : 
                       (N2718)? 1'b0 : 1'b0;
  assign N279 = N2589;
  assign valid_n[96] = (N280)? N2622 : 
                       (N2719)? 1'b0 : 1'b0;
  assign N280 = N2590;
  assign valid_n[97] = (N281)? N2622 : 
                       (N2720)? 1'b0 : 1'b0;
  assign N281 = N2591;
  assign valid_n[98] = (N282)? N2622 : 
                       (N2721)? 1'b0 : 1'b0;
  assign N282 = N2592;
  assign valid_n[99] = (N283)? N2622 : 
                       (N2722)? 1'b0 : 1'b0;
  assign N283 = N2593;
  assign valid_n[100] = (N284)? N2622 : 
                        (N2723)? 1'b0 : 1'b0;
  assign N284 = N2594;
  assign valid_n[101] = (N285)? N2622 : 
                        (N2724)? 1'b0 : 1'b0;
  assign N285 = N2595;
  assign valid_n[102] = (N286)? N2622 : 
                        (N2725)? 1'b0 : 1'b0;
  assign N286 = N2596;
  assign valid_n[103] = (N287)? N2622 : 
                        (N2726)? 1'b0 : 1'b0;
  assign N287 = N2597;
  assign valid_n[104] = (N288)? N2622 : 
                        (N2727)? 1'b0 : 1'b0;
  assign N288 = N2598;
  assign valid_n[105] = (N289)? N2622 : 
                        (N2728)? 1'b0 : 1'b0;
  assign N289 = N2599;
  assign valid_n[106] = (N290)? N2622 : 
                        (N2729)? 1'b0 : 1'b0;
  assign N290 = N2600;
  assign valid_n[107] = (N291)? N2622 : 
                        (N2730)? 1'b0 : 1'b0;
  assign N291 = N2601;
  assign valid_n[108] = (N292)? N2622 : 
                        (N2731)? 1'b0 : 1'b0;
  assign N292 = N2602;
  assign valid_n[109] = (N293)? N2622 : 
                        (N2732)? 1'b0 : 1'b0;
  assign N293 = N2603;
  assign valid_n[110] = (N294)? N2622 : 
                        (N2733)? 1'b0 : 1'b0;
  assign N294 = N2604;
  assign valid_n[111] = (N295)? N2622 : 
                        (N2734)? 1'b0 : 1'b0;
  assign N295 = N2605;
  assign valid_n[112] = (N296)? N2622 : 
                        (N2735)? 1'b0 : 1'b0;
  assign N296 = N2606;
  assign valid_n[113] = (N297)? N2622 : 
                        (N2736)? 1'b0 : 1'b0;
  assign N297 = N2607;
  assign valid_n[114] = (N298)? N2622 : 
                        (N2737)? 1'b0 : 1'b0;
  assign N298 = N2608;
  assign valid_n[115] = (N299)? N2622 : 
                        (N2738)? 1'b0 : 1'b0;
  assign N299 = N2609;
  assign valid_n[116] = (N300)? N2622 : 
                        (N2739)? 1'b0 : 1'b0;
  assign N300 = N2610;
  assign valid_n[117] = (N301)? N2622 : 
                        (N2740)? 1'b0 : 1'b0;
  assign N301 = N2611;
  assign valid_n[118] = (N302)? N2622 : 
                        (N2741)? 1'b0 : 1'b0;
  assign N302 = N2612;
  assign valid_n[119] = (N303)? N2622 : 
                        (N2742)? 1'b0 : 1'b0;
  assign N303 = N2613;
  assign valid_n[120] = (N304)? N2622 : 
                        (N2743)? 1'b0 : 1'b0;
  assign N304 = N2614;
  assign valid_n[121] = (N305)? N2622 : 
                        (N2744)? 1'b0 : 1'b0;
  assign N305 = N2615;
  assign valid_n[122] = (N306)? N2622 : 
                        (N2745)? 1'b0 : 1'b0;
  assign N306 = N2616;
  assign valid_n[123] = (N307)? N2622 : 
                        (N2746)? 1'b0 : 1'b0;
  assign N307 = N2617;
  assign valid_n[124] = (N308)? N2622 : 
                        (N2747)? 1'b0 : 1'b0;
  assign N308 = N2618;
  assign valid_n[125] = (N309)? N2622 : 
                        (N2748)? 1'b0 : 1'b0;
  assign N309 = N2619;
  assign valid_n[126] = (N310)? N2622 : 
                        (N2749)? 1'b0 : 1'b0;
  assign N310 = N2620;
  assign valid_n[127] = (N311)? N2622 : 
                        (N2750)? 1'b0 : 1'b0;
  assign N311 = N2621;
  assign data_nn[63:32] = (N312)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                          (N313)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                          (N314)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                          (N315)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                          (N316)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                          (N317)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                          (N318)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                          (N319)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                          (N320)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                          (N321)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                          (N322)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                          (N323)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                          (N324)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                          (N325)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                          (N326)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                          (N327)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                          (N328)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                          (N329)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                          (N330)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                          (N331)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                          (N332)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                          (N333)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                          (N334)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                          (N335)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                          (N336)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                          (N337)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                          (N338)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                          (N339)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                          (N340)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                          (N341)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                          (N342)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                          (N343)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                          (N344)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                          (N345)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                          (N346)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                          (N347)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                          (N348)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                          (N349)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                          (N350)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                          (N351)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                          (N352)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                          (N353)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                          (N354)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                          (N355)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                          (N356)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                          (N357)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                          (N358)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                          (N359)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                          (N360)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                          (N361)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                          (N362)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                          (N363)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                          (N364)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                          (N365)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                          (N366)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                          (N367)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                          (N368)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                          (N369)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                          (N370)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                          (N371)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                          (N372)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                          (N373)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                          (N374)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                          (N375)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                          (N376)? data_o[2047:2016] : 
                          (N377)? data_o[2015:1984] : 
                          (N378)? data_o[1983:1952] : 
                          (N379)? data_o[1951:1920] : 
                          (N380)? data_o[1919:1888] : 
                          (N381)? data_o[1887:1856] : 
                          (N382)? data_o[1855:1824] : 
                          (N383)? data_o[1823:1792] : 
                          (N384)? data_o[1791:1760] : 
                          (N385)? data_o[1759:1728] : 
                          (N386)? data_o[1727:1696] : 
                          (N387)? data_o[1695:1664] : 
                          (N388)? data_o[1663:1632] : 
                          (N389)? data_o[1631:1600] : 
                          (N390)? data_o[1599:1568] : 
                          (N391)? data_o[1567:1536] : 
                          (N392)? data_o[1535:1504] : 
                          (N393)? data_o[1503:1472] : 
                          (N394)? data_o[1471:1440] : 
                          (N395)? data_o[1439:1408] : 
                          (N396)? data_o[1407:1376] : 
                          (N397)? data_o[1375:1344] : 
                          (N398)? data_o[1343:1312] : 
                          (N399)? data_o[1311:1280] : 
                          (N400)? data_o[1279:1248] : 
                          (N401)? data_o[1247:1216] : 
                          (N402)? data_o[1215:1184] : 
                          (N403)? data_o[1183:1152] : 
                          (N404)? data_o[1151:1120] : 
                          (N405)? data_o[1119:1088] : 
                          (N406)? data_o[1087:1056] : 
                          (N407)? data_o[1055:1024] : 
                          (N408)? data_o[1023:992] : 
                          (N409)? data_o[991:960] : 
                          (N410)? data_o[959:928] : 
                          (N411)? data_o[927:896] : 
                          (N412)? data_o[895:864] : 
                          (N413)? data_o[863:832] : 
                          (N414)? data_o[831:800] : 
                          (N415)? data_o[799:768] : 
                          (N416)? data_o[767:736] : 
                          (N417)? data_o[735:704] : 
                          (N418)? data_o[703:672] : 
                          (N419)? data_o[671:640] : 
                          (N420)? data_o[639:608] : 
                          (N421)? data_o[607:576] : 
                          (N422)? data_o[575:544] : 
                          (N423)? data_o[543:512] : 
                          (N424)? data_o[511:480] : 
                          (N425)? data_o[479:448] : 
                          (N426)? data_o[447:416] : 
                          (N427)? data_o[415:384] : 
                          (N428)? data_o[383:352] : 
                          (N429)? data_o[351:320] : 
                          (N430)? data_o[319:288] : 
                          (N431)? data_o[287:256] : 
                          (N432)? data_o[255:224] : 
                          (N433)? data_o[223:192] : 
                          (N434)? data_o[191:160] : 
                          (N435)? data_o[159:128] : 
                          (N436)? data_o[127:96] : 
                          (N437)? data_o[95:64] : 
                          (N438)? data_o[63:32] : 1'b0;
  assign N312 = N5522;
  assign N313 = N5523;
  assign N314 = N5524;
  assign N315 = N5525;
  assign N316 = N5526;
  assign N317 = N5527;
  assign N318 = N5528;
  assign N319 = N5529;
  assign N320 = N5530;
  assign N321 = N5531;
  assign N322 = N5532;
  assign N323 = N5533;
  assign N324 = N3475;
  assign N325 = N3474;
  assign N326 = N3473;
  assign N327 = N3472;
  assign N328 = N3471;
  assign N329 = N3470;
  assign N330 = N3469;
  assign N331 = N3468;
  assign N332 = N3467;
  assign N333 = N3466;
  assign N334 = N3465;
  assign N335 = N3464;
  assign N336 = N3463;
  assign N337 = N3462;
  assign N338 = N3461;
  assign N339 = N3460;
  assign N340 = N3459;
  assign N341 = N3458;
  assign N342 = N3457;
  assign N343 = N3456;
  assign N344 = N3455;
  assign N345 = N3454;
  assign N346 = N3453;
  assign N347 = N3452;
  assign N348 = N3451;
  assign N349 = N3450;
  assign N350 = N3449;
  assign N351 = N3448;
  assign N352 = N3447;
  assign N353 = N3446;
  assign N354 = N3445;
  assign N355 = N3444;
  assign N356 = N3443;
  assign N357 = N3442;
  assign N358 = N3441;
  assign N359 = N3440;
  assign N360 = N3439;
  assign N361 = N3438;
  assign N362 = N3437;
  assign N363 = N3436;
  assign N364 = N3435;
  assign N365 = N3434;
  assign N366 = N3433;
  assign N367 = N3432;
  assign N368 = N3431;
  assign N369 = N3430;
  assign N370 = N3429;
  assign N371 = N3428;
  assign N372 = N3427;
  assign N373 = N3426;
  assign N374 = N3425;
  assign N375 = N3424;
  assign N376 = N3423;
  assign N377 = N3422;
  assign N378 = N3421;
  assign N379 = N3420;
  assign N380 = N3419;
  assign N381 = N3418;
  assign N382 = N3417;
  assign N383 = N3416;
  assign N384 = N3415;
  assign N385 = N3414;
  assign N386 = N3413;
  assign N387 = N3412;
  assign N388 = N3411;
  assign N389 = N3410;
  assign N390 = N3409;
  assign N391 = N3408;
  assign N392 = N3407;
  assign N393 = N3406;
  assign N394 = N3405;
  assign N395 = N3404;
  assign N396 = N3403;
  assign N397 = N3402;
  assign N398 = N3401;
  assign N399 = N3400;
  assign N400 = N3399;
  assign N401 = N3398;
  assign N402 = N3397;
  assign N403 = N3396;
  assign N404 = N3395;
  assign N405 = N3394;
  assign N406 = N3393;
  assign N407 = N3392;
  assign N408 = N3391;
  assign N409 = N3390;
  assign N410 = N3389;
  assign N411 = N3388;
  assign N412 = N3387;
  assign N413 = N3386;
  assign N414 = N3385;
  assign N415 = N3384;
  assign N416 = N3383;
  assign N417 = N3382;
  assign N418 = N3381;
  assign N419 = N3380;
  assign N420 = N3379;
  assign N421 = N3378;
  assign N422 = N3377;
  assign N423 = N3376;
  assign N424 = N3375;
  assign N425 = N3374;
  assign N426 = N3373;
  assign N427 = N3372;
  assign N428 = N3371;
  assign N429 = N3370;
  assign N430 = N3369;
  assign N431 = N3368;
  assign N432 = N3367;
  assign N433 = N3366;
  assign N434 = N3365;
  assign N435 = N3364;
  assign N436 = N3363;
  assign N437 = N3362;
  assign N438 = N3361;
  assign data_nn[95:64] = (N313)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                          (N314)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                          (N315)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                          (N316)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                          (N317)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                          (N318)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                          (N319)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                          (N320)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                          (N321)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                          (N322)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                          (N323)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                          (N324)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                          (N325)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                          (N326)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                          (N327)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                          (N328)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                          (N329)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                          (N330)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                          (N331)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                          (N332)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                          (N333)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                          (N334)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                          (N335)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                          (N336)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                          (N337)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                          (N338)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                          (N339)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                          (N340)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                          (N341)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                          (N342)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                          (N343)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                          (N344)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                          (N345)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                          (N346)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                          (N347)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                          (N348)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                          (N349)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                          (N350)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                          (N351)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                          (N352)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                          (N353)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                          (N354)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                          (N355)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                          (N356)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                          (N357)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                          (N358)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                          (N359)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                          (N360)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                          (N361)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                          (N362)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                          (N363)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                          (N364)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                          (N365)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                          (N366)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                          (N367)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                          (N368)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                          (N369)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                          (N370)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                          (N371)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                          (N372)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                          (N373)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                          (N374)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                          (N375)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                          (N376)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                          (N377)? data_o[2047:2016] : 
                          (N378)? data_o[2015:1984] : 
                          (N379)? data_o[1983:1952] : 
                          (N380)? data_o[1951:1920] : 
                          (N381)? data_o[1919:1888] : 
                          (N382)? data_o[1887:1856] : 
                          (N383)? data_o[1855:1824] : 
                          (N384)? data_o[1823:1792] : 
                          (N385)? data_o[1791:1760] : 
                          (N386)? data_o[1759:1728] : 
                          (N387)? data_o[1727:1696] : 
                          (N388)? data_o[1695:1664] : 
                          (N389)? data_o[1663:1632] : 
                          (N390)? data_o[1631:1600] : 
                          (N391)? data_o[1599:1568] : 
                          (N392)? data_o[1567:1536] : 
                          (N393)? data_o[1535:1504] : 
                          (N394)? data_o[1503:1472] : 
                          (N395)? data_o[1471:1440] : 
                          (N396)? data_o[1439:1408] : 
                          (N397)? data_o[1407:1376] : 
                          (N398)? data_o[1375:1344] : 
                          (N399)? data_o[1343:1312] : 
                          (N400)? data_o[1311:1280] : 
                          (N401)? data_o[1279:1248] : 
                          (N402)? data_o[1247:1216] : 
                          (N403)? data_o[1215:1184] : 
                          (N404)? data_o[1183:1152] : 
                          (N405)? data_o[1151:1120] : 
                          (N406)? data_o[1119:1088] : 
                          (N407)? data_o[1087:1056] : 
                          (N408)? data_o[1055:1024] : 
                          (N409)? data_o[1023:992] : 
                          (N410)? data_o[991:960] : 
                          (N411)? data_o[959:928] : 
                          (N412)? data_o[927:896] : 
                          (N413)? data_o[895:864] : 
                          (N414)? data_o[863:832] : 
                          (N415)? data_o[831:800] : 
                          (N416)? data_o[799:768] : 
                          (N417)? data_o[767:736] : 
                          (N418)? data_o[735:704] : 
                          (N419)? data_o[703:672] : 
                          (N420)? data_o[671:640] : 
                          (N421)? data_o[639:608] : 
                          (N422)? data_o[607:576] : 
                          (N423)? data_o[575:544] : 
                          (N424)? data_o[543:512] : 
                          (N425)? data_o[511:480] : 
                          (N426)? data_o[479:448] : 
                          (N427)? data_o[447:416] : 
                          (N428)? data_o[415:384] : 
                          (N429)? data_o[383:352] : 
                          (N430)? data_o[351:320] : 
                          (N431)? data_o[319:288] : 
                          (N432)? data_o[287:256] : 
                          (N433)? data_o[255:224] : 
                          (N434)? data_o[223:192] : 
                          (N435)? data_o[191:160] : 
                          (N436)? data_o[159:128] : 
                          (N437)? data_o[127:96] : 
                          (N438)? data_o[95:64] : 1'b0;
  assign data_nn[127:96] = (N314)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                           (N315)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                           (N316)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                           (N317)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                           (N318)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                           (N319)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                           (N320)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                           (N321)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                           (N322)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                           (N323)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                           (N324)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                           (N325)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                           (N326)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                           (N327)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                           (N328)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                           (N329)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                           (N330)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                           (N331)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                           (N332)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                           (N333)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                           (N334)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                           (N335)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                           (N336)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                           (N337)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                           (N338)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                           (N339)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                           (N340)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                           (N341)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                           (N342)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                           (N343)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                           (N344)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                           (N345)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                           (N346)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                           (N347)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                           (N348)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                           (N349)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                           (N350)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                           (N351)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                           (N352)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                           (N353)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                           (N354)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                           (N355)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                           (N356)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                           (N357)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                           (N358)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                           (N359)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                           (N360)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                           (N361)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                           (N362)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                           (N363)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                           (N364)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                           (N365)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                           (N366)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                           (N367)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                           (N368)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                           (N369)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                           (N370)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                           (N371)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                           (N372)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                           (N373)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                           (N374)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                           (N375)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                           (N376)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                           (N377)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                           (N378)? data_o[2047:2016] : 
                           (N379)? data_o[2015:1984] : 
                           (N380)? data_o[1983:1952] : 
                           (N381)? data_o[1951:1920] : 
                           (N382)? data_o[1919:1888] : 
                           (N383)? data_o[1887:1856] : 
                           (N384)? data_o[1855:1824] : 
                           (N385)? data_o[1823:1792] : 
                           (N386)? data_o[1791:1760] : 
                           (N387)? data_o[1759:1728] : 
                           (N388)? data_o[1727:1696] : 
                           (N389)? data_o[1695:1664] : 
                           (N390)? data_o[1663:1632] : 
                           (N391)? data_o[1631:1600] : 
                           (N392)? data_o[1599:1568] : 
                           (N393)? data_o[1567:1536] : 
                           (N394)? data_o[1535:1504] : 
                           (N395)? data_o[1503:1472] : 
                           (N396)? data_o[1471:1440] : 
                           (N397)? data_o[1439:1408] : 
                           (N398)? data_o[1407:1376] : 
                           (N399)? data_o[1375:1344] : 
                           (N400)? data_o[1343:1312] : 
                           (N401)? data_o[1311:1280] : 
                           (N402)? data_o[1279:1248] : 
                           (N403)? data_o[1247:1216] : 
                           (N404)? data_o[1215:1184] : 
                           (N405)? data_o[1183:1152] : 
                           (N406)? data_o[1151:1120] : 
                           (N407)? data_o[1119:1088] : 
                           (N408)? data_o[1087:1056] : 
                           (N409)? data_o[1055:1024] : 
                           (N410)? data_o[1023:992] : 
                           (N411)? data_o[991:960] : 
                           (N412)? data_o[959:928] : 
                           (N413)? data_o[927:896] : 
                           (N414)? data_o[895:864] : 
                           (N415)? data_o[863:832] : 
                           (N416)? data_o[831:800] : 
                           (N417)? data_o[799:768] : 
                           (N418)? data_o[767:736] : 
                           (N419)? data_o[735:704] : 
                           (N420)? data_o[703:672] : 
                           (N421)? data_o[671:640] : 
                           (N422)? data_o[639:608] : 
                           (N423)? data_o[607:576] : 
                           (N424)? data_o[575:544] : 
                           (N425)? data_o[543:512] : 
                           (N426)? data_o[511:480] : 
                           (N427)? data_o[479:448] : 
                           (N428)? data_o[447:416] : 
                           (N429)? data_o[415:384] : 
                           (N430)? data_o[383:352] : 
                           (N431)? data_o[351:320] : 
                           (N432)? data_o[319:288] : 
                           (N433)? data_o[287:256] : 
                           (N434)? data_o[255:224] : 
                           (N435)? data_o[223:192] : 
                           (N436)? data_o[191:160] : 
                           (N437)? data_o[159:128] : 
                           (N438)? data_o[127:96] : 1'b0;
  assign data_nn[159:128] = (N315)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N316)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N317)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N318)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N319)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N320)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N321)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N322)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N323)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N324)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N325)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N326)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N327)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N328)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N329)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N330)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N331)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N332)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N333)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N334)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N335)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N336)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N337)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N338)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N339)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N340)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N341)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N342)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N343)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N344)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N345)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N346)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N347)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N348)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N349)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N350)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N351)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N352)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N353)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N354)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N355)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N356)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N357)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N358)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N359)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N360)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N361)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N362)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N363)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N364)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N365)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N366)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N367)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N368)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N369)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N370)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N371)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N372)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N373)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N374)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N375)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N376)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N377)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N378)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N379)? data_o[2047:2016] : 
                            (N380)? data_o[2015:1984] : 
                            (N381)? data_o[1983:1952] : 
                            (N382)? data_o[1951:1920] : 
                            (N383)? data_o[1919:1888] : 
                            (N384)? data_o[1887:1856] : 
                            (N385)? data_o[1855:1824] : 
                            (N386)? data_o[1823:1792] : 
                            (N387)? data_o[1791:1760] : 
                            (N388)? data_o[1759:1728] : 
                            (N389)? data_o[1727:1696] : 
                            (N390)? data_o[1695:1664] : 
                            (N391)? data_o[1663:1632] : 
                            (N392)? data_o[1631:1600] : 
                            (N393)? data_o[1599:1568] : 
                            (N394)? data_o[1567:1536] : 
                            (N395)? data_o[1535:1504] : 
                            (N396)? data_o[1503:1472] : 
                            (N397)? data_o[1471:1440] : 
                            (N398)? data_o[1439:1408] : 
                            (N399)? data_o[1407:1376] : 
                            (N400)? data_o[1375:1344] : 
                            (N401)? data_o[1343:1312] : 
                            (N402)? data_o[1311:1280] : 
                            (N403)? data_o[1279:1248] : 
                            (N404)? data_o[1247:1216] : 
                            (N405)? data_o[1215:1184] : 
                            (N406)? data_o[1183:1152] : 
                            (N407)? data_o[1151:1120] : 
                            (N408)? data_o[1119:1088] : 
                            (N409)? data_o[1087:1056] : 
                            (N410)? data_o[1055:1024] : 
                            (N411)? data_o[1023:992] : 
                            (N412)? data_o[991:960] : 
                            (N413)? data_o[959:928] : 
                            (N414)? data_o[927:896] : 
                            (N415)? data_o[895:864] : 
                            (N416)? data_o[863:832] : 
                            (N417)? data_o[831:800] : 
                            (N418)? data_o[799:768] : 
                            (N419)? data_o[767:736] : 
                            (N420)? data_o[735:704] : 
                            (N421)? data_o[703:672] : 
                            (N422)? data_o[671:640] : 
                            (N423)? data_o[639:608] : 
                            (N424)? data_o[607:576] : 
                            (N425)? data_o[575:544] : 
                            (N426)? data_o[543:512] : 
                            (N427)? data_o[511:480] : 
                            (N428)? data_o[479:448] : 
                            (N429)? data_o[447:416] : 
                            (N430)? data_o[415:384] : 
                            (N431)? data_o[383:352] : 
                            (N432)? data_o[351:320] : 
                            (N433)? data_o[319:288] : 
                            (N434)? data_o[287:256] : 
                            (N435)? data_o[255:224] : 
                            (N436)? data_o[223:192] : 
                            (N437)? data_o[191:160] : 
                            (N438)? data_o[159:128] : 1'b0;
  assign data_nn[191:160] = (N316)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N317)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N318)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N319)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N320)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N321)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N322)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N323)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N324)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N325)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N326)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N327)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N328)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N329)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N330)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N331)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N332)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N333)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N334)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N335)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N336)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N337)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N338)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N339)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N340)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N341)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N342)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N343)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N344)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N345)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N346)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N347)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N348)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N349)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N350)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N351)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N352)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N353)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N354)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N355)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N356)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N357)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N358)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N359)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N360)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N361)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N362)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N363)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N364)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N365)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N366)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N367)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N368)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N369)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N370)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N371)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N372)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N373)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N374)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N375)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N376)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N377)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N378)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N379)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N380)? data_o[2047:2016] : 
                            (N381)? data_o[2015:1984] : 
                            (N382)? data_o[1983:1952] : 
                            (N383)? data_o[1951:1920] : 
                            (N384)? data_o[1919:1888] : 
                            (N385)? data_o[1887:1856] : 
                            (N386)? data_o[1855:1824] : 
                            (N387)? data_o[1823:1792] : 
                            (N388)? data_o[1791:1760] : 
                            (N389)? data_o[1759:1728] : 
                            (N390)? data_o[1727:1696] : 
                            (N391)? data_o[1695:1664] : 
                            (N392)? data_o[1663:1632] : 
                            (N393)? data_o[1631:1600] : 
                            (N394)? data_o[1599:1568] : 
                            (N395)? data_o[1567:1536] : 
                            (N396)? data_o[1535:1504] : 
                            (N397)? data_o[1503:1472] : 
                            (N398)? data_o[1471:1440] : 
                            (N399)? data_o[1439:1408] : 
                            (N400)? data_o[1407:1376] : 
                            (N401)? data_o[1375:1344] : 
                            (N402)? data_o[1343:1312] : 
                            (N403)? data_o[1311:1280] : 
                            (N404)? data_o[1279:1248] : 
                            (N405)? data_o[1247:1216] : 
                            (N406)? data_o[1215:1184] : 
                            (N407)? data_o[1183:1152] : 
                            (N408)? data_o[1151:1120] : 
                            (N409)? data_o[1119:1088] : 
                            (N410)? data_o[1087:1056] : 
                            (N411)? data_o[1055:1024] : 
                            (N412)? data_o[1023:992] : 
                            (N413)? data_o[991:960] : 
                            (N414)? data_o[959:928] : 
                            (N415)? data_o[927:896] : 
                            (N416)? data_o[895:864] : 
                            (N417)? data_o[863:832] : 
                            (N418)? data_o[831:800] : 
                            (N419)? data_o[799:768] : 
                            (N420)? data_o[767:736] : 
                            (N421)? data_o[735:704] : 
                            (N422)? data_o[703:672] : 
                            (N423)? data_o[671:640] : 
                            (N424)? data_o[639:608] : 
                            (N425)? data_o[607:576] : 
                            (N426)? data_o[575:544] : 
                            (N427)? data_o[543:512] : 
                            (N428)? data_o[511:480] : 
                            (N429)? data_o[479:448] : 
                            (N430)? data_o[447:416] : 
                            (N431)? data_o[415:384] : 
                            (N432)? data_o[383:352] : 
                            (N433)? data_o[351:320] : 
                            (N434)? data_o[319:288] : 
                            (N435)? data_o[287:256] : 
                            (N436)? data_o[255:224] : 
                            (N437)? data_o[223:192] : 
                            (N438)? data_o[191:160] : 1'b0;
  assign data_nn[223:192] = (N439)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N440)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N441)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N442)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N443)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N444)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N445)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N446)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N447)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N448)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N449)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N450)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N451)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N452)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N453)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N454)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N455)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N456)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N457)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N458)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N459)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N460)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N461)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N462)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N463)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N464)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N465)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N466)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N467)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N468)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N469)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N470)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N471)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N472)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N473)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N474)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N475)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N476)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N477)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N478)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N479)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N480)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N481)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N482)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N483)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N484)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N485)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N486)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N487)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N488)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N489)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N490)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N491)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N492)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N493)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N494)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N495)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N496)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N497)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N498)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N499)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N500)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N501)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N502)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N503)? data_o[2047:2016] : 
                            (N504)? data_o[2015:1984] : 
                            (N505)? data_o[1983:1952] : 
                            (N506)? data_o[1951:1920] : 
                            (N507)? data_o[1919:1888] : 
                            (N508)? data_o[1887:1856] : 
                            (N509)? data_o[1855:1824] : 
                            (N510)? data_o[1823:1792] : 
                            (N511)? data_o[1791:1760] : 
                            (N512)? data_o[1759:1728] : 
                            (N513)? data_o[1727:1696] : 
                            (N514)? data_o[1695:1664] : 
                            (N515)? data_o[1663:1632] : 
                            (N516)? data_o[1631:1600] : 
                            (N517)? data_o[1599:1568] : 
                            (N518)? data_o[1567:1536] : 
                            (N519)? data_o[1535:1504] : 
                            (N520)? data_o[1503:1472] : 
                            (N521)? data_o[1471:1440] : 
                            (N522)? data_o[1439:1408] : 
                            (N523)? data_o[1407:1376] : 
                            (N524)? data_o[1375:1344] : 
                            (N525)? data_o[1343:1312] : 
                            (N526)? data_o[1311:1280] : 
                            (N527)? data_o[1279:1248] : 
                            (N528)? data_o[1247:1216] : 
                            (N529)? data_o[1215:1184] : 
                            (N530)? data_o[1183:1152] : 
                            (N531)? data_o[1151:1120] : 
                            (N532)? data_o[1119:1088] : 
                            (N533)? data_o[1087:1056] : 
                            (N534)? data_o[1055:1024] : 
                            (N535)? data_o[1023:992] : 
                            (N536)? data_o[991:960] : 
                            (N537)? data_o[959:928] : 
                            (N538)? data_o[927:896] : 
                            (N539)? data_o[895:864] : 
                            (N540)? data_o[863:832] : 
                            (N541)? data_o[831:800] : 
                            (N542)? data_o[799:768] : 
                            (N543)? data_o[767:736] : 
                            (N544)? data_o[735:704] : 
                            (N545)? data_o[703:672] : 
                            (N546)? data_o[671:640] : 
                            (N547)? data_o[639:608] : 
                            (N548)? data_o[607:576] : 
                            (N549)? data_o[575:544] : 
                            (N550)? data_o[543:512] : 
                            (N551)? data_o[511:480] : 
                            (N552)? data_o[479:448] : 
                            (N553)? data_o[447:416] : 
                            (N554)? data_o[415:384] : 
                            (N555)? data_o[383:352] : 
                            (N556)? data_o[351:320] : 
                            (N557)? data_o[319:288] : 
                            (N558)? data_o[287:256] : 
                            (N559)? data_o[255:224] : 
                            (N560)? data_o[223:192] : 1'b0;
  assign N439 = N5449;
  assign N440 = N5450;
  assign N441 = N5451;
  assign N442 = N5452;
  assign N443 = N3127;
  assign N444 = N3126;
  assign N445 = N3125;
  assign N446 = N3124;
  assign N447 = N3123;
  assign N448 = N3122;
  assign N449 = N3121;
  assign N450 = N3120;
  assign N451 = N3119;
  assign N452 = N3118;
  assign N453 = N3117;
  assign N454 = N3116;
  assign N455 = N3115;
  assign N456 = N3114;
  assign N457 = N3113;
  assign N458 = N3112;
  assign N459 = N3111;
  assign N460 = N3110;
  assign N461 = N3109;
  assign N462 = N3108;
  assign N463 = N3107;
  assign N464 = N3106;
  assign N465 = N3105;
  assign N466 = N3104;
  assign N467 = N3103;
  assign N468 = N3102;
  assign N469 = N3101;
  assign N470 = N3100;
  assign N471 = N3099;
  assign N472 = N3098;
  assign N473 = N3097;
  assign N474 = N3096;
  assign N475 = N3095;
  assign N476 = N3094;
  assign N477 = N3093;
  assign N478 = N3092;
  assign N479 = N3091;
  assign N480 = N3090;
  assign N481 = N3089;
  assign N482 = N3088;
  assign N483 = N3087;
  assign N484 = N3086;
  assign N485 = N3085;
  assign N486 = N3084;
  assign N487 = N3083;
  assign N488 = N3082;
  assign N489 = N3081;
  assign N490 = N3080;
  assign N491 = N3079;
  assign N492 = N3078;
  assign N493 = N3077;
  assign N494 = N3076;
  assign N495 = N3075;
  assign N496 = N3074;
  assign N497 = N3073;
  assign N498 = N3072;
  assign N499 = N3071;
  assign N500 = N3070;
  assign N501 = N3069;
  assign N502 = N3068;
  assign N503 = N3067;
  assign N504 = N3066;
  assign N505 = N3065;
  assign N506 = N3064;
  assign N507 = N3063;
  assign N508 = N3062;
  assign N509 = N3061;
  assign N510 = N3060;
  assign N511 = N3059;
  assign N512 = N3058;
  assign N513 = N3057;
  assign N514 = N3056;
  assign N515 = N3055;
  assign N516 = N3054;
  assign N517 = N3053;
  assign N518 = N3052;
  assign N519 = N3051;
  assign N520 = N3050;
  assign N521 = N3049;
  assign N522 = N3048;
  assign N523 = N3047;
  assign N524 = N3046;
  assign N525 = N3045;
  assign N526 = N3044;
  assign N527 = N3043;
  assign N528 = N3042;
  assign N529 = N3041;
  assign N530 = N3040;
  assign N531 = N3039;
  assign N532 = N3038;
  assign N533 = N3037;
  assign N534 = N3036;
  assign N535 = N3035;
  assign N536 = N3034;
  assign N537 = N3033;
  assign N538 = N3032;
  assign N539 = N3031;
  assign N540 = N3030;
  assign N541 = N3029;
  assign N542 = N3028;
  assign N543 = N3027;
  assign N544 = N3026;
  assign N545 = N3025;
  assign N546 = N3024;
  assign N547 = N3023;
  assign N548 = N3022;
  assign N549 = N3021;
  assign N550 = N3020;
  assign N551 = N3019;
  assign N552 = N3018;
  assign N553 = N3017;
  assign N554 = N3016;
  assign N555 = N3015;
  assign N556 = N3014;
  assign N557 = N3013;
  assign N558 = N3012;
  assign N559 = N3011;
  assign N560 = N3010;
  assign data_nn[255:224] = (N440)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N441)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N442)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N443)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N444)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N445)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N446)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N447)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N448)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N449)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N450)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N451)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N452)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N453)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N454)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N455)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N456)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N457)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N458)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N459)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N460)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N461)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N462)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N463)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N464)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N465)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N466)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N467)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N468)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N469)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N470)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N471)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N472)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N473)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N474)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N475)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N476)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N477)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N478)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N479)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N480)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N481)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N482)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N483)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N484)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N485)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N486)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N487)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N488)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N489)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N490)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N491)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N492)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N493)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N494)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N495)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N496)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N497)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N498)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N499)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N500)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N501)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N502)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N503)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N504)? data_o[2047:2016] : 
                            (N505)? data_o[2015:1984] : 
                            (N506)? data_o[1983:1952] : 
                            (N507)? data_o[1951:1920] : 
                            (N508)? data_o[1919:1888] : 
                            (N509)? data_o[1887:1856] : 
                            (N510)? data_o[1855:1824] : 
                            (N511)? data_o[1823:1792] : 
                            (N512)? data_o[1791:1760] : 
                            (N513)? data_o[1759:1728] : 
                            (N514)? data_o[1727:1696] : 
                            (N515)? data_o[1695:1664] : 
                            (N516)? data_o[1663:1632] : 
                            (N517)? data_o[1631:1600] : 
                            (N518)? data_o[1599:1568] : 
                            (N519)? data_o[1567:1536] : 
                            (N520)? data_o[1535:1504] : 
                            (N521)? data_o[1503:1472] : 
                            (N522)? data_o[1471:1440] : 
                            (N523)? data_o[1439:1408] : 
                            (N524)? data_o[1407:1376] : 
                            (N525)? data_o[1375:1344] : 
                            (N526)? data_o[1343:1312] : 
                            (N527)? data_o[1311:1280] : 
                            (N528)? data_o[1279:1248] : 
                            (N529)? data_o[1247:1216] : 
                            (N530)? data_o[1215:1184] : 
                            (N531)? data_o[1183:1152] : 
                            (N532)? data_o[1151:1120] : 
                            (N533)? data_o[1119:1088] : 
                            (N534)? data_o[1087:1056] : 
                            (N535)? data_o[1055:1024] : 
                            (N536)? data_o[1023:992] : 
                            (N537)? data_o[991:960] : 
                            (N538)? data_o[959:928] : 
                            (N539)? data_o[927:896] : 
                            (N540)? data_o[895:864] : 
                            (N541)? data_o[863:832] : 
                            (N542)? data_o[831:800] : 
                            (N543)? data_o[799:768] : 
                            (N544)? data_o[767:736] : 
                            (N545)? data_o[735:704] : 
                            (N546)? data_o[703:672] : 
                            (N547)? data_o[671:640] : 
                            (N548)? data_o[639:608] : 
                            (N549)? data_o[607:576] : 
                            (N550)? data_o[575:544] : 
                            (N551)? data_o[543:512] : 
                            (N552)? data_o[511:480] : 
                            (N553)? data_o[479:448] : 
                            (N554)? data_o[447:416] : 
                            (N555)? data_o[415:384] : 
                            (N556)? data_o[383:352] : 
                            (N557)? data_o[351:320] : 
                            (N558)? data_o[319:288] : 
                            (N559)? data_o[287:256] : 
                            (N560)? data_o[255:224] : 1'b0;
  assign data_nn[287:256] = (N441)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N442)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N443)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N444)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N445)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N446)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N447)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N448)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N449)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N450)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N451)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N452)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N453)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N454)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N455)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N456)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N457)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N458)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N459)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N460)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N461)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N462)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N463)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N464)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N465)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N466)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N467)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N468)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N469)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N470)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N471)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N472)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N473)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N474)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N475)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N476)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N477)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N478)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N479)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N480)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N481)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N482)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N483)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N484)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N485)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N486)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N487)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N488)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N489)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N490)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N491)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N492)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N493)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N494)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N495)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N496)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N497)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N498)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N499)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N500)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N501)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N502)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N503)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N504)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N505)? data_o[2047:2016] : 
                            (N506)? data_o[2015:1984] : 
                            (N507)? data_o[1983:1952] : 
                            (N508)? data_o[1951:1920] : 
                            (N509)? data_o[1919:1888] : 
                            (N510)? data_o[1887:1856] : 
                            (N511)? data_o[1855:1824] : 
                            (N512)? data_o[1823:1792] : 
                            (N513)? data_o[1791:1760] : 
                            (N514)? data_o[1759:1728] : 
                            (N515)? data_o[1727:1696] : 
                            (N516)? data_o[1695:1664] : 
                            (N517)? data_o[1663:1632] : 
                            (N518)? data_o[1631:1600] : 
                            (N519)? data_o[1599:1568] : 
                            (N520)? data_o[1567:1536] : 
                            (N521)? data_o[1535:1504] : 
                            (N522)? data_o[1503:1472] : 
                            (N523)? data_o[1471:1440] : 
                            (N524)? data_o[1439:1408] : 
                            (N525)? data_o[1407:1376] : 
                            (N526)? data_o[1375:1344] : 
                            (N527)? data_o[1343:1312] : 
                            (N528)? data_o[1311:1280] : 
                            (N529)? data_o[1279:1248] : 
                            (N530)? data_o[1247:1216] : 
                            (N531)? data_o[1215:1184] : 
                            (N532)? data_o[1183:1152] : 
                            (N533)? data_o[1151:1120] : 
                            (N534)? data_o[1119:1088] : 
                            (N535)? data_o[1087:1056] : 
                            (N536)? data_o[1055:1024] : 
                            (N537)? data_o[1023:992] : 
                            (N538)? data_o[991:960] : 
                            (N539)? data_o[959:928] : 
                            (N540)? data_o[927:896] : 
                            (N541)? data_o[895:864] : 
                            (N542)? data_o[863:832] : 
                            (N543)? data_o[831:800] : 
                            (N544)? data_o[799:768] : 
                            (N545)? data_o[767:736] : 
                            (N546)? data_o[735:704] : 
                            (N547)? data_o[703:672] : 
                            (N548)? data_o[671:640] : 
                            (N549)? data_o[639:608] : 
                            (N550)? data_o[607:576] : 
                            (N551)? data_o[575:544] : 
                            (N552)? data_o[543:512] : 
                            (N553)? data_o[511:480] : 
                            (N554)? data_o[479:448] : 
                            (N555)? data_o[447:416] : 
                            (N556)? data_o[415:384] : 
                            (N557)? data_o[383:352] : 
                            (N558)? data_o[351:320] : 
                            (N559)? data_o[319:288] : 
                            (N560)? data_o[287:256] : 1'b0;
  assign data_nn[319:288] = (N442)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N443)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N444)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N445)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N446)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N447)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N448)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N449)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N450)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N451)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N452)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N453)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N454)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N455)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N456)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N457)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N458)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N459)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N460)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N461)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N462)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N463)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N464)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N465)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N466)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N467)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N468)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N469)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N470)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N471)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N472)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N473)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N474)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N475)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N476)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N477)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N478)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N479)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N480)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N481)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N482)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N483)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N484)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N485)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N486)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N487)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N488)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N489)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N490)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N491)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N492)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N493)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N494)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N495)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N496)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N497)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N498)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N499)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N500)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N501)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N502)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N503)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N504)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N505)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N506)? data_o[2047:2016] : 
                            (N507)? data_o[2015:1984] : 
                            (N508)? data_o[1983:1952] : 
                            (N509)? data_o[1951:1920] : 
                            (N510)? data_o[1919:1888] : 
                            (N511)? data_o[1887:1856] : 
                            (N512)? data_o[1855:1824] : 
                            (N513)? data_o[1823:1792] : 
                            (N514)? data_o[1791:1760] : 
                            (N515)? data_o[1759:1728] : 
                            (N516)? data_o[1727:1696] : 
                            (N517)? data_o[1695:1664] : 
                            (N518)? data_o[1663:1632] : 
                            (N519)? data_o[1631:1600] : 
                            (N520)? data_o[1599:1568] : 
                            (N521)? data_o[1567:1536] : 
                            (N522)? data_o[1535:1504] : 
                            (N523)? data_o[1503:1472] : 
                            (N524)? data_o[1471:1440] : 
                            (N525)? data_o[1439:1408] : 
                            (N526)? data_o[1407:1376] : 
                            (N527)? data_o[1375:1344] : 
                            (N528)? data_o[1343:1312] : 
                            (N529)? data_o[1311:1280] : 
                            (N530)? data_o[1279:1248] : 
                            (N531)? data_o[1247:1216] : 
                            (N532)? data_o[1215:1184] : 
                            (N533)? data_o[1183:1152] : 
                            (N534)? data_o[1151:1120] : 
                            (N535)? data_o[1119:1088] : 
                            (N536)? data_o[1087:1056] : 
                            (N537)? data_o[1055:1024] : 
                            (N538)? data_o[1023:992] : 
                            (N539)? data_o[991:960] : 
                            (N540)? data_o[959:928] : 
                            (N541)? data_o[927:896] : 
                            (N542)? data_o[895:864] : 
                            (N543)? data_o[863:832] : 
                            (N544)? data_o[831:800] : 
                            (N545)? data_o[799:768] : 
                            (N546)? data_o[767:736] : 
                            (N547)? data_o[735:704] : 
                            (N548)? data_o[703:672] : 
                            (N549)? data_o[671:640] : 
                            (N550)? data_o[639:608] : 
                            (N551)? data_o[607:576] : 
                            (N552)? data_o[575:544] : 
                            (N553)? data_o[543:512] : 
                            (N554)? data_o[511:480] : 
                            (N555)? data_o[479:448] : 
                            (N556)? data_o[447:416] : 
                            (N557)? data_o[415:384] : 
                            (N558)? data_o[383:352] : 
                            (N559)? data_o[351:320] : 
                            (N560)? data_o[319:288] : 1'b0;
  assign data_nn[351:320] = (N443)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N444)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N445)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N446)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N447)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N448)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N449)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N450)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N451)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N452)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N453)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N454)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N455)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N456)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N457)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N458)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N459)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N460)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N461)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N462)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N463)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N464)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N465)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N466)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N467)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N468)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N469)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N470)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N471)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N472)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N473)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N474)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N475)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N476)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N477)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N478)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N479)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N480)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N481)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N482)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N483)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N484)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N485)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N486)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N487)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N488)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N489)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N490)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N491)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N492)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N493)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N494)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N495)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N496)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N497)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N498)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N499)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N500)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N501)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N502)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N503)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N504)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N505)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N506)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N507)? data_o[2047:2016] : 
                            (N508)? data_o[2015:1984] : 
                            (N509)? data_o[1983:1952] : 
                            (N510)? data_o[1951:1920] : 
                            (N511)? data_o[1919:1888] : 
                            (N512)? data_o[1887:1856] : 
                            (N513)? data_o[1855:1824] : 
                            (N514)? data_o[1823:1792] : 
                            (N515)? data_o[1791:1760] : 
                            (N516)? data_o[1759:1728] : 
                            (N517)? data_o[1727:1696] : 
                            (N518)? data_o[1695:1664] : 
                            (N519)? data_o[1663:1632] : 
                            (N520)? data_o[1631:1600] : 
                            (N521)? data_o[1599:1568] : 
                            (N522)? data_o[1567:1536] : 
                            (N523)? data_o[1535:1504] : 
                            (N524)? data_o[1503:1472] : 
                            (N525)? data_o[1471:1440] : 
                            (N526)? data_o[1439:1408] : 
                            (N527)? data_o[1407:1376] : 
                            (N528)? data_o[1375:1344] : 
                            (N529)? data_o[1343:1312] : 
                            (N530)? data_o[1311:1280] : 
                            (N531)? data_o[1279:1248] : 
                            (N532)? data_o[1247:1216] : 
                            (N533)? data_o[1215:1184] : 
                            (N534)? data_o[1183:1152] : 
                            (N535)? data_o[1151:1120] : 
                            (N536)? data_o[1119:1088] : 
                            (N537)? data_o[1087:1056] : 
                            (N538)? data_o[1055:1024] : 
                            (N539)? data_o[1023:992] : 
                            (N540)? data_o[991:960] : 
                            (N541)? data_o[959:928] : 
                            (N542)? data_o[927:896] : 
                            (N543)? data_o[895:864] : 
                            (N544)? data_o[863:832] : 
                            (N545)? data_o[831:800] : 
                            (N546)? data_o[799:768] : 
                            (N547)? data_o[767:736] : 
                            (N548)? data_o[735:704] : 
                            (N549)? data_o[703:672] : 
                            (N550)? data_o[671:640] : 
                            (N551)? data_o[639:608] : 
                            (N552)? data_o[607:576] : 
                            (N553)? data_o[575:544] : 
                            (N554)? data_o[543:512] : 
                            (N555)? data_o[511:480] : 
                            (N556)? data_o[479:448] : 
                            (N557)? data_o[447:416] : 
                            (N558)? data_o[415:384] : 
                            (N559)? data_o[383:352] : 
                            (N560)? data_o[351:320] : 1'b0;
  assign data_nn[383:352] = (N561)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N562)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N563)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N564)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N565)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N566)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N567)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N568)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N569)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N570)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N571)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N572)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N573)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N574)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N575)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N576)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N577)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N578)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N579)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N580)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N581)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N582)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N583)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N584)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N585)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N586)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N587)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N588)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N589)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N590)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N591)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N592)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N593)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N594)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N595)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N596)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N597)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N598)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N599)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N600)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N601)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N602)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N603)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N604)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N605)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N606)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N607)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N608)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N609)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N610)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N611)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N612)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N613)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N614)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N615)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N616)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N617)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N618)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N619)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N620)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N621)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N622)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N623)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N624)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N625)? data_o[2047:2016] : 
                            (N626)? data_o[2015:1984] : 
                            (N627)? data_o[1983:1952] : 
                            (N628)? data_o[1951:1920] : 
                            (N629)? data_o[1919:1888] : 
                            (N630)? data_o[1887:1856] : 
                            (N631)? data_o[1855:1824] : 
                            (N632)? data_o[1823:1792] : 
                            (N633)? data_o[1791:1760] : 
                            (N634)? data_o[1759:1728] : 
                            (N635)? data_o[1727:1696] : 
                            (N636)? data_o[1695:1664] : 
                            (N637)? data_o[1663:1632] : 
                            (N638)? data_o[1631:1600] : 
                            (N639)? data_o[1599:1568] : 
                            (N640)? data_o[1567:1536] : 
                            (N641)? data_o[1535:1504] : 
                            (N642)? data_o[1503:1472] : 
                            (N643)? data_o[1471:1440] : 
                            (N644)? data_o[1439:1408] : 
                            (N645)? data_o[1407:1376] : 
                            (N646)? data_o[1375:1344] : 
                            (N647)? data_o[1343:1312] : 
                            (N648)? data_o[1311:1280] : 
                            (N649)? data_o[1279:1248] : 
                            (N650)? data_o[1247:1216] : 
                            (N651)? data_o[1215:1184] : 
                            (N652)? data_o[1183:1152] : 
                            (N653)? data_o[1151:1120] : 
                            (N654)? data_o[1119:1088] : 
                            (N655)? data_o[1087:1056] : 
                            (N656)? data_o[1055:1024] : 
                            (N657)? data_o[1023:992] : 
                            (N658)? data_o[991:960] : 
                            (N659)? data_o[959:928] : 
                            (N660)? data_o[927:896] : 
                            (N661)? data_o[895:864] : 
                            (N662)? data_o[863:832] : 
                            (N663)? data_o[831:800] : 
                            (N664)? data_o[799:768] : 
                            (N665)? data_o[767:736] : 
                            (N666)? data_o[735:704] : 
                            (N667)? data_o[703:672] : 
                            (N668)? data_o[671:640] : 
                            (N669)? data_o[639:608] : 
                            (N670)? data_o[607:576] : 
                            (N671)? data_o[575:544] : 
                            (N672)? data_o[543:512] : 
                            (N673)? data_o[511:480] : 
                            (N674)? data_o[479:448] : 
                            (N675)? data_o[447:416] : 
                            (N676)? data_o[415:384] : 
                            (N677)? data_o[383:352] : 1'b0;
  assign N561 = N3244;
  assign N562 = N3243;
  assign N563 = N3242;
  assign N564 = N3241;
  assign N565 = N3240;
  assign N566 = N3239;
  assign N567 = N3238;
  assign N568 = N3237;
  assign N569 = N3236;
  assign N570 = N3235;
  assign N571 = N3234;
  assign N572 = N3233;
  assign N573 = N3232;
  assign N574 = N3231;
  assign N575 = N3230;
  assign N576 = N3229;
  assign N577 = N3228;
  assign N578 = N3227;
  assign N579 = N3226;
  assign N580 = N3225;
  assign N581 = N3224;
  assign N582 = N3223;
  assign N583 = N3222;
  assign N584 = N3221;
  assign N585 = N3220;
  assign N586 = N3219;
  assign N587 = N3218;
  assign N588 = N3217;
  assign N589 = N3216;
  assign N590 = N3215;
  assign N591 = N3214;
  assign N592 = N3213;
  assign N593 = N3212;
  assign N594 = N3211;
  assign N595 = N3210;
  assign N596 = N3209;
  assign N597 = N3208;
  assign N598 = N3207;
  assign N599 = N3206;
  assign N600 = N3205;
  assign N601 = N3204;
  assign N602 = N3203;
  assign N603 = N3202;
  assign N604 = N3201;
  assign N605 = N3200;
  assign N606 = N3199;
  assign N607 = N3198;
  assign N608 = N3197;
  assign N609 = N3196;
  assign N610 = N3195;
  assign N611 = N3194;
  assign N612 = N3193;
  assign N613 = N3192;
  assign N614 = N3191;
  assign N615 = N3190;
  assign N616 = N3189;
  assign N617 = N3188;
  assign N618 = N3187;
  assign N619 = N3186;
  assign N620 = N3185;
  assign N621 = N3184;
  assign N622 = N3183;
  assign N623 = N3182;
  assign N624 = N3181;
  assign N625 = N3180;
  assign N626 = N3179;
  assign N627 = N3178;
  assign N628 = N3177;
  assign N629 = N3176;
  assign N630 = N3175;
  assign N631 = N3174;
  assign N632 = N3173;
  assign N633 = N3172;
  assign N634 = N3171;
  assign N635 = N3170;
  assign N636 = N3169;
  assign N637 = N3168;
  assign N638 = N3167;
  assign N639 = N3166;
  assign N640 = N3165;
  assign N641 = N3164;
  assign N642 = N3163;
  assign N643 = N3162;
  assign N644 = N3161;
  assign N645 = N3160;
  assign N646 = N3159;
  assign N647 = N3158;
  assign N648 = N3157;
  assign N649 = N3156;
  assign N650 = N3155;
  assign N651 = N3154;
  assign N652 = N3153;
  assign N653 = N3152;
  assign N654 = N3151;
  assign N655 = N3150;
  assign N656 = N3149;
  assign N657 = N3148;
  assign N658 = N3147;
  assign N659 = N3146;
  assign N660 = N3145;
  assign N661 = N3144;
  assign N662 = N3143;
  assign N663 = N3142;
  assign N664 = N3141;
  assign N665 = N3140;
  assign N666 = N3139;
  assign N667 = N3138;
  assign N668 = N3137;
  assign N669 = N3136;
  assign N670 = N3135;
  assign N671 = N3134;
  assign N672 = N3133;
  assign N673 = N3132;
  assign N674 = N3131;
  assign N675 = N3130;
  assign N676 = N3129;
  assign N677 = N3128;
  assign data_nn[415:384] = (N678)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N679)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N680)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N681)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N682)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N683)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N684)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N685)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N686)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N687)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N688)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N689)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N690)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N691)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N692)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N693)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N694)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N695)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N696)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N697)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N698)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N699)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N700)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N701)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N702)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N703)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N704)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N705)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N706)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N707)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N708)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N709)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N710)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N711)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N712)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N713)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N714)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N715)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N716)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N717)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N718)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N719)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N720)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N721)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N722)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N723)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N724)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N725)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N726)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N727)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N728)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N729)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N730)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N731)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N732)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N733)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N734)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N735)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N736)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N737)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N738)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N739)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N740)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N741)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N742)? data_o[2047:2016] : 
                            (N743)? data_o[2015:1984] : 
                            (N744)? data_o[1983:1952] : 
                            (N745)? data_o[1951:1920] : 
                            (N746)? data_o[1919:1888] : 
                            (N747)? data_o[1887:1856] : 
                            (N748)? data_o[1855:1824] : 
                            (N749)? data_o[1823:1792] : 
                            (N750)? data_o[1791:1760] : 
                            (N751)? data_o[1759:1728] : 
                            (N752)? data_o[1727:1696] : 
                            (N753)? data_o[1695:1664] : 
                            (N754)? data_o[1663:1632] : 
                            (N755)? data_o[1631:1600] : 
                            (N756)? data_o[1599:1568] : 
                            (N757)? data_o[1567:1536] : 
                            (N758)? data_o[1535:1504] : 
                            (N759)? data_o[1503:1472] : 
                            (N760)? data_o[1471:1440] : 
                            (N761)? data_o[1439:1408] : 
                            (N762)? data_o[1407:1376] : 
                            (N763)? data_o[1375:1344] : 
                            (N764)? data_o[1343:1312] : 
                            (N765)? data_o[1311:1280] : 
                            (N766)? data_o[1279:1248] : 
                            (N767)? data_o[1247:1216] : 
                            (N768)? data_o[1215:1184] : 
                            (N769)? data_o[1183:1152] : 
                            (N770)? data_o[1151:1120] : 
                            (N771)? data_o[1119:1088] : 
                            (N772)? data_o[1087:1056] : 
                            (N773)? data_o[1055:1024] : 
                            (N774)? data_o[1023:992] : 
                            (N775)? data_o[991:960] : 
                            (N776)? data_o[959:928] : 
                            (N777)? data_o[927:896] : 
                            (N778)? data_o[895:864] : 
                            (N779)? data_o[863:832] : 
                            (N780)? data_o[831:800] : 
                            (N781)? data_o[799:768] : 
                            (N782)? data_o[767:736] : 
                            (N783)? data_o[735:704] : 
                            (N784)? data_o[703:672] : 
                            (N785)? data_o[671:640] : 
                            (N786)? data_o[639:608] : 
                            (N787)? data_o[607:576] : 
                            (N788)? data_o[575:544] : 
                            (N789)? data_o[543:512] : 
                            (N790)? data_o[511:480] : 
                            (N791)? data_o[479:448] : 
                            (N792)? data_o[447:416] : 
                            (N793)? data_o[415:384] : 1'b0;
  assign N678 = N3360;
  assign N679 = N3359;
  assign N680 = N3358;
  assign N681 = N3357;
  assign N682 = N3356;
  assign N683 = N3355;
  assign N684 = N3354;
  assign N685 = N3353;
  assign N686 = N3352;
  assign N687 = N3351;
  assign N688 = N3350;
  assign N689 = N3349;
  assign N690 = N3348;
  assign N691 = N3347;
  assign N692 = N3346;
  assign N693 = N3345;
  assign N694 = N3344;
  assign N695 = N3343;
  assign N696 = N3342;
  assign N697 = N3341;
  assign N698 = N3340;
  assign N699 = N3339;
  assign N700 = N3338;
  assign N701 = N3337;
  assign N702 = N3336;
  assign N703 = N3335;
  assign N704 = N3334;
  assign N705 = N3333;
  assign N706 = N3332;
  assign N707 = N3331;
  assign N708 = N3330;
  assign N709 = N3329;
  assign N710 = N3328;
  assign N711 = N3327;
  assign N712 = N3326;
  assign N713 = N3325;
  assign N714 = N3324;
  assign N715 = N3323;
  assign N716 = N3322;
  assign N717 = N3321;
  assign N718 = N3320;
  assign N719 = N3319;
  assign N720 = N3318;
  assign N721 = N3317;
  assign N722 = N3316;
  assign N723 = N3315;
  assign N724 = N3314;
  assign N725 = N3313;
  assign N726 = N3312;
  assign N727 = N3311;
  assign N728 = N3310;
  assign N729 = N3309;
  assign N730 = N3308;
  assign N731 = N3307;
  assign N732 = N3306;
  assign N733 = N3305;
  assign N734 = N3304;
  assign N735 = N3303;
  assign N736 = N3302;
  assign N737 = N3301;
  assign N738 = N3300;
  assign N739 = N3299;
  assign N740 = N3298;
  assign N741 = N3297;
  assign N742 = N3296;
  assign N743 = N3295;
  assign N744 = N3294;
  assign N745 = N3293;
  assign N746 = N3292;
  assign N747 = N3291;
  assign N748 = N3290;
  assign N749 = N3289;
  assign N750 = N3288;
  assign N751 = N3287;
  assign N752 = N3286;
  assign N753 = N3285;
  assign N754 = N3284;
  assign N755 = N3283;
  assign N756 = N3282;
  assign N757 = N3281;
  assign N758 = N3280;
  assign N759 = N3279;
  assign N760 = N3278;
  assign N761 = N3277;
  assign N762 = N3276;
  assign N763 = N3275;
  assign N764 = N3274;
  assign N765 = N3273;
  assign N766 = N3272;
  assign N767 = N3271;
  assign N768 = N3270;
  assign N769 = N3269;
  assign N770 = N3268;
  assign N771 = N3267;
  assign N772 = N3266;
  assign N773 = N3265;
  assign N774 = N3264;
  assign N775 = N3263;
  assign N776 = N3262;
  assign N777 = N3261;
  assign N778 = N3260;
  assign N779 = N3259;
  assign N780 = N3258;
  assign N781 = N3257;
  assign N782 = N3256;
  assign N783 = N3255;
  assign N784 = N3254;
  assign N785 = N3253;
  assign N786 = N3252;
  assign N787 = N3251;
  assign N788 = N3250;
  assign N789 = N3249;
  assign N790 = N3248;
  assign N791 = N3247;
  assign N792 = N3246;
  assign N793 = N3245;
  assign data_nn[447:416] = (N324)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N325)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N326)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N327)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N328)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N329)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N330)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N331)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N332)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N333)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N334)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N335)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N336)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N337)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N338)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N339)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N340)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N341)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N342)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N343)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N344)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N345)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N346)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N347)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N348)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N349)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N350)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N351)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N352)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N353)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N354)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N355)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N356)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N357)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N358)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N359)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N360)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N361)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N362)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N363)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N364)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N365)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N366)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N367)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N368)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N369)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N370)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N371)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N372)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N373)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N374)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N375)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N376)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N377)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N378)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N379)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N380)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N381)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N382)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N383)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N384)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N385)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N386)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N387)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N388)? data_o[2047:2016] : 
                            (N389)? data_o[2015:1984] : 
                            (N390)? data_o[1983:1952] : 
                            (N391)? data_o[1951:1920] : 
                            (N392)? data_o[1919:1888] : 
                            (N393)? data_o[1887:1856] : 
                            (N394)? data_o[1855:1824] : 
                            (N395)? data_o[1823:1792] : 
                            (N396)? data_o[1791:1760] : 
                            (N397)? data_o[1759:1728] : 
                            (N398)? data_o[1727:1696] : 
                            (N399)? data_o[1695:1664] : 
                            (N400)? data_o[1663:1632] : 
                            (N401)? data_o[1631:1600] : 
                            (N402)? data_o[1599:1568] : 
                            (N403)? data_o[1567:1536] : 
                            (N404)? data_o[1535:1504] : 
                            (N405)? data_o[1503:1472] : 
                            (N406)? data_o[1471:1440] : 
                            (N407)? data_o[1439:1408] : 
                            (N408)? data_o[1407:1376] : 
                            (N409)? data_o[1375:1344] : 
                            (N410)? data_o[1343:1312] : 
                            (N411)? data_o[1311:1280] : 
                            (N412)? data_o[1279:1248] : 
                            (N413)? data_o[1247:1216] : 
                            (N414)? data_o[1215:1184] : 
                            (N415)? data_o[1183:1152] : 
                            (N416)? data_o[1151:1120] : 
                            (N417)? data_o[1119:1088] : 
                            (N418)? data_o[1087:1056] : 
                            (N419)? data_o[1055:1024] : 
                            (N420)? data_o[1023:992] : 
                            (N421)? data_o[991:960] : 
                            (N422)? data_o[959:928] : 
                            (N423)? data_o[927:896] : 
                            (N424)? data_o[895:864] : 
                            (N425)? data_o[863:832] : 
                            (N426)? data_o[831:800] : 
                            (N427)? data_o[799:768] : 
                            (N428)? data_o[767:736] : 
                            (N429)? data_o[735:704] : 
                            (N430)? data_o[703:672] : 
                            (N431)? data_o[671:640] : 
                            (N432)? data_o[639:608] : 
                            (N433)? data_o[607:576] : 
                            (N434)? data_o[575:544] : 
                            (N435)? data_o[543:512] : 
                            (N436)? data_o[511:480] : 
                            (N437)? data_o[479:448] : 
                            (N438)? data_o[447:416] : 1'b0;
  assign data_nn[479:448] = (N794)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N795)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N796)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N797)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N798)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N799)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N800)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N801)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N802)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N803)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N804)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N805)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N806)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N807)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N808)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N809)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N810)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N811)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N812)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N813)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N814)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N815)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N816)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N817)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N818)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N819)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N820)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N821)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N822)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N823)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N824)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N825)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N826)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N827)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N828)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N829)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N830)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N831)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N832)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N833)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N834)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N835)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N836)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N837)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N838)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N839)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N840)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N841)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N842)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N843)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N844)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N845)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N846)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N847)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N848)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N849)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N850)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N851)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N852)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N853)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N854)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N855)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N856)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N857)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N858)? data_o[2047:2016] : 
                            (N859)? data_o[2015:1984] : 
                            (N860)? data_o[1983:1952] : 
                            (N861)? data_o[1951:1920] : 
                            (N862)? data_o[1919:1888] : 
                            (N863)? data_o[1887:1856] : 
                            (N864)? data_o[1855:1824] : 
                            (N865)? data_o[1823:1792] : 
                            (N866)? data_o[1791:1760] : 
                            (N867)? data_o[1759:1728] : 
                            (N868)? data_o[1727:1696] : 
                            (N869)? data_o[1695:1664] : 
                            (N870)? data_o[1663:1632] : 
                            (N871)? data_o[1631:1600] : 
                            (N872)? data_o[1599:1568] : 
                            (N873)? data_o[1567:1536] : 
                            (N874)? data_o[1535:1504] : 
                            (N875)? data_o[1503:1472] : 
                            (N876)? data_o[1471:1440] : 
                            (N877)? data_o[1439:1408] : 
                            (N878)? data_o[1407:1376] : 
                            (N879)? data_o[1375:1344] : 
                            (N880)? data_o[1343:1312] : 
                            (N881)? data_o[1311:1280] : 
                            (N882)? data_o[1279:1248] : 
                            (N883)? data_o[1247:1216] : 
                            (N884)? data_o[1215:1184] : 
                            (N885)? data_o[1183:1152] : 
                            (N886)? data_o[1151:1120] : 
                            (N887)? data_o[1119:1088] : 
                            (N888)? data_o[1087:1056] : 
                            (N889)? data_o[1055:1024] : 
                            (N890)? data_o[1023:992] : 
                            (N891)? data_o[991:960] : 
                            (N892)? data_o[959:928] : 
                            (N893)? data_o[927:896] : 
                            (N894)? data_o[895:864] : 
                            (N895)? data_o[863:832] : 
                            (N896)? data_o[831:800] : 
                            (N897)? data_o[799:768] : 
                            (N898)? data_o[767:736] : 
                            (N899)? data_o[735:704] : 
                            (N900)? data_o[703:672] : 
                            (N901)? data_o[671:640] : 
                            (N902)? data_o[639:608] : 
                            (N903)? data_o[607:576] : 
                            (N904)? data_o[575:544] : 
                            (N905)? data_o[543:512] : 
                            (N906)? data_o[511:480] : 
                            (N907)? data_o[479:448] : 1'b0;
  assign N794 = N5534;
  assign N795 = N5535;
  assign N796 = N5536;
  assign N797 = N5537;
  assign N798 = N3521;
  assign N799 = N3520;
  assign N800 = N3519;
  assign N801 = N3518;
  assign N802 = N3517;
  assign N803 = N3516;
  assign N804 = N3515;
  assign N805 = N3514;
  assign N806 = N3513;
  assign N807 = N3512;
  assign N808 = N3511;
  assign N809 = N3510;
  assign N810 = N3509;
  assign N811 = N3508;
  assign N812 = N3507;
  assign N813 = N3506;
  assign N814 = N3505;
  assign N815 = N3504;
  assign N816 = N3503;
  assign N817 = N3502;
  assign N818 = N3501;
  assign N819 = N3500;
  assign N820 = N3499;
  assign N821 = N3498;
  assign N822 = N3497;
  assign N823 = N3496;
  assign N824 = N3495;
  assign N825 = N3494;
  assign N826 = N3493;
  assign N827 = N3492;
  assign N828 = N3491;
  assign N829 = N3490;
  assign N830 = N3489;
  assign N831 = N3488;
  assign N832 = N3487;
  assign N833 = N3486;
  assign N834 = N3485;
  assign N835 = N3484;
  assign N836 = N3483;
  assign N837 = N3482;
  assign N838 = N3481;
  assign N839 = N3480;
  assign N840 = N3479;
  assign N841 = N3478;
  assign N842 = N3477;
  assign N843 = N3476;
  assign N844 = N4236;
  assign N845 = N4235;
  assign N846 = N4234;
  assign N847 = N4233;
  assign N848 = N4232;
  assign N849 = N4231;
  assign N850 = N4230;
  assign N851 = N4229;
  assign N852 = N4228;
  assign N853 = N4227;
  assign N854 = N4226;
  assign N855 = N4225;
  assign N856 = N4224;
  assign N857 = N4223;
  assign N858 = N4222;
  assign N859 = N4221;
  assign N860 = N4220;
  assign N861 = N4219;
  assign N862 = N4218;
  assign N863 = N4217;
  assign N864 = N4216;
  assign N865 = N4215;
  assign N866 = N4214;
  assign N867 = N4213;
  assign N868 = N4212;
  assign N869 = N4211;
  assign N870 = N4210;
  assign N871 = N4209;
  assign N872 = N4208;
  assign N873 = N4207;
  assign N874 = N4206;
  assign N875 = N4205;
  assign N876 = N4204;
  assign N877 = N4203;
  assign N878 = N4202;
  assign N879 = N4201;
  assign N880 = N4200;
  assign N881 = N4199;
  assign N882 = N4198;
  assign N883 = N4197;
  assign N884 = N4196;
  assign N885 = N4195;
  assign N886 = N4194;
  assign N887 = N4193;
  assign N888 = N4192;
  assign N889 = N4191;
  assign N890 = N4190;
  assign N891 = N4189;
  assign N892 = N4188;
  assign N893 = N4187;
  assign N894 = N4186;
  assign N895 = N4185;
  assign N896 = N4184;
  assign N897 = N4183;
  assign N898 = N4182;
  assign N899 = N4181;
  assign N900 = N4180;
  assign N901 = N4179;
  assign N902 = N4178;
  assign N903 = N4177;
  assign N904 = N4176;
  assign N905 = N4175;
  assign N906 = N4174;
  assign N907 = N4173;
  assign data_nn[511:480] = (N795)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N796)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N797)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N798)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N799)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N800)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N801)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N802)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N803)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N804)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N805)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N806)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N807)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N808)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N809)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N810)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N811)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N812)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N813)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N814)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N815)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N816)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N817)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N818)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N819)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N820)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N821)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N822)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N823)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N824)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N825)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N826)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N827)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N828)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N829)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N830)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N831)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N832)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N833)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N834)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N835)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N836)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N837)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N838)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N839)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N840)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N841)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N842)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N843)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N844)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N845)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N846)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N847)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N848)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N849)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N850)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N851)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N852)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N853)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N854)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N855)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N856)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N857)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N858)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N859)? data_o[2047:2016] : 
                            (N860)? data_o[2015:1984] : 
                            (N861)? data_o[1983:1952] : 
                            (N862)? data_o[1951:1920] : 
                            (N863)? data_o[1919:1888] : 
                            (N864)? data_o[1887:1856] : 
                            (N865)? data_o[1855:1824] : 
                            (N866)? data_o[1823:1792] : 
                            (N867)? data_o[1791:1760] : 
                            (N868)? data_o[1759:1728] : 
                            (N869)? data_o[1727:1696] : 
                            (N870)? data_o[1695:1664] : 
                            (N871)? data_o[1663:1632] : 
                            (N872)? data_o[1631:1600] : 
                            (N873)? data_o[1599:1568] : 
                            (N874)? data_o[1567:1536] : 
                            (N875)? data_o[1535:1504] : 
                            (N876)? data_o[1503:1472] : 
                            (N877)? data_o[1471:1440] : 
                            (N878)? data_o[1439:1408] : 
                            (N879)? data_o[1407:1376] : 
                            (N880)? data_o[1375:1344] : 
                            (N881)? data_o[1343:1312] : 
                            (N882)? data_o[1311:1280] : 
                            (N883)? data_o[1279:1248] : 
                            (N884)? data_o[1247:1216] : 
                            (N885)? data_o[1215:1184] : 
                            (N886)? data_o[1183:1152] : 
                            (N887)? data_o[1151:1120] : 
                            (N888)? data_o[1119:1088] : 
                            (N889)? data_o[1087:1056] : 
                            (N890)? data_o[1055:1024] : 
                            (N891)? data_o[1023:992] : 
                            (N892)? data_o[991:960] : 
                            (N893)? data_o[959:928] : 
                            (N894)? data_o[927:896] : 
                            (N895)? data_o[895:864] : 
                            (N896)? data_o[863:832] : 
                            (N897)? data_o[831:800] : 
                            (N898)? data_o[799:768] : 
                            (N899)? data_o[767:736] : 
                            (N900)? data_o[735:704] : 
                            (N901)? data_o[703:672] : 
                            (N902)? data_o[671:640] : 
                            (N903)? data_o[639:608] : 
                            (N904)? data_o[607:576] : 
                            (N905)? data_o[575:544] : 
                            (N906)? data_o[543:512] : 
                            (N907)? data_o[511:480] : 1'b0;
  assign data_nn[543:512] = (N796)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N797)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N798)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N799)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N800)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N801)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N802)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N803)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N804)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N805)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N806)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N807)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N808)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N809)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N810)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N811)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N812)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N813)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N814)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N815)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N816)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N817)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N818)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N819)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N820)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N821)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N822)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N823)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N824)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N825)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N826)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N827)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N828)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N829)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N830)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N831)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N832)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N833)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N834)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N835)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N836)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N837)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N838)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N839)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N840)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N841)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N842)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N843)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N844)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N845)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N846)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N847)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N848)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N849)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N850)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N851)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N852)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N853)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N854)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N855)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N856)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N857)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N858)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N859)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N860)? data_o[2047:2016] : 
                            (N861)? data_o[2015:1984] : 
                            (N862)? data_o[1983:1952] : 
                            (N863)? data_o[1951:1920] : 
                            (N864)? data_o[1919:1888] : 
                            (N865)? data_o[1887:1856] : 
                            (N866)? data_o[1855:1824] : 
                            (N867)? data_o[1823:1792] : 
                            (N868)? data_o[1791:1760] : 
                            (N869)? data_o[1759:1728] : 
                            (N870)? data_o[1727:1696] : 
                            (N871)? data_o[1695:1664] : 
                            (N872)? data_o[1663:1632] : 
                            (N873)? data_o[1631:1600] : 
                            (N874)? data_o[1599:1568] : 
                            (N875)? data_o[1567:1536] : 
                            (N876)? data_o[1535:1504] : 
                            (N877)? data_o[1503:1472] : 
                            (N878)? data_o[1471:1440] : 
                            (N879)? data_o[1439:1408] : 
                            (N880)? data_o[1407:1376] : 
                            (N881)? data_o[1375:1344] : 
                            (N882)? data_o[1343:1312] : 
                            (N883)? data_o[1311:1280] : 
                            (N884)? data_o[1279:1248] : 
                            (N885)? data_o[1247:1216] : 
                            (N886)? data_o[1215:1184] : 
                            (N887)? data_o[1183:1152] : 
                            (N888)? data_o[1151:1120] : 
                            (N889)? data_o[1119:1088] : 
                            (N890)? data_o[1087:1056] : 
                            (N891)? data_o[1055:1024] : 
                            (N892)? data_o[1023:992] : 
                            (N893)? data_o[991:960] : 
                            (N894)? data_o[959:928] : 
                            (N895)? data_o[927:896] : 
                            (N896)? data_o[895:864] : 
                            (N897)? data_o[863:832] : 
                            (N898)? data_o[831:800] : 
                            (N899)? data_o[799:768] : 
                            (N900)? data_o[767:736] : 
                            (N901)? data_o[735:704] : 
                            (N902)? data_o[703:672] : 
                            (N903)? data_o[671:640] : 
                            (N904)? data_o[639:608] : 
                            (N905)? data_o[607:576] : 
                            (N906)? data_o[575:544] : 
                            (N907)? data_o[543:512] : 1'b0;
  assign data_nn[575:544] = (N797)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N798)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N799)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N800)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N801)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N802)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N803)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N804)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N805)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N806)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N807)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N808)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N809)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N810)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N811)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N812)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N813)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N814)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N815)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N816)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N817)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N818)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N819)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N820)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N821)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N822)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N823)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N824)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N825)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N826)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N827)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N828)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N829)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N830)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N831)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N832)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N833)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N834)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N835)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N836)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N837)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N838)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N839)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N840)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N841)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N842)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N843)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N844)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N845)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N846)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N847)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N848)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N849)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N850)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N851)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N852)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N853)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N854)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N855)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N856)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N857)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N858)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N859)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N860)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N861)? data_o[2047:2016] : 
                            (N862)? data_o[2015:1984] : 
                            (N863)? data_o[1983:1952] : 
                            (N864)? data_o[1951:1920] : 
                            (N865)? data_o[1919:1888] : 
                            (N866)? data_o[1887:1856] : 
                            (N867)? data_o[1855:1824] : 
                            (N868)? data_o[1823:1792] : 
                            (N869)? data_o[1791:1760] : 
                            (N870)? data_o[1759:1728] : 
                            (N871)? data_o[1727:1696] : 
                            (N872)? data_o[1695:1664] : 
                            (N873)? data_o[1663:1632] : 
                            (N874)? data_o[1631:1600] : 
                            (N875)? data_o[1599:1568] : 
                            (N876)? data_o[1567:1536] : 
                            (N877)? data_o[1535:1504] : 
                            (N878)? data_o[1503:1472] : 
                            (N879)? data_o[1471:1440] : 
                            (N880)? data_o[1439:1408] : 
                            (N881)? data_o[1407:1376] : 
                            (N882)? data_o[1375:1344] : 
                            (N883)? data_o[1343:1312] : 
                            (N884)? data_o[1311:1280] : 
                            (N885)? data_o[1279:1248] : 
                            (N886)? data_o[1247:1216] : 
                            (N887)? data_o[1215:1184] : 
                            (N888)? data_o[1183:1152] : 
                            (N889)? data_o[1151:1120] : 
                            (N890)? data_o[1119:1088] : 
                            (N891)? data_o[1087:1056] : 
                            (N892)? data_o[1055:1024] : 
                            (N893)? data_o[1023:992] : 
                            (N894)? data_o[991:960] : 
                            (N895)? data_o[959:928] : 
                            (N896)? data_o[927:896] : 
                            (N897)? data_o[895:864] : 
                            (N898)? data_o[863:832] : 
                            (N899)? data_o[831:800] : 
                            (N900)? data_o[799:768] : 
                            (N901)? data_o[767:736] : 
                            (N902)? data_o[735:704] : 
                            (N903)? data_o[703:672] : 
                            (N904)? data_o[671:640] : 
                            (N905)? data_o[639:608] : 
                            (N906)? data_o[607:576] : 
                            (N907)? data_o[575:544] : 1'b0;
  assign data_nn[607:576] = (N798)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N799)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N800)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N801)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N802)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N803)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N804)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N805)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N806)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N807)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N808)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N809)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N810)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N811)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N812)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N813)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N814)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N815)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N816)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N817)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N818)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N819)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N820)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N821)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N822)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N823)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N824)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N825)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N826)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N827)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N828)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N829)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N830)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N831)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N832)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N833)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N834)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N835)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N836)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N837)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N838)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N839)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N840)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N841)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N842)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N843)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N844)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N845)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N846)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N847)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N848)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N849)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N850)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N851)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N852)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N853)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N854)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N855)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N856)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N857)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N858)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N859)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N860)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N861)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N862)? data_o[2047:2016] : 
                            (N863)? data_o[2015:1984] : 
                            (N864)? data_o[1983:1952] : 
                            (N865)? data_o[1951:1920] : 
                            (N866)? data_o[1919:1888] : 
                            (N867)? data_o[1887:1856] : 
                            (N868)? data_o[1855:1824] : 
                            (N869)? data_o[1823:1792] : 
                            (N870)? data_o[1791:1760] : 
                            (N871)? data_o[1759:1728] : 
                            (N872)? data_o[1727:1696] : 
                            (N873)? data_o[1695:1664] : 
                            (N874)? data_o[1663:1632] : 
                            (N875)? data_o[1631:1600] : 
                            (N876)? data_o[1599:1568] : 
                            (N877)? data_o[1567:1536] : 
                            (N878)? data_o[1535:1504] : 
                            (N879)? data_o[1503:1472] : 
                            (N880)? data_o[1471:1440] : 
                            (N881)? data_o[1439:1408] : 
                            (N882)? data_o[1407:1376] : 
                            (N883)? data_o[1375:1344] : 
                            (N884)? data_o[1343:1312] : 
                            (N885)? data_o[1311:1280] : 
                            (N886)? data_o[1279:1248] : 
                            (N887)? data_o[1247:1216] : 
                            (N888)? data_o[1215:1184] : 
                            (N889)? data_o[1183:1152] : 
                            (N890)? data_o[1151:1120] : 
                            (N891)? data_o[1119:1088] : 
                            (N892)? data_o[1087:1056] : 
                            (N893)? data_o[1055:1024] : 
                            (N894)? data_o[1023:992] : 
                            (N895)? data_o[991:960] : 
                            (N896)? data_o[959:928] : 
                            (N897)? data_o[927:896] : 
                            (N898)? data_o[895:864] : 
                            (N899)? data_o[863:832] : 
                            (N900)? data_o[831:800] : 
                            (N901)? data_o[799:768] : 
                            (N902)? data_o[767:736] : 
                            (N903)? data_o[735:704] : 
                            (N904)? data_o[703:672] : 
                            (N905)? data_o[671:640] : 
                            (N906)? data_o[639:608] : 
                            (N907)? data_o[607:576] : 1'b0;
  assign data_nn[639:608] = (N908)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N909)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N910)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N911)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N912)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N913)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N914)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N915)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N916)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N917)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N918)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N919)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N920)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N921)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N922)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N923)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N924)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N925)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N926)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N927)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N928)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N929)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N930)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N931)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N932)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N933)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N934)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N935)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N936)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N937)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N938)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N939)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N940)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N941)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N942)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N943)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N944)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N945)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N946)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N947)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N948)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N949)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N950)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N951)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N952)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N953)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N954)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N955)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N956)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N957)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N958)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N959)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N960)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N961)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N962)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N963)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N964)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N965)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N966)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N967)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N968)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N969)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N970)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N971)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N972)? data_o[2047:2016] : 
                            (N973)? data_o[2015:1984] : 
                            (N974)? data_o[1983:1952] : 
                            (N975)? data_o[1951:1920] : 
                            (N976)? data_o[1919:1888] : 
                            (N977)? data_o[1887:1856] : 
                            (N978)? data_o[1855:1824] : 
                            (N979)? data_o[1823:1792] : 
                            (N980)? data_o[1791:1760] : 
                            (N981)? data_o[1759:1728] : 
                            (N982)? data_o[1727:1696] : 
                            (N983)? data_o[1695:1664] : 
                            (N984)? data_o[1663:1632] : 
                            (N985)? data_o[1631:1600] : 
                            (N986)? data_o[1599:1568] : 
                            (N987)? data_o[1567:1536] : 
                            (N988)? data_o[1535:1504] : 
                            (N989)? data_o[1503:1472] : 
                            (N990)? data_o[1471:1440] : 
                            (N991)? data_o[1439:1408] : 
                            (N992)? data_o[1407:1376] : 
                            (N993)? data_o[1375:1344] : 
                            (N994)? data_o[1343:1312] : 
                            (N995)? data_o[1311:1280] : 
                            (N996)? data_o[1279:1248] : 
                            (N997)? data_o[1247:1216] : 
                            (N998)? data_o[1215:1184] : 
                            (N999)? data_o[1183:1152] : 
                            (N1000)? data_o[1151:1120] : 
                            (N1001)? data_o[1119:1088] : 
                            (N1002)? data_o[1087:1056] : 
                            (N1003)? data_o[1055:1024] : 
                            (N1004)? data_o[1023:992] : 
                            (N1005)? data_o[991:960] : 
                            (N1006)? data_o[959:928] : 
                            (N1007)? data_o[927:896] : 
                            (N1008)? data_o[895:864] : 
                            (N1009)? data_o[863:832] : 
                            (N1010)? data_o[831:800] : 
                            (N1011)? data_o[799:768] : 
                            (N1012)? data_o[767:736] : 
                            (N1013)? data_o[735:704] : 
                            (N1014)? data_o[703:672] : 
                            (N1015)? data_o[671:640] : 
                            (N1016)? data_o[639:608] : 1'b0;
  assign N908 = N5538;
  assign N909 = N5539;
  assign N910 = N5540;
  assign N911 = N5541;
  assign N912 = N3626;
  assign N913 = N3625;
  assign N914 = N3624;
  assign N915 = N3623;
  assign N916 = N3622;
  assign N917 = N3621;
  assign N918 = N3620;
  assign N919 = N3619;
  assign N920 = N3618;
  assign N921 = N3617;
  assign N922 = N3616;
  assign N923 = N3615;
  assign N924 = N3614;
  assign N925 = N3613;
  assign N926 = N3612;
  assign N927 = N3611;
  assign N928 = N3610;
  assign N929 = N3609;
  assign N930 = N3608;
  assign N931 = N3607;
  assign N932 = N3606;
  assign N933 = N3605;
  assign N934 = N3604;
  assign N935 = N3603;
  assign N936 = N3602;
  assign N937 = N3601;
  assign N938 = N3600;
  assign N939 = N3599;
  assign N940 = N3598;
  assign N941 = N3597;
  assign N942 = N3596;
  assign N943 = N3595;
  assign N944 = N3594;
  assign N945 = N3593;
  assign N946 = N3592;
  assign N947 = N3591;
  assign N948 = N3590;
  assign N949 = N3589;
  assign N950 = N3588;
  assign N951 = N3587;
  assign N952 = N3586;
  assign N953 = N3585;
  assign N954 = N3584;
  assign N955 = N3583;
  assign N956 = N3582;
  assign N957 = N3581;
  assign N958 = N3580;
  assign N959 = N3579;
  assign N960 = N3578;
  assign N961 = N3577;
  assign N962 = N3576;
  assign N963 = N3575;
  assign N964 = N3574;
  assign N965 = N3573;
  assign N966 = N3572;
  assign N967 = N3571;
  assign N968 = N3570;
  assign N969 = N3569;
  assign N970 = N3568;
  assign N971 = N3567;
  assign N972 = N3566;
  assign N973 = N3565;
  assign N974 = N3564;
  assign N975 = N3563;
  assign N976 = N3562;
  assign N977 = N3561;
  assign N978 = N3560;
  assign N979 = N3559;
  assign N980 = N3558;
  assign N981 = N3557;
  assign N982 = N3556;
  assign N983 = N3555;
  assign N984 = N3554;
  assign N985 = N3553;
  assign N986 = N3552;
  assign N987 = N3551;
  assign N988 = N3550;
  assign N989 = N3549;
  assign N990 = N3548;
  assign N991 = N3547;
  assign N992 = N3546;
  assign N993 = N3545;
  assign N994 = N3544;
  assign N995 = N3543;
  assign N996 = N3542;
  assign N997 = N3541;
  assign N998 = N3540;
  assign N999 = N3539;
  assign N1000 = N3538;
  assign N1001 = N3537;
  assign N1002 = N3536;
  assign N1003 = N3535;
  assign N1004 = N3534;
  assign N1005 = N3533;
  assign N1006 = N3532;
  assign N1007 = N3531;
  assign N1008 = N3530;
  assign N1009 = N3529;
  assign N1010 = N3528;
  assign N1011 = N3527;
  assign N1012 = N3526;
  assign N1013 = N3525;
  assign N1014 = N3524;
  assign N1015 = N3523;
  assign N1016 = N3522;
  assign data_nn[671:640] = (N909)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N910)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N911)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N912)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N913)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N914)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N915)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N916)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N917)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N918)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N919)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N920)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N921)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N922)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N923)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N924)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N925)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N926)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N927)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N928)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N929)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N930)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N931)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N932)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N933)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N934)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N935)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N936)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N937)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N938)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N939)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N940)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N941)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N942)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N943)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N944)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N945)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N946)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N947)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N948)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N949)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N950)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N951)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N952)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N953)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N954)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N955)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N956)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N957)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N958)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N959)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N960)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N961)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N962)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N963)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N964)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N965)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N966)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N967)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N968)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N969)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N970)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N971)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N972)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N973)? data_o[2047:2016] : 
                            (N974)? data_o[2015:1984] : 
                            (N975)? data_o[1983:1952] : 
                            (N976)? data_o[1951:1920] : 
                            (N977)? data_o[1919:1888] : 
                            (N978)? data_o[1887:1856] : 
                            (N979)? data_o[1855:1824] : 
                            (N980)? data_o[1823:1792] : 
                            (N981)? data_o[1791:1760] : 
                            (N982)? data_o[1759:1728] : 
                            (N983)? data_o[1727:1696] : 
                            (N984)? data_o[1695:1664] : 
                            (N985)? data_o[1663:1632] : 
                            (N986)? data_o[1631:1600] : 
                            (N987)? data_o[1599:1568] : 
                            (N988)? data_o[1567:1536] : 
                            (N989)? data_o[1535:1504] : 
                            (N990)? data_o[1503:1472] : 
                            (N991)? data_o[1471:1440] : 
                            (N992)? data_o[1439:1408] : 
                            (N993)? data_o[1407:1376] : 
                            (N994)? data_o[1375:1344] : 
                            (N995)? data_o[1343:1312] : 
                            (N996)? data_o[1311:1280] : 
                            (N997)? data_o[1279:1248] : 
                            (N998)? data_o[1247:1216] : 
                            (N999)? data_o[1215:1184] : 
                            (N1000)? data_o[1183:1152] : 
                            (N1001)? data_o[1151:1120] : 
                            (N1002)? data_o[1119:1088] : 
                            (N1003)? data_o[1087:1056] : 
                            (N1004)? data_o[1055:1024] : 
                            (N1005)? data_o[1023:992] : 
                            (N1006)? data_o[991:960] : 
                            (N1007)? data_o[959:928] : 
                            (N1008)? data_o[927:896] : 
                            (N1009)? data_o[895:864] : 
                            (N1010)? data_o[863:832] : 
                            (N1011)? data_o[831:800] : 
                            (N1012)? data_o[799:768] : 
                            (N1013)? data_o[767:736] : 
                            (N1014)? data_o[735:704] : 
                            (N1015)? data_o[703:672] : 
                            (N1016)? data_o[671:640] : 1'b0;
  assign data_nn[703:672] = (N910)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N911)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N912)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N913)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N914)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N915)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N916)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N917)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N918)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N919)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N920)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N921)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N922)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N923)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N924)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N925)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N926)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N927)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N928)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N929)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N930)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N931)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N932)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N933)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N934)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N935)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N936)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N937)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N938)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N939)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N940)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N941)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N942)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N943)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N944)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N945)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N946)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N947)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N948)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N949)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N950)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N951)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N952)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N953)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N954)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N955)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N956)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N957)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N958)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N959)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N960)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N961)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N962)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N963)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N964)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N965)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N966)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N967)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N968)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N969)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N970)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N971)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N972)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N973)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N974)? data_o[2047:2016] : 
                            (N975)? data_o[2015:1984] : 
                            (N976)? data_o[1983:1952] : 
                            (N977)? data_o[1951:1920] : 
                            (N978)? data_o[1919:1888] : 
                            (N979)? data_o[1887:1856] : 
                            (N980)? data_o[1855:1824] : 
                            (N981)? data_o[1823:1792] : 
                            (N982)? data_o[1791:1760] : 
                            (N983)? data_o[1759:1728] : 
                            (N984)? data_o[1727:1696] : 
                            (N985)? data_o[1695:1664] : 
                            (N986)? data_o[1663:1632] : 
                            (N987)? data_o[1631:1600] : 
                            (N988)? data_o[1599:1568] : 
                            (N989)? data_o[1567:1536] : 
                            (N990)? data_o[1535:1504] : 
                            (N991)? data_o[1503:1472] : 
                            (N992)? data_o[1471:1440] : 
                            (N993)? data_o[1439:1408] : 
                            (N994)? data_o[1407:1376] : 
                            (N995)? data_o[1375:1344] : 
                            (N996)? data_o[1343:1312] : 
                            (N997)? data_o[1311:1280] : 
                            (N998)? data_o[1279:1248] : 
                            (N999)? data_o[1247:1216] : 
                            (N1000)? data_o[1215:1184] : 
                            (N1001)? data_o[1183:1152] : 
                            (N1002)? data_o[1151:1120] : 
                            (N1003)? data_o[1119:1088] : 
                            (N1004)? data_o[1087:1056] : 
                            (N1005)? data_o[1055:1024] : 
                            (N1006)? data_o[1023:992] : 
                            (N1007)? data_o[991:960] : 
                            (N1008)? data_o[959:928] : 
                            (N1009)? data_o[927:896] : 
                            (N1010)? data_o[895:864] : 
                            (N1011)? data_o[863:832] : 
                            (N1012)? data_o[831:800] : 
                            (N1013)? data_o[799:768] : 
                            (N1014)? data_o[767:736] : 
                            (N1015)? data_o[735:704] : 
                            (N1016)? data_o[703:672] : 1'b0;
  assign data_nn[735:704] = (N911)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N912)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N913)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N914)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N915)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N916)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N917)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N918)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N919)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N920)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N921)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N922)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N923)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N924)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N925)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N926)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N927)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N928)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N929)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N930)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N931)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N932)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N933)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N934)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N935)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N936)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N937)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N938)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N939)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N940)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N941)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N942)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N943)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N944)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N945)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N946)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N947)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N948)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N949)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N950)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N951)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N952)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N953)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N954)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N955)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N956)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N957)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N958)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N959)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N960)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N961)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N962)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N963)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N964)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N965)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N966)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N967)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N968)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N969)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N970)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N971)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N972)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N973)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N974)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N975)? data_o[2047:2016] : 
                            (N976)? data_o[2015:1984] : 
                            (N977)? data_o[1983:1952] : 
                            (N978)? data_o[1951:1920] : 
                            (N979)? data_o[1919:1888] : 
                            (N980)? data_o[1887:1856] : 
                            (N981)? data_o[1855:1824] : 
                            (N982)? data_o[1823:1792] : 
                            (N983)? data_o[1791:1760] : 
                            (N984)? data_o[1759:1728] : 
                            (N985)? data_o[1727:1696] : 
                            (N986)? data_o[1695:1664] : 
                            (N987)? data_o[1663:1632] : 
                            (N988)? data_o[1631:1600] : 
                            (N989)? data_o[1599:1568] : 
                            (N990)? data_o[1567:1536] : 
                            (N991)? data_o[1535:1504] : 
                            (N992)? data_o[1503:1472] : 
                            (N993)? data_o[1471:1440] : 
                            (N994)? data_o[1439:1408] : 
                            (N995)? data_o[1407:1376] : 
                            (N996)? data_o[1375:1344] : 
                            (N997)? data_o[1343:1312] : 
                            (N998)? data_o[1311:1280] : 
                            (N999)? data_o[1279:1248] : 
                            (N1000)? data_o[1247:1216] : 
                            (N1001)? data_o[1215:1184] : 
                            (N1002)? data_o[1183:1152] : 
                            (N1003)? data_o[1151:1120] : 
                            (N1004)? data_o[1119:1088] : 
                            (N1005)? data_o[1087:1056] : 
                            (N1006)? data_o[1055:1024] : 
                            (N1007)? data_o[1023:992] : 
                            (N1008)? data_o[991:960] : 
                            (N1009)? data_o[959:928] : 
                            (N1010)? data_o[927:896] : 
                            (N1011)? data_o[895:864] : 
                            (N1012)? data_o[863:832] : 
                            (N1013)? data_o[831:800] : 
                            (N1014)? data_o[799:768] : 
                            (N1015)? data_o[767:736] : 
                            (N1016)? data_o[735:704] : 1'b0;
  assign data_nn[767:736] = (N912)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N913)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N914)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N915)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N916)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N917)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N918)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N919)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N920)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N921)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N922)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N923)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N924)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N925)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N926)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N927)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N928)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N929)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N930)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N931)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N932)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N933)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N934)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N935)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N936)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N937)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N938)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N939)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N940)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N941)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N942)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N943)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N944)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N945)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N946)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N947)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N948)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N949)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N950)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N951)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N952)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N953)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N954)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N955)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N956)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N957)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N958)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N959)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N960)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N961)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N962)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N963)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N964)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N965)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N966)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N967)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N968)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N969)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N970)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N971)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N972)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N973)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N974)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N975)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N976)? data_o[2047:2016] : 
                            (N977)? data_o[2015:1984] : 
                            (N978)? data_o[1983:1952] : 
                            (N979)? data_o[1951:1920] : 
                            (N980)? data_o[1919:1888] : 
                            (N981)? data_o[1887:1856] : 
                            (N982)? data_o[1855:1824] : 
                            (N983)? data_o[1823:1792] : 
                            (N984)? data_o[1791:1760] : 
                            (N985)? data_o[1759:1728] : 
                            (N986)? data_o[1727:1696] : 
                            (N987)? data_o[1695:1664] : 
                            (N988)? data_o[1663:1632] : 
                            (N989)? data_o[1631:1600] : 
                            (N990)? data_o[1599:1568] : 
                            (N991)? data_o[1567:1536] : 
                            (N992)? data_o[1535:1504] : 
                            (N993)? data_o[1503:1472] : 
                            (N994)? data_o[1471:1440] : 
                            (N995)? data_o[1439:1408] : 
                            (N996)? data_o[1407:1376] : 
                            (N997)? data_o[1375:1344] : 
                            (N998)? data_o[1343:1312] : 
                            (N999)? data_o[1311:1280] : 
                            (N1000)? data_o[1279:1248] : 
                            (N1001)? data_o[1247:1216] : 
                            (N1002)? data_o[1215:1184] : 
                            (N1003)? data_o[1183:1152] : 
                            (N1004)? data_o[1151:1120] : 
                            (N1005)? data_o[1119:1088] : 
                            (N1006)? data_o[1087:1056] : 
                            (N1007)? data_o[1055:1024] : 
                            (N1008)? data_o[1023:992] : 
                            (N1009)? data_o[991:960] : 
                            (N1010)? data_o[959:928] : 
                            (N1011)? data_o[927:896] : 
                            (N1012)? data_o[895:864] : 
                            (N1013)? data_o[863:832] : 
                            (N1014)? data_o[831:800] : 
                            (N1015)? data_o[799:768] : 
                            (N1016)? data_o[767:736] : 1'b0;
  assign data_nn[799:768] = (N1017)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N1018)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N1019)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N1020)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N1021)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N1022)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N1023)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N1024)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N1025)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N1026)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N1027)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N1028)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N1029)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N1030)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N1031)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N1032)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N1033)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N1034)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N1035)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N1036)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N1037)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N1038)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N1039)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N1040)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N1041)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N1042)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N1043)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N1044)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N1045)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N1046)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N1047)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N1048)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N1049)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N1050)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N1051)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N1052)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N1053)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N1054)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N1055)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N1056)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N1057)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N1058)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N1059)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N1060)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N1061)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N1062)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N1063)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N1064)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N1065)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N1066)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N1067)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N1068)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N1069)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N1070)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N1071)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N1072)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N1073)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N1074)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N1075)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N1076)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N1077)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N1078)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N1079)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N1080)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N1081)? data_o[2047:2016] : 
                            (N1082)? data_o[2015:1984] : 
                            (N1083)? data_o[1983:1952] : 
                            (N1084)? data_o[1951:1920] : 
                            (N1085)? data_o[1919:1888] : 
                            (N1086)? data_o[1887:1856] : 
                            (N1087)? data_o[1855:1824] : 
                            (N1088)? data_o[1823:1792] : 
                            (N1089)? data_o[1791:1760] : 
                            (N1090)? data_o[1759:1728] : 
                            (N1091)? data_o[1727:1696] : 
                            (N1092)? data_o[1695:1664] : 
                            (N1093)? data_o[1663:1632] : 
                            (N1094)? data_o[1631:1600] : 
                            (N1095)? data_o[1599:1568] : 
                            (N1096)? data_o[1567:1536] : 
                            (N1097)? data_o[1535:1504] : 
                            (N1098)? data_o[1503:1472] : 
                            (N1099)? data_o[1471:1440] : 
                            (N1100)? data_o[1439:1408] : 
                            (N1101)? data_o[1407:1376] : 
                            (N1102)? data_o[1375:1344] : 
                            (N1103)? data_o[1343:1312] : 
                            (N1104)? data_o[1311:1280] : 
                            (N1105)? data_o[1279:1248] : 
                            (N1106)? data_o[1247:1216] : 
                            (N1107)? data_o[1215:1184] : 
                            (N1108)? data_o[1183:1152] : 
                            (N1109)? data_o[1151:1120] : 
                            (N1110)? data_o[1119:1088] : 
                            (N1111)? data_o[1087:1056] : 
                            (N1112)? data_o[1055:1024] : 
                            (N1113)? data_o[1023:992] : 
                            (N1114)? data_o[991:960] : 
                            (N1115)? data_o[959:928] : 
                            (N1116)? data_o[927:896] : 
                            (N1117)? data_o[895:864] : 
                            (N1118)? data_o[863:832] : 
                            (N1119)? data_o[831:800] : 
                            (N1120)? data_o[799:768] : 1'b0;
  assign N1017 = N3730;
  assign N1018 = N3729;
  assign N1019 = N3728;
  assign N1020 = N3727;
  assign N1021 = N3726;
  assign N1022 = N3725;
  assign N1023 = N3724;
  assign N1024 = N3723;
  assign N1025 = N3722;
  assign N1026 = N3721;
  assign N1027 = N3720;
  assign N1028 = N3719;
  assign N1029 = N3718;
  assign N1030 = N3717;
  assign N1031 = N3716;
  assign N1032 = N3715;
  assign N1033 = N3714;
  assign N1034 = N3713;
  assign N1035 = N3712;
  assign N1036 = N3711;
  assign N1037 = N3710;
  assign N1038 = N3709;
  assign N1039 = N3708;
  assign N1040 = N3707;
  assign N1041 = N3706;
  assign N1042 = N3705;
  assign N1043 = N3704;
  assign N1044 = N3703;
  assign N1045 = N3702;
  assign N1046 = N3701;
  assign N1047 = N3700;
  assign N1048 = N3699;
  assign N1049 = N3698;
  assign N1050 = N3697;
  assign N1051 = N3696;
  assign N1052 = N3695;
  assign N1053 = N3694;
  assign N1054 = N3693;
  assign N1055 = N3692;
  assign N1056 = N3691;
  assign N1057 = N3690;
  assign N1058 = N3689;
  assign N1059 = N3688;
  assign N1060 = N3687;
  assign N1061 = N3686;
  assign N1062 = N3685;
  assign N1063 = N3684;
  assign N1064 = N3683;
  assign N1065 = N3682;
  assign N1066 = N3681;
  assign N1067 = N3680;
  assign N1068 = N3679;
  assign N1069 = N3678;
  assign N1070 = N3677;
  assign N1071 = N3676;
  assign N1072 = N3675;
  assign N1073 = N3674;
  assign N1074 = N3673;
  assign N1075 = N3672;
  assign N1076 = N3671;
  assign N1077 = N3670;
  assign N1078 = N3669;
  assign N1079 = N3668;
  assign N1080 = N3667;
  assign N1081 = N3666;
  assign N1082 = N3665;
  assign N1083 = N3664;
  assign N1084 = N3663;
  assign N1085 = N3662;
  assign N1086 = N3661;
  assign N1087 = N3660;
  assign N1088 = N3659;
  assign N1089 = N3658;
  assign N1090 = N3657;
  assign N1091 = N3656;
  assign N1092 = N3655;
  assign N1093 = N3654;
  assign N1094 = N3653;
  assign N1095 = N3652;
  assign N1096 = N3651;
  assign N1097 = N3650;
  assign N1098 = N3649;
  assign N1099 = N3648;
  assign N1100 = N3647;
  assign N1101 = N3646;
  assign N1102 = N3645;
  assign N1103 = N3644;
  assign N1104 = N3643;
  assign N1105 = N3642;
  assign N1106 = N3641;
  assign N1107 = N3640;
  assign N1108 = N3639;
  assign N1109 = N3638;
  assign N1110 = N3637;
  assign N1111 = N3636;
  assign N1112 = N3635;
  assign N1113 = N3634;
  assign N1114 = N3633;
  assign N1115 = N3632;
  assign N1116 = N3631;
  assign N1117 = N3630;
  assign N1118 = N3629;
  assign N1119 = N3628;
  assign N1120 = N3627;
  assign data_nn[831:800] = (N1121)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N1122)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N1123)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N1124)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N1125)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N1126)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N1127)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N1128)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N1129)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N1130)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N1131)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N1132)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N1133)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N1134)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N1135)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N1136)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N1137)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N1138)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N1139)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N1140)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N1141)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N1142)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N1143)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N1144)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N1145)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N1146)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N1147)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N1148)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N1149)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N1150)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N1151)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N1152)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N1153)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N1154)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N1155)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N1156)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N1157)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N1158)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N1159)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N1160)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N1161)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N1162)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N1163)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N1164)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N1165)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N1166)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N1167)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N1168)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N1169)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N1170)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N1171)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N1172)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N1173)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N1174)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N1175)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N1176)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N1177)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N1178)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N1179)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N1180)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N1181)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N1182)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N1183)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N1184)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N1185)? data_o[2047:2016] : 
                            (N1186)? data_o[2015:1984] : 
                            (N1187)? data_o[1983:1952] : 
                            (N1188)? data_o[1951:1920] : 
                            (N1189)? data_o[1919:1888] : 
                            (N1190)? data_o[1887:1856] : 
                            (N1191)? data_o[1855:1824] : 
                            (N1192)? data_o[1823:1792] : 
                            (N1193)? data_o[1791:1760] : 
                            (N1194)? data_o[1759:1728] : 
                            (N1195)? data_o[1727:1696] : 
                            (N1196)? data_o[1695:1664] : 
                            (N1197)? data_o[1663:1632] : 
                            (N1198)? data_o[1631:1600] : 
                            (N1199)? data_o[1599:1568] : 
                            (N1200)? data_o[1567:1536] : 
                            (N1201)? data_o[1535:1504] : 
                            (N1202)? data_o[1503:1472] : 
                            (N1203)? data_o[1471:1440] : 
                            (N1204)? data_o[1439:1408] : 
                            (N1205)? data_o[1407:1376] : 
                            (N1206)? data_o[1375:1344] : 
                            (N1207)? data_o[1343:1312] : 
                            (N1208)? data_o[1311:1280] : 
                            (N1209)? data_o[1279:1248] : 
                            (N1210)? data_o[1247:1216] : 
                            (N1211)? data_o[1215:1184] : 
                            (N1212)? data_o[1183:1152] : 
                            (N1213)? data_o[1151:1120] : 
                            (N1214)? data_o[1119:1088] : 
                            (N1215)? data_o[1087:1056] : 
                            (N1216)? data_o[1055:1024] : 
                            (N1217)? data_o[1023:992] : 
                            (N1218)? data_o[991:960] : 
                            (N1219)? data_o[959:928] : 
                            (N1220)? data_o[927:896] : 
                            (N1221)? data_o[895:864] : 
                            (N1222)? data_o[863:832] : 
                            (N1223)? data_o[831:800] : 1'b0;
  assign N1121 = N5542;
  assign N1122 = N5543;
  assign N1123 = N5544;
  assign N1124 = N3830;
  assign N1125 = N3829;
  assign N1126 = N3828;
  assign N1127 = N3827;
  assign N1128 = N3826;
  assign N1129 = N3825;
  assign N1130 = N3824;
  assign N1131 = N3823;
  assign N1132 = N3822;
  assign N1133 = N3821;
  assign N1134 = N3820;
  assign N1135 = N3819;
  assign N1136 = N3818;
  assign N1137 = N3817;
  assign N1138 = N3816;
  assign N1139 = N3815;
  assign N1140 = N3814;
  assign N1141 = N3813;
  assign N1142 = N3812;
  assign N1143 = N3811;
  assign N1144 = N3810;
  assign N1145 = N3809;
  assign N1146 = N3808;
  assign N1147 = N3807;
  assign N1148 = N3806;
  assign N1149 = N3805;
  assign N1150 = N3804;
  assign N1151 = N3803;
  assign N1152 = N3802;
  assign N1153 = N3801;
  assign N1154 = N3800;
  assign N1155 = N3799;
  assign N1156 = N3798;
  assign N1157 = N3797;
  assign N1158 = N3796;
  assign N1159 = N3795;
  assign N1160 = N3794;
  assign N1161 = N3793;
  assign N1162 = N3792;
  assign N1163 = N3791;
  assign N1164 = N3790;
  assign N1165 = N3789;
  assign N1166 = N3788;
  assign N1167 = N3787;
  assign N1168 = N3786;
  assign N1169 = N3785;
  assign N1170 = N3784;
  assign N1171 = N3783;
  assign N1172 = N3782;
  assign N1173 = N3781;
  assign N1174 = N3780;
  assign N1175 = N3779;
  assign N1176 = N3778;
  assign N1177 = N3777;
  assign N1178 = N3776;
  assign N1179 = N3775;
  assign N1180 = N3774;
  assign N1181 = N3773;
  assign N1182 = N3772;
  assign N1183 = N3771;
  assign N1184 = N3770;
  assign N1185 = N3769;
  assign N1186 = N3768;
  assign N1187 = N3767;
  assign N1188 = N3766;
  assign N1189 = N3765;
  assign N1190 = N3764;
  assign N1191 = N3763;
  assign N1192 = N3762;
  assign N1193 = N3761;
  assign N1194 = N3760;
  assign N1195 = N3759;
  assign N1196 = N3758;
  assign N1197 = N3757;
  assign N1198 = N3756;
  assign N1199 = N3755;
  assign N1200 = N3754;
  assign N1201 = N3753;
  assign N1202 = N3752;
  assign N1203 = N3751;
  assign N1204 = N3750;
  assign N1205 = N3749;
  assign N1206 = N3748;
  assign N1207 = N3747;
  assign N1208 = N3746;
  assign N1209 = N3745;
  assign N1210 = N3744;
  assign N1211 = N3743;
  assign N1212 = N3742;
  assign N1213 = N3741;
  assign N1214 = N3740;
  assign N1215 = N3739;
  assign N1216 = N3738;
  assign N1217 = N3737;
  assign N1218 = N3736;
  assign N1219 = N3735;
  assign N1220 = N3734;
  assign N1221 = N3733;
  assign N1222 = N3732;
  assign N1223 = N3731;
  assign data_nn[863:832] = (N1122)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N1123)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N1124)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N1125)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N1126)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N1127)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N1128)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N1129)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N1130)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N1131)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N1132)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N1133)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N1134)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N1135)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N1136)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N1137)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N1138)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N1139)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N1140)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N1141)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N1142)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N1143)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N1144)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N1145)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N1146)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N1147)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N1148)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N1149)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N1150)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N1151)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N1152)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N1153)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N1154)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N1155)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N1156)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N1157)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N1158)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N1159)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N1160)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N1161)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N1162)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N1163)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N1164)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N1165)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N1166)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N1167)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N1168)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N1169)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N1170)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N1171)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N1172)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N1173)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N1174)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N1175)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N1176)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N1177)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N1178)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N1179)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N1180)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N1181)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N1182)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N1183)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N1184)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N1185)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N1186)? data_o[2047:2016] : 
                            (N1187)? data_o[2015:1984] : 
                            (N1188)? data_o[1983:1952] : 
                            (N1189)? data_o[1951:1920] : 
                            (N1190)? data_o[1919:1888] : 
                            (N1191)? data_o[1887:1856] : 
                            (N1192)? data_o[1855:1824] : 
                            (N1193)? data_o[1823:1792] : 
                            (N1194)? data_o[1791:1760] : 
                            (N1195)? data_o[1759:1728] : 
                            (N1196)? data_o[1727:1696] : 
                            (N1197)? data_o[1695:1664] : 
                            (N1198)? data_o[1663:1632] : 
                            (N1199)? data_o[1631:1600] : 
                            (N1200)? data_o[1599:1568] : 
                            (N1201)? data_o[1567:1536] : 
                            (N1202)? data_o[1535:1504] : 
                            (N1203)? data_o[1503:1472] : 
                            (N1204)? data_o[1471:1440] : 
                            (N1205)? data_o[1439:1408] : 
                            (N1206)? data_o[1407:1376] : 
                            (N1207)? data_o[1375:1344] : 
                            (N1208)? data_o[1343:1312] : 
                            (N1209)? data_o[1311:1280] : 
                            (N1210)? data_o[1279:1248] : 
                            (N1211)? data_o[1247:1216] : 
                            (N1212)? data_o[1215:1184] : 
                            (N1213)? data_o[1183:1152] : 
                            (N1214)? data_o[1151:1120] : 
                            (N1215)? data_o[1119:1088] : 
                            (N1216)? data_o[1087:1056] : 
                            (N1217)? data_o[1055:1024] : 
                            (N1218)? data_o[1023:992] : 
                            (N1219)? data_o[991:960] : 
                            (N1220)? data_o[959:928] : 
                            (N1221)? data_o[927:896] : 
                            (N1222)? data_o[895:864] : 
                            (N1223)? data_o[863:832] : 1'b0;
  assign data_nn[895:864] = (N1123)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N1124)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N1125)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N1126)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N1127)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N1128)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N1129)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N1130)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N1131)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N1132)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N1133)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N1134)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N1135)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N1136)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N1137)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N1138)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N1139)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N1140)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N1141)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N1142)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N1143)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N1144)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N1145)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N1146)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N1147)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N1148)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N1149)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N1150)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N1151)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N1152)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N1153)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N1154)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N1155)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N1156)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N1157)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N1158)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N1159)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N1160)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N1161)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N1162)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N1163)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N1164)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N1165)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N1166)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N1167)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N1168)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N1169)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N1170)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N1171)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N1172)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N1173)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N1174)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N1175)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N1176)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N1177)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N1178)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N1179)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N1180)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N1181)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N1182)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N1183)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N1184)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N1185)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N1186)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N1187)? data_o[2047:2016] : 
                            (N1188)? data_o[2015:1984] : 
                            (N1189)? data_o[1983:1952] : 
                            (N1190)? data_o[1951:1920] : 
                            (N1191)? data_o[1919:1888] : 
                            (N1192)? data_o[1887:1856] : 
                            (N1193)? data_o[1855:1824] : 
                            (N1194)? data_o[1823:1792] : 
                            (N1195)? data_o[1791:1760] : 
                            (N1196)? data_o[1759:1728] : 
                            (N1197)? data_o[1727:1696] : 
                            (N1198)? data_o[1695:1664] : 
                            (N1199)? data_o[1663:1632] : 
                            (N1200)? data_o[1631:1600] : 
                            (N1201)? data_o[1599:1568] : 
                            (N1202)? data_o[1567:1536] : 
                            (N1203)? data_o[1535:1504] : 
                            (N1204)? data_o[1503:1472] : 
                            (N1205)? data_o[1471:1440] : 
                            (N1206)? data_o[1439:1408] : 
                            (N1207)? data_o[1407:1376] : 
                            (N1208)? data_o[1375:1344] : 
                            (N1209)? data_o[1343:1312] : 
                            (N1210)? data_o[1311:1280] : 
                            (N1211)? data_o[1279:1248] : 
                            (N1212)? data_o[1247:1216] : 
                            (N1213)? data_o[1215:1184] : 
                            (N1214)? data_o[1183:1152] : 
                            (N1215)? data_o[1151:1120] : 
                            (N1216)? data_o[1119:1088] : 
                            (N1217)? data_o[1087:1056] : 
                            (N1218)? data_o[1055:1024] : 
                            (N1219)? data_o[1023:992] : 
                            (N1220)? data_o[991:960] : 
                            (N1221)? data_o[959:928] : 
                            (N1222)? data_o[927:896] : 
                            (N1223)? data_o[895:864] : 1'b0;
  assign data_nn[927:896] = (N1124)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N1125)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N1126)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N1127)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N1128)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N1129)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N1130)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N1131)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N1132)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N1133)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N1134)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N1135)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N1136)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N1137)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N1138)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N1139)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N1140)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N1141)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N1142)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N1143)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N1144)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N1145)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N1146)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N1147)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N1148)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N1149)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N1150)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N1151)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N1152)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N1153)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N1154)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N1155)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N1156)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N1157)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N1158)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N1159)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N1160)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N1161)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N1162)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N1163)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N1164)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N1165)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N1166)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N1167)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N1168)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N1169)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N1170)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N1171)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N1172)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N1173)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N1174)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N1175)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N1176)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N1177)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N1178)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N1179)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N1180)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N1181)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N1182)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N1183)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N1184)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N1185)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N1186)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N1187)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N1188)? data_o[2047:2016] : 
                            (N1189)? data_o[2015:1984] : 
                            (N1190)? data_o[1983:1952] : 
                            (N1191)? data_o[1951:1920] : 
                            (N1192)? data_o[1919:1888] : 
                            (N1193)? data_o[1887:1856] : 
                            (N1194)? data_o[1855:1824] : 
                            (N1195)? data_o[1823:1792] : 
                            (N1196)? data_o[1791:1760] : 
                            (N1197)? data_o[1759:1728] : 
                            (N1198)? data_o[1727:1696] : 
                            (N1199)? data_o[1695:1664] : 
                            (N1200)? data_o[1663:1632] : 
                            (N1201)? data_o[1631:1600] : 
                            (N1202)? data_o[1599:1568] : 
                            (N1203)? data_o[1567:1536] : 
                            (N1204)? data_o[1535:1504] : 
                            (N1205)? data_o[1503:1472] : 
                            (N1206)? data_o[1471:1440] : 
                            (N1207)? data_o[1439:1408] : 
                            (N1208)? data_o[1407:1376] : 
                            (N1209)? data_o[1375:1344] : 
                            (N1210)? data_o[1343:1312] : 
                            (N1211)? data_o[1311:1280] : 
                            (N1212)? data_o[1279:1248] : 
                            (N1213)? data_o[1247:1216] : 
                            (N1214)? data_o[1215:1184] : 
                            (N1215)? data_o[1183:1152] : 
                            (N1216)? data_o[1151:1120] : 
                            (N1217)? data_o[1119:1088] : 
                            (N1218)? data_o[1087:1056] : 
                            (N1219)? data_o[1055:1024] : 
                            (N1220)? data_o[1023:992] : 
                            (N1221)? data_o[991:960] : 
                            (N1222)? data_o[959:928] : 
                            (N1223)? data_o[927:896] : 1'b0;
  assign data_nn[959:928] = (N1224)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N1225)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N1226)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N1227)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N1228)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N1229)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N1230)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N1231)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N1232)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N1233)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N1234)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N1235)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N1236)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N1237)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N1238)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N1239)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N1240)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N1241)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N1242)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N1243)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N1244)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N1245)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N1246)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N1247)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N1248)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N1249)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N1250)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N1251)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N1252)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N1253)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N1254)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N1255)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N1256)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N1257)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N1258)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N1259)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N1260)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N1261)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N1262)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N1263)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N1264)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N1265)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N1266)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N1267)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N1268)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N1269)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N1270)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N1271)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N1272)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N1273)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N1274)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N1275)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N1276)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N1277)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N1278)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N1279)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N1280)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N1281)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N1282)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N1283)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N1284)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N1285)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N1286)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N1287)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N1288)? data_o[2047:2016] : 
                            (N1289)? data_o[2015:1984] : 
                            (N1290)? data_o[1983:1952] : 
                            (N1291)? data_o[1951:1920] : 
                            (N1292)? data_o[1919:1888] : 
                            (N1293)? data_o[1887:1856] : 
                            (N1294)? data_o[1855:1824] : 
                            (N1295)? data_o[1823:1792] : 
                            (N1296)? data_o[1791:1760] : 
                            (N1297)? data_o[1759:1728] : 
                            (N1298)? data_o[1727:1696] : 
                            (N1299)? data_o[1695:1664] : 
                            (N1300)? data_o[1663:1632] : 
                            (N1301)? data_o[1631:1600] : 
                            (N1302)? data_o[1599:1568] : 
                            (N1303)? data_o[1567:1536] : 
                            (N1304)? data_o[1535:1504] : 
                            (N1305)? data_o[1503:1472] : 
                            (N1306)? data_o[1471:1440] : 
                            (N1307)? data_o[1439:1408] : 
                            (N1308)? data_o[1407:1376] : 
                            (N1309)? data_o[1375:1344] : 
                            (N1310)? data_o[1343:1312] : 
                            (N1311)? data_o[1311:1280] : 
                            (N1312)? data_o[1279:1248] : 
                            (N1313)? data_o[1247:1216] : 
                            (N1314)? data_o[1215:1184] : 
                            (N1315)? data_o[1183:1152] : 
                            (N1316)? data_o[1151:1120] : 
                            (N1317)? data_o[1119:1088] : 
                            (N1318)? data_o[1087:1056] : 
                            (N1319)? data_o[1055:1024] : 
                            (N1320)? data_o[1023:992] : 
                            (N1321)? data_o[991:960] : 
                            (N1322)? data_o[959:928] : 1'b0;
  assign N1224 = N5545;
  assign N1225 = N5546;
  assign N1226 = N5547;
  assign N1227 = N5548;
  assign N1228 = N3861;
  assign N1229 = N3860;
  assign N1230 = N3859;
  assign N1231 = N3858;
  assign N1232 = N3857;
  assign N1233 = N3856;
  assign N1234 = N3855;
  assign N1235 = N3854;
  assign N1236 = N3853;
  assign N1237 = N3852;
  assign N1238 = N3851;
  assign N1239 = N3850;
  assign N1240 = N3849;
  assign N1241 = N3848;
  assign N1242 = N3847;
  assign N1243 = N3846;
  assign N1244 = N3845;
  assign N1245 = N3844;
  assign N1246 = N3843;
  assign N1247 = N3842;
  assign N1248 = N3841;
  assign N1249 = N3840;
  assign N1250 = N3839;
  assign N1251 = N3838;
  assign N1252 = N3837;
  assign N1253 = N3836;
  assign N1254 = N3835;
  assign N1255 = N3834;
  assign N1256 = N3833;
  assign N1257 = N3832;
  assign N1258 = N3831;
  assign N1259 = N3989;
  assign N1260 = N3988;
  assign N1261 = N3987;
  assign N1262 = N3986;
  assign N1263 = N3985;
  assign N1264 = N3984;
  assign N1265 = N3983;
  assign N1266 = N3982;
  assign N1267 = N3981;
  assign N1268 = N3980;
  assign N1269 = N3979;
  assign N1270 = N3978;
  assign N1271 = N3977;
  assign N1272 = N3976;
  assign N1273 = N3975;
  assign N1274 = N3974;
  assign N1275 = N3973;
  assign N1276 = N3972;
  assign N1277 = N3971;
  assign N1278 = N3970;
  assign N1279 = N3969;
  assign N1280 = N3968;
  assign N1281 = N3967;
  assign N1282 = N3966;
  assign N1283 = N3965;
  assign N1284 = N3964;
  assign N1285 = N3963;
  assign N1286 = N3962;
  assign N1287 = N3961;
  assign N1288 = N3960;
  assign N1289 = N3959;
  assign N1290 = N3958;
  assign N1291 = N3957;
  assign N1292 = N3956;
  assign N1293 = N3955;
  assign N1294 = N3954;
  assign N1295 = N3953;
  assign N1296 = N3952;
  assign N1297 = N3951;
  assign N1298 = N3950;
  assign N1299 = N3949;
  assign N1300 = N3948;
  assign N1301 = N3947;
  assign N1302 = N3946;
  assign N1303 = N3945;
  assign N1304 = N3944;
  assign N1305 = N3943;
  assign N1306 = N3942;
  assign N1307 = N3941;
  assign N1308 = N3940;
  assign N1309 = N3939;
  assign N1310 = N3938;
  assign N1311 = N3937;
  assign N1312 = N3936;
  assign N1313 = N3935;
  assign N1314 = N3934;
  assign N1315 = N3933;
  assign N1316 = N3932;
  assign N1317 = N3931;
  assign N1318 = N3930;
  assign N1319 = N3929;
  assign N1320 = N3928;
  assign N1321 = N3927;
  assign N1322 = N3926;
  assign data_nn[991:960] = (N1225)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                            (N1226)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                            (N1227)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                            (N1228)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                            (N1229)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                            (N1230)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                            (N1231)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                            (N1232)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                            (N1233)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                            (N1234)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                            (N1235)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                            (N1236)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                            (N1237)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                            (N1238)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                            (N1239)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                            (N1240)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                            (N1241)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                            (N1242)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                            (N1243)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                            (N1244)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                            (N1245)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                            (N1246)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                            (N1247)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                            (N1248)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                            (N1249)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                            (N1250)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                            (N1251)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                            (N1252)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                            (N1253)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                            (N1254)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                            (N1255)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                            (N1256)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                            (N1257)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                            (N1258)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                            (N1259)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                            (N1260)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                            (N1261)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                            (N1262)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                            (N1263)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                            (N1264)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                            (N1265)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                            (N1266)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                            (N1267)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                            (N1268)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                            (N1269)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                            (N1270)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                            (N1271)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                            (N1272)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                            (N1273)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                            (N1274)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                            (N1275)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                            (N1276)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                            (N1277)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                            (N1278)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                            (N1279)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                            (N1280)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                            (N1281)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                            (N1282)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                            (N1283)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                            (N1284)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                            (N1285)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                            (N1286)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                            (N1287)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                            (N1288)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                            (N1289)? data_o[2047:2016] : 
                            (N1290)? data_o[2015:1984] : 
                            (N1291)? data_o[1983:1952] : 
                            (N1292)? data_o[1951:1920] : 
                            (N1293)? data_o[1919:1888] : 
                            (N1294)? data_o[1887:1856] : 
                            (N1295)? data_o[1855:1824] : 
                            (N1296)? data_o[1823:1792] : 
                            (N1297)? data_o[1791:1760] : 
                            (N1298)? data_o[1759:1728] : 
                            (N1299)? data_o[1727:1696] : 
                            (N1300)? data_o[1695:1664] : 
                            (N1301)? data_o[1663:1632] : 
                            (N1302)? data_o[1631:1600] : 
                            (N1303)? data_o[1599:1568] : 
                            (N1304)? data_o[1567:1536] : 
                            (N1305)? data_o[1535:1504] : 
                            (N1306)? data_o[1503:1472] : 
                            (N1307)? data_o[1471:1440] : 
                            (N1308)? data_o[1439:1408] : 
                            (N1309)? data_o[1407:1376] : 
                            (N1310)? data_o[1375:1344] : 
                            (N1311)? data_o[1343:1312] : 
                            (N1312)? data_o[1311:1280] : 
                            (N1313)? data_o[1279:1248] : 
                            (N1314)? data_o[1247:1216] : 
                            (N1315)? data_o[1215:1184] : 
                            (N1316)? data_o[1183:1152] : 
                            (N1317)? data_o[1151:1120] : 
                            (N1318)? data_o[1119:1088] : 
                            (N1319)? data_o[1087:1056] : 
                            (N1320)? data_o[1055:1024] : 
                            (N1321)? data_o[1023:992] : 
                            (N1322)? data_o[991:960] : 1'b0;
  assign data_nn[1023:992] = (N1226)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                             (N1227)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                             (N1228)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                             (N1229)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                             (N1230)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                             (N1231)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                             (N1232)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                             (N1233)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                             (N1234)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                             (N1235)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                             (N1236)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                             (N1237)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                             (N1238)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                             (N1239)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                             (N1240)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                             (N1241)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                             (N1242)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                             (N1243)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                             (N1244)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                             (N1245)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                             (N1246)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                             (N1247)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                             (N1248)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                             (N1249)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                             (N1250)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                             (N1251)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                             (N1252)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                             (N1253)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                             (N1254)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                             (N1255)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                             (N1256)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                             (N1257)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                             (N1258)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                             (N1259)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                             (N1260)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                             (N1261)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                             (N1262)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                             (N1263)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                             (N1264)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                             (N1265)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                             (N1266)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                             (N1267)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                             (N1268)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                             (N1269)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                             (N1270)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                             (N1271)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                             (N1272)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                             (N1273)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                             (N1274)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                             (N1275)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                             (N1276)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                             (N1277)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                             (N1278)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                             (N1279)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                             (N1280)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                             (N1281)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                             (N1282)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                             (N1283)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                             (N1284)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                             (N1285)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                             (N1286)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                             (N1287)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                             (N1288)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                             (N1289)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                             (N1290)? data_o[2047:2016] : 
                             (N1291)? data_o[2015:1984] : 
                             (N1292)? data_o[1983:1952] : 
                             (N1293)? data_o[1951:1920] : 
                             (N1294)? data_o[1919:1888] : 
                             (N1295)? data_o[1887:1856] : 
                             (N1296)? data_o[1855:1824] : 
                             (N1297)? data_o[1823:1792] : 
                             (N1298)? data_o[1791:1760] : 
                             (N1299)? data_o[1759:1728] : 
                             (N1300)? data_o[1727:1696] : 
                             (N1301)? data_o[1695:1664] : 
                             (N1302)? data_o[1663:1632] : 
                             (N1303)? data_o[1631:1600] : 
                             (N1304)? data_o[1599:1568] : 
                             (N1305)? data_o[1567:1536] : 
                             (N1306)? data_o[1535:1504] : 
                             (N1307)? data_o[1503:1472] : 
                             (N1308)? data_o[1471:1440] : 
                             (N1309)? data_o[1439:1408] : 
                             (N1310)? data_o[1407:1376] : 
                             (N1311)? data_o[1375:1344] : 
                             (N1312)? data_o[1343:1312] : 
                             (N1313)? data_o[1311:1280] : 
                             (N1314)? data_o[1279:1248] : 
                             (N1315)? data_o[1247:1216] : 
                             (N1316)? data_o[1215:1184] : 
                             (N1317)? data_o[1183:1152] : 
                             (N1318)? data_o[1151:1120] : 
                             (N1319)? data_o[1119:1088] : 
                             (N1320)? data_o[1087:1056] : 
                             (N1321)? data_o[1055:1024] : 
                             (N1322)? data_o[1023:992] : 1'b0;
  assign data_nn[1055:1024] = (N1227)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1228)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1229)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1230)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1231)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1232)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1233)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1234)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1235)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1236)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1237)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1238)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1239)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1240)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1241)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1242)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1243)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1244)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1245)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1246)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1247)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1248)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1249)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1250)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1251)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1252)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1253)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1254)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1255)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1256)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1257)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1258)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1259)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1260)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1261)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1262)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1263)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1264)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1265)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1266)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1267)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1268)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1269)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1270)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1271)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1272)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1273)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1274)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1275)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1276)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1277)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1278)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1279)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1280)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1281)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1282)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1283)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1284)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1285)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1286)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1287)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1288)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1289)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1290)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1291)? data_o[2047:2016] : 
                              (N1292)? data_o[2015:1984] : 
                              (N1293)? data_o[1983:1952] : 
                              (N1294)? data_o[1951:1920] : 
                              (N1295)? data_o[1919:1888] : 
                              (N1296)? data_o[1887:1856] : 
                              (N1297)? data_o[1855:1824] : 
                              (N1298)? data_o[1823:1792] : 
                              (N1299)? data_o[1791:1760] : 
                              (N1300)? data_o[1759:1728] : 
                              (N1301)? data_o[1727:1696] : 
                              (N1302)? data_o[1695:1664] : 
                              (N1303)? data_o[1663:1632] : 
                              (N1304)? data_o[1631:1600] : 
                              (N1305)? data_o[1599:1568] : 
                              (N1306)? data_o[1567:1536] : 
                              (N1307)? data_o[1535:1504] : 
                              (N1308)? data_o[1503:1472] : 
                              (N1309)? data_o[1471:1440] : 
                              (N1310)? data_o[1439:1408] : 
                              (N1311)? data_o[1407:1376] : 
                              (N1312)? data_o[1375:1344] : 
                              (N1313)? data_o[1343:1312] : 
                              (N1314)? data_o[1311:1280] : 
                              (N1315)? data_o[1279:1248] : 
                              (N1316)? data_o[1247:1216] : 
                              (N1317)? data_o[1215:1184] : 
                              (N1318)? data_o[1183:1152] : 
                              (N1319)? data_o[1151:1120] : 
                              (N1320)? data_o[1119:1088] : 
                              (N1321)? data_o[1087:1056] : 
                              (N1322)? data_o[1055:1024] : 1'b0;
  assign data_nn[1087:1056] = (N1228)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1229)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1230)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1231)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1232)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1233)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1234)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1235)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1236)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1237)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1238)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1239)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1240)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1241)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1242)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1243)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1244)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1245)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1246)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1247)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1248)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1249)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1250)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1251)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1252)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1253)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1254)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1255)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1256)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1257)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1258)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1259)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1260)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1261)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1262)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1263)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1264)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1265)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1266)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1267)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1268)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1269)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1270)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1271)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1272)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1273)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1274)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1275)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1276)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1277)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1278)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1279)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1280)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1281)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1282)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1283)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1284)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1285)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1286)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1287)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1288)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1289)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1290)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1291)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1292)? data_o[2047:2016] : 
                              (N1293)? data_o[2015:1984] : 
                              (N1294)? data_o[1983:1952] : 
                              (N1295)? data_o[1951:1920] : 
                              (N1296)? data_o[1919:1888] : 
                              (N1297)? data_o[1887:1856] : 
                              (N1298)? data_o[1855:1824] : 
                              (N1299)? data_o[1823:1792] : 
                              (N1300)? data_o[1791:1760] : 
                              (N1301)? data_o[1759:1728] : 
                              (N1302)? data_o[1727:1696] : 
                              (N1303)? data_o[1695:1664] : 
                              (N1304)? data_o[1663:1632] : 
                              (N1305)? data_o[1631:1600] : 
                              (N1306)? data_o[1599:1568] : 
                              (N1307)? data_o[1567:1536] : 
                              (N1308)? data_o[1535:1504] : 
                              (N1309)? data_o[1503:1472] : 
                              (N1310)? data_o[1471:1440] : 
                              (N1311)? data_o[1439:1408] : 
                              (N1312)? data_o[1407:1376] : 
                              (N1313)? data_o[1375:1344] : 
                              (N1314)? data_o[1343:1312] : 
                              (N1315)? data_o[1311:1280] : 
                              (N1316)? data_o[1279:1248] : 
                              (N1317)? data_o[1247:1216] : 
                              (N1318)? data_o[1215:1184] : 
                              (N1319)? data_o[1183:1152] : 
                              (N1320)? data_o[1151:1120] : 
                              (N1321)? data_o[1119:1088] : 
                              (N1322)? data_o[1087:1056] : 1'b0;
  assign data_nn[1119:1088] = (N1323)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1324)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1325)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1326)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1327)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1328)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1329)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1330)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1331)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1332)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1333)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1334)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1335)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1336)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1337)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1338)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1339)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1340)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1341)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1342)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1343)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1344)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1345)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1346)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1347)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1348)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1349)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1350)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1351)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1352)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1353)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1354)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1355)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1356)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1357)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1358)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1359)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1360)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1361)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1362)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1363)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1364)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1365)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1366)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1367)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1368)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1369)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1370)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1371)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1372)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1373)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1374)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1375)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1376)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1377)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1378)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1379)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1380)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1381)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1382)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1383)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1384)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1385)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1386)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1387)? data_o[2047:2016] : 
                              (N1388)? data_o[2015:1984] : 
                              (N1389)? data_o[1983:1952] : 
                              (N1390)? data_o[1951:1920] : 
                              (N1391)? data_o[1919:1888] : 
                              (N1392)? data_o[1887:1856] : 
                              (N1393)? data_o[1855:1824] : 
                              (N1394)? data_o[1823:1792] : 
                              (N1395)? data_o[1791:1760] : 
                              (N1396)? data_o[1759:1728] : 
                              (N1397)? data_o[1727:1696] : 
                              (N1398)? data_o[1695:1664] : 
                              (N1399)? data_o[1663:1632] : 
                              (N1400)? data_o[1631:1600] : 
                              (N1401)? data_o[1599:1568] : 
                              (N1402)? data_o[1567:1536] : 
                              (N1403)? data_o[1535:1504] : 
                              (N1404)? data_o[1503:1472] : 
                              (N1405)? data_o[1471:1440] : 
                              (N1406)? data_o[1439:1408] : 
                              (N1407)? data_o[1407:1376] : 
                              (N1408)? data_o[1375:1344] : 
                              (N1409)? data_o[1343:1312] : 
                              (N1410)? data_o[1311:1280] : 
                              (N1411)? data_o[1279:1248] : 
                              (N1412)? data_o[1247:1216] : 
                              (N1413)? data_o[1215:1184] : 
                              (N1414)? data_o[1183:1152] : 
                              (N1415)? data_o[1151:1120] : 
                              (N1416)? data_o[1119:1088] : 1'b0;
  assign N1323 = N5597;
  assign N1324 = N5598;
  assign N1325 = N5599;
  assign N1326 = N4172;
  assign N1327 = N4171;
  assign N1328 = N4170;
  assign N1329 = N4169;
  assign N1330 = N4168;
  assign N1331 = N4167;
  assign N1332 = N4166;
  assign N1333 = N4165;
  assign N1334 = N4164;
  assign N1335 = N4163;
  assign N1336 = N4162;
  assign N1337 = N4161;
  assign N1338 = N4160;
  assign N1339 = N4159;
  assign N1340 = N4158;
  assign N1341 = N4157;
  assign N1342 = N4156;
  assign N1343 = N4155;
  assign N1344 = N4154;
  assign N1345 = N4153;
  assign N1346 = N4152;
  assign N1347 = N4151;
  assign N1348 = N4150;
  assign N1349 = N4149;
  assign N1350 = N4148;
  assign N1351 = N4147;
  assign N1352 = N4146;
  assign N1353 = N3925;
  assign N1354 = N3924;
  assign N1355 = N3923;
  assign N1356 = N3922;
  assign N1357 = N3921;
  assign N1358 = N3920;
  assign N1359 = N3919;
  assign N1360 = N3918;
  assign N1361 = N3917;
  assign N1362 = N3916;
  assign N1363 = N3915;
  assign N1364 = N3914;
  assign N1365 = N3913;
  assign N1366 = N3912;
  assign N1367 = N3911;
  assign N1368 = N3910;
  assign N1369 = N3909;
  assign N1370 = N3908;
  assign N1371 = N3907;
  assign N1372 = N3906;
  assign N1373 = N3905;
  assign N1374 = N3904;
  assign N1375 = N3903;
  assign N1376 = N3902;
  assign N1377 = N3901;
  assign N1378 = N3900;
  assign N1379 = N3899;
  assign N1380 = N3898;
  assign N1381 = N3897;
  assign N1382 = N3896;
  assign N1383 = N3895;
  assign N1384 = N3894;
  assign N1385 = N3893;
  assign N1386 = N3892;
  assign N1387 = N3891;
  assign N1388 = N3890;
  assign N1389 = N3889;
  assign N1390 = N3888;
  assign N1391 = N3887;
  assign N1392 = N3886;
  assign N1393 = N3885;
  assign N1394 = N3884;
  assign N1395 = N3883;
  assign N1396 = N3882;
  assign N1397 = N3881;
  assign N1398 = N3880;
  assign N1399 = N3879;
  assign N1400 = N3878;
  assign N1401 = N3877;
  assign N1402 = N3876;
  assign N1403 = N3875;
  assign N1404 = N3874;
  assign N1405 = N3873;
  assign N1406 = N3872;
  assign N1407 = N3871;
  assign N1408 = N3870;
  assign N1409 = N3869;
  assign N1410 = N3868;
  assign N1411 = N3867;
  assign N1412 = N3866;
  assign N1413 = N3865;
  assign N1414 = N3864;
  assign N1415 = N3863;
  assign N1416 = N3862;
  assign data_nn[1151:1120] = (N1324)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1325)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1326)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1327)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1328)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1329)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1330)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1331)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1332)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1333)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1334)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1335)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1336)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1337)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1338)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1339)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1340)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1341)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1342)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1343)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1344)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1345)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1346)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1347)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1348)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1349)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1350)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1351)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1352)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1259)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1260)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1261)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1262)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1263)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1264)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1265)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1266)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1267)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1268)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1269)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1270)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1271)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1272)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1273)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1274)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1275)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1276)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1277)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1278)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1279)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1280)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1281)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1282)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1283)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1284)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1285)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1286)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1287)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1288)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1289)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1290)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1291)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1292)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1293)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1294)? data_o[2047:2016] : 
                              (N1295)? data_o[2015:1984] : 
                              (N1296)? data_o[1983:1952] : 
                              (N1297)? data_o[1951:1920] : 
                              (N1298)? data_o[1919:1888] : 
                              (N1299)? data_o[1887:1856] : 
                              (N1300)? data_o[1855:1824] : 
                              (N1301)? data_o[1823:1792] : 
                              (N1302)? data_o[1791:1760] : 
                              (N1303)? data_o[1759:1728] : 
                              (N1304)? data_o[1727:1696] : 
                              (N1305)? data_o[1695:1664] : 
                              (N1306)? data_o[1663:1632] : 
                              (N1307)? data_o[1631:1600] : 
                              (N1308)? data_o[1599:1568] : 
                              (N1309)? data_o[1567:1536] : 
                              (N1310)? data_o[1535:1504] : 
                              (N1311)? data_o[1503:1472] : 
                              (N1312)? data_o[1471:1440] : 
                              (N1313)? data_o[1439:1408] : 
                              (N1314)? data_o[1407:1376] : 
                              (N1315)? data_o[1375:1344] : 
                              (N1316)? data_o[1343:1312] : 
                              (N1317)? data_o[1311:1280] : 
                              (N1318)? data_o[1279:1248] : 
                              (N1319)? data_o[1247:1216] : 
                              (N1320)? data_o[1215:1184] : 
                              (N1321)? data_o[1183:1152] : 
                              (N1322)? data_o[1151:1120] : 1'b0;
  assign data_nn[1183:1152] = (N1417)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1418)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1419)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1420)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1421)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1422)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1423)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1424)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1425)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1426)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1427)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1428)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1429)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1430)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1431)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1432)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1433)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1434)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1435)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1436)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1437)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1438)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1439)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1440)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1441)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1442)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1443)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1444)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1445)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1446)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1447)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1448)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1449)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1450)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1451)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1452)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1453)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1454)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1455)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1456)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1457)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1458)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1459)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1460)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1461)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1462)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1463)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1464)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1465)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1466)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1467)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1468)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1469)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1470)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1471)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1472)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1473)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1474)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1475)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1476)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1477)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1478)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1479)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1480)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1481)? data_o[2047:2016] : 
                              (N1482)? data_o[2015:1984] : 
                              (N1483)? data_o[1983:1952] : 
                              (N1484)? data_o[1951:1920] : 
                              (N1485)? data_o[1919:1888] : 
                              (N1486)? data_o[1887:1856] : 
                              (N1487)? data_o[1855:1824] : 
                              (N1488)? data_o[1823:1792] : 
                              (N1489)? data_o[1791:1760] : 
                              (N1490)? data_o[1759:1728] : 
                              (N1491)? data_o[1727:1696] : 
                              (N1492)? data_o[1695:1664] : 
                              (N1493)? data_o[1663:1632] : 
                              (N1494)? data_o[1631:1600] : 
                              (N1495)? data_o[1599:1568] : 
                              (N1496)? data_o[1567:1536] : 
                              (N1497)? data_o[1535:1504] : 
                              (N1498)? data_o[1503:1472] : 
                              (N1499)? data_o[1471:1440] : 
                              (N1500)? data_o[1439:1408] : 
                              (N1501)? data_o[1407:1376] : 
                              (N1502)? data_o[1375:1344] : 
                              (N1503)? data_o[1343:1312] : 
                              (N1504)? data_o[1311:1280] : 
                              (N1505)? data_o[1279:1248] : 
                              (N1506)? data_o[1247:1216] : 
                              (N1507)? data_o[1215:1184] : 
                              (N1508)? data_o[1183:1152] : 1'b0;
  assign N1417 = N4081;
  assign N1418 = N4080;
  assign N1419 = N4079;
  assign N1420 = N4078;
  assign N1421 = N4077;
  assign N1422 = N4076;
  assign N1423 = N4075;
  assign N1424 = N4074;
  assign N1425 = N4073;
  assign N1426 = N4072;
  assign N1427 = N4071;
  assign N1428 = N4070;
  assign N1429 = N4069;
  assign N1430 = N4068;
  assign N1431 = N4067;
  assign N1432 = N4066;
  assign N1433 = N4065;
  assign N1434 = N4064;
  assign N1435 = N4063;
  assign N1436 = N4062;
  assign N1437 = N4061;
  assign N1438 = N4060;
  assign N1439 = N4059;
  assign N1440 = N4058;
  assign N1441 = N4057;
  assign N1442 = N4056;
  assign N1443 = N4055;
  assign N1444 = N4054;
  assign N1445 = N4053;
  assign N1446 = N4052;
  assign N1447 = N4051;
  assign N1448 = N4050;
  assign N1449 = N4049;
  assign N1450 = N4048;
  assign N1451 = N4047;
  assign N1452 = N4046;
  assign N1453 = N4045;
  assign N1454 = N4044;
  assign N1455 = N4043;
  assign N1456 = N4042;
  assign N1457 = N4041;
  assign N1458 = N4040;
  assign N1459 = N4039;
  assign N1460 = N4038;
  assign N1461 = N4037;
  assign N1462 = N4036;
  assign N1463 = N4035;
  assign N1464 = N4034;
  assign N1465 = N4033;
  assign N1466 = N4032;
  assign N1467 = N4031;
  assign N1468 = N4030;
  assign N1469 = N4029;
  assign N1470 = N4028;
  assign N1471 = N4027;
  assign N1472 = N4026;
  assign N1473 = N4025;
  assign N1474 = N4024;
  assign N1475 = N4023;
  assign N1476 = N4022;
  assign N1477 = N4021;
  assign N1478 = N4020;
  assign N1479 = N4019;
  assign N1480 = N4018;
  assign N1481 = N4017;
  assign N1482 = N4016;
  assign N1483 = N4015;
  assign N1484 = N4014;
  assign N1485 = N4013;
  assign N1486 = N4012;
  assign N1487 = N4011;
  assign N1488 = N4010;
  assign N1489 = N4009;
  assign N1490 = N4008;
  assign N1491 = N4007;
  assign N1492 = N4006;
  assign N1493 = N4005;
  assign N1494 = N4004;
  assign N1495 = N4003;
  assign N1496 = N4002;
  assign N1497 = N4001;
  assign N1498 = N4000;
  assign N1499 = N3999;
  assign N1500 = N3998;
  assign N1501 = N3997;
  assign N1502 = N3996;
  assign N1503 = N3995;
  assign N1504 = N3994;
  assign N1505 = N3993;
  assign N1506 = N3992;
  assign N1507 = N3991;
  assign N1508 = N3990;
  assign data_nn[1215:1184] = (N1326)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1327)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1328)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1329)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1330)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1331)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1332)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1333)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1334)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1335)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1336)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1337)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1338)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1339)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1340)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1341)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1342)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1343)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1344)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1345)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1346)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1347)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1348)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1349)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1350)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1351)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1352)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1509)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1510)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1511)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1512)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1513)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1514)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1515)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1516)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1517)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1518)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1519)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1520)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1521)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1522)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1523)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1524)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1525)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1526)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1527)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1528)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1529)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1530)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1531)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1532)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1533)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1534)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1535)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1536)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1537)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1538)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1539)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1540)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1541)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1542)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1543)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1544)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1545)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1546)? data_o[2047:2016] : 
                              (N1547)? data_o[2015:1984] : 
                              (N1548)? data_o[1983:1952] : 
                              (N1549)? data_o[1951:1920] : 
                              (N1550)? data_o[1919:1888] : 
                              (N1551)? data_o[1887:1856] : 
                              (N1552)? data_o[1855:1824] : 
                              (N1553)? data_o[1823:1792] : 
                              (N1554)? data_o[1791:1760] : 
                              (N1555)? data_o[1759:1728] : 
                              (N1556)? data_o[1727:1696] : 
                              (N1557)? data_o[1695:1664] : 
                              (N1558)? data_o[1663:1632] : 
                              (N1559)? data_o[1631:1600] : 
                              (N1560)? data_o[1599:1568] : 
                              (N1561)? data_o[1567:1536] : 
                              (N1562)? data_o[1535:1504] : 
                              (N1563)? data_o[1503:1472] : 
                              (N1564)? data_o[1471:1440] : 
                              (N1565)? data_o[1439:1408] : 
                              (N1566)? data_o[1407:1376] : 
                              (N1567)? data_o[1375:1344] : 
                              (N1568)? data_o[1343:1312] : 
                              (N1569)? data_o[1311:1280] : 
                              (N1570)? data_o[1279:1248] : 
                              (N1571)? data_o[1247:1216] : 
                              (N1572)? data_o[1215:1184] : 1'b0;
  assign N1509 = N4145;
  assign N1510 = N4144;
  assign N1511 = N4143;
  assign N1512 = N4142;
  assign N1513 = N4141;
  assign N1514 = N4140;
  assign N1515 = N4139;
  assign N1516 = N4138;
  assign N1517 = N4137;
  assign N1518 = N4136;
  assign N1519 = N4135;
  assign N1520 = N4134;
  assign N1521 = N4133;
  assign N1522 = N4132;
  assign N1523 = N4131;
  assign N1524 = N4130;
  assign N1525 = N4129;
  assign N1526 = N4128;
  assign N1527 = N4127;
  assign N1528 = N4126;
  assign N1529 = N4125;
  assign N1530 = N4124;
  assign N1531 = N4123;
  assign N1532 = N4122;
  assign N1533 = N4121;
  assign N1534 = N4120;
  assign N1535 = N4119;
  assign N1536 = N4118;
  assign N1537 = N4117;
  assign N1538 = N4116;
  assign N1539 = N4115;
  assign N1540 = N4114;
  assign N1541 = N4113;
  assign N1542 = N4112;
  assign N1543 = N4111;
  assign N1544 = N4110;
  assign N1545 = N4109;
  assign N1546 = N4108;
  assign N1547 = N4107;
  assign N1548 = N4106;
  assign N1549 = N4105;
  assign N1550 = N4104;
  assign N1551 = N4103;
  assign N1552 = N4102;
  assign N1553 = N4101;
  assign N1554 = N4100;
  assign N1555 = N4099;
  assign N1556 = N4098;
  assign N1557 = N4097;
  assign N1558 = N4096;
  assign N1559 = N4095;
  assign N1560 = N4094;
  assign N1561 = N4093;
  assign N1562 = N4092;
  assign N1563 = N4091;
  assign N1564 = N4090;
  assign N1565 = N4089;
  assign N1566 = N4088;
  assign N1567 = N4087;
  assign N1568 = N4086;
  assign N1569 = N4085;
  assign N1570 = N4084;
  assign N1571 = N4083;
  assign N1572 = N4082;
  assign data_nn[1247:1216] = (N1573)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1574)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1575)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1576)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1577)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1578)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1579)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1580)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1581)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1582)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1583)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1584)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1585)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1586)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1587)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1588)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1589)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1590)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1591)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1592)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1593)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1594)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1595)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1596)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1597)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1598)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N844)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N845)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N846)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N847)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N848)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N849)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N850)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N851)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N852)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N853)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N854)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N855)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N856)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N857)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N858)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N859)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N860)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N861)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N862)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N863)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N864)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N865)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N866)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N867)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N868)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N869)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N870)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N871)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N872)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N873)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N874)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N875)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N876)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N877)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N878)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N879)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N880)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N881)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N882)? data_o[2047:2016] : 
                              (N883)? data_o[2015:1984] : 
                              (N884)? data_o[1983:1952] : 
                              (N885)? data_o[1951:1920] : 
                              (N886)? data_o[1919:1888] : 
                              (N887)? data_o[1887:1856] : 
                              (N888)? data_o[1855:1824] : 
                              (N889)? data_o[1823:1792] : 
                              (N890)? data_o[1791:1760] : 
                              (N891)? data_o[1759:1728] : 
                              (N892)? data_o[1727:1696] : 
                              (N893)? data_o[1695:1664] : 
                              (N894)? data_o[1663:1632] : 
                              (N895)? data_o[1631:1600] : 
                              (N896)? data_o[1599:1568] : 
                              (N897)? data_o[1567:1536] : 
                              (N898)? data_o[1535:1504] : 
                              (N899)? data_o[1503:1472] : 
                              (N900)? data_o[1471:1440] : 
                              (N901)? data_o[1439:1408] : 
                              (N902)? data_o[1407:1376] : 
                              (N903)? data_o[1375:1344] : 
                              (N904)? data_o[1343:1312] : 
                              (N905)? data_o[1311:1280] : 
                              (N906)? data_o[1279:1248] : 
                              (N907)? data_o[1247:1216] : 1'b0;
  assign N1573 = N4262;
  assign N1574 = N4261;
  assign N1575 = N4260;
  assign N1576 = N4259;
  assign N1577 = N4258;
  assign N1578 = N4257;
  assign N1579 = N4256;
  assign N1580 = N4255;
  assign N1581 = N4254;
  assign N1582 = N4253;
  assign N1583 = N4252;
  assign N1584 = N4251;
  assign N1585 = N4250;
  assign N1586 = N4249;
  assign N1587 = N4248;
  assign N1588 = N4247;
  assign N1589 = N4246;
  assign N1590 = N4245;
  assign N1591 = N4244;
  assign N1592 = N4243;
  assign N1593 = N4242;
  assign N1594 = N4241;
  assign N1595 = N4240;
  assign N1596 = N4239;
  assign N1597 = N4238;
  assign N1598 = N4237;
  assign data_nn[1279:1248] = (N1599)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1600)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1601)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1602)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1603)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1604)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1605)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1606)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1607)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1608)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1609)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1610)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1611)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1612)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1613)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1614)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1615)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1616)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1617)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1618)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1619)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1620)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1621)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1622)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1623)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1624)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1625)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1626)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1627)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1628)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1629)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1630)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1631)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1632)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1633)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1634)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1635)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1636)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1637)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1638)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1639)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1640)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1641)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1642)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1643)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1644)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1645)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1646)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1647)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1648)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1649)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1650)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1651)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1652)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1653)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1654)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1655)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1656)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1657)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1658)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1659)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1660)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1661)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1662)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1663)? data_o[2047:2016] : 
                              (N1664)? data_o[2015:1984] : 
                              (N1665)? data_o[1983:1952] : 
                              (N1666)? data_o[1951:1920] : 
                              (N1667)? data_o[1919:1888] : 
                              (N1668)? data_o[1887:1856] : 
                              (N1669)? data_o[1855:1824] : 
                              (N1670)? data_o[1823:1792] : 
                              (N1671)? data_o[1791:1760] : 
                              (N1672)? data_o[1759:1728] : 
                              (N1673)? data_o[1727:1696] : 
                              (N1674)? data_o[1695:1664] : 
                              (N1675)? data_o[1663:1632] : 
                              (N1676)? data_o[1631:1600] : 
                              (N1677)? data_o[1599:1568] : 
                              (N1678)? data_o[1567:1536] : 
                              (N1679)? data_o[1535:1504] : 
                              (N1680)? data_o[1503:1472] : 
                              (N1681)? data_o[1471:1440] : 
                              (N1682)? data_o[1439:1408] : 
                              (N1683)? data_o[1407:1376] : 
                              (N1684)? data_o[1375:1344] : 
                              (N1685)? data_o[1343:1312] : 
                              (N1686)? data_o[1311:1280] : 
                              (N1687)? data_o[1279:1248] : 1'b0;
  assign N1599 = N5628;
  assign N1600 = N5629;
  assign N1601 = N5630;
  assign N1602 = N5631;
  assign N1603 = N4283;
  assign N1604 = N4282;
  assign N1605 = N4281;
  assign N1606 = N4280;
  assign N1607 = N4279;
  assign N1608 = N4278;
  assign N1609 = N4277;
  assign N1610 = N4276;
  assign N1611 = N4275;
  assign N1612 = N4274;
  assign N1613 = N4273;
  assign N1614 = N4272;
  assign N1615 = N4271;
  assign N1616 = N4270;
  assign N1617 = N4269;
  assign N1618 = N4268;
  assign N1619 = N4267;
  assign N1620 = N4266;
  assign N1621 = N4265;
  assign N1622 = N4264;
  assign N1623 = N4263;
  assign N1624 = N4870;
  assign N1625 = N4869;
  assign N1626 = N4868;
  assign N1627 = N4867;
  assign N1628 = N4866;
  assign N1629 = N4865;
  assign N1630 = N4864;
  assign N1631 = N4863;
  assign N1632 = N4862;
  assign N1633 = N4861;
  assign N1634 = N4860;
  assign N1635 = N4859;
  assign N1636 = N4858;
  assign N1637 = N4857;
  assign N1638 = N4856;
  assign N1639 = N4855;
  assign N1640 = N4854;
  assign N1641 = N4853;
  assign N1642 = N4852;
  assign N1643 = N4851;
  assign N1644 = N4850;
  assign N1645 = N4849;
  assign N1646 = N4848;
  assign N1647 = N4847;
  assign N1648 = N4846;
  assign N1649 = N4845;
  assign N1650 = N4844;
  assign N1651 = N4843;
  assign N1652 = N4842;
  assign N1653 = N4841;
  assign N1654 = N4840;
  assign N1655 = N4839;
  assign N1656 = N4838;
  assign N1657 = N4837;
  assign N1658 = N4836;
  assign N1659 = N4835;
  assign N1660 = N4834;
  assign N1661 = N4833;
  assign N1662 = N4832;
  assign N1663 = N4831;
  assign N1664 = N4830;
  assign N1665 = N4829;
  assign N1666 = N4828;
  assign N1667 = N4827;
  assign N1668 = N4826;
  assign N1669 = N4825;
  assign N1670 = N4824;
  assign N1671 = N4823;
  assign N1672 = N4822;
  assign N1673 = N4821;
  assign N1674 = N4820;
  assign N1675 = N4819;
  assign N1676 = N4818;
  assign N1677 = N4817;
  assign N1678 = N4816;
  assign N1679 = N4815;
  assign N1680 = N4814;
  assign N1681 = N4813;
  assign N1682 = N4812;
  assign N1683 = N4811;
  assign N1684 = N4810;
  assign N1685 = N4809;
  assign N1686 = N4808;
  assign N1687 = N4807;
  assign data_nn[1311:1280] = (N1600)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1601)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1602)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1603)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1604)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1605)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1606)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1607)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1608)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1609)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1610)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1611)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1612)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1613)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1614)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1615)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1616)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1617)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1618)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1619)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1620)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1621)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1622)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1623)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1624)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1625)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1626)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1627)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1628)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1629)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1630)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1631)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1632)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1633)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1634)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1635)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1636)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1637)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1638)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1639)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1640)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1641)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1642)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1643)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1644)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1645)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1646)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1647)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1648)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1649)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1650)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1651)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1652)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1653)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1654)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1655)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1656)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1657)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1658)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1659)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1660)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1661)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1662)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1663)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1664)? data_o[2047:2016] : 
                              (N1665)? data_o[2015:1984] : 
                              (N1666)? data_o[1983:1952] : 
                              (N1667)? data_o[1951:1920] : 
                              (N1668)? data_o[1919:1888] : 
                              (N1669)? data_o[1887:1856] : 
                              (N1670)? data_o[1855:1824] : 
                              (N1671)? data_o[1823:1792] : 
                              (N1672)? data_o[1791:1760] : 
                              (N1673)? data_o[1759:1728] : 
                              (N1674)? data_o[1727:1696] : 
                              (N1675)? data_o[1695:1664] : 
                              (N1676)? data_o[1663:1632] : 
                              (N1677)? data_o[1631:1600] : 
                              (N1678)? data_o[1599:1568] : 
                              (N1679)? data_o[1567:1536] : 
                              (N1680)? data_o[1535:1504] : 
                              (N1681)? data_o[1503:1472] : 
                              (N1682)? data_o[1471:1440] : 
                              (N1683)? data_o[1439:1408] : 
                              (N1684)? data_o[1407:1376] : 
                              (N1685)? data_o[1375:1344] : 
                              (N1686)? data_o[1343:1312] : 
                              (N1687)? data_o[1311:1280] : 1'b0;
  assign data_nn[1343:1312] = (N1601)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1602)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1603)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1604)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1605)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1606)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1607)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1608)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1609)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1610)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1611)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1612)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1613)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1614)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1615)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1616)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1617)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1618)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1619)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1620)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1621)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1622)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1623)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1624)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1625)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1626)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1627)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1628)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1629)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1630)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1631)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1632)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1633)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1634)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1635)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1636)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1637)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1638)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1639)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1640)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1641)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1642)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1643)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1644)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1645)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1646)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1647)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1648)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1649)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1650)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1651)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1652)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1653)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1654)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1655)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1656)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1657)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1658)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1659)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1660)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1661)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1662)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1663)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1664)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1665)? data_o[2047:2016] : 
                              (N1666)? data_o[2015:1984] : 
                              (N1667)? data_o[1983:1952] : 
                              (N1668)? data_o[1951:1920] : 
                              (N1669)? data_o[1919:1888] : 
                              (N1670)? data_o[1887:1856] : 
                              (N1671)? data_o[1855:1824] : 
                              (N1672)? data_o[1823:1792] : 
                              (N1673)? data_o[1791:1760] : 
                              (N1674)? data_o[1759:1728] : 
                              (N1675)? data_o[1727:1696] : 
                              (N1676)? data_o[1695:1664] : 
                              (N1677)? data_o[1663:1632] : 
                              (N1678)? data_o[1631:1600] : 
                              (N1679)? data_o[1599:1568] : 
                              (N1680)? data_o[1567:1536] : 
                              (N1681)? data_o[1535:1504] : 
                              (N1682)? data_o[1503:1472] : 
                              (N1683)? data_o[1471:1440] : 
                              (N1684)? data_o[1439:1408] : 
                              (N1685)? data_o[1407:1376] : 
                              (N1686)? data_o[1375:1344] : 
                              (N1687)? data_o[1343:1312] : 1'b0;
  assign data_nn[1375:1344] = (N1602)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1603)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1604)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1605)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1606)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1607)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1608)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1609)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1610)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1611)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1612)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1613)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1614)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1615)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1616)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1617)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1618)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1619)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1620)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1621)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1622)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1623)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1624)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1625)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1626)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1627)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1628)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1629)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1630)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1631)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1632)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1633)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1634)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1635)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1636)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1637)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1638)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1639)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1640)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1641)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1642)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1643)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1644)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1645)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1646)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1647)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1648)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1649)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1650)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1651)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1652)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1653)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1654)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1655)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1656)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1657)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1658)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1659)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1660)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1661)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1662)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1663)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1664)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1665)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1666)? data_o[2047:2016] : 
                              (N1667)? data_o[2015:1984] : 
                              (N1668)? data_o[1983:1952] : 
                              (N1669)? data_o[1951:1920] : 
                              (N1670)? data_o[1919:1888] : 
                              (N1671)? data_o[1887:1856] : 
                              (N1672)? data_o[1855:1824] : 
                              (N1673)? data_o[1823:1792] : 
                              (N1674)? data_o[1791:1760] : 
                              (N1675)? data_o[1759:1728] : 
                              (N1676)? data_o[1727:1696] : 
                              (N1677)? data_o[1695:1664] : 
                              (N1678)? data_o[1663:1632] : 
                              (N1679)? data_o[1631:1600] : 
                              (N1680)? data_o[1599:1568] : 
                              (N1681)? data_o[1567:1536] : 
                              (N1682)? data_o[1535:1504] : 
                              (N1683)? data_o[1503:1472] : 
                              (N1684)? data_o[1471:1440] : 
                              (N1685)? data_o[1439:1408] : 
                              (N1686)? data_o[1407:1376] : 
                              (N1687)? data_o[1375:1344] : 1'b0;
  assign data_nn[1407:1376] = (N1603)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1604)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1605)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1606)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1607)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1608)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1609)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1610)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1611)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1612)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1613)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1614)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1615)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1616)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1617)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1618)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1619)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1620)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1621)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1622)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1623)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1624)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1625)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1626)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1627)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1628)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1629)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1630)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1631)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1632)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1633)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1634)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1635)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1636)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1637)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1638)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1639)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1640)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1641)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1642)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1643)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1644)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1645)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1646)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1647)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1648)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1649)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1650)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1651)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1652)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1653)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1654)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1655)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1656)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1657)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1658)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1659)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1660)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1661)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1662)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1663)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1664)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1665)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1666)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1667)? data_o[2047:2016] : 
                              (N1668)? data_o[2015:1984] : 
                              (N1669)? data_o[1983:1952] : 
                              (N1670)? data_o[1951:1920] : 
                              (N1671)? data_o[1919:1888] : 
                              (N1672)? data_o[1887:1856] : 
                              (N1673)? data_o[1855:1824] : 
                              (N1674)? data_o[1823:1792] : 
                              (N1675)? data_o[1791:1760] : 
                              (N1676)? data_o[1759:1728] : 
                              (N1677)? data_o[1727:1696] : 
                              (N1678)? data_o[1695:1664] : 
                              (N1679)? data_o[1663:1632] : 
                              (N1680)? data_o[1631:1600] : 
                              (N1681)? data_o[1599:1568] : 
                              (N1682)? data_o[1567:1536] : 
                              (N1683)? data_o[1535:1504] : 
                              (N1684)? data_o[1503:1472] : 
                              (N1685)? data_o[1471:1440] : 
                              (N1686)? data_o[1439:1408] : 
                              (N1687)? data_o[1407:1376] : 1'b0;
  assign data_nn[1439:1408] = (N1688)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1689)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1690)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1691)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1692)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1693)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1694)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1695)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1696)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1697)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1698)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1699)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1700)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1701)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1702)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1703)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1704)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1705)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1706)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1707)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1708)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1709)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1710)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1711)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1712)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1713)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1714)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1715)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1716)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1717)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1718)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1719)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1720)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1721)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1722)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1723)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1724)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1725)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1726)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1727)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1728)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1729)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1730)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1731)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1732)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1733)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1734)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1735)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1736)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1737)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1738)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1739)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1740)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1741)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1742)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1743)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1744)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1745)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1746)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1747)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1748)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1749)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1750)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1751)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1752)? data_o[2047:2016] : 
                              (N1753)? data_o[2015:1984] : 
                              (N1754)? data_o[1983:1952] : 
                              (N1755)? data_o[1951:1920] : 
                              (N1756)? data_o[1919:1888] : 
                              (N1757)? data_o[1887:1856] : 
                              (N1758)? data_o[1855:1824] : 
                              (N1759)? data_o[1823:1792] : 
                              (N1760)? data_o[1791:1760] : 
                              (N1761)? data_o[1759:1728] : 
                              (N1762)? data_o[1727:1696] : 
                              (N1763)? data_o[1695:1664] : 
                              (N1764)? data_o[1663:1632] : 
                              (N1765)? data_o[1631:1600] : 
                              (N1766)? data_o[1599:1568] : 
                              (N1767)? data_o[1567:1536] : 
                              (N1768)? data_o[1535:1504] : 
                              (N1769)? data_o[1503:1472] : 
                              (N1770)? data_o[1471:1440] : 
                              (N1771)? data_o[1439:1408] : 1'b0;
  assign N1688 = N5632;
  assign N1689 = N5633;
  assign N1690 = N5634;
  assign N1691 = N5635;
  assign N1692 = N4363;
  assign N1693 = N4362;
  assign N1694 = N4361;
  assign N1695 = N4360;
  assign N1696 = N4359;
  assign N1697 = N4358;
  assign N1698 = N4357;
  assign N1699 = N4356;
  assign N1700 = N4355;
  assign N1701 = N4354;
  assign N1702 = N4353;
  assign N1703 = N4352;
  assign N1704 = N4351;
  assign N1705 = N4350;
  assign N1706 = N4349;
  assign N1707 = N4348;
  assign N1708 = N4347;
  assign N1709 = N4346;
  assign N1710 = N4345;
  assign N1711 = N4344;
  assign N1712 = N4343;
  assign N1713 = N4342;
  assign N1714 = N4341;
  assign N1715 = N4340;
  assign N1716 = N4339;
  assign N1717 = N4338;
  assign N1718 = N4337;
  assign N1719 = N4336;
  assign N1720 = N4335;
  assign N1721 = N4334;
  assign N1722 = N4333;
  assign N1723 = N4332;
  assign N1724 = N4331;
  assign N1725 = N4330;
  assign N1726 = N4329;
  assign N1727 = N4328;
  assign N1728 = N4327;
  assign N1729 = N4326;
  assign N1730 = N4325;
  assign N1731 = N4324;
  assign N1732 = N4323;
  assign N1733 = N4322;
  assign N1734 = N4321;
  assign N1735 = N4320;
  assign N1736 = N4319;
  assign N1737 = N4318;
  assign N1738 = N4317;
  assign N1739 = N4316;
  assign N1740 = N4315;
  assign N1741 = N4314;
  assign N1742 = N4313;
  assign N1743 = N4312;
  assign N1744 = N4311;
  assign N1745 = N4310;
  assign N1746 = N4309;
  assign N1747 = N4308;
  assign N1748 = N4307;
  assign N1749 = N4306;
  assign N1750 = N4305;
  assign N1751 = N4304;
  assign N1752 = N4303;
  assign N1753 = N4302;
  assign N1754 = N4301;
  assign N1755 = N4300;
  assign N1756 = N4299;
  assign N1757 = N4298;
  assign N1758 = N4297;
  assign N1759 = N4296;
  assign N1760 = N4295;
  assign N1761 = N4294;
  assign N1762 = N4293;
  assign N1763 = N4292;
  assign N1764 = N4291;
  assign N1765 = N4290;
  assign N1766 = N4289;
  assign N1767 = N4288;
  assign N1768 = N4287;
  assign N1769 = N4286;
  assign N1770 = N4285;
  assign N1771 = N4284;
  assign data_nn[1471:1440] = (N1689)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1690)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1691)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1692)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1693)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1694)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1695)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1696)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1697)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1698)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1699)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1700)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1701)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1702)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1703)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1704)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1705)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1706)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1707)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1708)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1709)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1710)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1711)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1712)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1713)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1714)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1715)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1716)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1717)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1718)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1719)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1720)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1721)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1722)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1723)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1724)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1725)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1726)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1727)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1728)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1729)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1730)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1731)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1732)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1733)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1734)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1735)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1736)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1737)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1738)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1739)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1740)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1741)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1742)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1743)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1744)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1745)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1746)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1747)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1748)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1749)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1750)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1751)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1752)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1753)? data_o[2047:2016] : 
                              (N1754)? data_o[2015:1984] : 
                              (N1755)? data_o[1983:1952] : 
                              (N1756)? data_o[1951:1920] : 
                              (N1757)? data_o[1919:1888] : 
                              (N1758)? data_o[1887:1856] : 
                              (N1759)? data_o[1855:1824] : 
                              (N1760)? data_o[1823:1792] : 
                              (N1761)? data_o[1791:1760] : 
                              (N1762)? data_o[1759:1728] : 
                              (N1763)? data_o[1727:1696] : 
                              (N1764)? data_o[1695:1664] : 
                              (N1765)? data_o[1663:1632] : 
                              (N1766)? data_o[1631:1600] : 
                              (N1767)? data_o[1599:1568] : 
                              (N1768)? data_o[1567:1536] : 
                              (N1769)? data_o[1535:1504] : 
                              (N1770)? data_o[1503:1472] : 
                              (N1771)? data_o[1471:1440] : 1'b0;
  assign data_nn[1503:1472] = (N1690)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1691)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1692)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1693)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1694)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1695)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1696)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1697)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1698)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1699)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1700)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1701)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1702)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1703)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1704)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1705)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1706)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1707)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1708)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1709)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1710)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1711)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1712)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1713)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1714)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1715)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1716)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1717)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1718)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1719)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1720)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1721)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1722)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1723)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1724)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1725)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1726)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1727)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1728)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1729)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1730)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1731)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1732)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1733)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1734)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1735)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1736)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1737)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1738)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1739)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1740)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1741)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1742)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1743)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1744)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1745)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1746)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1747)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1748)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1749)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1750)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1751)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1752)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1753)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1754)? data_o[2047:2016] : 
                              (N1755)? data_o[2015:1984] : 
                              (N1756)? data_o[1983:1952] : 
                              (N1757)? data_o[1951:1920] : 
                              (N1758)? data_o[1919:1888] : 
                              (N1759)? data_o[1887:1856] : 
                              (N1760)? data_o[1855:1824] : 
                              (N1761)? data_o[1823:1792] : 
                              (N1762)? data_o[1791:1760] : 
                              (N1763)? data_o[1759:1728] : 
                              (N1764)? data_o[1727:1696] : 
                              (N1765)? data_o[1695:1664] : 
                              (N1766)? data_o[1663:1632] : 
                              (N1767)? data_o[1631:1600] : 
                              (N1768)? data_o[1599:1568] : 
                              (N1769)? data_o[1567:1536] : 
                              (N1770)? data_o[1535:1504] : 
                              (N1771)? data_o[1503:1472] : 1'b0;
  assign data_nn[1535:1504] = (N1691)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1692)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1693)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1694)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1695)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1696)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1697)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1698)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1699)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1700)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1701)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1702)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1703)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1704)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1705)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1706)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1707)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1708)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1709)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1710)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1711)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1712)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1713)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1714)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1715)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1716)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1717)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1718)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1719)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1720)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1721)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1722)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1723)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1724)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1725)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1726)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1727)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1728)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1729)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1730)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1731)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1732)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1733)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1734)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1735)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1736)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1737)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1738)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1739)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1740)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1741)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1742)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1743)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1744)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1745)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1746)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1747)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1748)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1749)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1750)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1751)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1752)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1753)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1754)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1755)? data_o[2047:2016] : 
                              (N1756)? data_o[2015:1984] : 
                              (N1757)? data_o[1983:1952] : 
                              (N1758)? data_o[1951:1920] : 
                              (N1759)? data_o[1919:1888] : 
                              (N1760)? data_o[1887:1856] : 
                              (N1761)? data_o[1855:1824] : 
                              (N1762)? data_o[1823:1792] : 
                              (N1763)? data_o[1791:1760] : 
                              (N1764)? data_o[1759:1728] : 
                              (N1765)? data_o[1727:1696] : 
                              (N1766)? data_o[1695:1664] : 
                              (N1767)? data_o[1663:1632] : 
                              (N1768)? data_o[1631:1600] : 
                              (N1769)? data_o[1599:1568] : 
                              (N1770)? data_o[1567:1536] : 
                              (N1771)? data_o[1535:1504] : 1'b0;
  assign data_nn[1567:1536] = (N1692)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1693)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1694)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1695)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1696)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1697)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1698)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1699)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1700)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1701)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1702)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1703)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1704)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1705)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1706)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1707)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1708)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1709)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1710)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1711)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1712)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1713)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1714)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1715)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1716)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1717)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1718)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1719)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1720)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1721)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1722)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1723)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1724)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1725)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1726)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1727)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1728)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1729)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1730)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1731)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1732)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1733)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1734)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1735)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1736)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1737)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1738)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1739)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1740)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1741)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1742)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1743)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1744)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1745)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1746)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1747)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1748)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1749)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1750)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1751)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1752)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1753)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1754)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1755)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1756)? data_o[2047:2016] : 
                              (N1757)? data_o[2015:1984] : 
                              (N1758)? data_o[1983:1952] : 
                              (N1759)? data_o[1951:1920] : 
                              (N1760)? data_o[1919:1888] : 
                              (N1761)? data_o[1887:1856] : 
                              (N1762)? data_o[1855:1824] : 
                              (N1763)? data_o[1823:1792] : 
                              (N1764)? data_o[1791:1760] : 
                              (N1765)? data_o[1759:1728] : 
                              (N1766)? data_o[1727:1696] : 
                              (N1767)? data_o[1695:1664] : 
                              (N1768)? data_o[1663:1632] : 
                              (N1769)? data_o[1631:1600] : 
                              (N1770)? data_o[1599:1568] : 
                              (N1771)? data_o[1567:1536] : 1'b0;
  assign data_nn[1599:1568] = (N1772)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1773)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1774)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1775)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1776)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1777)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1778)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1779)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1780)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1781)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1782)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1783)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1784)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1785)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1786)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1787)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1788)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1789)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1790)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1791)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1792)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1793)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1794)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1795)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1796)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1797)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1798)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1799)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1800)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1801)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1802)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1803)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1804)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1805)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1806)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1807)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1808)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1809)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1810)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1811)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1812)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1813)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1814)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1815)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1816)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1817)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1818)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1819)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1820)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1821)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1822)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1823)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1824)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1825)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1826)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1827)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1828)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1829)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1830)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1831)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1832)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1833)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1834)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1835)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1836)? data_o[2047:2016] : 
                              (N1837)? data_o[2015:1984] : 
                              (N1838)? data_o[1983:1952] : 
                              (N1839)? data_o[1951:1920] : 
                              (N1840)? data_o[1919:1888] : 
                              (N1841)? data_o[1887:1856] : 
                              (N1842)? data_o[1855:1824] : 
                              (N1843)? data_o[1823:1792] : 
                              (N1844)? data_o[1791:1760] : 
                              (N1845)? data_o[1759:1728] : 
                              (N1846)? data_o[1727:1696] : 
                              (N1847)? data_o[1695:1664] : 
                              (N1848)? data_o[1663:1632] : 
                              (N1849)? data_o[1631:1600] : 
                              (N1850)? data_o[1599:1568] : 1'b0;
  assign N1772 = N4442;
  assign N1773 = N4441;
  assign N1774 = N4440;
  assign N1775 = N4439;
  assign N1776 = N4438;
  assign N1777 = N4437;
  assign N1778 = N4436;
  assign N1779 = N4435;
  assign N1780 = N4434;
  assign N1781 = N4433;
  assign N1782 = N4432;
  assign N1783 = N4431;
  assign N1784 = N4430;
  assign N1785 = N4429;
  assign N1786 = N4428;
  assign N1787 = N4427;
  assign N1788 = N4426;
  assign N1789 = N4425;
  assign N1790 = N4424;
  assign N1791 = N4423;
  assign N1792 = N4422;
  assign N1793 = N4421;
  assign N1794 = N4420;
  assign N1795 = N4419;
  assign N1796 = N4418;
  assign N1797 = N4417;
  assign N1798 = N4416;
  assign N1799 = N4415;
  assign N1800 = N4414;
  assign N1801 = N4413;
  assign N1802 = N4412;
  assign N1803 = N4411;
  assign N1804 = N4410;
  assign N1805 = N4409;
  assign N1806 = N4408;
  assign N1807 = N4407;
  assign N1808 = N4406;
  assign N1809 = N4405;
  assign N1810 = N4404;
  assign N1811 = N4403;
  assign N1812 = N4402;
  assign N1813 = N4401;
  assign N1814 = N4400;
  assign N1815 = N4399;
  assign N1816 = N4398;
  assign N1817 = N4397;
  assign N1818 = N4396;
  assign N1819 = N4395;
  assign N1820 = N4394;
  assign N1821 = N4393;
  assign N1822 = N4392;
  assign N1823 = N4391;
  assign N1824 = N4390;
  assign N1825 = N4389;
  assign N1826 = N4388;
  assign N1827 = N4387;
  assign N1828 = N4386;
  assign N1829 = N4385;
  assign N1830 = N4384;
  assign N1831 = N4383;
  assign N1832 = N4382;
  assign N1833 = N4381;
  assign N1834 = N4380;
  assign N1835 = N4379;
  assign N1836 = N4378;
  assign N1837 = N4377;
  assign N1838 = N4376;
  assign N1839 = N4375;
  assign N1840 = N4374;
  assign N1841 = N4373;
  assign N1842 = N4372;
  assign N1843 = N4371;
  assign N1844 = N4370;
  assign N1845 = N4369;
  assign N1846 = N4368;
  assign N1847 = N4367;
  assign N1848 = N4366;
  assign N1849 = N4365;
  assign N1850 = N4364;
  assign data_nn[1631:1600] = (N1851)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1852)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1853)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1854)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1855)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1856)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1857)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1858)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1859)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1860)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1861)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1862)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1863)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1864)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1865)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1866)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1867)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1868)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1869)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1870)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1871)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1872)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1873)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1874)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1875)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1876)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1877)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1878)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1879)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1880)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1881)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1882)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1883)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1884)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1885)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1886)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1887)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1888)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1889)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1890)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1891)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1892)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1893)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1894)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1895)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1896)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1897)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1898)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1899)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1900)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1901)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1902)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1903)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1904)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1905)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1906)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1907)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1908)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1909)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1910)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1911)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1912)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1913)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1914)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1915)? data_o[2047:2016] : 
                              (N1916)? data_o[2015:1984] : 
                              (N1917)? data_o[1983:1952] : 
                              (N1918)? data_o[1951:1920] : 
                              (N1919)? data_o[1919:1888] : 
                              (N1920)? data_o[1887:1856] : 
                              (N1921)? data_o[1855:1824] : 
                              (N1922)? data_o[1823:1792] : 
                              (N1923)? data_o[1791:1760] : 
                              (N1924)? data_o[1759:1728] : 
                              (N1925)? data_o[1727:1696] : 
                              (N1926)? data_o[1695:1664] : 
                              (N1927)? data_o[1663:1632] : 
                              (N1928)? data_o[1631:1600] : 1'b0;
  assign N1851 = N5639;
  assign N1852 = N5640;
  assign N1853 = N5641;
  assign N1854 = N5642;
  assign N1855 = N5643;
  assign N1856 = N5644;
  assign N1857 = N4523;
  assign N1858 = N4522;
  assign N1859 = N4521;
  assign N1860 = N4520;
  assign N1861 = N4519;
  assign N1862 = N4518;
  assign N1863 = N4517;
  assign N1864 = N4516;
  assign N1865 = N4506;
  assign N1866 = N4505;
  assign N1867 = N4504;
  assign N1868 = N4503;
  assign N1869 = N4502;
  assign N1870 = N4501;
  assign N1871 = N4500;
  assign N1872 = N4499;
  assign N1873 = N4498;
  assign N1874 = N4497;
  assign N1875 = N4496;
  assign N1876 = N4495;
  assign N1877 = N4494;
  assign N1878 = N4493;
  assign N1879 = N4492;
  assign N1880 = N4491;
  assign N1881 = N4490;
  assign N1882 = N4489;
  assign N1883 = N4488;
  assign N1884 = N4487;
  assign N1885 = N4486;
  assign N1886 = N4485;
  assign N1887 = N4484;
  assign N1888 = N4483;
  assign N1889 = N4482;
  assign N1890 = N4481;
  assign N1891 = N4480;
  assign N1892 = N4479;
  assign N1893 = N4478;
  assign N1894 = N4477;
  assign N1895 = N4476;
  assign N1896 = N4475;
  assign N1897 = N4474;
  assign N1898 = N4473;
  assign N1899 = N4472;
  assign N1900 = N4471;
  assign N1901 = N4470;
  assign N1902 = N4469;
  assign N1903 = N4468;
  assign N1904 = N4467;
  assign N1905 = N4466;
  assign N1906 = N4465;
  assign N1907 = N4464;
  assign N1908 = N4463;
  assign N1909 = N4462;
  assign N1910 = N4461;
  assign N1911 = N4460;
  assign N1912 = N4459;
  assign N1913 = N4458;
  assign N1914 = N4457;
  assign N1915 = N4456;
  assign N1916 = N4455;
  assign N1917 = N4454;
  assign N1918 = N4453;
  assign N1919 = N4452;
  assign N1920 = N4451;
  assign N1921 = N4450;
  assign N1922 = N4449;
  assign N1923 = N4448;
  assign N1924 = N4447;
  assign N1925 = N4446;
  assign N1926 = N4445;
  assign N1927 = N4444;
  assign N1928 = N4443;
  assign data_nn[1663:1632] = (N1852)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1853)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1854)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1855)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1856)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1857)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1858)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1859)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1860)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1861)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1862)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1863)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1864)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1865)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1866)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1867)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1868)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1869)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1870)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1871)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1872)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1873)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1874)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1875)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1876)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1877)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1878)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1879)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1880)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1881)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1882)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1883)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1884)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1885)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1886)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1887)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1888)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1889)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1890)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1891)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1892)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1893)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1894)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1895)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1896)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1897)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1898)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1899)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1900)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1901)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1902)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1903)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1904)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1905)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1906)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1907)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1908)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1909)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1910)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1911)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1912)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1913)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1914)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1915)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1916)? data_o[2047:2016] : 
                              (N1917)? data_o[2015:1984] : 
                              (N1918)? data_o[1983:1952] : 
                              (N1919)? data_o[1951:1920] : 
                              (N1920)? data_o[1919:1888] : 
                              (N1921)? data_o[1887:1856] : 
                              (N1922)? data_o[1855:1824] : 
                              (N1923)? data_o[1823:1792] : 
                              (N1924)? data_o[1791:1760] : 
                              (N1925)? data_o[1759:1728] : 
                              (N1926)? data_o[1727:1696] : 
                              (N1927)? data_o[1695:1664] : 
                              (N1928)? data_o[1663:1632] : 1'b0;
  assign data_nn[1695:1664] = (N1853)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1854)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1855)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1856)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1857)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1858)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1859)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1860)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1861)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1862)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1863)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1864)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1865)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1866)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1867)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1868)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1869)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1870)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1871)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1872)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1873)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1874)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1875)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1876)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1877)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1878)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1879)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1880)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1881)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1882)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1883)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1884)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1885)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1886)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1887)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1888)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1889)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1890)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1891)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1892)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1893)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1894)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1895)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1896)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1897)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1898)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1899)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1900)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1901)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1902)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1903)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1904)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1905)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1906)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1907)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1908)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1909)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1910)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1911)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1912)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1913)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1914)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1915)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1916)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1917)? data_o[2047:2016] : 
                              (N1918)? data_o[2015:1984] : 
                              (N1919)? data_o[1983:1952] : 
                              (N1920)? data_o[1951:1920] : 
                              (N1921)? data_o[1919:1888] : 
                              (N1922)? data_o[1887:1856] : 
                              (N1923)? data_o[1855:1824] : 
                              (N1924)? data_o[1823:1792] : 
                              (N1925)? data_o[1791:1760] : 
                              (N1926)? data_o[1759:1728] : 
                              (N1927)? data_o[1727:1696] : 
                              (N1928)? data_o[1695:1664] : 1'b0;
  assign data_nn[1727:1696] = (N1854)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1855)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1856)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1857)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1858)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1859)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1860)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1861)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1862)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1863)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1864)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1865)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1866)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1867)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1868)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1869)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1870)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1871)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1872)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1873)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1874)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1875)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1876)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1877)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1878)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1879)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1880)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1881)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1882)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1883)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1884)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1885)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1886)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1887)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1888)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1889)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1890)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1891)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1892)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1893)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1894)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1895)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1896)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1897)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1898)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1899)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1900)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1901)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1902)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1903)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1904)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1905)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1906)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1907)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1908)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1909)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1910)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1911)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1912)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1913)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1914)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1915)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1916)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1917)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1918)? data_o[2047:2016] : 
                              (N1919)? data_o[2015:1984] : 
                              (N1920)? data_o[1983:1952] : 
                              (N1921)? data_o[1951:1920] : 
                              (N1922)? data_o[1919:1888] : 
                              (N1923)? data_o[1887:1856] : 
                              (N1924)? data_o[1855:1824] : 
                              (N1925)? data_o[1823:1792] : 
                              (N1926)? data_o[1791:1760] : 
                              (N1927)? data_o[1759:1728] : 
                              (N1928)? data_o[1727:1696] : 1'b0;
  assign data_nn[1759:1728] = (N1929)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1930)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1931)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1932)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1933)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1934)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1935)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1936)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1937)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1938)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1939)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1940)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1941)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1942)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1943)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1944)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1945)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1946)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1947)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1948)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1949)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1950)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1951)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1952)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1953)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1954)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1955)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1956)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1957)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1958)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1959)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1960)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1961)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1962)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1963)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1964)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1965)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1966)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1967)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1968)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1969)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1970)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1971)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1972)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1973)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1974)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1975)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1976)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1977)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1978)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1979)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1980)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1981)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1982)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1983)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1984)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1985)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1986)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1987)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1988)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1989)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1990)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1991)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1992)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1993)? data_o[2047:2016] : 
                              (N1994)? data_o[2015:1984] : 
                              (N1995)? data_o[1983:1952] : 
                              (N1996)? data_o[1951:1920] : 
                              (N1997)? data_o[1919:1888] : 
                              (N1998)? data_o[1887:1856] : 
                              (N1999)? data_o[1855:1824] : 
                              (N2000)? data_o[1823:1792] : 
                              (N2001)? data_o[1791:1760] : 
                              (N2002)? data_o[1759:1728] : 1'b0;
  assign N1929 = N5637;
  assign N1930 = N4515;
  assign N1931 = N4514;
  assign N1932 = N4513;
  assign N1933 = N4512;
  assign N1934 = N4511;
  assign N1935 = N4510;
  assign N1936 = N4509;
  assign N1937 = N4508;
  assign N1938 = N4507;
  assign N1939 = N4669;
  assign N1940 = N4668;
  assign N1941 = N4667;
  assign N1942 = N4666;
  assign N1943 = N4665;
  assign N1944 = N4664;
  assign N1945 = N4663;
  assign N1946 = N4662;
  assign N1947 = N4661;
  assign N1948 = N4660;
  assign N1949 = N4659;
  assign N1950 = N4658;
  assign N1951 = N4657;
  assign N1952 = N4656;
  assign N1953 = N4655;
  assign N1954 = N4654;
  assign N1955 = N4653;
  assign N1956 = N4652;
  assign N1957 = N4651;
  assign N1958 = N4650;
  assign N1959 = N4649;
  assign N1960 = N4648;
  assign N1961 = N4647;
  assign N1962 = N4646;
  assign N1963 = N4645;
  assign N1964 = N4644;
  assign N1965 = N4643;
  assign N1966 = N4642;
  assign N1967 = N4641;
  assign N1968 = N4640;
  assign N1969 = N4639;
  assign N1970 = N4638;
  assign N1971 = N4637;
  assign N1972 = N4636;
  assign N1973 = N4635;
  assign N1974 = N4634;
  assign N1975 = N4633;
  assign N1976 = N4632;
  assign N1977 = N4631;
  assign N1978 = N4630;
  assign N1979 = N4629;
  assign N1980 = N4628;
  assign N1981 = N4627;
  assign N1982 = N4626;
  assign N1983 = N4625;
  assign N1984 = N4624;
  assign N1985 = N4623;
  assign N1986 = N4622;
  assign N1987 = N4621;
  assign N1988 = N4620;
  assign N1989 = N4619;
  assign N1990 = N4618;
  assign N1991 = N4617;
  assign N1992 = N4616;
  assign N1993 = N4615;
  assign N1994 = N4614;
  assign N1995 = N4613;
  assign N1996 = N4612;
  assign N1997 = N4611;
  assign N1998 = N4610;
  assign N1999 = N4609;
  assign N2000 = N4608;
  assign N2001 = N4607;
  assign N2002 = N4606;
  assign data_nn[1791:1760] = (N1930)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1931)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1932)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1933)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1934)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1935)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1936)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1937)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1938)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1939)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1940)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1941)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1942)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1943)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1944)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1945)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1946)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1947)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1948)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1949)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1950)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1951)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1952)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1953)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1954)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1955)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1956)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1957)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1958)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1959)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1960)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1961)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1962)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1963)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1964)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1965)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1966)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1967)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1968)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1969)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1970)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1971)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1972)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1973)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1974)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1975)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1976)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1977)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1978)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1979)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1980)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1981)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1982)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1983)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1984)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1985)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1986)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1987)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1988)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1989)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1990)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1991)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1992)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1993)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1994)? data_o[2047:2016] : 
                              (N1995)? data_o[2015:1984] : 
                              (N1996)? data_o[1983:1952] : 
                              (N1997)? data_o[1951:1920] : 
                              (N1998)? data_o[1919:1888] : 
                              (N1999)? data_o[1887:1856] : 
                              (N2000)? data_o[1855:1824] : 
                              (N2001)? data_o[1823:1792] : 
                              (N2002)? data_o[1791:1760] : 1'b0;
  assign data_nn[1823:1792] = (N1857)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1858)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1859)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1860)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1861)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1862)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1863)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1864)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1939)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1940)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1941)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1942)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1943)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1944)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1945)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1946)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1947)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1948)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1949)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1950)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1951)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1952)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1953)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1954)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1955)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1956)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1957)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1958)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1959)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1960)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1961)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1962)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1963)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1964)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1965)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1966)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1967)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1968)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1969)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1970)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1971)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1972)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1973)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1974)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1975)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1976)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1977)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1978)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1979)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1980)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1981)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1982)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1983)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1984)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1985)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1986)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1987)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1988)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1989)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1990)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1991)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1992)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1993)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1994)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1995)? data_o[2047:2016] : 
                              (N1996)? data_o[2015:1984] : 
                              (N1997)? data_o[1983:1952] : 
                              (N1998)? data_o[1951:1920] : 
                              (N1999)? data_o[1919:1888] : 
                              (N2000)? data_o[1887:1856] : 
                              (N2001)? data_o[1855:1824] : 
                              (N2002)? data_o[1823:1792] : 1'b0;
  assign data_nn[1855:1824] = (N2003)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N2004)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N2005)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N2006)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N2007)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N2008)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N2009)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1939)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1940)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1941)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1942)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1943)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1944)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1945)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1946)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1947)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1948)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1949)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1950)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1951)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1952)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1953)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1954)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1955)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1956)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1957)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1958)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1959)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1960)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1961)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1962)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1963)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1964)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1965)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1966)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1967)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1968)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1969)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1970)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1971)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1972)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1973)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1974)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1975)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1976)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1977)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1978)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1979)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1980)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1981)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1982)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1983)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1984)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1985)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1986)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1987)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1988)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1989)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1990)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1991)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1992)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1993)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1994)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1995)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1996)? data_o[2047:2016] : 
                              (N1997)? data_o[2015:1984] : 
                              (N1998)? data_o[1983:1952] : 
                              (N1999)? data_o[1951:1920] : 
                              (N2000)? data_o[1919:1888] : 
                              (N2001)? data_o[1887:1856] : 
                              (N2002)? data_o[1855:1824] : 1'b0;
  assign N2003 = N4530;
  assign N2004 = N4529;
  assign N2005 = N4528;
  assign N2006 = N4527;
  assign N2007 = N4526;
  assign N2008 = N4525;
  assign N2009 = N4524;
  assign data_nn[1887:1856] = (N2010)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N2011)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N2012)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N2013)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N2014)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N2015)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1939)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1940)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1941)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1942)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1943)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1944)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1945)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1946)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1947)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1948)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1949)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1950)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1951)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1952)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1953)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1954)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1955)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1956)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1957)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1958)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1959)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1960)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1961)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1962)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1963)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1964)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1965)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1966)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1967)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1968)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1969)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1970)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1971)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1972)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1973)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1974)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1975)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1976)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1977)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1978)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1979)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1980)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1981)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1982)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1983)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1984)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1985)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1986)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1987)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1988)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1989)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1990)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1991)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1992)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1993)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1994)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1995)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1996)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1997)? data_o[2047:2016] : 
                              (N1998)? data_o[2015:1984] : 
                              (N1999)? data_o[1983:1952] : 
                              (N2000)? data_o[1951:1920] : 
                              (N2001)? data_o[1919:1888] : 
                              (N2002)? data_o[1887:1856] : 1'b0;
  assign N2010 = N4536;
  assign N2011 = N4535;
  assign N2012 = N4534;
  assign N2013 = N4533;
  assign N2014 = N4532;
  assign N2015 = N4531;
  assign data_nn[1919:1888] = (N2016)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N2017)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N2018)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N2019)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N2020)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N2021)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N2022)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N2023)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N2024)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N2025)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N2026)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N2027)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N2028)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N2029)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N2030)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N2031)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N2032)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N2033)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N2034)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N2035)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N2036)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N2037)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N2038)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N2039)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N2040)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N2041)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N2042)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N2043)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N2044)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N2045)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N2046)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N2047)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N2048)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N2049)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N2050)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N2051)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N2052)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N2053)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N2054)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N2055)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N2056)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N2057)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N2058)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N2059)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N2060)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N2061)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N2062)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N2063)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N2064)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N2065)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N2066)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N2067)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N2068)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N2069)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N2070)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N2071)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N2072)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N2073)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N2074)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N2075)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N2076)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N2077)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N2078)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N2079)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N2080)? data_o[2047:2016] : 
                              (N2081)? data_o[2015:1984] : 
                              (N2082)? data_o[1983:1952] : 
                              (N2083)? data_o[1951:1920] : 
                              (N2084)? data_o[1919:1888] : 1'b0;
  assign N2016 = N4605;
  assign N2017 = N4604;
  assign N2018 = N4603;
  assign N2019 = N4602;
  assign N2020 = N4601;
  assign N2021 = N4600;
  assign N2022 = N4599;
  assign N2023 = N4598;
  assign N2024 = N4597;
  assign N2025 = N4596;
  assign N2026 = N4595;
  assign N2027 = N4594;
  assign N2028 = N4593;
  assign N2029 = N4592;
  assign N2030 = N4591;
  assign N2031 = N4590;
  assign N2032 = N4589;
  assign N2033 = N4588;
  assign N2034 = N4587;
  assign N2035 = N4586;
  assign N2036 = N4585;
  assign N2037 = N4584;
  assign N2038 = N4583;
  assign N2039 = N4582;
  assign N2040 = N4581;
  assign N2041 = N4580;
  assign N2042 = N4579;
  assign N2043 = N4578;
  assign N2044 = N4577;
  assign N2045 = N4576;
  assign N2046 = N4575;
  assign N2047 = N4574;
  assign N2048 = N4573;
  assign N2049 = N4572;
  assign N2050 = N4571;
  assign N2051 = N4570;
  assign N2052 = N4569;
  assign N2053 = N4568;
  assign N2054 = N4567;
  assign N2055 = N4566;
  assign N2056 = N4565;
  assign N2057 = N4564;
  assign N2058 = N4563;
  assign N2059 = N4562;
  assign N2060 = N4561;
  assign N2061 = N4560;
  assign N2062 = N4559;
  assign N2063 = N4558;
  assign N2064 = N4557;
  assign N2065 = N4556;
  assign N2066 = N4555;
  assign N2067 = N4554;
  assign N2068 = N4553;
  assign N2069 = N4552;
  assign N2070 = N4551;
  assign N2071 = N4550;
  assign N2072 = N4549;
  assign N2073 = N4548;
  assign N2074 = N4547;
  assign N2075 = N4546;
  assign N2076 = N4545;
  assign N2077 = N4544;
  assign N2078 = N4543;
  assign N2079 = N4542;
  assign N2080 = N4541;
  assign N2081 = N4540;
  assign N2082 = N4539;
  assign N2083 = N4538;
  assign N2084 = N4537;
  assign data_nn[1951:1920] = (N2085)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N2086)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N2087)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N2088)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1939)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1940)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1941)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1942)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1943)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1944)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1945)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1946)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1947)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1948)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1949)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1950)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1951)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1952)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1953)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1954)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1955)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1956)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1957)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1958)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1959)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1960)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1961)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1962)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1963)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1964)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1965)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1966)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1967)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1968)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1969)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1970)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1971)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1972)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1973)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1974)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1975)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1976)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1977)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1978)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1979)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1980)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1981)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1982)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1983)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1984)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1985)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1986)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1987)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1988)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1989)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1990)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1991)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1992)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1993)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1994)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1995)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1996)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1997)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1998)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1999)? data_o[2047:2016] : 
                              (N2000)? data_o[2015:1984] : 
                              (N2001)? data_o[1983:1952] : 
                              (N2002)? data_o[1951:1920] : 1'b0;
  assign N2085 = N4673;
  assign N2086 = N4672;
  assign N2087 = N4671;
  assign N2088 = N4670;
  assign data_nn[1983:1952] = (N2089)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N2090)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N2091)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N2092)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N2093)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N2094)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N2095)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N2096)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N2097)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N2098)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N2099)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N2100)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N2101)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N2102)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N2103)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N2104)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N2105)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N2106)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N2107)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N2108)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N2109)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N2110)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N2111)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N2112)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N2113)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N2114)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N2115)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N2116)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N2117)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N2118)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N2119)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N2120)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N2121)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N2122)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N2123)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N2124)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N2125)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N2126)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N2127)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N2128)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N2129)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N2130)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N2131)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N2132)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N2133)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N2134)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N2135)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N2136)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N2137)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N2138)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N2139)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N2140)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N2141)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N2142)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N2143)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N2144)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N2145)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N2146)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N2147)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N2148)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N2149)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N2150)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N2151)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N2152)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N2153)? data_o[2047:2016] : 
                              (N2154)? data_o[2015:1984] : 
                              (N2155)? data_o[1983:1952] : 1'b0;
  assign N2089 = N4740;
  assign N2090 = N4739;
  assign N2091 = N4738;
  assign N2092 = N4737;
  assign N2093 = N4736;
  assign N2094 = N4735;
  assign N2095 = N4734;
  assign N2096 = N4733;
  assign N2097 = N4732;
  assign N2098 = N4731;
  assign N2099 = N4730;
  assign N2100 = N4729;
  assign N2101 = N4728;
  assign N2102 = N4727;
  assign N2103 = N4726;
  assign N2104 = N4725;
  assign N2105 = N4724;
  assign N2106 = N4723;
  assign N2107 = N4722;
  assign N2108 = N4721;
  assign N2109 = N4720;
  assign N2110 = N4719;
  assign N2111 = N4718;
  assign N2112 = N4717;
  assign N2113 = N4716;
  assign N2114 = N4715;
  assign N2115 = N4714;
  assign N2116 = N4713;
  assign N2117 = N4712;
  assign N2118 = N4711;
  assign N2119 = N4710;
  assign N2120 = N4709;
  assign N2121 = N4708;
  assign N2122 = N4707;
  assign N2123 = N4706;
  assign N2124 = N4705;
  assign N2125 = N4704;
  assign N2126 = N4703;
  assign N2127 = N4702;
  assign N2128 = N4701;
  assign N2129 = N4700;
  assign N2130 = N4699;
  assign N2131 = N4698;
  assign N2132 = N4697;
  assign N2133 = N4696;
  assign N2134 = N4695;
  assign N2135 = N4694;
  assign N2136 = N4693;
  assign N2137 = N4692;
  assign N2138 = N4691;
  assign N2139 = N4690;
  assign N2140 = N4689;
  assign N2141 = N4688;
  assign N2142 = N4687;
  assign N2143 = N4686;
  assign N2144 = N4685;
  assign N2145 = N4684;
  assign N2146 = N4683;
  assign N2147 = N4682;
  assign N2148 = N4681;
  assign N2149 = N4680;
  assign N2150 = N4679;
  assign N2151 = N4678;
  assign N2152 = N4677;
  assign N2153 = N4676;
  assign N2154 = N4675;
  assign N2155 = N4674;
  assign data_nn[2015:1984] = (N2156)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N2157)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N2158)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N2159)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N2160)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N2161)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N2162)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N2163)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N2164)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N2165)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N2166)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N2167)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N2168)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N2169)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N2170)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N2171)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N2172)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N2173)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N2174)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N2175)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N2176)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N2177)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N2178)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N2179)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N2180)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N2181)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N2182)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N2183)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N2184)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N2185)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N2186)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N2187)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N2188)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N2189)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N2190)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N2191)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N2192)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N2193)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N2194)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N2195)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N2196)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N2197)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N2198)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N2199)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N2200)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N2201)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N2202)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N2203)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N2204)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N2205)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N2206)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N2207)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N2208)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N2209)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N2210)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N2211)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N2212)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N2213)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N2214)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N2215)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N2216)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N2217)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N2218)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N2219)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N2220)? data_o[2047:2016] : 
                              (N2221)? data_o[2015:1984] : 1'b0;
  assign N2156 = N4806;
  assign N2157 = N4805;
  assign N2158 = N4804;
  assign N2159 = N4803;
  assign N2160 = N4802;
  assign N2161 = N4801;
  assign N2162 = N4800;
  assign N2163 = N4799;
  assign N2164 = N4798;
  assign N2165 = N4797;
  assign N2166 = N4796;
  assign N2167 = N4795;
  assign N2168 = N4794;
  assign N2169 = N4793;
  assign N2170 = N4792;
  assign N2171 = N4791;
  assign N2172 = N4790;
  assign N2173 = N4789;
  assign N2174 = N4788;
  assign N2175 = N4787;
  assign N2176 = N4786;
  assign N2177 = N4785;
  assign N2178 = N4784;
  assign N2179 = N4783;
  assign N2180 = N4782;
  assign N2181 = N4781;
  assign N2182 = N4780;
  assign N2183 = N4779;
  assign N2184 = N4778;
  assign N2185 = N4777;
  assign N2186 = N4776;
  assign N2187 = N4775;
  assign N2188 = N4774;
  assign N2189 = N4773;
  assign N2190 = N4772;
  assign N2191 = N4771;
  assign N2192 = N4770;
  assign N2193 = N4769;
  assign N2194 = N4768;
  assign N2195 = N4767;
  assign N2196 = N4766;
  assign N2197 = N4765;
  assign N2198 = N4764;
  assign N2199 = N4763;
  assign N2200 = N4762;
  assign N2201 = N4761;
  assign N2202 = N4760;
  assign N2203 = N4759;
  assign N2204 = N4758;
  assign N2205 = N4757;
  assign N2206 = N4756;
  assign N2207 = N4755;
  assign N2208 = N4754;
  assign N2209 = N4753;
  assign N2210 = N4752;
  assign N2211 = N4751;
  assign N2212 = N4750;
  assign N2213 = N4749;
  assign N2214 = N4748;
  assign N2215 = N4747;
  assign N2216 = N4746;
  assign N2217 = N4745;
  assign N2218 = N4744;
  assign N2219 = N4743;
  assign N2220 = N4742;
  assign N2221 = N4741;
  assign data_nn[2047:2016] = (N2222)? { data_n_127__31_, data_n_127__30_, data_n_127__29_, data_n_127__28_, data_n_127__27_, data_n_127__26_, data_n_127__25_, data_n_127__24_, data_n_127__23_, data_n_127__22_, data_n_127__21_, data_n_127__20_, data_n_127__19_, data_n_127__18_, data_n_127__17_, data_n_127__16_, data_n_127__15_, data_n_127__14_, data_n_127__13_, data_n_127__12_, data_n_127__11_, data_n_127__10_, data_n_127__9_, data_n_127__8_, data_n_127__7_, data_n_127__6_, data_n_127__5_, data_n_127__4_, data_n_127__3_, data_n_127__2_, data_n_127__1_, data_n_127__0_ } : 
                              (N1624)? { data_n_126__31_, data_n_126__30_, data_n_126__29_, data_n_126__28_, data_n_126__27_, data_n_126__26_, data_n_126__25_, data_n_126__24_, data_n_126__23_, data_n_126__22_, data_n_126__21_, data_n_126__20_, data_n_126__19_, data_n_126__18_, data_n_126__17_, data_n_126__16_, data_n_126__15_, data_n_126__14_, data_n_126__13_, data_n_126__12_, data_n_126__11_, data_n_126__10_, data_n_126__9_, data_n_126__8_, data_n_126__7_, data_n_126__6_, data_n_126__5_, data_n_126__4_, data_n_126__3_, data_n_126__2_, data_n_126__1_, data_n_126__0_ } : 
                              (N1625)? { data_n_125__31_, data_n_125__30_, data_n_125__29_, data_n_125__28_, data_n_125__27_, data_n_125__26_, data_n_125__25_, data_n_125__24_, data_n_125__23_, data_n_125__22_, data_n_125__21_, data_n_125__20_, data_n_125__19_, data_n_125__18_, data_n_125__17_, data_n_125__16_, data_n_125__15_, data_n_125__14_, data_n_125__13_, data_n_125__12_, data_n_125__11_, data_n_125__10_, data_n_125__9_, data_n_125__8_, data_n_125__7_, data_n_125__6_, data_n_125__5_, data_n_125__4_, data_n_125__3_, data_n_125__2_, data_n_125__1_, data_n_125__0_ } : 
                              (N1626)? { data_n_124__31_, data_n_124__30_, data_n_124__29_, data_n_124__28_, data_n_124__27_, data_n_124__26_, data_n_124__25_, data_n_124__24_, data_n_124__23_, data_n_124__22_, data_n_124__21_, data_n_124__20_, data_n_124__19_, data_n_124__18_, data_n_124__17_, data_n_124__16_, data_n_124__15_, data_n_124__14_, data_n_124__13_, data_n_124__12_, data_n_124__11_, data_n_124__10_, data_n_124__9_, data_n_124__8_, data_n_124__7_, data_n_124__6_, data_n_124__5_, data_n_124__4_, data_n_124__3_, data_n_124__2_, data_n_124__1_, data_n_124__0_ } : 
                              (N1627)? { data_n_123__31_, data_n_123__30_, data_n_123__29_, data_n_123__28_, data_n_123__27_, data_n_123__26_, data_n_123__25_, data_n_123__24_, data_n_123__23_, data_n_123__22_, data_n_123__21_, data_n_123__20_, data_n_123__19_, data_n_123__18_, data_n_123__17_, data_n_123__16_, data_n_123__15_, data_n_123__14_, data_n_123__13_, data_n_123__12_, data_n_123__11_, data_n_123__10_, data_n_123__9_, data_n_123__8_, data_n_123__7_, data_n_123__6_, data_n_123__5_, data_n_123__4_, data_n_123__3_, data_n_123__2_, data_n_123__1_, data_n_123__0_ } : 
                              (N1628)? { data_n_122__31_, data_n_122__30_, data_n_122__29_, data_n_122__28_, data_n_122__27_, data_n_122__26_, data_n_122__25_, data_n_122__24_, data_n_122__23_, data_n_122__22_, data_n_122__21_, data_n_122__20_, data_n_122__19_, data_n_122__18_, data_n_122__17_, data_n_122__16_, data_n_122__15_, data_n_122__14_, data_n_122__13_, data_n_122__12_, data_n_122__11_, data_n_122__10_, data_n_122__9_, data_n_122__8_, data_n_122__7_, data_n_122__6_, data_n_122__5_, data_n_122__4_, data_n_122__3_, data_n_122__2_, data_n_122__1_, data_n_122__0_ } : 
                              (N1629)? { data_n_121__31_, data_n_121__30_, data_n_121__29_, data_n_121__28_, data_n_121__27_, data_n_121__26_, data_n_121__25_, data_n_121__24_, data_n_121__23_, data_n_121__22_, data_n_121__21_, data_n_121__20_, data_n_121__19_, data_n_121__18_, data_n_121__17_, data_n_121__16_, data_n_121__15_, data_n_121__14_, data_n_121__13_, data_n_121__12_, data_n_121__11_, data_n_121__10_, data_n_121__9_, data_n_121__8_, data_n_121__7_, data_n_121__6_, data_n_121__5_, data_n_121__4_, data_n_121__3_, data_n_121__2_, data_n_121__1_, data_n_121__0_ } : 
                              (N1630)? { data_n_120__31_, data_n_120__30_, data_n_120__29_, data_n_120__28_, data_n_120__27_, data_n_120__26_, data_n_120__25_, data_n_120__24_, data_n_120__23_, data_n_120__22_, data_n_120__21_, data_n_120__20_, data_n_120__19_, data_n_120__18_, data_n_120__17_, data_n_120__16_, data_n_120__15_, data_n_120__14_, data_n_120__13_, data_n_120__12_, data_n_120__11_, data_n_120__10_, data_n_120__9_, data_n_120__8_, data_n_120__7_, data_n_120__6_, data_n_120__5_, data_n_120__4_, data_n_120__3_, data_n_120__2_, data_n_120__1_, data_n_120__0_ } : 
                              (N1631)? { data_n_119__31_, data_n_119__30_, data_n_119__29_, data_n_119__28_, data_n_119__27_, data_n_119__26_, data_n_119__25_, data_n_119__24_, data_n_119__23_, data_n_119__22_, data_n_119__21_, data_n_119__20_, data_n_119__19_, data_n_119__18_, data_n_119__17_, data_n_119__16_, data_n_119__15_, data_n_119__14_, data_n_119__13_, data_n_119__12_, data_n_119__11_, data_n_119__10_, data_n_119__9_, data_n_119__8_, data_n_119__7_, data_n_119__6_, data_n_119__5_, data_n_119__4_, data_n_119__3_, data_n_119__2_, data_n_119__1_, data_n_119__0_ } : 
                              (N1632)? { data_n_118__31_, data_n_118__30_, data_n_118__29_, data_n_118__28_, data_n_118__27_, data_n_118__26_, data_n_118__25_, data_n_118__24_, data_n_118__23_, data_n_118__22_, data_n_118__21_, data_n_118__20_, data_n_118__19_, data_n_118__18_, data_n_118__17_, data_n_118__16_, data_n_118__15_, data_n_118__14_, data_n_118__13_, data_n_118__12_, data_n_118__11_, data_n_118__10_, data_n_118__9_, data_n_118__8_, data_n_118__7_, data_n_118__6_, data_n_118__5_, data_n_118__4_, data_n_118__3_, data_n_118__2_, data_n_118__1_, data_n_118__0_ } : 
                              (N1633)? { data_n_117__31_, data_n_117__30_, data_n_117__29_, data_n_117__28_, data_n_117__27_, data_n_117__26_, data_n_117__25_, data_n_117__24_, data_n_117__23_, data_n_117__22_, data_n_117__21_, data_n_117__20_, data_n_117__19_, data_n_117__18_, data_n_117__17_, data_n_117__16_, data_n_117__15_, data_n_117__14_, data_n_117__13_, data_n_117__12_, data_n_117__11_, data_n_117__10_, data_n_117__9_, data_n_117__8_, data_n_117__7_, data_n_117__6_, data_n_117__5_, data_n_117__4_, data_n_117__3_, data_n_117__2_, data_n_117__1_, data_n_117__0_ } : 
                              (N1634)? { data_n_116__31_, data_n_116__30_, data_n_116__29_, data_n_116__28_, data_n_116__27_, data_n_116__26_, data_n_116__25_, data_n_116__24_, data_n_116__23_, data_n_116__22_, data_n_116__21_, data_n_116__20_, data_n_116__19_, data_n_116__18_, data_n_116__17_, data_n_116__16_, data_n_116__15_, data_n_116__14_, data_n_116__13_, data_n_116__12_, data_n_116__11_, data_n_116__10_, data_n_116__9_, data_n_116__8_, data_n_116__7_, data_n_116__6_, data_n_116__5_, data_n_116__4_, data_n_116__3_, data_n_116__2_, data_n_116__1_, data_n_116__0_ } : 
                              (N1635)? { data_n_115__31_, data_n_115__30_, data_n_115__29_, data_n_115__28_, data_n_115__27_, data_n_115__26_, data_n_115__25_, data_n_115__24_, data_n_115__23_, data_n_115__22_, data_n_115__21_, data_n_115__20_, data_n_115__19_, data_n_115__18_, data_n_115__17_, data_n_115__16_, data_n_115__15_, data_n_115__14_, data_n_115__13_, data_n_115__12_, data_n_115__11_, data_n_115__10_, data_n_115__9_, data_n_115__8_, data_n_115__7_, data_n_115__6_, data_n_115__5_, data_n_115__4_, data_n_115__3_, data_n_115__2_, data_n_115__1_, data_n_115__0_ } : 
                              (N1636)? { data_n_114__31_, data_n_114__30_, data_n_114__29_, data_n_114__28_, data_n_114__27_, data_n_114__26_, data_n_114__25_, data_n_114__24_, data_n_114__23_, data_n_114__22_, data_n_114__21_, data_n_114__20_, data_n_114__19_, data_n_114__18_, data_n_114__17_, data_n_114__16_, data_n_114__15_, data_n_114__14_, data_n_114__13_, data_n_114__12_, data_n_114__11_, data_n_114__10_, data_n_114__9_, data_n_114__8_, data_n_114__7_, data_n_114__6_, data_n_114__5_, data_n_114__4_, data_n_114__3_, data_n_114__2_, data_n_114__1_, data_n_114__0_ } : 
                              (N1637)? { data_n_113__31_, data_n_113__30_, data_n_113__29_, data_n_113__28_, data_n_113__27_, data_n_113__26_, data_n_113__25_, data_n_113__24_, data_n_113__23_, data_n_113__22_, data_n_113__21_, data_n_113__20_, data_n_113__19_, data_n_113__18_, data_n_113__17_, data_n_113__16_, data_n_113__15_, data_n_113__14_, data_n_113__13_, data_n_113__12_, data_n_113__11_, data_n_113__10_, data_n_113__9_, data_n_113__8_, data_n_113__7_, data_n_113__6_, data_n_113__5_, data_n_113__4_, data_n_113__3_, data_n_113__2_, data_n_113__1_, data_n_113__0_ } : 
                              (N1638)? { data_n_112__31_, data_n_112__30_, data_n_112__29_, data_n_112__28_, data_n_112__27_, data_n_112__26_, data_n_112__25_, data_n_112__24_, data_n_112__23_, data_n_112__22_, data_n_112__21_, data_n_112__20_, data_n_112__19_, data_n_112__18_, data_n_112__17_, data_n_112__16_, data_n_112__15_, data_n_112__14_, data_n_112__13_, data_n_112__12_, data_n_112__11_, data_n_112__10_, data_n_112__9_, data_n_112__8_, data_n_112__7_, data_n_112__6_, data_n_112__5_, data_n_112__4_, data_n_112__3_, data_n_112__2_, data_n_112__1_, data_n_112__0_ } : 
                              (N1639)? { data_n_111__31_, data_n_111__30_, data_n_111__29_, data_n_111__28_, data_n_111__27_, data_n_111__26_, data_n_111__25_, data_n_111__24_, data_n_111__23_, data_n_111__22_, data_n_111__21_, data_n_111__20_, data_n_111__19_, data_n_111__18_, data_n_111__17_, data_n_111__16_, data_n_111__15_, data_n_111__14_, data_n_111__13_, data_n_111__12_, data_n_111__11_, data_n_111__10_, data_n_111__9_, data_n_111__8_, data_n_111__7_, data_n_111__6_, data_n_111__5_, data_n_111__4_, data_n_111__3_, data_n_111__2_, data_n_111__1_, data_n_111__0_ } : 
                              (N1640)? { data_n_110__31_, data_n_110__30_, data_n_110__29_, data_n_110__28_, data_n_110__27_, data_n_110__26_, data_n_110__25_, data_n_110__24_, data_n_110__23_, data_n_110__22_, data_n_110__21_, data_n_110__20_, data_n_110__19_, data_n_110__18_, data_n_110__17_, data_n_110__16_, data_n_110__15_, data_n_110__14_, data_n_110__13_, data_n_110__12_, data_n_110__11_, data_n_110__10_, data_n_110__9_, data_n_110__8_, data_n_110__7_, data_n_110__6_, data_n_110__5_, data_n_110__4_, data_n_110__3_, data_n_110__2_, data_n_110__1_, data_n_110__0_ } : 
                              (N1641)? { data_n_109__31_, data_n_109__30_, data_n_109__29_, data_n_109__28_, data_n_109__27_, data_n_109__26_, data_n_109__25_, data_n_109__24_, data_n_109__23_, data_n_109__22_, data_n_109__21_, data_n_109__20_, data_n_109__19_, data_n_109__18_, data_n_109__17_, data_n_109__16_, data_n_109__15_, data_n_109__14_, data_n_109__13_, data_n_109__12_, data_n_109__11_, data_n_109__10_, data_n_109__9_, data_n_109__8_, data_n_109__7_, data_n_109__6_, data_n_109__5_, data_n_109__4_, data_n_109__3_, data_n_109__2_, data_n_109__1_, data_n_109__0_ } : 
                              (N1642)? { data_n_108__31_, data_n_108__30_, data_n_108__29_, data_n_108__28_, data_n_108__27_, data_n_108__26_, data_n_108__25_, data_n_108__24_, data_n_108__23_, data_n_108__22_, data_n_108__21_, data_n_108__20_, data_n_108__19_, data_n_108__18_, data_n_108__17_, data_n_108__16_, data_n_108__15_, data_n_108__14_, data_n_108__13_, data_n_108__12_, data_n_108__11_, data_n_108__10_, data_n_108__9_, data_n_108__8_, data_n_108__7_, data_n_108__6_, data_n_108__5_, data_n_108__4_, data_n_108__3_, data_n_108__2_, data_n_108__1_, data_n_108__0_ } : 
                              (N1643)? { data_n_107__31_, data_n_107__30_, data_n_107__29_, data_n_107__28_, data_n_107__27_, data_n_107__26_, data_n_107__25_, data_n_107__24_, data_n_107__23_, data_n_107__22_, data_n_107__21_, data_n_107__20_, data_n_107__19_, data_n_107__18_, data_n_107__17_, data_n_107__16_, data_n_107__15_, data_n_107__14_, data_n_107__13_, data_n_107__12_, data_n_107__11_, data_n_107__10_, data_n_107__9_, data_n_107__8_, data_n_107__7_, data_n_107__6_, data_n_107__5_, data_n_107__4_, data_n_107__3_, data_n_107__2_, data_n_107__1_, data_n_107__0_ } : 
                              (N1644)? { data_n_106__31_, data_n_106__30_, data_n_106__29_, data_n_106__28_, data_n_106__27_, data_n_106__26_, data_n_106__25_, data_n_106__24_, data_n_106__23_, data_n_106__22_, data_n_106__21_, data_n_106__20_, data_n_106__19_, data_n_106__18_, data_n_106__17_, data_n_106__16_, data_n_106__15_, data_n_106__14_, data_n_106__13_, data_n_106__12_, data_n_106__11_, data_n_106__10_, data_n_106__9_, data_n_106__8_, data_n_106__7_, data_n_106__6_, data_n_106__5_, data_n_106__4_, data_n_106__3_, data_n_106__2_, data_n_106__1_, data_n_106__0_ } : 
                              (N1645)? { data_n_105__31_, data_n_105__30_, data_n_105__29_, data_n_105__28_, data_n_105__27_, data_n_105__26_, data_n_105__25_, data_n_105__24_, data_n_105__23_, data_n_105__22_, data_n_105__21_, data_n_105__20_, data_n_105__19_, data_n_105__18_, data_n_105__17_, data_n_105__16_, data_n_105__15_, data_n_105__14_, data_n_105__13_, data_n_105__12_, data_n_105__11_, data_n_105__10_, data_n_105__9_, data_n_105__8_, data_n_105__7_, data_n_105__6_, data_n_105__5_, data_n_105__4_, data_n_105__3_, data_n_105__2_, data_n_105__1_, data_n_105__0_ } : 
                              (N1646)? { data_n_104__31_, data_n_104__30_, data_n_104__29_, data_n_104__28_, data_n_104__27_, data_n_104__26_, data_n_104__25_, data_n_104__24_, data_n_104__23_, data_n_104__22_, data_n_104__21_, data_n_104__20_, data_n_104__19_, data_n_104__18_, data_n_104__17_, data_n_104__16_, data_n_104__15_, data_n_104__14_, data_n_104__13_, data_n_104__12_, data_n_104__11_, data_n_104__10_, data_n_104__9_, data_n_104__8_, data_n_104__7_, data_n_104__6_, data_n_104__5_, data_n_104__4_, data_n_104__3_, data_n_104__2_, data_n_104__1_, data_n_104__0_ } : 
                              (N1647)? { data_n_103__31_, data_n_103__30_, data_n_103__29_, data_n_103__28_, data_n_103__27_, data_n_103__26_, data_n_103__25_, data_n_103__24_, data_n_103__23_, data_n_103__22_, data_n_103__21_, data_n_103__20_, data_n_103__19_, data_n_103__18_, data_n_103__17_, data_n_103__16_, data_n_103__15_, data_n_103__14_, data_n_103__13_, data_n_103__12_, data_n_103__11_, data_n_103__10_, data_n_103__9_, data_n_103__8_, data_n_103__7_, data_n_103__6_, data_n_103__5_, data_n_103__4_, data_n_103__3_, data_n_103__2_, data_n_103__1_, data_n_103__0_ } : 
                              (N1648)? { data_n_102__31_, data_n_102__30_, data_n_102__29_, data_n_102__28_, data_n_102__27_, data_n_102__26_, data_n_102__25_, data_n_102__24_, data_n_102__23_, data_n_102__22_, data_n_102__21_, data_n_102__20_, data_n_102__19_, data_n_102__18_, data_n_102__17_, data_n_102__16_, data_n_102__15_, data_n_102__14_, data_n_102__13_, data_n_102__12_, data_n_102__11_, data_n_102__10_, data_n_102__9_, data_n_102__8_, data_n_102__7_, data_n_102__6_, data_n_102__5_, data_n_102__4_, data_n_102__3_, data_n_102__2_, data_n_102__1_, data_n_102__0_ } : 
                              (N1649)? { data_n_101__31_, data_n_101__30_, data_n_101__29_, data_n_101__28_, data_n_101__27_, data_n_101__26_, data_n_101__25_, data_n_101__24_, data_n_101__23_, data_n_101__22_, data_n_101__21_, data_n_101__20_, data_n_101__19_, data_n_101__18_, data_n_101__17_, data_n_101__16_, data_n_101__15_, data_n_101__14_, data_n_101__13_, data_n_101__12_, data_n_101__11_, data_n_101__10_, data_n_101__9_, data_n_101__8_, data_n_101__7_, data_n_101__6_, data_n_101__5_, data_n_101__4_, data_n_101__3_, data_n_101__2_, data_n_101__1_, data_n_101__0_ } : 
                              (N1650)? { data_n_100__31_, data_n_100__30_, data_n_100__29_, data_n_100__28_, data_n_100__27_, data_n_100__26_, data_n_100__25_, data_n_100__24_, data_n_100__23_, data_n_100__22_, data_n_100__21_, data_n_100__20_, data_n_100__19_, data_n_100__18_, data_n_100__17_, data_n_100__16_, data_n_100__15_, data_n_100__14_, data_n_100__13_, data_n_100__12_, data_n_100__11_, data_n_100__10_, data_n_100__9_, data_n_100__8_, data_n_100__7_, data_n_100__6_, data_n_100__5_, data_n_100__4_, data_n_100__3_, data_n_100__2_, data_n_100__1_, data_n_100__0_ } : 
                              (N1651)? { data_n_99__31_, data_n_99__30_, data_n_99__29_, data_n_99__28_, data_n_99__27_, data_n_99__26_, data_n_99__25_, data_n_99__24_, data_n_99__23_, data_n_99__22_, data_n_99__21_, data_n_99__20_, data_n_99__19_, data_n_99__18_, data_n_99__17_, data_n_99__16_, data_n_99__15_, data_n_99__14_, data_n_99__13_, data_n_99__12_, data_n_99__11_, data_n_99__10_, data_n_99__9_, data_n_99__8_, data_n_99__7_, data_n_99__6_, data_n_99__5_, data_n_99__4_, data_n_99__3_, data_n_99__2_, data_n_99__1_, data_n_99__0_ } : 
                              (N1652)? { data_n_98__31_, data_n_98__30_, data_n_98__29_, data_n_98__28_, data_n_98__27_, data_n_98__26_, data_n_98__25_, data_n_98__24_, data_n_98__23_, data_n_98__22_, data_n_98__21_, data_n_98__20_, data_n_98__19_, data_n_98__18_, data_n_98__17_, data_n_98__16_, data_n_98__15_, data_n_98__14_, data_n_98__13_, data_n_98__12_, data_n_98__11_, data_n_98__10_, data_n_98__9_, data_n_98__8_, data_n_98__7_, data_n_98__6_, data_n_98__5_, data_n_98__4_, data_n_98__3_, data_n_98__2_, data_n_98__1_, data_n_98__0_ } : 
                              (N1653)? { data_n_97__31_, data_n_97__30_, data_n_97__29_, data_n_97__28_, data_n_97__27_, data_n_97__26_, data_n_97__25_, data_n_97__24_, data_n_97__23_, data_n_97__22_, data_n_97__21_, data_n_97__20_, data_n_97__19_, data_n_97__18_, data_n_97__17_, data_n_97__16_, data_n_97__15_, data_n_97__14_, data_n_97__13_, data_n_97__12_, data_n_97__11_, data_n_97__10_, data_n_97__9_, data_n_97__8_, data_n_97__7_, data_n_97__6_, data_n_97__5_, data_n_97__4_, data_n_97__3_, data_n_97__2_, data_n_97__1_, data_n_97__0_ } : 
                              (N1654)? { data_n_96__31_, data_n_96__30_, data_n_96__29_, data_n_96__28_, data_n_96__27_, data_n_96__26_, data_n_96__25_, data_n_96__24_, data_n_96__23_, data_n_96__22_, data_n_96__21_, data_n_96__20_, data_n_96__19_, data_n_96__18_, data_n_96__17_, data_n_96__16_, data_n_96__15_, data_n_96__14_, data_n_96__13_, data_n_96__12_, data_n_96__11_, data_n_96__10_, data_n_96__9_, data_n_96__8_, data_n_96__7_, data_n_96__6_, data_n_96__5_, data_n_96__4_, data_n_96__3_, data_n_96__2_, data_n_96__1_, data_n_96__0_ } : 
                              (N1655)? { data_n_95__31_, data_n_95__30_, data_n_95__29_, data_n_95__28_, data_n_95__27_, data_n_95__26_, data_n_95__25_, data_n_95__24_, data_n_95__23_, data_n_95__22_, data_n_95__21_, data_n_95__20_, data_n_95__19_, data_n_95__18_, data_n_95__17_, data_n_95__16_, data_n_95__15_, data_n_95__14_, data_n_95__13_, data_n_95__12_, data_n_95__11_, data_n_95__10_, data_n_95__9_, data_n_95__8_, data_n_95__7_, data_n_95__6_, data_n_95__5_, data_n_95__4_, data_n_95__3_, data_n_95__2_, data_n_95__1_, data_n_95__0_ } : 
                              (N1656)? { data_n_94__31_, data_n_94__30_, data_n_94__29_, data_n_94__28_, data_n_94__27_, data_n_94__26_, data_n_94__25_, data_n_94__24_, data_n_94__23_, data_n_94__22_, data_n_94__21_, data_n_94__20_, data_n_94__19_, data_n_94__18_, data_n_94__17_, data_n_94__16_, data_n_94__15_, data_n_94__14_, data_n_94__13_, data_n_94__12_, data_n_94__11_, data_n_94__10_, data_n_94__9_, data_n_94__8_, data_n_94__7_, data_n_94__6_, data_n_94__5_, data_n_94__4_, data_n_94__3_, data_n_94__2_, data_n_94__1_, data_n_94__0_ } : 
                              (N1657)? { data_n_93__31_, data_n_93__30_, data_n_93__29_, data_n_93__28_, data_n_93__27_, data_n_93__26_, data_n_93__25_, data_n_93__24_, data_n_93__23_, data_n_93__22_, data_n_93__21_, data_n_93__20_, data_n_93__19_, data_n_93__18_, data_n_93__17_, data_n_93__16_, data_n_93__15_, data_n_93__14_, data_n_93__13_, data_n_93__12_, data_n_93__11_, data_n_93__10_, data_n_93__9_, data_n_93__8_, data_n_93__7_, data_n_93__6_, data_n_93__5_, data_n_93__4_, data_n_93__3_, data_n_93__2_, data_n_93__1_, data_n_93__0_ } : 
                              (N1658)? { data_n_92__31_, data_n_92__30_, data_n_92__29_, data_n_92__28_, data_n_92__27_, data_n_92__26_, data_n_92__25_, data_n_92__24_, data_n_92__23_, data_n_92__22_, data_n_92__21_, data_n_92__20_, data_n_92__19_, data_n_92__18_, data_n_92__17_, data_n_92__16_, data_n_92__15_, data_n_92__14_, data_n_92__13_, data_n_92__12_, data_n_92__11_, data_n_92__10_, data_n_92__9_, data_n_92__8_, data_n_92__7_, data_n_92__6_, data_n_92__5_, data_n_92__4_, data_n_92__3_, data_n_92__2_, data_n_92__1_, data_n_92__0_ } : 
                              (N1659)? { data_n_91__31_, data_n_91__30_, data_n_91__29_, data_n_91__28_, data_n_91__27_, data_n_91__26_, data_n_91__25_, data_n_91__24_, data_n_91__23_, data_n_91__22_, data_n_91__21_, data_n_91__20_, data_n_91__19_, data_n_91__18_, data_n_91__17_, data_n_91__16_, data_n_91__15_, data_n_91__14_, data_n_91__13_, data_n_91__12_, data_n_91__11_, data_n_91__10_, data_n_91__9_, data_n_91__8_, data_n_91__7_, data_n_91__6_, data_n_91__5_, data_n_91__4_, data_n_91__3_, data_n_91__2_, data_n_91__1_, data_n_91__0_ } : 
                              (N1660)? { data_n_90__31_, data_n_90__30_, data_n_90__29_, data_n_90__28_, data_n_90__27_, data_n_90__26_, data_n_90__25_, data_n_90__24_, data_n_90__23_, data_n_90__22_, data_n_90__21_, data_n_90__20_, data_n_90__19_, data_n_90__18_, data_n_90__17_, data_n_90__16_, data_n_90__15_, data_n_90__14_, data_n_90__13_, data_n_90__12_, data_n_90__11_, data_n_90__10_, data_n_90__9_, data_n_90__8_, data_n_90__7_, data_n_90__6_, data_n_90__5_, data_n_90__4_, data_n_90__3_, data_n_90__2_, data_n_90__1_, data_n_90__0_ } : 
                              (N1661)? { data_n_89__31_, data_n_89__30_, data_n_89__29_, data_n_89__28_, data_n_89__27_, data_n_89__26_, data_n_89__25_, data_n_89__24_, data_n_89__23_, data_n_89__22_, data_n_89__21_, data_n_89__20_, data_n_89__19_, data_n_89__18_, data_n_89__17_, data_n_89__16_, data_n_89__15_, data_n_89__14_, data_n_89__13_, data_n_89__12_, data_n_89__11_, data_n_89__10_, data_n_89__9_, data_n_89__8_, data_n_89__7_, data_n_89__6_, data_n_89__5_, data_n_89__4_, data_n_89__3_, data_n_89__2_, data_n_89__1_, data_n_89__0_ } : 
                              (N1662)? { data_n_88__31_, data_n_88__30_, data_n_88__29_, data_n_88__28_, data_n_88__27_, data_n_88__26_, data_n_88__25_, data_n_88__24_, data_n_88__23_, data_n_88__22_, data_n_88__21_, data_n_88__20_, data_n_88__19_, data_n_88__18_, data_n_88__17_, data_n_88__16_, data_n_88__15_, data_n_88__14_, data_n_88__13_, data_n_88__12_, data_n_88__11_, data_n_88__10_, data_n_88__9_, data_n_88__8_, data_n_88__7_, data_n_88__6_, data_n_88__5_, data_n_88__4_, data_n_88__3_, data_n_88__2_, data_n_88__1_, data_n_88__0_ } : 
                              (N1663)? { data_n_87__31_, data_n_87__30_, data_n_87__29_, data_n_87__28_, data_n_87__27_, data_n_87__26_, data_n_87__25_, data_n_87__24_, data_n_87__23_, data_n_87__22_, data_n_87__21_, data_n_87__20_, data_n_87__19_, data_n_87__18_, data_n_87__17_, data_n_87__16_, data_n_87__15_, data_n_87__14_, data_n_87__13_, data_n_87__12_, data_n_87__11_, data_n_87__10_, data_n_87__9_, data_n_87__8_, data_n_87__7_, data_n_87__6_, data_n_87__5_, data_n_87__4_, data_n_87__3_, data_n_87__2_, data_n_87__1_, data_n_87__0_ } : 
                              (N1664)? { data_n_86__31_, data_n_86__30_, data_n_86__29_, data_n_86__28_, data_n_86__27_, data_n_86__26_, data_n_86__25_, data_n_86__24_, data_n_86__23_, data_n_86__22_, data_n_86__21_, data_n_86__20_, data_n_86__19_, data_n_86__18_, data_n_86__17_, data_n_86__16_, data_n_86__15_, data_n_86__14_, data_n_86__13_, data_n_86__12_, data_n_86__11_, data_n_86__10_, data_n_86__9_, data_n_86__8_, data_n_86__7_, data_n_86__6_, data_n_86__5_, data_n_86__4_, data_n_86__3_, data_n_86__2_, data_n_86__1_, data_n_86__0_ } : 
                              (N1665)? { data_n_85__31_, data_n_85__30_, data_n_85__29_, data_n_85__28_, data_n_85__27_, data_n_85__26_, data_n_85__25_, data_n_85__24_, data_n_85__23_, data_n_85__22_, data_n_85__21_, data_n_85__20_, data_n_85__19_, data_n_85__18_, data_n_85__17_, data_n_85__16_, data_n_85__15_, data_n_85__14_, data_n_85__13_, data_n_85__12_, data_n_85__11_, data_n_85__10_, data_n_85__9_, data_n_85__8_, data_n_85__7_, data_n_85__6_, data_n_85__5_, data_n_85__4_, data_n_85__3_, data_n_85__2_, data_n_85__1_, data_n_85__0_ } : 
                              (N1666)? { data_n_84__31_, data_n_84__30_, data_n_84__29_, data_n_84__28_, data_n_84__27_, data_n_84__26_, data_n_84__25_, data_n_84__24_, data_n_84__23_, data_n_84__22_, data_n_84__21_, data_n_84__20_, data_n_84__19_, data_n_84__18_, data_n_84__17_, data_n_84__16_, data_n_84__15_, data_n_84__14_, data_n_84__13_, data_n_84__12_, data_n_84__11_, data_n_84__10_, data_n_84__9_, data_n_84__8_, data_n_84__7_, data_n_84__6_, data_n_84__5_, data_n_84__4_, data_n_84__3_, data_n_84__2_, data_n_84__1_, data_n_84__0_ } : 
                              (N1667)? { data_n_83__31_, data_n_83__30_, data_n_83__29_, data_n_83__28_, data_n_83__27_, data_n_83__26_, data_n_83__25_, data_n_83__24_, data_n_83__23_, data_n_83__22_, data_n_83__21_, data_n_83__20_, data_n_83__19_, data_n_83__18_, data_n_83__17_, data_n_83__16_, data_n_83__15_, data_n_83__14_, data_n_83__13_, data_n_83__12_, data_n_83__11_, data_n_83__10_, data_n_83__9_, data_n_83__8_, data_n_83__7_, data_n_83__6_, data_n_83__5_, data_n_83__4_, data_n_83__3_, data_n_83__2_, data_n_83__1_, data_n_83__0_ } : 
                              (N1668)? { data_n_82__31_, data_n_82__30_, data_n_82__29_, data_n_82__28_, data_n_82__27_, data_n_82__26_, data_n_82__25_, data_n_82__24_, data_n_82__23_, data_n_82__22_, data_n_82__21_, data_n_82__20_, data_n_82__19_, data_n_82__18_, data_n_82__17_, data_n_82__16_, data_n_82__15_, data_n_82__14_, data_n_82__13_, data_n_82__12_, data_n_82__11_, data_n_82__10_, data_n_82__9_, data_n_82__8_, data_n_82__7_, data_n_82__6_, data_n_82__5_, data_n_82__4_, data_n_82__3_, data_n_82__2_, data_n_82__1_, data_n_82__0_ } : 
                              (N1669)? { data_n_81__31_, data_n_81__30_, data_n_81__29_, data_n_81__28_, data_n_81__27_, data_n_81__26_, data_n_81__25_, data_n_81__24_, data_n_81__23_, data_n_81__22_, data_n_81__21_, data_n_81__20_, data_n_81__19_, data_n_81__18_, data_n_81__17_, data_n_81__16_, data_n_81__15_, data_n_81__14_, data_n_81__13_, data_n_81__12_, data_n_81__11_, data_n_81__10_, data_n_81__9_, data_n_81__8_, data_n_81__7_, data_n_81__6_, data_n_81__5_, data_n_81__4_, data_n_81__3_, data_n_81__2_, data_n_81__1_, data_n_81__0_ } : 
                              (N1670)? { data_n_80__31_, data_n_80__30_, data_n_80__29_, data_n_80__28_, data_n_80__27_, data_n_80__26_, data_n_80__25_, data_n_80__24_, data_n_80__23_, data_n_80__22_, data_n_80__21_, data_n_80__20_, data_n_80__19_, data_n_80__18_, data_n_80__17_, data_n_80__16_, data_n_80__15_, data_n_80__14_, data_n_80__13_, data_n_80__12_, data_n_80__11_, data_n_80__10_, data_n_80__9_, data_n_80__8_, data_n_80__7_, data_n_80__6_, data_n_80__5_, data_n_80__4_, data_n_80__3_, data_n_80__2_, data_n_80__1_, data_n_80__0_ } : 
                              (N1671)? { data_n_79__31_, data_n_79__30_, data_n_79__29_, data_n_79__28_, data_n_79__27_, data_n_79__26_, data_n_79__25_, data_n_79__24_, data_n_79__23_, data_n_79__22_, data_n_79__21_, data_n_79__20_, data_n_79__19_, data_n_79__18_, data_n_79__17_, data_n_79__16_, data_n_79__15_, data_n_79__14_, data_n_79__13_, data_n_79__12_, data_n_79__11_, data_n_79__10_, data_n_79__9_, data_n_79__8_, data_n_79__7_, data_n_79__6_, data_n_79__5_, data_n_79__4_, data_n_79__3_, data_n_79__2_, data_n_79__1_, data_n_79__0_ } : 
                              (N1672)? { data_n_78__31_, data_n_78__30_, data_n_78__29_, data_n_78__28_, data_n_78__27_, data_n_78__26_, data_n_78__25_, data_n_78__24_, data_n_78__23_, data_n_78__22_, data_n_78__21_, data_n_78__20_, data_n_78__19_, data_n_78__18_, data_n_78__17_, data_n_78__16_, data_n_78__15_, data_n_78__14_, data_n_78__13_, data_n_78__12_, data_n_78__11_, data_n_78__10_, data_n_78__9_, data_n_78__8_, data_n_78__7_, data_n_78__6_, data_n_78__5_, data_n_78__4_, data_n_78__3_, data_n_78__2_, data_n_78__1_, data_n_78__0_ } : 
                              (N1673)? { data_n_77__31_, data_n_77__30_, data_n_77__29_, data_n_77__28_, data_n_77__27_, data_n_77__26_, data_n_77__25_, data_n_77__24_, data_n_77__23_, data_n_77__22_, data_n_77__21_, data_n_77__20_, data_n_77__19_, data_n_77__18_, data_n_77__17_, data_n_77__16_, data_n_77__15_, data_n_77__14_, data_n_77__13_, data_n_77__12_, data_n_77__11_, data_n_77__10_, data_n_77__9_, data_n_77__8_, data_n_77__7_, data_n_77__6_, data_n_77__5_, data_n_77__4_, data_n_77__3_, data_n_77__2_, data_n_77__1_, data_n_77__0_ } : 
                              (N1674)? { data_n_76__31_, data_n_76__30_, data_n_76__29_, data_n_76__28_, data_n_76__27_, data_n_76__26_, data_n_76__25_, data_n_76__24_, data_n_76__23_, data_n_76__22_, data_n_76__21_, data_n_76__20_, data_n_76__19_, data_n_76__18_, data_n_76__17_, data_n_76__16_, data_n_76__15_, data_n_76__14_, data_n_76__13_, data_n_76__12_, data_n_76__11_, data_n_76__10_, data_n_76__9_, data_n_76__8_, data_n_76__7_, data_n_76__6_, data_n_76__5_, data_n_76__4_, data_n_76__3_, data_n_76__2_, data_n_76__1_, data_n_76__0_ } : 
                              (N1675)? { data_n_75__31_, data_n_75__30_, data_n_75__29_, data_n_75__28_, data_n_75__27_, data_n_75__26_, data_n_75__25_, data_n_75__24_, data_n_75__23_, data_n_75__22_, data_n_75__21_, data_n_75__20_, data_n_75__19_, data_n_75__18_, data_n_75__17_, data_n_75__16_, data_n_75__15_, data_n_75__14_, data_n_75__13_, data_n_75__12_, data_n_75__11_, data_n_75__10_, data_n_75__9_, data_n_75__8_, data_n_75__7_, data_n_75__6_, data_n_75__5_, data_n_75__4_, data_n_75__3_, data_n_75__2_, data_n_75__1_, data_n_75__0_ } : 
                              (N1676)? { data_n_74__31_, data_n_74__30_, data_n_74__29_, data_n_74__28_, data_n_74__27_, data_n_74__26_, data_n_74__25_, data_n_74__24_, data_n_74__23_, data_n_74__22_, data_n_74__21_, data_n_74__20_, data_n_74__19_, data_n_74__18_, data_n_74__17_, data_n_74__16_, data_n_74__15_, data_n_74__14_, data_n_74__13_, data_n_74__12_, data_n_74__11_, data_n_74__10_, data_n_74__9_, data_n_74__8_, data_n_74__7_, data_n_74__6_, data_n_74__5_, data_n_74__4_, data_n_74__3_, data_n_74__2_, data_n_74__1_, data_n_74__0_ } : 
                              (N1677)? { data_n_73__31_, data_n_73__30_, data_n_73__29_, data_n_73__28_, data_n_73__27_, data_n_73__26_, data_n_73__25_, data_n_73__24_, data_n_73__23_, data_n_73__22_, data_n_73__21_, data_n_73__20_, data_n_73__19_, data_n_73__18_, data_n_73__17_, data_n_73__16_, data_n_73__15_, data_n_73__14_, data_n_73__13_, data_n_73__12_, data_n_73__11_, data_n_73__10_, data_n_73__9_, data_n_73__8_, data_n_73__7_, data_n_73__6_, data_n_73__5_, data_n_73__4_, data_n_73__3_, data_n_73__2_, data_n_73__1_, data_n_73__0_ } : 
                              (N1678)? { data_n_72__31_, data_n_72__30_, data_n_72__29_, data_n_72__28_, data_n_72__27_, data_n_72__26_, data_n_72__25_, data_n_72__24_, data_n_72__23_, data_n_72__22_, data_n_72__21_, data_n_72__20_, data_n_72__19_, data_n_72__18_, data_n_72__17_, data_n_72__16_, data_n_72__15_, data_n_72__14_, data_n_72__13_, data_n_72__12_, data_n_72__11_, data_n_72__10_, data_n_72__9_, data_n_72__8_, data_n_72__7_, data_n_72__6_, data_n_72__5_, data_n_72__4_, data_n_72__3_, data_n_72__2_, data_n_72__1_, data_n_72__0_ } : 
                              (N1679)? { data_n_71__31_, data_n_71__30_, data_n_71__29_, data_n_71__28_, data_n_71__27_, data_n_71__26_, data_n_71__25_, data_n_71__24_, data_n_71__23_, data_n_71__22_, data_n_71__21_, data_n_71__20_, data_n_71__19_, data_n_71__18_, data_n_71__17_, data_n_71__16_, data_n_71__15_, data_n_71__14_, data_n_71__13_, data_n_71__12_, data_n_71__11_, data_n_71__10_, data_n_71__9_, data_n_71__8_, data_n_71__7_, data_n_71__6_, data_n_71__5_, data_n_71__4_, data_n_71__3_, data_n_71__2_, data_n_71__1_, data_n_71__0_ } : 
                              (N1680)? { data_n_70__31_, data_n_70__30_, data_n_70__29_, data_n_70__28_, data_n_70__27_, data_n_70__26_, data_n_70__25_, data_n_70__24_, data_n_70__23_, data_n_70__22_, data_n_70__21_, data_n_70__20_, data_n_70__19_, data_n_70__18_, data_n_70__17_, data_n_70__16_, data_n_70__15_, data_n_70__14_, data_n_70__13_, data_n_70__12_, data_n_70__11_, data_n_70__10_, data_n_70__9_, data_n_70__8_, data_n_70__7_, data_n_70__6_, data_n_70__5_, data_n_70__4_, data_n_70__3_, data_n_70__2_, data_n_70__1_, data_n_70__0_ } : 
                              (N1681)? { data_n_69__31_, data_n_69__30_, data_n_69__29_, data_n_69__28_, data_n_69__27_, data_n_69__26_, data_n_69__25_, data_n_69__24_, data_n_69__23_, data_n_69__22_, data_n_69__21_, data_n_69__20_, data_n_69__19_, data_n_69__18_, data_n_69__17_, data_n_69__16_, data_n_69__15_, data_n_69__14_, data_n_69__13_, data_n_69__12_, data_n_69__11_, data_n_69__10_, data_n_69__9_, data_n_69__8_, data_n_69__7_, data_n_69__6_, data_n_69__5_, data_n_69__4_, data_n_69__3_, data_n_69__2_, data_n_69__1_, data_n_69__0_ } : 
                              (N1682)? { data_n_68__31_, data_n_68__30_, data_n_68__29_, data_n_68__28_, data_n_68__27_, data_n_68__26_, data_n_68__25_, data_n_68__24_, data_n_68__23_, data_n_68__22_, data_n_68__21_, data_n_68__20_, data_n_68__19_, data_n_68__18_, data_n_68__17_, data_n_68__16_, data_n_68__15_, data_n_68__14_, data_n_68__13_, data_n_68__12_, data_n_68__11_, data_n_68__10_, data_n_68__9_, data_n_68__8_, data_n_68__7_, data_n_68__6_, data_n_68__5_, data_n_68__4_, data_n_68__3_, data_n_68__2_, data_n_68__1_, data_n_68__0_ } : 
                              (N1683)? { data_n_67__31_, data_n_67__30_, data_n_67__29_, data_n_67__28_, data_n_67__27_, data_n_67__26_, data_n_67__25_, data_n_67__24_, data_n_67__23_, data_n_67__22_, data_n_67__21_, data_n_67__20_, data_n_67__19_, data_n_67__18_, data_n_67__17_, data_n_67__16_, data_n_67__15_, data_n_67__14_, data_n_67__13_, data_n_67__12_, data_n_67__11_, data_n_67__10_, data_n_67__9_, data_n_67__8_, data_n_67__7_, data_n_67__6_, data_n_67__5_, data_n_67__4_, data_n_67__3_, data_n_67__2_, data_n_67__1_, data_n_67__0_ } : 
                              (N1684)? { data_n_66__31_, data_n_66__30_, data_n_66__29_, data_n_66__28_, data_n_66__27_, data_n_66__26_, data_n_66__25_, data_n_66__24_, data_n_66__23_, data_n_66__22_, data_n_66__21_, data_n_66__20_, data_n_66__19_, data_n_66__18_, data_n_66__17_, data_n_66__16_, data_n_66__15_, data_n_66__14_, data_n_66__13_, data_n_66__12_, data_n_66__11_, data_n_66__10_, data_n_66__9_, data_n_66__8_, data_n_66__7_, data_n_66__6_, data_n_66__5_, data_n_66__4_, data_n_66__3_, data_n_66__2_, data_n_66__1_, data_n_66__0_ } : 
                              (N1685)? { data_n_65__31_, data_n_65__30_, data_n_65__29_, data_n_65__28_, data_n_65__27_, data_n_65__26_, data_n_65__25_, data_n_65__24_, data_n_65__23_, data_n_65__22_, data_n_65__21_, data_n_65__20_, data_n_65__19_, data_n_65__18_, data_n_65__17_, data_n_65__16_, data_n_65__15_, data_n_65__14_, data_n_65__13_, data_n_65__12_, data_n_65__11_, data_n_65__10_, data_n_65__9_, data_n_65__8_, data_n_65__7_, data_n_65__6_, data_n_65__5_, data_n_65__4_, data_n_65__3_, data_n_65__2_, data_n_65__1_, data_n_65__0_ } : 
                              (N1686)? { data_n_64__31_, data_n_64__30_, data_n_64__29_, data_n_64__28_, data_n_64__27_, data_n_64__26_, data_n_64__25_, data_n_64__24_, data_n_64__23_, data_n_64__22_, data_n_64__21_, data_n_64__20_, data_n_64__19_, data_n_64__18_, data_n_64__17_, data_n_64__16_, data_n_64__15_, data_n_64__14_, data_n_64__13_, data_n_64__12_, data_n_64__11_, data_n_64__10_, data_n_64__9_, data_n_64__8_, data_n_64__7_, data_n_64__6_, data_n_64__5_, data_n_64__4_, data_n_64__3_, data_n_64__2_, data_n_64__1_, data_n_64__0_ } : 
                              (N1687)? data_o[2047:2016] : 1'b0;
  assign N2222 = N4871;
  assign { N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872 } = (N2223)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, valid_n } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       (N2881)? { valid_n[126:64], valid_o } : 1'b0;
  assign N2223 = yumi_cnt_i[6];
  assign { N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999 } = (N2224)? { N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       (N2816)? { N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872 } : 1'b0;
  assign N2224 = yumi_cnt_i[5];
  assign { N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094 } = (N2225)? { N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       (N2783)? { N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999 } : 1'b0;
  assign N2225 = yumi_cnt_i[4];
  assign { N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173 } = (N2226)? { N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               (N2766)? { N5164, N5163, N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094 } : 1'b0;
  assign N2226 = yumi_cnt_i[3];
  assign { N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244 } = (N2227)? { N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (N2757)? { N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173 } : 1'b0;
  assign N2227 = yumi_cnt_i[2];
  assign { N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311 } = (N2228)? { N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N2752)? { N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244 } : 1'b0;
  assign N2228 = yumi_cnt_i[1];
  assign valid_nn = (N2229)? { N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312 } : 
                    (N2751)? { N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311 } : 1'b0;
  assign N2229 = yumi_cnt_i[0];
  assign ready_o = ~valid_r[63];
  assign N2230 = valid_i & ready_o;
  assign N2366 = ~N2238;
  assign N2367 = ~N2239;
  assign N2368 = ~N2240;
  assign N2369 = ~N2241;
  assign N2370 = ~N2242;
  assign N2371 = ~N2243;
  assign N2372 = ~N2244;
  assign N2373 = ~N2245;
  assign N2374 = ~N2246;
  assign N2375 = ~N2247;
  assign N2376 = ~N2248;
  assign N2377 = ~N2249;
  assign N2378 = ~N2250;
  assign N2379 = ~N2251;
  assign N2380 = ~N2252;
  assign N2381 = ~N2253;
  assign N2382 = ~N2254;
  assign N2383 = ~N2255;
  assign N2384 = ~N2256;
  assign N2385 = ~N2257;
  assign N2386 = ~N2258;
  assign N2387 = ~N2259;
  assign N2388 = ~N2260;
  assign N2389 = ~N2261;
  assign N2390 = ~N2262;
  assign N2391 = ~N2263;
  assign N2392 = ~N2264;
  assign N2393 = ~N2265;
  assign N2394 = ~N2266;
  assign N2395 = ~N2267;
  assign N2396 = ~N2268;
  assign N2397 = ~N2269;
  assign N2398 = ~N2270;
  assign N2399 = ~N2271;
  assign N2400 = ~N2272;
  assign N2401 = ~N2273;
  assign N2402 = ~N2274;
  assign N2403 = ~N2275;
  assign N2404 = ~N2276;
  assign N2405 = ~N2277;
  assign N2406 = ~N2278;
  assign N2407 = ~N2279;
  assign N2408 = ~N2280;
  assign N2409 = ~N2281;
  assign N2410 = ~N2282;
  assign N2411 = ~N2283;
  assign N2412 = ~N2284;
  assign N2413 = ~N2285;
  assign N2414 = ~N2286;
  assign N2415 = ~N2287;
  assign N2416 = ~N2288;
  assign N2417 = ~N2289;
  assign N2418 = ~N2290;
  assign N2419 = ~N2291;
  assign N2420 = ~N2292;
  assign N2421 = ~N2293;
  assign N2422 = ~N2294;
  assign N2423 = ~N2295;
  assign N2424 = ~N2296;
  assign N2425 = ~N2297;
  assign N2426 = ~N2298;
  assign N2427 = ~N2299;
  assign N2428 = ~N2300;
  assign N2429 = ~N2301;
  assign N2430 = ~N2302;
  assign N2431 = ~N2303;
  assign N2432 = ~N2304;
  assign N2433 = ~N2305;
  assign N2434 = ~N2306;
  assign N2435 = ~N2307;
  assign N2436 = ~N2308;
  assign N2437 = ~N2309;
  assign N2438 = ~N2310;
  assign N2439 = ~N2311;
  assign N2440 = ~N2312;
  assign N2441 = ~N2313;
  assign N2442 = ~N2314;
  assign N2443 = ~N2315;
  assign N2444 = ~N2316;
  assign N2445 = ~N2317;
  assign N2446 = ~N2318;
  assign N2447 = ~N2319;
  assign N2448 = ~N2320;
  assign N2449 = ~N2321;
  assign N2450 = ~N2322;
  assign N2451 = ~N2323;
  assign N2452 = ~N2324;
  assign N2453 = ~N2325;
  assign N2454 = ~N2326;
  assign N2455 = ~N2327;
  assign N2456 = ~N2328;
  assign N2457 = ~N2329;
  assign N2458 = ~N2330;
  assign N2459 = ~N2331;
  assign N2460 = ~N2332;
  assign N2461 = ~N2333;
  assign N2462 = ~N2334;
  assign N2463 = ~N2335;
  assign N2464 = ~N2336;
  assign N2465 = ~N2337;
  assign N2466 = ~N2338;
  assign N2467 = ~N2339;
  assign N2468 = ~N2340;
  assign N2469 = ~N2341;
  assign N2470 = ~N2342;
  assign N2471 = ~N2343;
  assign N2472 = ~N2344;
  assign N2473 = ~N2345;
  assign N2474 = ~N2346;
  assign N2475 = ~N2347;
  assign N2476 = ~N2348;
  assign N2477 = ~N2349;
  assign N2478 = ~N2350;
  assign N2479 = ~N2351;
  assign N2480 = ~N2352;
  assign N2481 = ~N2353;
  assign N2482 = ~N2354;
  assign N2483 = ~N2355;
  assign N2484 = ~N2356;
  assign N2485 = ~N2357;
  assign N2486 = ~N2358;
  assign N2487 = ~N2359;
  assign N2488 = ~N2360;
  assign N2489 = ~N2361;
  assign N2490 = ~N2362;
  assign N2491 = ~N2363;
  assign N2492 = ~N2364;
  assign N2493 = ~N2365;
  assign N2622 = valid_i & ready_o;
  assign N2623 = ~N2494;
  assign N2624 = ~N2495;
  assign N2625 = ~N2496;
  assign N2626 = ~N2497;
  assign N2627 = ~N2498;
  assign N2628 = ~N2499;
  assign N2629 = ~N2500;
  assign N2630 = ~N2501;
  assign N2631 = ~N2502;
  assign N2632 = ~N2503;
  assign N2633 = ~N2504;
  assign N2634 = ~N2505;
  assign N2635 = ~N2506;
  assign N2636 = ~N2507;
  assign N2637 = ~N2508;
  assign N2638 = ~N2509;
  assign N2639 = ~N2510;
  assign N2640 = ~N2511;
  assign N2641 = ~N2512;
  assign N2642 = ~N2513;
  assign N2643 = ~N2514;
  assign N2644 = ~N2515;
  assign N2645 = ~N2516;
  assign N2646 = ~N2517;
  assign N2647 = ~N2518;
  assign N2648 = ~N2519;
  assign N2649 = ~N2520;
  assign N2650 = ~N2521;
  assign N2651 = ~N2522;
  assign N2652 = ~N2523;
  assign N2653 = ~N2524;
  assign N2654 = ~N2525;
  assign N2655 = ~N2526;
  assign N2656 = ~N2527;
  assign N2657 = ~N2528;
  assign N2658 = ~N2529;
  assign N2659 = ~N2530;
  assign N2660 = ~N2531;
  assign N2661 = ~N2532;
  assign N2662 = ~N2533;
  assign N2663 = ~N2534;
  assign N2664 = ~N2535;
  assign N2665 = ~N2536;
  assign N2666 = ~N2537;
  assign N2667 = ~N2538;
  assign N2668 = ~N2539;
  assign N2669 = ~N2540;
  assign N2670 = ~N2541;
  assign N2671 = ~N2542;
  assign N2672 = ~N2543;
  assign N2673 = ~N2544;
  assign N2674 = ~N2545;
  assign N2675 = ~N2546;
  assign N2676 = ~N2547;
  assign N2677 = ~N2548;
  assign N2678 = ~N2549;
  assign N2679 = ~N2550;
  assign N2680 = ~N2551;
  assign N2681 = ~N2552;
  assign N2682 = ~N2553;
  assign N2683 = ~N2554;
  assign N2684 = ~N2555;
  assign N2685 = ~N2556;
  assign N2686 = ~N2557;
  assign N2687 = ~N2558;
  assign N2688 = ~N2559;
  assign N2689 = ~N2560;
  assign N2690 = ~N2561;
  assign N2691 = ~N2562;
  assign N2692 = ~N2563;
  assign N2693 = ~N2564;
  assign N2694 = ~N2565;
  assign N2695 = ~N2566;
  assign N2696 = ~N2567;
  assign N2697 = ~N2568;
  assign N2698 = ~N2569;
  assign N2699 = ~N2570;
  assign N2700 = ~N2571;
  assign N2701 = ~N2572;
  assign N2702 = ~N2573;
  assign N2703 = ~N2574;
  assign N2704 = ~N2575;
  assign N2705 = ~N2576;
  assign N2706 = ~N2577;
  assign N2707 = ~N2578;
  assign N2708 = ~N2579;
  assign N2709 = ~N2580;
  assign N2710 = ~N2581;
  assign N2711 = ~N2582;
  assign N2712 = ~N2583;
  assign N2713 = ~N2584;
  assign N2714 = ~N2585;
  assign N2715 = ~N2586;
  assign N2716 = ~N2587;
  assign N2717 = ~N2588;
  assign N2718 = ~N2589;
  assign N2719 = ~N2590;
  assign N2720 = ~N2591;
  assign N2721 = ~N2592;
  assign N2722 = ~N2593;
  assign N2723 = ~N2594;
  assign N2724 = ~N2595;
  assign N2725 = ~N2596;
  assign N2726 = ~N2597;
  assign N2727 = ~N2598;
  assign N2728 = ~N2599;
  assign N2729 = ~N2600;
  assign N2730 = ~N2601;
  assign N2731 = ~N2602;
  assign N2732 = ~N2603;
  assign N2733 = ~N2604;
  assign N2734 = ~N2605;
  assign N2735 = ~N2606;
  assign N2736 = ~N2607;
  assign N2737 = ~N2608;
  assign N2738 = ~N2609;
  assign N2739 = ~N2610;
  assign N2740 = ~N2611;
  assign N2741 = ~N2612;
  assign N2742 = ~N2613;
  assign N2743 = ~N2614;
  assign N2744 = ~N2615;
  assign N2745 = ~N2616;
  assign N2746 = ~N2617;
  assign N2747 = ~N2618;
  assign N2748 = ~N2619;
  assign N2749 = ~N2620;
  assign N2750 = ~N2621;
  assign N2751 = ~yumi_cnt_i[0];
  assign N2752 = ~yumi_cnt_i[1];
  assign N2753 = N2751 & N2752;
  assign N2754 = N2751 & yumi_cnt_i[1];
  assign N2755 = yumi_cnt_i[0] & N2752;
  assign N2756 = yumi_cnt_i[0] & yumi_cnt_i[1];
  assign N2757 = ~yumi_cnt_i[2];
  assign N2758 = N2753 & N2757;
  assign N2759 = N2753 & yumi_cnt_i[2];
  assign N2760 = N2755 & N2757;
  assign N2761 = N2755 & yumi_cnt_i[2];
  assign N2762 = N2754 & N2757;
  assign N2763 = N2754 & yumi_cnt_i[2];
  assign N2764 = N2756 & N2757;
  assign N2765 = N2756 & yumi_cnt_i[2];
  assign N2766 = ~yumi_cnt_i[3];
  assign N2767 = N2758 & N2766;
  assign N2768 = N2758 & yumi_cnt_i[3];
  assign N2769 = N2760 & N2766;
  assign N2770 = N2760 & yumi_cnt_i[3];
  assign N2771 = N2762 & N2766;
  assign N2772 = N2762 & yumi_cnt_i[3];
  assign N2773 = N2764 & N2766;
  assign N2774 = N2764 & yumi_cnt_i[3];
  assign N2775 = N2759 & N2766;
  assign N2776 = N2759 & yumi_cnt_i[3];
  assign N2777 = N2761 & N2766;
  assign N2778 = N2761 & yumi_cnt_i[3];
  assign N2779 = N2763 & N2766;
  assign N2780 = N2763 & yumi_cnt_i[3];
  assign N2781 = N2765 & N2766;
  assign N2782 = N2765 & yumi_cnt_i[3];
  assign N2783 = ~yumi_cnt_i[4];
  assign N2784 = N2767 & N2783;
  assign N2785 = N2767 & yumi_cnt_i[4];
  assign N2786 = N2769 & N2783;
  assign N2787 = N2769 & yumi_cnt_i[4];
  assign N2788 = N2771 & N2783;
  assign N2789 = N2771 & yumi_cnt_i[4];
  assign N2790 = N2773 & N2783;
  assign N2791 = N2773 & yumi_cnt_i[4];
  assign N2792 = N2775 & N2783;
  assign N2793 = N2775 & yumi_cnt_i[4];
  assign N2794 = N2777 & N2783;
  assign N2795 = N2777 & yumi_cnt_i[4];
  assign N2796 = N2779 & N2783;
  assign N2797 = N2779 & yumi_cnt_i[4];
  assign N2798 = N2781 & N2783;
  assign N2799 = N2781 & yumi_cnt_i[4];
  assign N2800 = N2768 & N2783;
  assign N2801 = N2768 & yumi_cnt_i[4];
  assign N2802 = N2770 & N2783;
  assign N2803 = N2770 & yumi_cnt_i[4];
  assign N2804 = N2772 & N2783;
  assign N2805 = N2772 & yumi_cnt_i[4];
  assign N2806 = N2774 & N2783;
  assign N2807 = N2774 & yumi_cnt_i[4];
  assign N2808 = N2776 & N2783;
  assign N2809 = N2776 & yumi_cnt_i[4];
  assign N2810 = N2778 & N2783;
  assign N2811 = N2778 & yumi_cnt_i[4];
  assign N2812 = N2780 & N2783;
  assign N2813 = N2780 & yumi_cnt_i[4];
  assign N2814 = N2782 & N2783;
  assign N2815 = N2782 & yumi_cnt_i[4];
  assign N2816 = ~yumi_cnt_i[5];
  assign N2817 = N2784 & N2816;
  assign N2818 = N2784 & yumi_cnt_i[5];
  assign N2819 = N2786 & N2816;
  assign N2820 = N2786 & yumi_cnt_i[5];
  assign N2821 = N2788 & N2816;
  assign N2822 = N2788 & yumi_cnt_i[5];
  assign N2823 = N2790 & N2816;
  assign N2824 = N2790 & yumi_cnt_i[5];
  assign N2825 = N2792 & N2816;
  assign N2826 = N2792 & yumi_cnt_i[5];
  assign N2827 = N2794 & N2816;
  assign N2828 = N2794 & yumi_cnt_i[5];
  assign N2829 = N2796 & N2816;
  assign N2830 = N2796 & yumi_cnt_i[5];
  assign N2831 = N2798 & N2816;
  assign N2832 = N2798 & yumi_cnt_i[5];
  assign N2833 = N2800 & N2816;
  assign N2834 = N2800 & yumi_cnt_i[5];
  assign N2835 = N2802 & N2816;
  assign N2836 = N2802 & yumi_cnt_i[5];
  assign N2837 = N2804 & N2816;
  assign N2838 = N2804 & yumi_cnt_i[5];
  assign N2839 = N2806 & N2816;
  assign N2840 = N2806 & yumi_cnt_i[5];
  assign N2841 = N2808 & N2816;
  assign N2842 = N2808 & yumi_cnt_i[5];
  assign N2843 = N2810 & N2816;
  assign N2844 = N2810 & yumi_cnt_i[5];
  assign N2845 = N2812 & N2816;
  assign N2846 = N2812 & yumi_cnt_i[5];
  assign N2847 = N2814 & N2816;
  assign N2848 = N2814 & yumi_cnt_i[5];
  assign N2849 = N2785 & N2816;
  assign N2850 = N2785 & yumi_cnt_i[5];
  assign N2851 = N2787 & N2816;
  assign N2852 = N2787 & yumi_cnt_i[5];
  assign N2853 = N2789 & N2816;
  assign N2854 = N2789 & yumi_cnt_i[5];
  assign N2855 = N2791 & N2816;
  assign N2856 = N2791 & yumi_cnt_i[5];
  assign N2857 = N2793 & N2816;
  assign N2858 = N2793 & yumi_cnt_i[5];
  assign N2859 = N2795 & N2816;
  assign N2860 = N2795 & yumi_cnt_i[5];
  assign N2861 = N2797 & N2816;
  assign N2862 = N2797 & yumi_cnt_i[5];
  assign N2863 = N2799 & N2816;
  assign N2864 = N2799 & yumi_cnt_i[5];
  assign N2865 = N2801 & N2816;
  assign N2866 = N2801 & yumi_cnt_i[5];
  assign N2867 = N2803 & N2816;
  assign N2868 = N2803 & yumi_cnt_i[5];
  assign N2869 = N2805 & N2816;
  assign N2870 = N2805 & yumi_cnt_i[5];
  assign N2871 = N2807 & N2816;
  assign N2872 = N2807 & yumi_cnt_i[5];
  assign N2873 = N2809 & N2816;
  assign N2874 = N2809 & yumi_cnt_i[5];
  assign N2875 = N2811 & N2816;
  assign N2876 = N2811 & yumi_cnt_i[5];
  assign N2877 = N2813 & N2816;
  assign N2878 = N2813 & yumi_cnt_i[5];
  assign N2879 = N2815 & N2816;
  assign N2880 = N2815 & yumi_cnt_i[5];
  assign N2881 = ~yumi_cnt_i[6];
  assign N2882 = N2817 & N2881;
  assign N2883 = N2817 & yumi_cnt_i[6];
  assign N2884 = N2819 & N2881;
  assign N2885 = N2819 & yumi_cnt_i[6];
  assign N2886 = N2821 & N2881;
  assign N2887 = N2821 & yumi_cnt_i[6];
  assign N2888 = N2823 & N2881;
  assign N2889 = N2823 & yumi_cnt_i[6];
  assign N2890 = N2825 & N2881;
  assign N2891 = N2825 & yumi_cnt_i[6];
  assign N2892 = N2827 & N2881;
  assign N2893 = N2827 & yumi_cnt_i[6];
  assign N2894 = N2829 & N2881;
  assign N2895 = N2829 & yumi_cnt_i[6];
  assign N2896 = N2831 & N2881;
  assign N2897 = N2831 & yumi_cnt_i[6];
  assign N2898 = N2833 & N2881;
  assign N2899 = N2833 & yumi_cnt_i[6];
  assign N2900 = N2835 & N2881;
  assign N2901 = N2835 & yumi_cnt_i[6];
  assign N2902 = N2837 & N2881;
  assign N2903 = N2837 & yumi_cnt_i[6];
  assign N2904 = N2839 & N2881;
  assign N2905 = N2839 & yumi_cnt_i[6];
  assign N2906 = N2841 & N2881;
  assign N2907 = N2841 & yumi_cnt_i[6];
  assign N2908 = N2843 & N2881;
  assign N2909 = N2843 & yumi_cnt_i[6];
  assign N2910 = N2845 & N2881;
  assign N2911 = N2845 & yumi_cnt_i[6];
  assign N2912 = N2847 & N2881;
  assign N2913 = N2847 & yumi_cnt_i[6];
  assign N2914 = N2849 & N2881;
  assign N2915 = N2849 & yumi_cnt_i[6];
  assign N2916 = N2851 & N2881;
  assign N2917 = N2851 & yumi_cnt_i[6];
  assign N2918 = N2853 & N2881;
  assign N2919 = N2853 & yumi_cnt_i[6];
  assign N2920 = N2855 & N2881;
  assign N2921 = N2855 & yumi_cnt_i[6];
  assign N2922 = N2857 & N2881;
  assign N2923 = N2857 & yumi_cnt_i[6];
  assign N2924 = N2859 & N2881;
  assign N2925 = N2859 & yumi_cnt_i[6];
  assign N2926 = N2861 & N2881;
  assign N2927 = N2861 & yumi_cnt_i[6];
  assign N2928 = N2863 & N2881;
  assign N2929 = N2863 & yumi_cnt_i[6];
  assign N2930 = N2865 & N2881;
  assign N2931 = N2865 & yumi_cnt_i[6];
  assign N2932 = N2867 & N2881;
  assign N2933 = N2867 & yumi_cnt_i[6];
  assign N2934 = N2869 & N2881;
  assign N2935 = N2869 & yumi_cnt_i[6];
  assign N2936 = N2871 & N2881;
  assign N2937 = N2871 & yumi_cnt_i[6];
  assign N2938 = N2873 & N2881;
  assign N2939 = N2873 & yumi_cnt_i[6];
  assign N2940 = N2875 & N2881;
  assign N2941 = N2875 & yumi_cnt_i[6];
  assign N2942 = N2877 & N2881;
  assign N2943 = N2877 & yumi_cnt_i[6];
  assign N2944 = N2879 & N2881;
  assign N2945 = N2879 & yumi_cnt_i[6];
  assign N2946 = N2818 & N2881;
  assign N2947 = N2818 & yumi_cnt_i[6];
  assign N2948 = N2820 & N2881;
  assign N2949 = N2820 & yumi_cnt_i[6];
  assign N2950 = N2822 & N2881;
  assign N2951 = N2822 & yumi_cnt_i[6];
  assign N2952 = N2824 & N2881;
  assign N2953 = N2824 & yumi_cnt_i[6];
  assign N2954 = N2826 & N2881;
  assign N2955 = N2826 & yumi_cnt_i[6];
  assign N2956 = N2828 & N2881;
  assign N2957 = N2828 & yumi_cnt_i[6];
  assign N2958 = N2830 & N2881;
  assign N2959 = N2830 & yumi_cnt_i[6];
  assign N2960 = N2832 & N2881;
  assign N2961 = N2832 & yumi_cnt_i[6];
  assign N2962 = N2834 & N2881;
  assign N2963 = N2834 & yumi_cnt_i[6];
  assign N2964 = N2836 & N2881;
  assign N2965 = N2836 & yumi_cnt_i[6];
  assign N2966 = N2838 & N2881;
  assign N2967 = N2838 & yumi_cnt_i[6];
  assign N2968 = N2840 & N2881;
  assign N2969 = N2840 & yumi_cnt_i[6];
  assign N2970 = N2842 & N2881;
  assign N2971 = N2842 & yumi_cnt_i[6];
  assign N2972 = N2844 & N2881;
  assign N2973 = N2844 & yumi_cnt_i[6];
  assign N2974 = N2846 & N2881;
  assign N2975 = N2846 & yumi_cnt_i[6];
  assign N2976 = N2848 & N2881;
  assign N2977 = N2848 & yumi_cnt_i[6];
  assign N2978 = N2850 & N2881;
  assign N2979 = N2850 & yumi_cnt_i[6];
  assign N2980 = N2852 & N2881;
  assign N2981 = N2852 & yumi_cnt_i[6];
  assign N2982 = N2854 & N2881;
  assign N2983 = N2854 & yumi_cnt_i[6];
  assign N2984 = N2856 & N2881;
  assign N2985 = N2856 & yumi_cnt_i[6];
  assign N2986 = N2858 & N2881;
  assign N2987 = N2858 & yumi_cnt_i[6];
  assign N2988 = N2860 & N2881;
  assign N2989 = N2860 & yumi_cnt_i[6];
  assign N2990 = N2862 & N2881;
  assign N2991 = N2862 & yumi_cnt_i[6];
  assign N2992 = N2864 & N2881;
  assign N2993 = N2864 & yumi_cnt_i[6];
  assign N2994 = N2866 & N2881;
  assign N2995 = N2866 & yumi_cnt_i[6];
  assign N2996 = N2868 & N2881;
  assign N2997 = N2868 & yumi_cnt_i[6];
  assign N2998 = N2870 & N2881;
  assign N2999 = N2870 & yumi_cnt_i[6];
  assign N3000 = N2872 & N2881;
  assign N3001 = N2872 & yumi_cnt_i[6];
  assign N3002 = N2874 & N2881;
  assign N3003 = N2874 & yumi_cnt_i[6];
  assign N3004 = N2876 & N2881;
  assign N3005 = N2876 & yumi_cnt_i[6];
  assign N3006 = N2878 & N2881;
  assign N3007 = N2878 & yumi_cnt_i[6];
  assign N3008 = N2880 & N2881;
  assign N3009 = N2880 & yumi_cnt_i[6];

  always @(posedge clk_i) begin
    if(reset_i) begin
      valid_r_63_sv2v_reg <= 1'b0;
      valid_r_62_sv2v_reg <= 1'b0;
      valid_r_61_sv2v_reg <= 1'b0;
      valid_r_60_sv2v_reg <= 1'b0;
      valid_r_59_sv2v_reg <= 1'b0;
      valid_r_58_sv2v_reg <= 1'b0;
      valid_r_57_sv2v_reg <= 1'b0;
      valid_r_56_sv2v_reg <= 1'b0;
      valid_r_55_sv2v_reg <= 1'b0;
      valid_r_54_sv2v_reg <= 1'b0;
      valid_r_53_sv2v_reg <= 1'b0;
      valid_r_52_sv2v_reg <= 1'b0;
      valid_r_51_sv2v_reg <= 1'b0;
      valid_r_50_sv2v_reg <= 1'b0;
      valid_r_49_sv2v_reg <= 1'b0;
      valid_r_48_sv2v_reg <= 1'b0;
      valid_r_47_sv2v_reg <= 1'b0;
      valid_r_46_sv2v_reg <= 1'b0;
      valid_r_45_sv2v_reg <= 1'b0;
      valid_r_44_sv2v_reg <= 1'b0;
      valid_r_43_sv2v_reg <= 1'b0;
      valid_r_42_sv2v_reg <= 1'b0;
      valid_r_41_sv2v_reg <= 1'b0;
      valid_r_40_sv2v_reg <= 1'b0;
      valid_r_39_sv2v_reg <= 1'b0;
      valid_r_38_sv2v_reg <= 1'b0;
      valid_r_37_sv2v_reg <= 1'b0;
      valid_r_36_sv2v_reg <= 1'b0;
      valid_r_35_sv2v_reg <= 1'b0;
      valid_r_34_sv2v_reg <= 1'b0;
      valid_r_33_sv2v_reg <= 1'b0;
      valid_r_32_sv2v_reg <= 1'b0;
      valid_r_31_sv2v_reg <= 1'b0;
      valid_r_30_sv2v_reg <= 1'b0;
      valid_r_29_sv2v_reg <= 1'b0;
      valid_r_28_sv2v_reg <= 1'b0;
      valid_r_27_sv2v_reg <= 1'b0;
      valid_r_26_sv2v_reg <= 1'b0;
      valid_r_25_sv2v_reg <= 1'b0;
      valid_r_24_sv2v_reg <= 1'b0;
      valid_r_23_sv2v_reg <= 1'b0;
      valid_r_22_sv2v_reg <= 1'b0;
      valid_r_21_sv2v_reg <= 1'b0;
      valid_r_20_sv2v_reg <= 1'b0;
      valid_r_19_sv2v_reg <= 1'b0;
      valid_r_18_sv2v_reg <= 1'b0;
      valid_r_17_sv2v_reg <= 1'b0;
      valid_r_16_sv2v_reg <= 1'b0;
      valid_r_15_sv2v_reg <= 1'b0;
      valid_r_14_sv2v_reg <= 1'b0;
      valid_r_13_sv2v_reg <= 1'b0;
      valid_r_12_sv2v_reg <= 1'b0;
      valid_r_11_sv2v_reg <= 1'b0;
      valid_r_10_sv2v_reg <= 1'b0;
      valid_r_9_sv2v_reg <= 1'b0;
      valid_r_8_sv2v_reg <= 1'b0;
      valid_r_7_sv2v_reg <= 1'b0;
      valid_r_6_sv2v_reg <= 1'b0;
      valid_r_5_sv2v_reg <= 1'b0;
      valid_r_4_sv2v_reg <= 1'b0;
      valid_r_3_sv2v_reg <= 1'b0;
      valid_r_2_sv2v_reg <= 1'b0;
      valid_r_1_sv2v_reg <= 1'b0;
      valid_r_0_sv2v_reg <= 1'b0;
      num_els_r_6_sv2v_reg <= 1'b0;
      num_els_r_5_sv2v_reg <= 1'b0;
      num_els_r_4_sv2v_reg <= 1'b0;
      num_els_r_3_sv2v_reg <= 1'b0;
      num_els_r_2_sv2v_reg <= 1'b0;
      num_els_r_1_sv2v_reg <= 1'b0;
      num_els_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      valid_r_63_sv2v_reg <= valid_nn[63];
      valid_r_62_sv2v_reg <= valid_nn[62];
      valid_r_61_sv2v_reg <= valid_nn[61];
      valid_r_60_sv2v_reg <= valid_nn[60];
      valid_r_59_sv2v_reg <= valid_nn[59];
      valid_r_58_sv2v_reg <= valid_nn[58];
      valid_r_57_sv2v_reg <= valid_nn[57];
      valid_r_56_sv2v_reg <= valid_nn[56];
      valid_r_55_sv2v_reg <= valid_nn[55];
      valid_r_54_sv2v_reg <= valid_nn[54];
      valid_r_53_sv2v_reg <= valid_nn[53];
      valid_r_52_sv2v_reg <= valid_nn[52];
      valid_r_51_sv2v_reg <= valid_nn[51];
      valid_r_50_sv2v_reg <= valid_nn[50];
      valid_r_49_sv2v_reg <= valid_nn[49];
      valid_r_48_sv2v_reg <= valid_nn[48];
      valid_r_47_sv2v_reg <= valid_nn[47];
      valid_r_46_sv2v_reg <= valid_nn[46];
      valid_r_45_sv2v_reg <= valid_nn[45];
      valid_r_44_sv2v_reg <= valid_nn[44];
      valid_r_43_sv2v_reg <= valid_nn[43];
      valid_r_42_sv2v_reg <= valid_nn[42];
      valid_r_41_sv2v_reg <= valid_nn[41];
      valid_r_40_sv2v_reg <= valid_nn[40];
      valid_r_39_sv2v_reg <= valid_nn[39];
      valid_r_38_sv2v_reg <= valid_nn[38];
      valid_r_37_sv2v_reg <= valid_nn[37];
      valid_r_36_sv2v_reg <= valid_nn[36];
      valid_r_35_sv2v_reg <= valid_nn[35];
      valid_r_34_sv2v_reg <= valid_nn[34];
      valid_r_33_sv2v_reg <= valid_nn[33];
      valid_r_32_sv2v_reg <= valid_nn[32];
      valid_r_31_sv2v_reg <= valid_nn[31];
      valid_r_30_sv2v_reg <= valid_nn[30];
      valid_r_29_sv2v_reg <= valid_nn[29];
      valid_r_28_sv2v_reg <= valid_nn[28];
      valid_r_27_sv2v_reg <= valid_nn[27];
      valid_r_26_sv2v_reg <= valid_nn[26];
      valid_r_25_sv2v_reg <= valid_nn[25];
      valid_r_24_sv2v_reg <= valid_nn[24];
      valid_r_23_sv2v_reg <= valid_nn[23];
      valid_r_22_sv2v_reg <= valid_nn[22];
      valid_r_21_sv2v_reg <= valid_nn[21];
      valid_r_20_sv2v_reg <= valid_nn[20];
      valid_r_19_sv2v_reg <= valid_nn[19];
      valid_r_18_sv2v_reg <= valid_nn[18];
      valid_r_17_sv2v_reg <= valid_nn[17];
      valid_r_16_sv2v_reg <= valid_nn[16];
      valid_r_15_sv2v_reg <= valid_nn[15];
      valid_r_14_sv2v_reg <= valid_nn[14];
      valid_r_13_sv2v_reg <= valid_nn[13];
      valid_r_12_sv2v_reg <= valid_nn[12];
      valid_r_11_sv2v_reg <= valid_nn[11];
      valid_r_10_sv2v_reg <= valid_nn[10];
      valid_r_9_sv2v_reg <= valid_nn[9];
      valid_r_8_sv2v_reg <= valid_nn[8];
      valid_r_7_sv2v_reg <= valid_nn[7];
      valid_r_6_sv2v_reg <= valid_nn[6];
      valid_r_5_sv2v_reg <= valid_nn[5];
      valid_r_4_sv2v_reg <= valid_nn[4];
      valid_r_3_sv2v_reg <= valid_nn[3];
      valid_r_2_sv2v_reg <= valid_nn[2];
      valid_r_1_sv2v_reg <= valid_nn[1];
      valid_r_0_sv2v_reg <= valid_nn[0];
      num_els_r_6_sv2v_reg <= num_els_n[6];
      num_els_r_5_sv2v_reg <= num_els_n[5];
      num_els_r_4_sv2v_reg <= num_els_n[4];
      num_els_r_3_sv2v_reg <= num_els_n[3];
      num_els_r_2_sv2v_reg <= num_els_n[2];
      num_els_r_1_sv2v_reg <= num_els_n[1];
      num_els_r_0_sv2v_reg <= num_els_n[0];
    end 
    if(1'b1) begin
      data_r_2047_sv2v_reg <= data_nn[2047];
      data_r_2046_sv2v_reg <= data_nn[2046];
      data_r_2045_sv2v_reg <= data_nn[2045];
      data_r_2044_sv2v_reg <= data_nn[2044];
      data_r_2043_sv2v_reg <= data_nn[2043];
      data_r_2042_sv2v_reg <= data_nn[2042];
      data_r_2041_sv2v_reg <= data_nn[2041];
      data_r_2040_sv2v_reg <= data_nn[2040];
      data_r_2039_sv2v_reg <= data_nn[2039];
      data_r_2038_sv2v_reg <= data_nn[2038];
      data_r_2037_sv2v_reg <= data_nn[2037];
      data_r_2036_sv2v_reg <= data_nn[2036];
      data_r_2035_sv2v_reg <= data_nn[2035];
      data_r_2034_sv2v_reg <= data_nn[2034];
      data_r_2033_sv2v_reg <= data_nn[2033];
      data_r_2032_sv2v_reg <= data_nn[2032];
      data_r_2031_sv2v_reg <= data_nn[2031];
      data_r_2030_sv2v_reg <= data_nn[2030];
      data_r_2029_sv2v_reg <= data_nn[2029];
      data_r_2028_sv2v_reg <= data_nn[2028];
      data_r_2027_sv2v_reg <= data_nn[2027];
      data_r_2026_sv2v_reg <= data_nn[2026];
      data_r_2025_sv2v_reg <= data_nn[2025];
      data_r_2024_sv2v_reg <= data_nn[2024];
      data_r_2023_sv2v_reg <= data_nn[2023];
      data_r_2022_sv2v_reg <= data_nn[2022];
      data_r_2021_sv2v_reg <= data_nn[2021];
      data_r_2020_sv2v_reg <= data_nn[2020];
      data_r_2019_sv2v_reg <= data_nn[2019];
      data_r_2018_sv2v_reg <= data_nn[2018];
      data_r_2017_sv2v_reg <= data_nn[2017];
      data_r_2016_sv2v_reg <= data_nn[2016];
      data_r_2015_sv2v_reg <= data_nn[2015];
      data_r_2014_sv2v_reg <= data_nn[2014];
      data_r_2013_sv2v_reg <= data_nn[2013];
      data_r_2012_sv2v_reg <= data_nn[2012];
      data_r_2011_sv2v_reg <= data_nn[2011];
      data_r_2010_sv2v_reg <= data_nn[2010];
      data_r_2009_sv2v_reg <= data_nn[2009];
      data_r_2008_sv2v_reg <= data_nn[2008];
      data_r_2007_sv2v_reg <= data_nn[2007];
      data_r_2006_sv2v_reg <= data_nn[2006];
      data_r_2005_sv2v_reg <= data_nn[2005];
      data_r_2004_sv2v_reg <= data_nn[2004];
      data_r_2003_sv2v_reg <= data_nn[2003];
      data_r_2002_sv2v_reg <= data_nn[2002];
      data_r_2001_sv2v_reg <= data_nn[2001];
      data_r_2000_sv2v_reg <= data_nn[2000];
      data_r_1999_sv2v_reg <= data_nn[1999];
      data_r_1998_sv2v_reg <= data_nn[1998];
      data_r_1997_sv2v_reg <= data_nn[1997];
      data_r_1996_sv2v_reg <= data_nn[1996];
      data_r_1995_sv2v_reg <= data_nn[1995];
      data_r_1994_sv2v_reg <= data_nn[1994];
      data_r_1993_sv2v_reg <= data_nn[1993];
      data_r_1992_sv2v_reg <= data_nn[1992];
      data_r_1991_sv2v_reg <= data_nn[1991];
      data_r_1990_sv2v_reg <= data_nn[1990];
      data_r_1989_sv2v_reg <= data_nn[1989];
      data_r_1988_sv2v_reg <= data_nn[1988];
      data_r_1987_sv2v_reg <= data_nn[1987];
      data_r_1986_sv2v_reg <= data_nn[1986];
      data_r_1985_sv2v_reg <= data_nn[1985];
      data_r_1984_sv2v_reg <= data_nn[1984];
      data_r_1983_sv2v_reg <= data_nn[1983];
      data_r_1982_sv2v_reg <= data_nn[1982];
      data_r_1981_sv2v_reg <= data_nn[1981];
      data_r_1980_sv2v_reg <= data_nn[1980];
      data_r_1979_sv2v_reg <= data_nn[1979];
      data_r_1978_sv2v_reg <= data_nn[1978];
      data_r_1977_sv2v_reg <= data_nn[1977];
      data_r_1976_sv2v_reg <= data_nn[1976];
      data_r_1975_sv2v_reg <= data_nn[1975];
      data_r_1974_sv2v_reg <= data_nn[1974];
      data_r_1973_sv2v_reg <= data_nn[1973];
      data_r_1972_sv2v_reg <= data_nn[1972];
      data_r_1971_sv2v_reg <= data_nn[1971];
      data_r_1970_sv2v_reg <= data_nn[1970];
      data_r_1969_sv2v_reg <= data_nn[1969];
      data_r_1968_sv2v_reg <= data_nn[1968];
      data_r_1967_sv2v_reg <= data_nn[1967];
      data_r_1966_sv2v_reg <= data_nn[1966];
      data_r_1965_sv2v_reg <= data_nn[1965];
      data_r_1964_sv2v_reg <= data_nn[1964];
      data_r_1963_sv2v_reg <= data_nn[1963];
      data_r_1962_sv2v_reg <= data_nn[1962];
      data_r_1961_sv2v_reg <= data_nn[1961];
      data_r_1960_sv2v_reg <= data_nn[1960];
      data_r_1959_sv2v_reg <= data_nn[1959];
      data_r_1958_sv2v_reg <= data_nn[1958];
      data_r_1957_sv2v_reg <= data_nn[1957];
      data_r_1956_sv2v_reg <= data_nn[1956];
      data_r_1955_sv2v_reg <= data_nn[1955];
      data_r_1954_sv2v_reg <= data_nn[1954];
      data_r_1953_sv2v_reg <= data_nn[1953];
      data_r_1952_sv2v_reg <= data_nn[1952];
      data_r_1951_sv2v_reg <= data_nn[1951];
      data_r_1950_sv2v_reg <= data_nn[1950];
      data_r_1949_sv2v_reg <= data_nn[1949];
      data_r_1948_sv2v_reg <= data_nn[1948];
      data_r_1947_sv2v_reg <= data_nn[1947];
      data_r_1946_sv2v_reg <= data_nn[1946];
      data_r_1945_sv2v_reg <= data_nn[1945];
      data_r_1944_sv2v_reg <= data_nn[1944];
      data_r_1943_sv2v_reg <= data_nn[1943];
      data_r_1942_sv2v_reg <= data_nn[1942];
      data_r_1941_sv2v_reg <= data_nn[1941];
      data_r_1940_sv2v_reg <= data_nn[1940];
      data_r_1939_sv2v_reg <= data_nn[1939];
      data_r_1938_sv2v_reg <= data_nn[1938];
      data_r_1937_sv2v_reg <= data_nn[1937];
      data_r_1936_sv2v_reg <= data_nn[1936];
      data_r_1935_sv2v_reg <= data_nn[1935];
      data_r_1934_sv2v_reg <= data_nn[1934];
      data_r_1933_sv2v_reg <= data_nn[1933];
      data_r_1932_sv2v_reg <= data_nn[1932];
      data_r_1931_sv2v_reg <= data_nn[1931];
      data_r_1930_sv2v_reg <= data_nn[1930];
      data_r_1929_sv2v_reg <= data_nn[1929];
      data_r_1928_sv2v_reg <= data_nn[1928];
      data_r_1927_sv2v_reg <= data_nn[1927];
      data_r_1926_sv2v_reg <= data_nn[1926];
      data_r_1925_sv2v_reg <= data_nn[1925];
      data_r_1924_sv2v_reg <= data_nn[1924];
      data_r_1923_sv2v_reg <= data_nn[1923];
      data_r_1922_sv2v_reg <= data_nn[1922];
      data_r_1921_sv2v_reg <= data_nn[1921];
      data_r_1920_sv2v_reg <= data_nn[1920];
      data_r_1919_sv2v_reg <= data_nn[1919];
      data_r_1918_sv2v_reg <= data_nn[1918];
      data_r_1917_sv2v_reg <= data_nn[1917];
      data_r_1916_sv2v_reg <= data_nn[1916];
      data_r_1915_sv2v_reg <= data_nn[1915];
      data_r_1914_sv2v_reg <= data_nn[1914];
      data_r_1913_sv2v_reg <= data_nn[1913];
      data_r_1912_sv2v_reg <= data_nn[1912];
      data_r_1911_sv2v_reg <= data_nn[1911];
      data_r_1910_sv2v_reg <= data_nn[1910];
      data_r_1909_sv2v_reg <= data_nn[1909];
      data_r_1908_sv2v_reg <= data_nn[1908];
      data_r_1907_sv2v_reg <= data_nn[1907];
      data_r_1906_sv2v_reg <= data_nn[1906];
      data_r_1905_sv2v_reg <= data_nn[1905];
      data_r_1904_sv2v_reg <= data_nn[1904];
      data_r_1903_sv2v_reg <= data_nn[1903];
      data_r_1902_sv2v_reg <= data_nn[1902];
      data_r_1901_sv2v_reg <= data_nn[1901];
      data_r_1900_sv2v_reg <= data_nn[1900];
      data_r_1899_sv2v_reg <= data_nn[1899];
      data_r_1898_sv2v_reg <= data_nn[1898];
      data_r_1897_sv2v_reg <= data_nn[1897];
      data_r_1896_sv2v_reg <= data_nn[1896];
      data_r_1895_sv2v_reg <= data_nn[1895];
      data_r_1894_sv2v_reg <= data_nn[1894];
      data_r_1893_sv2v_reg <= data_nn[1893];
      data_r_1892_sv2v_reg <= data_nn[1892];
      data_r_1891_sv2v_reg <= data_nn[1891];
      data_r_1890_sv2v_reg <= data_nn[1890];
      data_r_1889_sv2v_reg <= data_nn[1889];
      data_r_1888_sv2v_reg <= data_nn[1888];
      data_r_1887_sv2v_reg <= data_nn[1887];
      data_r_1886_sv2v_reg <= data_nn[1886];
      data_r_1885_sv2v_reg <= data_nn[1885];
      data_r_1884_sv2v_reg <= data_nn[1884];
      data_r_1883_sv2v_reg <= data_nn[1883];
      data_r_1882_sv2v_reg <= data_nn[1882];
      data_r_1881_sv2v_reg <= data_nn[1881];
      data_r_1880_sv2v_reg <= data_nn[1880];
      data_r_1879_sv2v_reg <= data_nn[1879];
      data_r_1878_sv2v_reg <= data_nn[1878];
      data_r_1877_sv2v_reg <= data_nn[1877];
      data_r_1876_sv2v_reg <= data_nn[1876];
      data_r_1875_sv2v_reg <= data_nn[1875];
      data_r_1874_sv2v_reg <= data_nn[1874];
      data_r_1873_sv2v_reg <= data_nn[1873];
      data_r_1872_sv2v_reg <= data_nn[1872];
      data_r_1871_sv2v_reg <= data_nn[1871];
      data_r_1870_sv2v_reg <= data_nn[1870];
      data_r_1869_sv2v_reg <= data_nn[1869];
      data_r_1868_sv2v_reg <= data_nn[1868];
      data_r_1867_sv2v_reg <= data_nn[1867];
      data_r_1866_sv2v_reg <= data_nn[1866];
      data_r_1865_sv2v_reg <= data_nn[1865];
      data_r_1864_sv2v_reg <= data_nn[1864];
      data_r_1863_sv2v_reg <= data_nn[1863];
      data_r_1862_sv2v_reg <= data_nn[1862];
      data_r_1861_sv2v_reg <= data_nn[1861];
      data_r_1860_sv2v_reg <= data_nn[1860];
      data_r_1859_sv2v_reg <= data_nn[1859];
      data_r_1858_sv2v_reg <= data_nn[1858];
      data_r_1857_sv2v_reg <= data_nn[1857];
      data_r_1856_sv2v_reg <= data_nn[1856];
      data_r_1855_sv2v_reg <= data_nn[1855];
      data_r_1854_sv2v_reg <= data_nn[1854];
      data_r_1853_sv2v_reg <= data_nn[1853];
      data_r_1852_sv2v_reg <= data_nn[1852];
      data_r_1851_sv2v_reg <= data_nn[1851];
      data_r_1850_sv2v_reg <= data_nn[1850];
      data_r_1849_sv2v_reg <= data_nn[1849];
      data_r_1848_sv2v_reg <= data_nn[1848];
      data_r_1847_sv2v_reg <= data_nn[1847];
      data_r_1846_sv2v_reg <= data_nn[1846];
      data_r_1845_sv2v_reg <= data_nn[1845];
      data_r_1844_sv2v_reg <= data_nn[1844];
      data_r_1843_sv2v_reg <= data_nn[1843];
      data_r_1842_sv2v_reg <= data_nn[1842];
      data_r_1841_sv2v_reg <= data_nn[1841];
      data_r_1840_sv2v_reg <= data_nn[1840];
      data_r_1839_sv2v_reg <= data_nn[1839];
      data_r_1838_sv2v_reg <= data_nn[1838];
      data_r_1837_sv2v_reg <= data_nn[1837];
      data_r_1836_sv2v_reg <= data_nn[1836];
      data_r_1835_sv2v_reg <= data_nn[1835];
      data_r_1834_sv2v_reg <= data_nn[1834];
      data_r_1833_sv2v_reg <= data_nn[1833];
      data_r_1832_sv2v_reg <= data_nn[1832];
      data_r_1831_sv2v_reg <= data_nn[1831];
      data_r_1830_sv2v_reg <= data_nn[1830];
      data_r_1829_sv2v_reg <= data_nn[1829];
      data_r_1828_sv2v_reg <= data_nn[1828];
      data_r_1827_sv2v_reg <= data_nn[1827];
      data_r_1826_sv2v_reg <= data_nn[1826];
      data_r_1825_sv2v_reg <= data_nn[1825];
      data_r_1824_sv2v_reg <= data_nn[1824];
      data_r_1823_sv2v_reg <= data_nn[1823];
      data_r_1822_sv2v_reg <= data_nn[1822];
      data_r_1821_sv2v_reg <= data_nn[1821];
      data_r_1820_sv2v_reg <= data_nn[1820];
      data_r_1819_sv2v_reg <= data_nn[1819];
      data_r_1818_sv2v_reg <= data_nn[1818];
      data_r_1817_sv2v_reg <= data_nn[1817];
      data_r_1816_sv2v_reg <= data_nn[1816];
      data_r_1815_sv2v_reg <= data_nn[1815];
      data_r_1814_sv2v_reg <= data_nn[1814];
      data_r_1813_sv2v_reg <= data_nn[1813];
      data_r_1812_sv2v_reg <= data_nn[1812];
      data_r_1811_sv2v_reg <= data_nn[1811];
      data_r_1810_sv2v_reg <= data_nn[1810];
      data_r_1809_sv2v_reg <= data_nn[1809];
      data_r_1808_sv2v_reg <= data_nn[1808];
      data_r_1807_sv2v_reg <= data_nn[1807];
      data_r_1806_sv2v_reg <= data_nn[1806];
      data_r_1805_sv2v_reg <= data_nn[1805];
      data_r_1804_sv2v_reg <= data_nn[1804];
      data_r_1803_sv2v_reg <= data_nn[1803];
      data_r_1802_sv2v_reg <= data_nn[1802];
      data_r_1801_sv2v_reg <= data_nn[1801];
      data_r_1800_sv2v_reg <= data_nn[1800];
      data_r_1799_sv2v_reg <= data_nn[1799];
      data_r_1798_sv2v_reg <= data_nn[1798];
      data_r_1797_sv2v_reg <= data_nn[1797];
      data_r_1796_sv2v_reg <= data_nn[1796];
      data_r_1795_sv2v_reg <= data_nn[1795];
      data_r_1794_sv2v_reg <= data_nn[1794];
      data_r_1793_sv2v_reg <= data_nn[1793];
      data_r_1792_sv2v_reg <= data_nn[1792];
      data_r_1791_sv2v_reg <= data_nn[1791];
      data_r_1790_sv2v_reg <= data_nn[1790];
      data_r_1789_sv2v_reg <= data_nn[1789];
      data_r_1788_sv2v_reg <= data_nn[1788];
      data_r_1787_sv2v_reg <= data_nn[1787];
      data_r_1786_sv2v_reg <= data_nn[1786];
      data_r_1785_sv2v_reg <= data_nn[1785];
      data_r_1784_sv2v_reg <= data_nn[1784];
      data_r_1783_sv2v_reg <= data_nn[1783];
      data_r_1782_sv2v_reg <= data_nn[1782];
      data_r_1781_sv2v_reg <= data_nn[1781];
      data_r_1780_sv2v_reg <= data_nn[1780];
      data_r_1779_sv2v_reg <= data_nn[1779];
      data_r_1778_sv2v_reg <= data_nn[1778];
      data_r_1777_sv2v_reg <= data_nn[1777];
      data_r_1776_sv2v_reg <= data_nn[1776];
      data_r_1775_sv2v_reg <= data_nn[1775];
      data_r_1774_sv2v_reg <= data_nn[1774];
      data_r_1773_sv2v_reg <= data_nn[1773];
      data_r_1772_sv2v_reg <= data_nn[1772];
      data_r_1771_sv2v_reg <= data_nn[1771];
      data_r_1770_sv2v_reg <= data_nn[1770];
      data_r_1769_sv2v_reg <= data_nn[1769];
      data_r_1768_sv2v_reg <= data_nn[1768];
      data_r_1767_sv2v_reg <= data_nn[1767];
      data_r_1766_sv2v_reg <= data_nn[1766];
      data_r_1765_sv2v_reg <= data_nn[1765];
      data_r_1764_sv2v_reg <= data_nn[1764];
      data_r_1763_sv2v_reg <= data_nn[1763];
      data_r_1762_sv2v_reg <= data_nn[1762];
      data_r_1761_sv2v_reg <= data_nn[1761];
      data_r_1760_sv2v_reg <= data_nn[1760];
      data_r_1759_sv2v_reg <= data_nn[1759];
      data_r_1758_sv2v_reg <= data_nn[1758];
      data_r_1757_sv2v_reg <= data_nn[1757];
      data_r_1756_sv2v_reg <= data_nn[1756];
      data_r_1755_sv2v_reg <= data_nn[1755];
      data_r_1754_sv2v_reg <= data_nn[1754];
      data_r_1753_sv2v_reg <= data_nn[1753];
      data_r_1752_sv2v_reg <= data_nn[1752];
      data_r_1751_sv2v_reg <= data_nn[1751];
      data_r_1750_sv2v_reg <= data_nn[1750];
      data_r_1749_sv2v_reg <= data_nn[1749];
      data_r_1748_sv2v_reg <= data_nn[1748];
      data_r_1747_sv2v_reg <= data_nn[1747];
      data_r_1746_sv2v_reg <= data_nn[1746];
      data_r_1745_sv2v_reg <= data_nn[1745];
      data_r_1744_sv2v_reg <= data_nn[1744];
      data_r_1743_sv2v_reg <= data_nn[1743];
      data_r_1742_sv2v_reg <= data_nn[1742];
      data_r_1741_sv2v_reg <= data_nn[1741];
      data_r_1740_sv2v_reg <= data_nn[1740];
      data_r_1739_sv2v_reg <= data_nn[1739];
      data_r_1738_sv2v_reg <= data_nn[1738];
      data_r_1737_sv2v_reg <= data_nn[1737];
      data_r_1736_sv2v_reg <= data_nn[1736];
      data_r_1735_sv2v_reg <= data_nn[1735];
      data_r_1734_sv2v_reg <= data_nn[1734];
      data_r_1733_sv2v_reg <= data_nn[1733];
      data_r_1732_sv2v_reg <= data_nn[1732];
      data_r_1731_sv2v_reg <= data_nn[1731];
      data_r_1730_sv2v_reg <= data_nn[1730];
      data_r_1729_sv2v_reg <= data_nn[1729];
      data_r_1728_sv2v_reg <= data_nn[1728];
      data_r_1727_sv2v_reg <= data_nn[1727];
      data_r_1726_sv2v_reg <= data_nn[1726];
      data_r_1725_sv2v_reg <= data_nn[1725];
      data_r_1724_sv2v_reg <= data_nn[1724];
      data_r_1723_sv2v_reg <= data_nn[1723];
      data_r_1722_sv2v_reg <= data_nn[1722];
      data_r_1721_sv2v_reg <= data_nn[1721];
      data_r_1720_sv2v_reg <= data_nn[1720];
      data_r_1719_sv2v_reg <= data_nn[1719];
      data_r_1718_sv2v_reg <= data_nn[1718];
      data_r_1717_sv2v_reg <= data_nn[1717];
      data_r_1716_sv2v_reg <= data_nn[1716];
      data_r_1715_sv2v_reg <= data_nn[1715];
      data_r_1714_sv2v_reg <= data_nn[1714];
      data_r_1713_sv2v_reg <= data_nn[1713];
      data_r_1712_sv2v_reg <= data_nn[1712];
      data_r_1711_sv2v_reg <= data_nn[1711];
      data_r_1710_sv2v_reg <= data_nn[1710];
      data_r_1709_sv2v_reg <= data_nn[1709];
      data_r_1708_sv2v_reg <= data_nn[1708];
      data_r_1707_sv2v_reg <= data_nn[1707];
      data_r_1706_sv2v_reg <= data_nn[1706];
      data_r_1705_sv2v_reg <= data_nn[1705];
      data_r_1704_sv2v_reg <= data_nn[1704];
      data_r_1703_sv2v_reg <= data_nn[1703];
      data_r_1702_sv2v_reg <= data_nn[1702];
      data_r_1701_sv2v_reg <= data_nn[1701];
      data_r_1700_sv2v_reg <= data_nn[1700];
      data_r_1699_sv2v_reg <= data_nn[1699];
      data_r_1698_sv2v_reg <= data_nn[1698];
      data_r_1697_sv2v_reg <= data_nn[1697];
      data_r_1696_sv2v_reg <= data_nn[1696];
      data_r_1695_sv2v_reg <= data_nn[1695];
      data_r_1694_sv2v_reg <= data_nn[1694];
      data_r_1693_sv2v_reg <= data_nn[1693];
      data_r_1692_sv2v_reg <= data_nn[1692];
      data_r_1691_sv2v_reg <= data_nn[1691];
      data_r_1690_sv2v_reg <= data_nn[1690];
      data_r_1689_sv2v_reg <= data_nn[1689];
      data_r_1688_sv2v_reg <= data_nn[1688];
      data_r_1687_sv2v_reg <= data_nn[1687];
      data_r_1686_sv2v_reg <= data_nn[1686];
      data_r_1685_sv2v_reg <= data_nn[1685];
      data_r_1684_sv2v_reg <= data_nn[1684];
      data_r_1683_sv2v_reg <= data_nn[1683];
      data_r_1682_sv2v_reg <= data_nn[1682];
      data_r_1681_sv2v_reg <= data_nn[1681];
      data_r_1680_sv2v_reg <= data_nn[1680];
      data_r_1679_sv2v_reg <= data_nn[1679];
      data_r_1678_sv2v_reg <= data_nn[1678];
      data_r_1677_sv2v_reg <= data_nn[1677];
      data_r_1676_sv2v_reg <= data_nn[1676];
      data_r_1675_sv2v_reg <= data_nn[1675];
      data_r_1674_sv2v_reg <= data_nn[1674];
      data_r_1673_sv2v_reg <= data_nn[1673];
      data_r_1672_sv2v_reg <= data_nn[1672];
      data_r_1671_sv2v_reg <= data_nn[1671];
      data_r_1670_sv2v_reg <= data_nn[1670];
      data_r_1669_sv2v_reg <= data_nn[1669];
      data_r_1668_sv2v_reg <= data_nn[1668];
      data_r_1667_sv2v_reg <= data_nn[1667];
      data_r_1666_sv2v_reg <= data_nn[1666];
      data_r_1665_sv2v_reg <= data_nn[1665];
      data_r_1664_sv2v_reg <= data_nn[1664];
      data_r_1663_sv2v_reg <= data_nn[1663];
      data_r_1662_sv2v_reg <= data_nn[1662];
      data_r_1661_sv2v_reg <= data_nn[1661];
      data_r_1660_sv2v_reg <= data_nn[1660];
      data_r_1659_sv2v_reg <= data_nn[1659];
      data_r_1658_sv2v_reg <= data_nn[1658];
      data_r_1657_sv2v_reg <= data_nn[1657];
      data_r_1656_sv2v_reg <= data_nn[1656];
      data_r_1655_sv2v_reg <= data_nn[1655];
      data_r_1654_sv2v_reg <= data_nn[1654];
      data_r_1653_sv2v_reg <= data_nn[1653];
      data_r_1652_sv2v_reg <= data_nn[1652];
      data_r_1651_sv2v_reg <= data_nn[1651];
      data_r_1650_sv2v_reg <= data_nn[1650];
      data_r_1649_sv2v_reg <= data_nn[1649];
      data_r_1648_sv2v_reg <= data_nn[1648];
      data_r_1647_sv2v_reg <= data_nn[1647];
      data_r_1646_sv2v_reg <= data_nn[1646];
      data_r_1645_sv2v_reg <= data_nn[1645];
      data_r_1644_sv2v_reg <= data_nn[1644];
      data_r_1643_sv2v_reg <= data_nn[1643];
      data_r_1642_sv2v_reg <= data_nn[1642];
      data_r_1641_sv2v_reg <= data_nn[1641];
      data_r_1640_sv2v_reg <= data_nn[1640];
      data_r_1639_sv2v_reg <= data_nn[1639];
      data_r_1638_sv2v_reg <= data_nn[1638];
      data_r_1637_sv2v_reg <= data_nn[1637];
      data_r_1636_sv2v_reg <= data_nn[1636];
      data_r_1635_sv2v_reg <= data_nn[1635];
      data_r_1634_sv2v_reg <= data_nn[1634];
      data_r_1633_sv2v_reg <= data_nn[1633];
      data_r_1632_sv2v_reg <= data_nn[1632];
      data_r_1631_sv2v_reg <= data_nn[1631];
      data_r_1630_sv2v_reg <= data_nn[1630];
      data_r_1629_sv2v_reg <= data_nn[1629];
      data_r_1628_sv2v_reg <= data_nn[1628];
      data_r_1627_sv2v_reg <= data_nn[1627];
      data_r_1626_sv2v_reg <= data_nn[1626];
      data_r_1625_sv2v_reg <= data_nn[1625];
      data_r_1624_sv2v_reg <= data_nn[1624];
      data_r_1623_sv2v_reg <= data_nn[1623];
      data_r_1622_sv2v_reg <= data_nn[1622];
      data_r_1621_sv2v_reg <= data_nn[1621];
      data_r_1620_sv2v_reg <= data_nn[1620];
      data_r_1619_sv2v_reg <= data_nn[1619];
      data_r_1618_sv2v_reg <= data_nn[1618];
      data_r_1617_sv2v_reg <= data_nn[1617];
      data_r_1616_sv2v_reg <= data_nn[1616];
      data_r_1615_sv2v_reg <= data_nn[1615];
      data_r_1614_sv2v_reg <= data_nn[1614];
      data_r_1613_sv2v_reg <= data_nn[1613];
      data_r_1612_sv2v_reg <= data_nn[1612];
      data_r_1611_sv2v_reg <= data_nn[1611];
      data_r_1610_sv2v_reg <= data_nn[1610];
      data_r_1609_sv2v_reg <= data_nn[1609];
      data_r_1608_sv2v_reg <= data_nn[1608];
      data_r_1607_sv2v_reg <= data_nn[1607];
      data_r_1606_sv2v_reg <= data_nn[1606];
      data_r_1605_sv2v_reg <= data_nn[1605];
      data_r_1604_sv2v_reg <= data_nn[1604];
      data_r_1603_sv2v_reg <= data_nn[1603];
      data_r_1602_sv2v_reg <= data_nn[1602];
      data_r_1601_sv2v_reg <= data_nn[1601];
      data_r_1600_sv2v_reg <= data_nn[1600];
      data_r_1599_sv2v_reg <= data_nn[1599];
      data_r_1598_sv2v_reg <= data_nn[1598];
      data_r_1597_sv2v_reg <= data_nn[1597];
      data_r_1596_sv2v_reg <= data_nn[1596];
      data_r_1595_sv2v_reg <= data_nn[1595];
      data_r_1594_sv2v_reg <= data_nn[1594];
      data_r_1593_sv2v_reg <= data_nn[1593];
      data_r_1592_sv2v_reg <= data_nn[1592];
      data_r_1591_sv2v_reg <= data_nn[1591];
      data_r_1590_sv2v_reg <= data_nn[1590];
      data_r_1589_sv2v_reg <= data_nn[1589];
      data_r_1588_sv2v_reg <= data_nn[1588];
      data_r_1587_sv2v_reg <= data_nn[1587];
      data_r_1586_sv2v_reg <= data_nn[1586];
      data_r_1585_sv2v_reg <= data_nn[1585];
      data_r_1584_sv2v_reg <= data_nn[1584];
      data_r_1583_sv2v_reg <= data_nn[1583];
      data_r_1582_sv2v_reg <= data_nn[1582];
      data_r_1581_sv2v_reg <= data_nn[1581];
      data_r_1580_sv2v_reg <= data_nn[1580];
      data_r_1579_sv2v_reg <= data_nn[1579];
      data_r_1578_sv2v_reg <= data_nn[1578];
      data_r_1577_sv2v_reg <= data_nn[1577];
      data_r_1576_sv2v_reg <= data_nn[1576];
      data_r_1575_sv2v_reg <= data_nn[1575];
      data_r_1574_sv2v_reg <= data_nn[1574];
      data_r_1573_sv2v_reg <= data_nn[1573];
      data_r_1572_sv2v_reg <= data_nn[1572];
      data_r_1571_sv2v_reg <= data_nn[1571];
      data_r_1570_sv2v_reg <= data_nn[1570];
      data_r_1569_sv2v_reg <= data_nn[1569];
      data_r_1568_sv2v_reg <= data_nn[1568];
      data_r_1567_sv2v_reg <= data_nn[1567];
      data_r_1566_sv2v_reg <= data_nn[1566];
      data_r_1565_sv2v_reg <= data_nn[1565];
      data_r_1564_sv2v_reg <= data_nn[1564];
      data_r_1563_sv2v_reg <= data_nn[1563];
      data_r_1562_sv2v_reg <= data_nn[1562];
      data_r_1561_sv2v_reg <= data_nn[1561];
      data_r_1560_sv2v_reg <= data_nn[1560];
      data_r_1559_sv2v_reg <= data_nn[1559];
      data_r_1558_sv2v_reg <= data_nn[1558];
      data_r_1557_sv2v_reg <= data_nn[1557];
      data_r_1556_sv2v_reg <= data_nn[1556];
      data_r_1555_sv2v_reg <= data_nn[1555];
      data_r_1554_sv2v_reg <= data_nn[1554];
      data_r_1553_sv2v_reg <= data_nn[1553];
      data_r_1552_sv2v_reg <= data_nn[1552];
      data_r_1551_sv2v_reg <= data_nn[1551];
      data_r_1550_sv2v_reg <= data_nn[1550];
      data_r_1549_sv2v_reg <= data_nn[1549];
      data_r_1548_sv2v_reg <= data_nn[1548];
      data_r_1547_sv2v_reg <= data_nn[1547];
      data_r_1546_sv2v_reg <= data_nn[1546];
      data_r_1545_sv2v_reg <= data_nn[1545];
      data_r_1544_sv2v_reg <= data_nn[1544];
      data_r_1543_sv2v_reg <= data_nn[1543];
      data_r_1542_sv2v_reg <= data_nn[1542];
      data_r_1541_sv2v_reg <= data_nn[1541];
      data_r_1540_sv2v_reg <= data_nn[1540];
      data_r_1539_sv2v_reg <= data_nn[1539];
      data_r_1538_sv2v_reg <= data_nn[1538];
      data_r_1537_sv2v_reg <= data_nn[1537];
      data_r_1536_sv2v_reg <= data_nn[1536];
      data_r_1535_sv2v_reg <= data_nn[1535];
      data_r_1534_sv2v_reg <= data_nn[1534];
      data_r_1533_sv2v_reg <= data_nn[1533];
      data_r_1532_sv2v_reg <= data_nn[1532];
      data_r_1531_sv2v_reg <= data_nn[1531];
      data_r_1530_sv2v_reg <= data_nn[1530];
      data_r_1529_sv2v_reg <= data_nn[1529];
      data_r_1528_sv2v_reg <= data_nn[1528];
      data_r_1527_sv2v_reg <= data_nn[1527];
      data_r_1526_sv2v_reg <= data_nn[1526];
      data_r_1525_sv2v_reg <= data_nn[1525];
      data_r_1524_sv2v_reg <= data_nn[1524];
      data_r_1523_sv2v_reg <= data_nn[1523];
      data_r_1522_sv2v_reg <= data_nn[1522];
      data_r_1521_sv2v_reg <= data_nn[1521];
      data_r_1520_sv2v_reg <= data_nn[1520];
      data_r_1519_sv2v_reg <= data_nn[1519];
      data_r_1518_sv2v_reg <= data_nn[1518];
      data_r_1517_sv2v_reg <= data_nn[1517];
      data_r_1516_sv2v_reg <= data_nn[1516];
      data_r_1515_sv2v_reg <= data_nn[1515];
      data_r_1514_sv2v_reg <= data_nn[1514];
      data_r_1513_sv2v_reg <= data_nn[1513];
      data_r_1512_sv2v_reg <= data_nn[1512];
      data_r_1511_sv2v_reg <= data_nn[1511];
      data_r_1510_sv2v_reg <= data_nn[1510];
      data_r_1509_sv2v_reg <= data_nn[1509];
      data_r_1508_sv2v_reg <= data_nn[1508];
      data_r_1507_sv2v_reg <= data_nn[1507];
      data_r_1506_sv2v_reg <= data_nn[1506];
      data_r_1505_sv2v_reg <= data_nn[1505];
      data_r_1504_sv2v_reg <= data_nn[1504];
      data_r_1503_sv2v_reg <= data_nn[1503];
      data_r_1502_sv2v_reg <= data_nn[1502];
      data_r_1501_sv2v_reg <= data_nn[1501];
      data_r_1500_sv2v_reg <= data_nn[1500];
      data_r_1499_sv2v_reg <= data_nn[1499];
      data_r_1498_sv2v_reg <= data_nn[1498];
      data_r_1497_sv2v_reg <= data_nn[1497];
      data_r_1496_sv2v_reg <= data_nn[1496];
      data_r_1495_sv2v_reg <= data_nn[1495];
      data_r_1494_sv2v_reg <= data_nn[1494];
      data_r_1493_sv2v_reg <= data_nn[1493];
      data_r_1492_sv2v_reg <= data_nn[1492];
      data_r_1491_sv2v_reg <= data_nn[1491];
      data_r_1490_sv2v_reg <= data_nn[1490];
      data_r_1489_sv2v_reg <= data_nn[1489];
      data_r_1488_sv2v_reg <= data_nn[1488];
      data_r_1487_sv2v_reg <= data_nn[1487];
      data_r_1486_sv2v_reg <= data_nn[1486];
      data_r_1485_sv2v_reg <= data_nn[1485];
      data_r_1484_sv2v_reg <= data_nn[1484];
      data_r_1483_sv2v_reg <= data_nn[1483];
      data_r_1482_sv2v_reg <= data_nn[1482];
      data_r_1481_sv2v_reg <= data_nn[1481];
      data_r_1480_sv2v_reg <= data_nn[1480];
      data_r_1479_sv2v_reg <= data_nn[1479];
      data_r_1478_sv2v_reg <= data_nn[1478];
      data_r_1477_sv2v_reg <= data_nn[1477];
      data_r_1476_sv2v_reg <= data_nn[1476];
      data_r_1475_sv2v_reg <= data_nn[1475];
      data_r_1474_sv2v_reg <= data_nn[1474];
      data_r_1473_sv2v_reg <= data_nn[1473];
      data_r_1472_sv2v_reg <= data_nn[1472];
      data_r_1471_sv2v_reg <= data_nn[1471];
      data_r_1470_sv2v_reg <= data_nn[1470];
      data_r_1469_sv2v_reg <= data_nn[1469];
      data_r_1468_sv2v_reg <= data_nn[1468];
      data_r_1467_sv2v_reg <= data_nn[1467];
      data_r_1466_sv2v_reg <= data_nn[1466];
      data_r_1465_sv2v_reg <= data_nn[1465];
      data_r_1464_sv2v_reg <= data_nn[1464];
      data_r_1463_sv2v_reg <= data_nn[1463];
      data_r_1462_sv2v_reg <= data_nn[1462];
      data_r_1461_sv2v_reg <= data_nn[1461];
      data_r_1460_sv2v_reg <= data_nn[1460];
      data_r_1459_sv2v_reg <= data_nn[1459];
      data_r_1458_sv2v_reg <= data_nn[1458];
      data_r_1457_sv2v_reg <= data_nn[1457];
      data_r_1456_sv2v_reg <= data_nn[1456];
      data_r_1455_sv2v_reg <= data_nn[1455];
      data_r_1454_sv2v_reg <= data_nn[1454];
      data_r_1453_sv2v_reg <= data_nn[1453];
      data_r_1452_sv2v_reg <= data_nn[1452];
      data_r_1451_sv2v_reg <= data_nn[1451];
      data_r_1450_sv2v_reg <= data_nn[1450];
      data_r_1449_sv2v_reg <= data_nn[1449];
      data_r_1448_sv2v_reg <= data_nn[1448];
      data_r_1447_sv2v_reg <= data_nn[1447];
      data_r_1446_sv2v_reg <= data_nn[1446];
      data_r_1445_sv2v_reg <= data_nn[1445];
      data_r_1444_sv2v_reg <= data_nn[1444];
      data_r_1443_sv2v_reg <= data_nn[1443];
      data_r_1442_sv2v_reg <= data_nn[1442];
      data_r_1441_sv2v_reg <= data_nn[1441];
      data_r_1440_sv2v_reg <= data_nn[1440];
      data_r_1439_sv2v_reg <= data_nn[1439];
      data_r_1438_sv2v_reg <= data_nn[1438];
      data_r_1437_sv2v_reg <= data_nn[1437];
      data_r_1436_sv2v_reg <= data_nn[1436];
      data_r_1435_sv2v_reg <= data_nn[1435];
      data_r_1434_sv2v_reg <= data_nn[1434];
      data_r_1433_sv2v_reg <= data_nn[1433];
      data_r_1432_sv2v_reg <= data_nn[1432];
      data_r_1431_sv2v_reg <= data_nn[1431];
      data_r_1430_sv2v_reg <= data_nn[1430];
      data_r_1429_sv2v_reg <= data_nn[1429];
      data_r_1428_sv2v_reg <= data_nn[1428];
      data_r_1427_sv2v_reg <= data_nn[1427];
      data_r_1426_sv2v_reg <= data_nn[1426];
      data_r_1425_sv2v_reg <= data_nn[1425];
      data_r_1424_sv2v_reg <= data_nn[1424];
      data_r_1423_sv2v_reg <= data_nn[1423];
      data_r_1422_sv2v_reg <= data_nn[1422];
      data_r_1421_sv2v_reg <= data_nn[1421];
      data_r_1420_sv2v_reg <= data_nn[1420];
      data_r_1419_sv2v_reg <= data_nn[1419];
      data_r_1418_sv2v_reg <= data_nn[1418];
      data_r_1417_sv2v_reg <= data_nn[1417];
      data_r_1416_sv2v_reg <= data_nn[1416];
      data_r_1415_sv2v_reg <= data_nn[1415];
      data_r_1414_sv2v_reg <= data_nn[1414];
      data_r_1413_sv2v_reg <= data_nn[1413];
      data_r_1412_sv2v_reg <= data_nn[1412];
      data_r_1411_sv2v_reg <= data_nn[1411];
      data_r_1410_sv2v_reg <= data_nn[1410];
      data_r_1409_sv2v_reg <= data_nn[1409];
      data_r_1408_sv2v_reg <= data_nn[1408];
      data_r_1407_sv2v_reg <= data_nn[1407];
      data_r_1406_sv2v_reg <= data_nn[1406];
      data_r_1405_sv2v_reg <= data_nn[1405];
      data_r_1404_sv2v_reg <= data_nn[1404];
      data_r_1403_sv2v_reg <= data_nn[1403];
      data_r_1402_sv2v_reg <= data_nn[1402];
      data_r_1401_sv2v_reg <= data_nn[1401];
      data_r_1400_sv2v_reg <= data_nn[1400];
      data_r_1399_sv2v_reg <= data_nn[1399];
      data_r_1398_sv2v_reg <= data_nn[1398];
      data_r_1397_sv2v_reg <= data_nn[1397];
      data_r_1396_sv2v_reg <= data_nn[1396];
      data_r_1395_sv2v_reg <= data_nn[1395];
      data_r_1394_sv2v_reg <= data_nn[1394];
      data_r_1393_sv2v_reg <= data_nn[1393];
      data_r_1392_sv2v_reg <= data_nn[1392];
      data_r_1391_sv2v_reg <= data_nn[1391];
      data_r_1390_sv2v_reg <= data_nn[1390];
      data_r_1389_sv2v_reg <= data_nn[1389];
      data_r_1388_sv2v_reg <= data_nn[1388];
      data_r_1387_sv2v_reg <= data_nn[1387];
      data_r_1386_sv2v_reg <= data_nn[1386];
      data_r_1385_sv2v_reg <= data_nn[1385];
      data_r_1384_sv2v_reg <= data_nn[1384];
      data_r_1383_sv2v_reg <= data_nn[1383];
      data_r_1382_sv2v_reg <= data_nn[1382];
      data_r_1381_sv2v_reg <= data_nn[1381];
      data_r_1380_sv2v_reg <= data_nn[1380];
      data_r_1379_sv2v_reg <= data_nn[1379];
      data_r_1378_sv2v_reg <= data_nn[1378];
      data_r_1377_sv2v_reg <= data_nn[1377];
      data_r_1376_sv2v_reg <= data_nn[1376];
      data_r_1375_sv2v_reg <= data_nn[1375];
      data_r_1374_sv2v_reg <= data_nn[1374];
      data_r_1373_sv2v_reg <= data_nn[1373];
      data_r_1372_sv2v_reg <= data_nn[1372];
      data_r_1371_sv2v_reg <= data_nn[1371];
      data_r_1370_sv2v_reg <= data_nn[1370];
      data_r_1369_sv2v_reg <= data_nn[1369];
      data_r_1368_sv2v_reg <= data_nn[1368];
      data_r_1367_sv2v_reg <= data_nn[1367];
      data_r_1366_sv2v_reg <= data_nn[1366];
      data_r_1365_sv2v_reg <= data_nn[1365];
      data_r_1364_sv2v_reg <= data_nn[1364];
      data_r_1363_sv2v_reg <= data_nn[1363];
      data_r_1362_sv2v_reg <= data_nn[1362];
      data_r_1361_sv2v_reg <= data_nn[1361];
      data_r_1360_sv2v_reg <= data_nn[1360];
      data_r_1359_sv2v_reg <= data_nn[1359];
      data_r_1358_sv2v_reg <= data_nn[1358];
      data_r_1357_sv2v_reg <= data_nn[1357];
      data_r_1356_sv2v_reg <= data_nn[1356];
      data_r_1355_sv2v_reg <= data_nn[1355];
      data_r_1354_sv2v_reg <= data_nn[1354];
      data_r_1353_sv2v_reg <= data_nn[1353];
      data_r_1352_sv2v_reg <= data_nn[1352];
      data_r_1351_sv2v_reg <= data_nn[1351];
      data_r_1350_sv2v_reg <= data_nn[1350];
      data_r_1349_sv2v_reg <= data_nn[1349];
      data_r_1348_sv2v_reg <= data_nn[1348];
      data_r_1347_sv2v_reg <= data_nn[1347];
      data_r_1346_sv2v_reg <= data_nn[1346];
      data_r_1345_sv2v_reg <= data_nn[1345];
      data_r_1344_sv2v_reg <= data_nn[1344];
      data_r_1343_sv2v_reg <= data_nn[1343];
      data_r_1342_sv2v_reg <= data_nn[1342];
      data_r_1341_sv2v_reg <= data_nn[1341];
      data_r_1340_sv2v_reg <= data_nn[1340];
      data_r_1339_sv2v_reg <= data_nn[1339];
      data_r_1338_sv2v_reg <= data_nn[1338];
      data_r_1337_sv2v_reg <= data_nn[1337];
      data_r_1336_sv2v_reg <= data_nn[1336];
      data_r_1335_sv2v_reg <= data_nn[1335];
      data_r_1334_sv2v_reg <= data_nn[1334];
      data_r_1333_sv2v_reg <= data_nn[1333];
      data_r_1332_sv2v_reg <= data_nn[1332];
      data_r_1331_sv2v_reg <= data_nn[1331];
      data_r_1330_sv2v_reg <= data_nn[1330];
      data_r_1329_sv2v_reg <= data_nn[1329];
      data_r_1328_sv2v_reg <= data_nn[1328];
      data_r_1327_sv2v_reg <= data_nn[1327];
      data_r_1326_sv2v_reg <= data_nn[1326];
      data_r_1325_sv2v_reg <= data_nn[1325];
      data_r_1324_sv2v_reg <= data_nn[1324];
      data_r_1323_sv2v_reg <= data_nn[1323];
      data_r_1322_sv2v_reg <= data_nn[1322];
      data_r_1321_sv2v_reg <= data_nn[1321];
      data_r_1320_sv2v_reg <= data_nn[1320];
      data_r_1319_sv2v_reg <= data_nn[1319];
      data_r_1318_sv2v_reg <= data_nn[1318];
      data_r_1317_sv2v_reg <= data_nn[1317];
      data_r_1316_sv2v_reg <= data_nn[1316];
      data_r_1315_sv2v_reg <= data_nn[1315];
      data_r_1314_sv2v_reg <= data_nn[1314];
      data_r_1313_sv2v_reg <= data_nn[1313];
      data_r_1312_sv2v_reg <= data_nn[1312];
      data_r_1311_sv2v_reg <= data_nn[1311];
      data_r_1310_sv2v_reg <= data_nn[1310];
      data_r_1309_sv2v_reg <= data_nn[1309];
      data_r_1308_sv2v_reg <= data_nn[1308];
      data_r_1307_sv2v_reg <= data_nn[1307];
      data_r_1306_sv2v_reg <= data_nn[1306];
      data_r_1305_sv2v_reg <= data_nn[1305];
      data_r_1304_sv2v_reg <= data_nn[1304];
      data_r_1303_sv2v_reg <= data_nn[1303];
      data_r_1302_sv2v_reg <= data_nn[1302];
      data_r_1301_sv2v_reg <= data_nn[1301];
      data_r_1300_sv2v_reg <= data_nn[1300];
      data_r_1299_sv2v_reg <= data_nn[1299];
      data_r_1298_sv2v_reg <= data_nn[1298];
      data_r_1297_sv2v_reg <= data_nn[1297];
      data_r_1296_sv2v_reg <= data_nn[1296];
      data_r_1295_sv2v_reg <= data_nn[1295];
      data_r_1294_sv2v_reg <= data_nn[1294];
      data_r_1293_sv2v_reg <= data_nn[1293];
      data_r_1292_sv2v_reg <= data_nn[1292];
      data_r_1291_sv2v_reg <= data_nn[1291];
      data_r_1290_sv2v_reg <= data_nn[1290];
      data_r_1289_sv2v_reg <= data_nn[1289];
      data_r_1288_sv2v_reg <= data_nn[1288];
      data_r_1287_sv2v_reg <= data_nn[1287];
      data_r_1286_sv2v_reg <= data_nn[1286];
      data_r_1285_sv2v_reg <= data_nn[1285];
      data_r_1284_sv2v_reg <= data_nn[1284];
      data_r_1283_sv2v_reg <= data_nn[1283];
      data_r_1282_sv2v_reg <= data_nn[1282];
      data_r_1281_sv2v_reg <= data_nn[1281];
      data_r_1280_sv2v_reg <= data_nn[1280];
      data_r_1279_sv2v_reg <= data_nn[1279];
      data_r_1278_sv2v_reg <= data_nn[1278];
      data_r_1277_sv2v_reg <= data_nn[1277];
      data_r_1276_sv2v_reg <= data_nn[1276];
      data_r_1275_sv2v_reg <= data_nn[1275];
      data_r_1274_sv2v_reg <= data_nn[1274];
      data_r_1273_sv2v_reg <= data_nn[1273];
      data_r_1272_sv2v_reg <= data_nn[1272];
      data_r_1271_sv2v_reg <= data_nn[1271];
      data_r_1270_sv2v_reg <= data_nn[1270];
      data_r_1269_sv2v_reg <= data_nn[1269];
      data_r_1268_sv2v_reg <= data_nn[1268];
      data_r_1267_sv2v_reg <= data_nn[1267];
      data_r_1266_sv2v_reg <= data_nn[1266];
      data_r_1265_sv2v_reg <= data_nn[1265];
      data_r_1264_sv2v_reg <= data_nn[1264];
      data_r_1263_sv2v_reg <= data_nn[1263];
      data_r_1262_sv2v_reg <= data_nn[1262];
      data_r_1261_sv2v_reg <= data_nn[1261];
      data_r_1260_sv2v_reg <= data_nn[1260];
      data_r_1259_sv2v_reg <= data_nn[1259];
      data_r_1258_sv2v_reg <= data_nn[1258];
      data_r_1257_sv2v_reg <= data_nn[1257];
      data_r_1256_sv2v_reg <= data_nn[1256];
      data_r_1255_sv2v_reg <= data_nn[1255];
      data_r_1254_sv2v_reg <= data_nn[1254];
      data_r_1253_sv2v_reg <= data_nn[1253];
      data_r_1252_sv2v_reg <= data_nn[1252];
      data_r_1251_sv2v_reg <= data_nn[1251];
      data_r_1250_sv2v_reg <= data_nn[1250];
      data_r_1249_sv2v_reg <= data_nn[1249];
      data_r_1248_sv2v_reg <= data_nn[1248];
      data_r_1247_sv2v_reg <= data_nn[1247];
      data_r_1246_sv2v_reg <= data_nn[1246];
      data_r_1245_sv2v_reg <= data_nn[1245];
      data_r_1244_sv2v_reg <= data_nn[1244];
      data_r_1243_sv2v_reg <= data_nn[1243];
      data_r_1242_sv2v_reg <= data_nn[1242];
      data_r_1241_sv2v_reg <= data_nn[1241];
      data_r_1240_sv2v_reg <= data_nn[1240];
      data_r_1239_sv2v_reg <= data_nn[1239];
      data_r_1238_sv2v_reg <= data_nn[1238];
      data_r_1237_sv2v_reg <= data_nn[1237];
      data_r_1236_sv2v_reg <= data_nn[1236];
      data_r_1235_sv2v_reg <= data_nn[1235];
      data_r_1234_sv2v_reg <= data_nn[1234];
      data_r_1233_sv2v_reg <= data_nn[1233];
      data_r_1232_sv2v_reg <= data_nn[1232];
      data_r_1231_sv2v_reg <= data_nn[1231];
      data_r_1230_sv2v_reg <= data_nn[1230];
      data_r_1229_sv2v_reg <= data_nn[1229];
      data_r_1228_sv2v_reg <= data_nn[1228];
      data_r_1227_sv2v_reg <= data_nn[1227];
      data_r_1226_sv2v_reg <= data_nn[1226];
      data_r_1225_sv2v_reg <= data_nn[1225];
      data_r_1224_sv2v_reg <= data_nn[1224];
      data_r_1223_sv2v_reg <= data_nn[1223];
      data_r_1222_sv2v_reg <= data_nn[1222];
      data_r_1221_sv2v_reg <= data_nn[1221];
      data_r_1220_sv2v_reg <= data_nn[1220];
      data_r_1219_sv2v_reg <= data_nn[1219];
      data_r_1218_sv2v_reg <= data_nn[1218];
      data_r_1217_sv2v_reg <= data_nn[1217];
      data_r_1216_sv2v_reg <= data_nn[1216];
      data_r_1215_sv2v_reg <= data_nn[1215];
      data_r_1214_sv2v_reg <= data_nn[1214];
      data_r_1213_sv2v_reg <= data_nn[1213];
      data_r_1212_sv2v_reg <= data_nn[1212];
      data_r_1211_sv2v_reg <= data_nn[1211];
      data_r_1210_sv2v_reg <= data_nn[1210];
      data_r_1209_sv2v_reg <= data_nn[1209];
      data_r_1208_sv2v_reg <= data_nn[1208];
      data_r_1207_sv2v_reg <= data_nn[1207];
      data_r_1206_sv2v_reg <= data_nn[1206];
      data_r_1205_sv2v_reg <= data_nn[1205];
      data_r_1204_sv2v_reg <= data_nn[1204];
      data_r_1203_sv2v_reg <= data_nn[1203];
      data_r_1202_sv2v_reg <= data_nn[1202];
      data_r_1201_sv2v_reg <= data_nn[1201];
      data_r_1200_sv2v_reg <= data_nn[1200];
      data_r_1199_sv2v_reg <= data_nn[1199];
      data_r_1198_sv2v_reg <= data_nn[1198];
      data_r_1197_sv2v_reg <= data_nn[1197];
      data_r_1196_sv2v_reg <= data_nn[1196];
      data_r_1195_sv2v_reg <= data_nn[1195];
      data_r_1194_sv2v_reg <= data_nn[1194];
      data_r_1193_sv2v_reg <= data_nn[1193];
      data_r_1192_sv2v_reg <= data_nn[1192];
      data_r_1191_sv2v_reg <= data_nn[1191];
      data_r_1190_sv2v_reg <= data_nn[1190];
      data_r_1189_sv2v_reg <= data_nn[1189];
      data_r_1188_sv2v_reg <= data_nn[1188];
      data_r_1187_sv2v_reg <= data_nn[1187];
      data_r_1186_sv2v_reg <= data_nn[1186];
      data_r_1185_sv2v_reg <= data_nn[1185];
      data_r_1184_sv2v_reg <= data_nn[1184];
      data_r_1183_sv2v_reg <= data_nn[1183];
      data_r_1182_sv2v_reg <= data_nn[1182];
      data_r_1181_sv2v_reg <= data_nn[1181];
      data_r_1180_sv2v_reg <= data_nn[1180];
      data_r_1179_sv2v_reg <= data_nn[1179];
      data_r_1178_sv2v_reg <= data_nn[1178];
      data_r_1177_sv2v_reg <= data_nn[1177];
      data_r_1176_sv2v_reg <= data_nn[1176];
      data_r_1175_sv2v_reg <= data_nn[1175];
      data_r_1174_sv2v_reg <= data_nn[1174];
      data_r_1173_sv2v_reg <= data_nn[1173];
      data_r_1172_sv2v_reg <= data_nn[1172];
      data_r_1171_sv2v_reg <= data_nn[1171];
      data_r_1170_sv2v_reg <= data_nn[1170];
      data_r_1169_sv2v_reg <= data_nn[1169];
      data_r_1168_sv2v_reg <= data_nn[1168];
      data_r_1167_sv2v_reg <= data_nn[1167];
      data_r_1166_sv2v_reg <= data_nn[1166];
      data_r_1165_sv2v_reg <= data_nn[1165];
      data_r_1164_sv2v_reg <= data_nn[1164];
      data_r_1163_sv2v_reg <= data_nn[1163];
      data_r_1162_sv2v_reg <= data_nn[1162];
      data_r_1161_sv2v_reg <= data_nn[1161];
      data_r_1160_sv2v_reg <= data_nn[1160];
      data_r_1159_sv2v_reg <= data_nn[1159];
      data_r_1158_sv2v_reg <= data_nn[1158];
      data_r_1157_sv2v_reg <= data_nn[1157];
      data_r_1156_sv2v_reg <= data_nn[1156];
      data_r_1155_sv2v_reg <= data_nn[1155];
      data_r_1154_sv2v_reg <= data_nn[1154];
      data_r_1153_sv2v_reg <= data_nn[1153];
      data_r_1152_sv2v_reg <= data_nn[1152];
      data_r_1151_sv2v_reg <= data_nn[1151];
      data_r_1150_sv2v_reg <= data_nn[1150];
      data_r_1149_sv2v_reg <= data_nn[1149];
      data_r_1148_sv2v_reg <= data_nn[1148];
      data_r_1147_sv2v_reg <= data_nn[1147];
      data_r_1146_sv2v_reg <= data_nn[1146];
      data_r_1145_sv2v_reg <= data_nn[1145];
      data_r_1144_sv2v_reg <= data_nn[1144];
      data_r_1143_sv2v_reg <= data_nn[1143];
      data_r_1142_sv2v_reg <= data_nn[1142];
      data_r_1141_sv2v_reg <= data_nn[1141];
      data_r_1140_sv2v_reg <= data_nn[1140];
      data_r_1139_sv2v_reg <= data_nn[1139];
      data_r_1138_sv2v_reg <= data_nn[1138];
      data_r_1137_sv2v_reg <= data_nn[1137];
      data_r_1136_sv2v_reg <= data_nn[1136];
      data_r_1135_sv2v_reg <= data_nn[1135];
      data_r_1134_sv2v_reg <= data_nn[1134];
      data_r_1133_sv2v_reg <= data_nn[1133];
      data_r_1132_sv2v_reg <= data_nn[1132];
      data_r_1131_sv2v_reg <= data_nn[1131];
      data_r_1130_sv2v_reg <= data_nn[1130];
      data_r_1129_sv2v_reg <= data_nn[1129];
      data_r_1128_sv2v_reg <= data_nn[1128];
      data_r_1127_sv2v_reg <= data_nn[1127];
      data_r_1126_sv2v_reg <= data_nn[1126];
      data_r_1125_sv2v_reg <= data_nn[1125];
      data_r_1124_sv2v_reg <= data_nn[1124];
      data_r_1123_sv2v_reg <= data_nn[1123];
      data_r_1122_sv2v_reg <= data_nn[1122];
      data_r_1121_sv2v_reg <= data_nn[1121];
      data_r_1120_sv2v_reg <= data_nn[1120];
      data_r_1119_sv2v_reg <= data_nn[1119];
      data_r_1118_sv2v_reg <= data_nn[1118];
      data_r_1117_sv2v_reg <= data_nn[1117];
      data_r_1116_sv2v_reg <= data_nn[1116];
      data_r_1115_sv2v_reg <= data_nn[1115];
      data_r_1114_sv2v_reg <= data_nn[1114];
      data_r_1113_sv2v_reg <= data_nn[1113];
      data_r_1112_sv2v_reg <= data_nn[1112];
      data_r_1111_sv2v_reg <= data_nn[1111];
      data_r_1110_sv2v_reg <= data_nn[1110];
      data_r_1109_sv2v_reg <= data_nn[1109];
      data_r_1108_sv2v_reg <= data_nn[1108];
      data_r_1107_sv2v_reg <= data_nn[1107];
      data_r_1106_sv2v_reg <= data_nn[1106];
      data_r_1105_sv2v_reg <= data_nn[1105];
      data_r_1104_sv2v_reg <= data_nn[1104];
      data_r_1103_sv2v_reg <= data_nn[1103];
      data_r_1102_sv2v_reg <= data_nn[1102];
      data_r_1101_sv2v_reg <= data_nn[1101];
      data_r_1100_sv2v_reg <= data_nn[1100];
      data_r_1099_sv2v_reg <= data_nn[1099];
      data_r_1098_sv2v_reg <= data_nn[1098];
      data_r_1097_sv2v_reg <= data_nn[1097];
      data_r_1096_sv2v_reg <= data_nn[1096];
      data_r_1095_sv2v_reg <= data_nn[1095];
      data_r_1094_sv2v_reg <= data_nn[1094];
      data_r_1093_sv2v_reg <= data_nn[1093];
      data_r_1092_sv2v_reg <= data_nn[1092];
      data_r_1091_sv2v_reg <= data_nn[1091];
      data_r_1090_sv2v_reg <= data_nn[1090];
      data_r_1089_sv2v_reg <= data_nn[1089];
      data_r_1088_sv2v_reg <= data_nn[1088];
      data_r_1087_sv2v_reg <= data_nn[1087];
      data_r_1086_sv2v_reg <= data_nn[1086];
      data_r_1085_sv2v_reg <= data_nn[1085];
      data_r_1084_sv2v_reg <= data_nn[1084];
      data_r_1083_sv2v_reg <= data_nn[1083];
      data_r_1082_sv2v_reg <= data_nn[1082];
      data_r_1081_sv2v_reg <= data_nn[1081];
      data_r_1080_sv2v_reg <= data_nn[1080];
      data_r_1079_sv2v_reg <= data_nn[1079];
      data_r_1078_sv2v_reg <= data_nn[1078];
      data_r_1077_sv2v_reg <= data_nn[1077];
      data_r_1076_sv2v_reg <= data_nn[1076];
      data_r_1075_sv2v_reg <= data_nn[1075];
      data_r_1074_sv2v_reg <= data_nn[1074];
      data_r_1073_sv2v_reg <= data_nn[1073];
      data_r_1072_sv2v_reg <= data_nn[1072];
      data_r_1071_sv2v_reg <= data_nn[1071];
      data_r_1070_sv2v_reg <= data_nn[1070];
      data_r_1069_sv2v_reg <= data_nn[1069];
      data_r_1068_sv2v_reg <= data_nn[1068];
      data_r_1067_sv2v_reg <= data_nn[1067];
      data_r_1066_sv2v_reg <= data_nn[1066];
      data_r_1065_sv2v_reg <= data_nn[1065];
      data_r_1064_sv2v_reg <= data_nn[1064];
      data_r_1063_sv2v_reg <= data_nn[1063];
      data_r_1062_sv2v_reg <= data_nn[1062];
      data_r_1061_sv2v_reg <= data_nn[1061];
      data_r_1060_sv2v_reg <= data_nn[1060];
      data_r_1059_sv2v_reg <= data_nn[1059];
      data_r_1058_sv2v_reg <= data_nn[1058];
      data_r_1057_sv2v_reg <= data_nn[1057];
      data_r_1056_sv2v_reg <= data_nn[1056];
      data_r_1055_sv2v_reg <= data_nn[1055];
      data_r_1054_sv2v_reg <= data_nn[1054];
      data_r_1053_sv2v_reg <= data_nn[1053];
      data_r_1052_sv2v_reg <= data_nn[1052];
      data_r_1051_sv2v_reg <= data_nn[1051];
      data_r_1050_sv2v_reg <= data_nn[1050];
      data_r_1049_sv2v_reg <= data_nn[1049];
      data_r_1048_sv2v_reg <= data_nn[1048];
      data_r_1047_sv2v_reg <= data_nn[1047];
      data_r_1046_sv2v_reg <= data_nn[1046];
      data_r_1045_sv2v_reg <= data_nn[1045];
      data_r_1044_sv2v_reg <= data_nn[1044];
      data_r_1043_sv2v_reg <= data_nn[1043];
      data_r_1042_sv2v_reg <= data_nn[1042];
      data_r_1041_sv2v_reg <= data_nn[1041];
      data_r_1040_sv2v_reg <= data_nn[1040];
      data_r_1039_sv2v_reg <= data_nn[1039];
      data_r_1038_sv2v_reg <= data_nn[1038];
      data_r_1037_sv2v_reg <= data_nn[1037];
      data_r_1036_sv2v_reg <= data_nn[1036];
      data_r_1035_sv2v_reg <= data_nn[1035];
      data_r_1034_sv2v_reg <= data_nn[1034];
      data_r_1033_sv2v_reg <= data_nn[1033];
      data_r_1032_sv2v_reg <= data_nn[1032];
      data_r_1031_sv2v_reg <= data_nn[1031];
      data_r_1030_sv2v_reg <= data_nn[1030];
      data_r_1029_sv2v_reg <= data_nn[1029];
      data_r_1028_sv2v_reg <= data_nn[1028];
      data_r_1027_sv2v_reg <= data_nn[1027];
      data_r_1026_sv2v_reg <= data_nn[1026];
      data_r_1025_sv2v_reg <= data_nn[1025];
      data_r_1024_sv2v_reg <= data_nn[1024];
      data_r_1023_sv2v_reg <= data_nn[1023];
      data_r_1022_sv2v_reg <= data_nn[1022];
      data_r_1021_sv2v_reg <= data_nn[1021];
      data_r_1020_sv2v_reg <= data_nn[1020];
      data_r_1019_sv2v_reg <= data_nn[1019];
      data_r_1018_sv2v_reg <= data_nn[1018];
      data_r_1017_sv2v_reg <= data_nn[1017];
      data_r_1016_sv2v_reg <= data_nn[1016];
      data_r_1015_sv2v_reg <= data_nn[1015];
      data_r_1014_sv2v_reg <= data_nn[1014];
      data_r_1013_sv2v_reg <= data_nn[1013];
      data_r_1012_sv2v_reg <= data_nn[1012];
      data_r_1011_sv2v_reg <= data_nn[1011];
      data_r_1010_sv2v_reg <= data_nn[1010];
      data_r_1009_sv2v_reg <= data_nn[1009];
      data_r_1008_sv2v_reg <= data_nn[1008];
      data_r_1007_sv2v_reg <= data_nn[1007];
      data_r_1006_sv2v_reg <= data_nn[1006];
      data_r_1005_sv2v_reg <= data_nn[1005];
      data_r_1004_sv2v_reg <= data_nn[1004];
      data_r_1003_sv2v_reg <= data_nn[1003];
      data_r_1002_sv2v_reg <= data_nn[1002];
      data_r_1001_sv2v_reg <= data_nn[1001];
      data_r_1000_sv2v_reg <= data_nn[1000];
      data_r_999_sv2v_reg <= data_nn[999];
      data_r_998_sv2v_reg <= data_nn[998];
      data_r_997_sv2v_reg <= data_nn[997];
      data_r_996_sv2v_reg <= data_nn[996];
      data_r_995_sv2v_reg <= data_nn[995];
      data_r_994_sv2v_reg <= data_nn[994];
      data_r_993_sv2v_reg <= data_nn[993];
      data_r_992_sv2v_reg <= data_nn[992];
      data_r_991_sv2v_reg <= data_nn[991];
      data_r_990_sv2v_reg <= data_nn[990];
      data_r_989_sv2v_reg <= data_nn[989];
      data_r_988_sv2v_reg <= data_nn[988];
      data_r_987_sv2v_reg <= data_nn[987];
      data_r_986_sv2v_reg <= data_nn[986];
      data_r_985_sv2v_reg <= data_nn[985];
      data_r_984_sv2v_reg <= data_nn[984];
      data_r_983_sv2v_reg <= data_nn[983];
      data_r_982_sv2v_reg <= data_nn[982];
      data_r_981_sv2v_reg <= data_nn[981];
      data_r_980_sv2v_reg <= data_nn[980];
      data_r_979_sv2v_reg <= data_nn[979];
      data_r_978_sv2v_reg <= data_nn[978];
      data_r_977_sv2v_reg <= data_nn[977];
      data_r_976_sv2v_reg <= data_nn[976];
      data_r_975_sv2v_reg <= data_nn[975];
      data_r_974_sv2v_reg <= data_nn[974];
      data_r_973_sv2v_reg <= data_nn[973];
      data_r_972_sv2v_reg <= data_nn[972];
      data_r_971_sv2v_reg <= data_nn[971];
      data_r_970_sv2v_reg <= data_nn[970];
      data_r_969_sv2v_reg <= data_nn[969];
      data_r_968_sv2v_reg <= data_nn[968];
      data_r_967_sv2v_reg <= data_nn[967];
      data_r_966_sv2v_reg <= data_nn[966];
      data_r_965_sv2v_reg <= data_nn[965];
      data_r_964_sv2v_reg <= data_nn[964];
      data_r_963_sv2v_reg <= data_nn[963];
      data_r_962_sv2v_reg <= data_nn[962];
      data_r_961_sv2v_reg <= data_nn[961];
      data_r_960_sv2v_reg <= data_nn[960];
      data_r_959_sv2v_reg <= data_nn[959];
      data_r_958_sv2v_reg <= data_nn[958];
      data_r_957_sv2v_reg <= data_nn[957];
      data_r_956_sv2v_reg <= data_nn[956];
      data_r_955_sv2v_reg <= data_nn[955];
      data_r_954_sv2v_reg <= data_nn[954];
      data_r_953_sv2v_reg <= data_nn[953];
      data_r_952_sv2v_reg <= data_nn[952];
      data_r_951_sv2v_reg <= data_nn[951];
      data_r_950_sv2v_reg <= data_nn[950];
      data_r_949_sv2v_reg <= data_nn[949];
      data_r_948_sv2v_reg <= data_nn[948];
      data_r_947_sv2v_reg <= data_nn[947];
      data_r_946_sv2v_reg <= data_nn[946];
      data_r_945_sv2v_reg <= data_nn[945];
      data_r_944_sv2v_reg <= data_nn[944];
      data_r_943_sv2v_reg <= data_nn[943];
      data_r_942_sv2v_reg <= data_nn[942];
      data_r_941_sv2v_reg <= data_nn[941];
      data_r_940_sv2v_reg <= data_nn[940];
      data_r_939_sv2v_reg <= data_nn[939];
      data_r_938_sv2v_reg <= data_nn[938];
      data_r_937_sv2v_reg <= data_nn[937];
      data_r_936_sv2v_reg <= data_nn[936];
      data_r_935_sv2v_reg <= data_nn[935];
      data_r_934_sv2v_reg <= data_nn[934];
      data_r_933_sv2v_reg <= data_nn[933];
      data_r_932_sv2v_reg <= data_nn[932];
      data_r_931_sv2v_reg <= data_nn[931];
      data_r_930_sv2v_reg <= data_nn[930];
      data_r_929_sv2v_reg <= data_nn[929];
      data_r_928_sv2v_reg <= data_nn[928];
      data_r_927_sv2v_reg <= data_nn[927];
      data_r_926_sv2v_reg <= data_nn[926];
      data_r_925_sv2v_reg <= data_nn[925];
      data_r_924_sv2v_reg <= data_nn[924];
      data_r_923_sv2v_reg <= data_nn[923];
      data_r_922_sv2v_reg <= data_nn[922];
      data_r_921_sv2v_reg <= data_nn[921];
      data_r_920_sv2v_reg <= data_nn[920];
      data_r_919_sv2v_reg <= data_nn[919];
      data_r_918_sv2v_reg <= data_nn[918];
      data_r_917_sv2v_reg <= data_nn[917];
      data_r_916_sv2v_reg <= data_nn[916];
      data_r_915_sv2v_reg <= data_nn[915];
      data_r_914_sv2v_reg <= data_nn[914];
      data_r_913_sv2v_reg <= data_nn[913];
      data_r_912_sv2v_reg <= data_nn[912];
      data_r_911_sv2v_reg <= data_nn[911];
      data_r_910_sv2v_reg <= data_nn[910];
      data_r_909_sv2v_reg <= data_nn[909];
      data_r_908_sv2v_reg <= data_nn[908];
      data_r_907_sv2v_reg <= data_nn[907];
      data_r_906_sv2v_reg <= data_nn[906];
      data_r_905_sv2v_reg <= data_nn[905];
      data_r_904_sv2v_reg <= data_nn[904];
      data_r_903_sv2v_reg <= data_nn[903];
      data_r_902_sv2v_reg <= data_nn[902];
      data_r_901_sv2v_reg <= data_nn[901];
      data_r_900_sv2v_reg <= data_nn[900];
      data_r_899_sv2v_reg <= data_nn[899];
      data_r_898_sv2v_reg <= data_nn[898];
      data_r_897_sv2v_reg <= data_nn[897];
      data_r_896_sv2v_reg <= data_nn[896];
      data_r_895_sv2v_reg <= data_nn[895];
      data_r_894_sv2v_reg <= data_nn[894];
      data_r_893_sv2v_reg <= data_nn[893];
      data_r_892_sv2v_reg <= data_nn[892];
      data_r_891_sv2v_reg <= data_nn[891];
      data_r_890_sv2v_reg <= data_nn[890];
      data_r_889_sv2v_reg <= data_nn[889];
      data_r_888_sv2v_reg <= data_nn[888];
      data_r_887_sv2v_reg <= data_nn[887];
      data_r_886_sv2v_reg <= data_nn[886];
      data_r_885_sv2v_reg <= data_nn[885];
      data_r_884_sv2v_reg <= data_nn[884];
      data_r_883_sv2v_reg <= data_nn[883];
      data_r_882_sv2v_reg <= data_nn[882];
      data_r_881_sv2v_reg <= data_nn[881];
      data_r_880_sv2v_reg <= data_nn[880];
      data_r_879_sv2v_reg <= data_nn[879];
      data_r_878_sv2v_reg <= data_nn[878];
      data_r_877_sv2v_reg <= data_nn[877];
      data_r_876_sv2v_reg <= data_nn[876];
      data_r_875_sv2v_reg <= data_nn[875];
      data_r_874_sv2v_reg <= data_nn[874];
      data_r_873_sv2v_reg <= data_nn[873];
      data_r_872_sv2v_reg <= data_nn[872];
      data_r_871_sv2v_reg <= data_nn[871];
      data_r_870_sv2v_reg <= data_nn[870];
      data_r_869_sv2v_reg <= data_nn[869];
      data_r_868_sv2v_reg <= data_nn[868];
      data_r_867_sv2v_reg <= data_nn[867];
      data_r_866_sv2v_reg <= data_nn[866];
      data_r_865_sv2v_reg <= data_nn[865];
      data_r_864_sv2v_reg <= data_nn[864];
      data_r_863_sv2v_reg <= data_nn[863];
      data_r_862_sv2v_reg <= data_nn[862];
      data_r_861_sv2v_reg <= data_nn[861];
      data_r_860_sv2v_reg <= data_nn[860];
      data_r_859_sv2v_reg <= data_nn[859];
      data_r_858_sv2v_reg <= data_nn[858];
      data_r_857_sv2v_reg <= data_nn[857];
      data_r_856_sv2v_reg <= data_nn[856];
      data_r_855_sv2v_reg <= data_nn[855];
      data_r_854_sv2v_reg <= data_nn[854];
      data_r_853_sv2v_reg <= data_nn[853];
      data_r_852_sv2v_reg <= data_nn[852];
      data_r_851_sv2v_reg <= data_nn[851];
      data_r_850_sv2v_reg <= data_nn[850];
      data_r_849_sv2v_reg <= data_nn[849];
      data_r_848_sv2v_reg <= data_nn[848];
      data_r_847_sv2v_reg <= data_nn[847];
      data_r_846_sv2v_reg <= data_nn[846];
      data_r_845_sv2v_reg <= data_nn[845];
      data_r_844_sv2v_reg <= data_nn[844];
      data_r_843_sv2v_reg <= data_nn[843];
      data_r_842_sv2v_reg <= data_nn[842];
      data_r_841_sv2v_reg <= data_nn[841];
      data_r_840_sv2v_reg <= data_nn[840];
      data_r_839_sv2v_reg <= data_nn[839];
      data_r_838_sv2v_reg <= data_nn[838];
      data_r_837_sv2v_reg <= data_nn[837];
      data_r_836_sv2v_reg <= data_nn[836];
      data_r_835_sv2v_reg <= data_nn[835];
      data_r_834_sv2v_reg <= data_nn[834];
      data_r_833_sv2v_reg <= data_nn[833];
      data_r_832_sv2v_reg <= data_nn[832];
      data_r_831_sv2v_reg <= data_nn[831];
      data_r_830_sv2v_reg <= data_nn[830];
      data_r_829_sv2v_reg <= data_nn[829];
      data_r_828_sv2v_reg <= data_nn[828];
      data_r_827_sv2v_reg <= data_nn[827];
      data_r_826_sv2v_reg <= data_nn[826];
      data_r_825_sv2v_reg <= data_nn[825];
      data_r_824_sv2v_reg <= data_nn[824];
      data_r_823_sv2v_reg <= data_nn[823];
      data_r_822_sv2v_reg <= data_nn[822];
      data_r_821_sv2v_reg <= data_nn[821];
      data_r_820_sv2v_reg <= data_nn[820];
      data_r_819_sv2v_reg <= data_nn[819];
      data_r_818_sv2v_reg <= data_nn[818];
      data_r_817_sv2v_reg <= data_nn[817];
      data_r_816_sv2v_reg <= data_nn[816];
      data_r_815_sv2v_reg <= data_nn[815];
      data_r_814_sv2v_reg <= data_nn[814];
      data_r_813_sv2v_reg <= data_nn[813];
      data_r_812_sv2v_reg <= data_nn[812];
      data_r_811_sv2v_reg <= data_nn[811];
      data_r_810_sv2v_reg <= data_nn[810];
      data_r_809_sv2v_reg <= data_nn[809];
      data_r_808_sv2v_reg <= data_nn[808];
      data_r_807_sv2v_reg <= data_nn[807];
      data_r_806_sv2v_reg <= data_nn[806];
      data_r_805_sv2v_reg <= data_nn[805];
      data_r_804_sv2v_reg <= data_nn[804];
      data_r_803_sv2v_reg <= data_nn[803];
      data_r_802_sv2v_reg <= data_nn[802];
      data_r_801_sv2v_reg <= data_nn[801];
      data_r_800_sv2v_reg <= data_nn[800];
      data_r_799_sv2v_reg <= data_nn[799];
      data_r_798_sv2v_reg <= data_nn[798];
      data_r_797_sv2v_reg <= data_nn[797];
      data_r_796_sv2v_reg <= data_nn[796];
      data_r_795_sv2v_reg <= data_nn[795];
      data_r_794_sv2v_reg <= data_nn[794];
      data_r_793_sv2v_reg <= data_nn[793];
      data_r_792_sv2v_reg <= data_nn[792];
      data_r_791_sv2v_reg <= data_nn[791];
      data_r_790_sv2v_reg <= data_nn[790];
      data_r_789_sv2v_reg <= data_nn[789];
      data_r_788_sv2v_reg <= data_nn[788];
      data_r_787_sv2v_reg <= data_nn[787];
      data_r_786_sv2v_reg <= data_nn[786];
      data_r_785_sv2v_reg <= data_nn[785];
      data_r_784_sv2v_reg <= data_nn[784];
      data_r_783_sv2v_reg <= data_nn[783];
      data_r_782_sv2v_reg <= data_nn[782];
      data_r_781_sv2v_reg <= data_nn[781];
      data_r_780_sv2v_reg <= data_nn[780];
      data_r_779_sv2v_reg <= data_nn[779];
      data_r_778_sv2v_reg <= data_nn[778];
      data_r_777_sv2v_reg <= data_nn[777];
      data_r_776_sv2v_reg <= data_nn[776];
      data_r_775_sv2v_reg <= data_nn[775];
      data_r_774_sv2v_reg <= data_nn[774];
      data_r_773_sv2v_reg <= data_nn[773];
      data_r_772_sv2v_reg <= data_nn[772];
      data_r_771_sv2v_reg <= data_nn[771];
      data_r_770_sv2v_reg <= data_nn[770];
      data_r_769_sv2v_reg <= data_nn[769];
      data_r_768_sv2v_reg <= data_nn[768];
      data_r_767_sv2v_reg <= data_nn[767];
      data_r_766_sv2v_reg <= data_nn[766];
      data_r_765_sv2v_reg <= data_nn[765];
      data_r_764_sv2v_reg <= data_nn[764];
      data_r_763_sv2v_reg <= data_nn[763];
      data_r_762_sv2v_reg <= data_nn[762];
      data_r_761_sv2v_reg <= data_nn[761];
      data_r_760_sv2v_reg <= data_nn[760];
      data_r_759_sv2v_reg <= data_nn[759];
      data_r_758_sv2v_reg <= data_nn[758];
      data_r_757_sv2v_reg <= data_nn[757];
      data_r_756_sv2v_reg <= data_nn[756];
      data_r_755_sv2v_reg <= data_nn[755];
      data_r_754_sv2v_reg <= data_nn[754];
      data_r_753_sv2v_reg <= data_nn[753];
      data_r_752_sv2v_reg <= data_nn[752];
      data_r_751_sv2v_reg <= data_nn[751];
      data_r_750_sv2v_reg <= data_nn[750];
      data_r_749_sv2v_reg <= data_nn[749];
      data_r_748_sv2v_reg <= data_nn[748];
      data_r_747_sv2v_reg <= data_nn[747];
      data_r_746_sv2v_reg <= data_nn[746];
      data_r_745_sv2v_reg <= data_nn[745];
      data_r_744_sv2v_reg <= data_nn[744];
      data_r_743_sv2v_reg <= data_nn[743];
      data_r_742_sv2v_reg <= data_nn[742];
      data_r_741_sv2v_reg <= data_nn[741];
      data_r_740_sv2v_reg <= data_nn[740];
      data_r_739_sv2v_reg <= data_nn[739];
      data_r_738_sv2v_reg <= data_nn[738];
      data_r_737_sv2v_reg <= data_nn[737];
      data_r_736_sv2v_reg <= data_nn[736];
      data_r_735_sv2v_reg <= data_nn[735];
      data_r_734_sv2v_reg <= data_nn[734];
      data_r_733_sv2v_reg <= data_nn[733];
      data_r_732_sv2v_reg <= data_nn[732];
      data_r_731_sv2v_reg <= data_nn[731];
      data_r_730_sv2v_reg <= data_nn[730];
      data_r_729_sv2v_reg <= data_nn[729];
      data_r_728_sv2v_reg <= data_nn[728];
      data_r_727_sv2v_reg <= data_nn[727];
      data_r_726_sv2v_reg <= data_nn[726];
      data_r_725_sv2v_reg <= data_nn[725];
      data_r_724_sv2v_reg <= data_nn[724];
      data_r_723_sv2v_reg <= data_nn[723];
      data_r_722_sv2v_reg <= data_nn[722];
      data_r_721_sv2v_reg <= data_nn[721];
      data_r_720_sv2v_reg <= data_nn[720];
      data_r_719_sv2v_reg <= data_nn[719];
      data_r_718_sv2v_reg <= data_nn[718];
      data_r_717_sv2v_reg <= data_nn[717];
      data_r_716_sv2v_reg <= data_nn[716];
      data_r_715_sv2v_reg <= data_nn[715];
      data_r_714_sv2v_reg <= data_nn[714];
      data_r_713_sv2v_reg <= data_nn[713];
      data_r_712_sv2v_reg <= data_nn[712];
      data_r_711_sv2v_reg <= data_nn[711];
      data_r_710_sv2v_reg <= data_nn[710];
      data_r_709_sv2v_reg <= data_nn[709];
      data_r_708_sv2v_reg <= data_nn[708];
      data_r_707_sv2v_reg <= data_nn[707];
      data_r_706_sv2v_reg <= data_nn[706];
      data_r_705_sv2v_reg <= data_nn[705];
      data_r_704_sv2v_reg <= data_nn[704];
      data_r_703_sv2v_reg <= data_nn[703];
      data_r_702_sv2v_reg <= data_nn[702];
      data_r_701_sv2v_reg <= data_nn[701];
      data_r_700_sv2v_reg <= data_nn[700];
      data_r_699_sv2v_reg <= data_nn[699];
      data_r_698_sv2v_reg <= data_nn[698];
      data_r_697_sv2v_reg <= data_nn[697];
      data_r_696_sv2v_reg <= data_nn[696];
      data_r_695_sv2v_reg <= data_nn[695];
      data_r_694_sv2v_reg <= data_nn[694];
      data_r_693_sv2v_reg <= data_nn[693];
      data_r_692_sv2v_reg <= data_nn[692];
      data_r_691_sv2v_reg <= data_nn[691];
      data_r_690_sv2v_reg <= data_nn[690];
      data_r_689_sv2v_reg <= data_nn[689];
      data_r_688_sv2v_reg <= data_nn[688];
      data_r_687_sv2v_reg <= data_nn[687];
      data_r_686_sv2v_reg <= data_nn[686];
      data_r_685_sv2v_reg <= data_nn[685];
      data_r_684_sv2v_reg <= data_nn[684];
      data_r_683_sv2v_reg <= data_nn[683];
      data_r_682_sv2v_reg <= data_nn[682];
      data_r_681_sv2v_reg <= data_nn[681];
      data_r_680_sv2v_reg <= data_nn[680];
      data_r_679_sv2v_reg <= data_nn[679];
      data_r_678_sv2v_reg <= data_nn[678];
      data_r_677_sv2v_reg <= data_nn[677];
      data_r_676_sv2v_reg <= data_nn[676];
      data_r_675_sv2v_reg <= data_nn[675];
      data_r_674_sv2v_reg <= data_nn[674];
      data_r_673_sv2v_reg <= data_nn[673];
      data_r_672_sv2v_reg <= data_nn[672];
      data_r_671_sv2v_reg <= data_nn[671];
      data_r_670_sv2v_reg <= data_nn[670];
      data_r_669_sv2v_reg <= data_nn[669];
      data_r_668_sv2v_reg <= data_nn[668];
      data_r_667_sv2v_reg <= data_nn[667];
      data_r_666_sv2v_reg <= data_nn[666];
      data_r_665_sv2v_reg <= data_nn[665];
      data_r_664_sv2v_reg <= data_nn[664];
      data_r_663_sv2v_reg <= data_nn[663];
      data_r_662_sv2v_reg <= data_nn[662];
      data_r_661_sv2v_reg <= data_nn[661];
      data_r_660_sv2v_reg <= data_nn[660];
      data_r_659_sv2v_reg <= data_nn[659];
      data_r_658_sv2v_reg <= data_nn[658];
      data_r_657_sv2v_reg <= data_nn[657];
      data_r_656_sv2v_reg <= data_nn[656];
      data_r_655_sv2v_reg <= data_nn[655];
      data_r_654_sv2v_reg <= data_nn[654];
      data_r_653_sv2v_reg <= data_nn[653];
      data_r_652_sv2v_reg <= data_nn[652];
      data_r_651_sv2v_reg <= data_nn[651];
      data_r_650_sv2v_reg <= data_nn[650];
      data_r_649_sv2v_reg <= data_nn[649];
      data_r_648_sv2v_reg <= data_nn[648];
      data_r_647_sv2v_reg <= data_nn[647];
      data_r_646_sv2v_reg <= data_nn[646];
      data_r_645_sv2v_reg <= data_nn[645];
      data_r_644_sv2v_reg <= data_nn[644];
      data_r_643_sv2v_reg <= data_nn[643];
      data_r_642_sv2v_reg <= data_nn[642];
      data_r_641_sv2v_reg <= data_nn[641];
      data_r_640_sv2v_reg <= data_nn[640];
      data_r_639_sv2v_reg <= data_nn[639];
      data_r_638_sv2v_reg <= data_nn[638];
      data_r_637_sv2v_reg <= data_nn[637];
      data_r_636_sv2v_reg <= data_nn[636];
      data_r_635_sv2v_reg <= data_nn[635];
      data_r_634_sv2v_reg <= data_nn[634];
      data_r_633_sv2v_reg <= data_nn[633];
      data_r_632_sv2v_reg <= data_nn[632];
      data_r_631_sv2v_reg <= data_nn[631];
      data_r_630_sv2v_reg <= data_nn[630];
      data_r_629_sv2v_reg <= data_nn[629];
      data_r_628_sv2v_reg <= data_nn[628];
      data_r_627_sv2v_reg <= data_nn[627];
      data_r_626_sv2v_reg <= data_nn[626];
      data_r_625_sv2v_reg <= data_nn[625];
      data_r_624_sv2v_reg <= data_nn[624];
      data_r_623_sv2v_reg <= data_nn[623];
      data_r_622_sv2v_reg <= data_nn[622];
      data_r_621_sv2v_reg <= data_nn[621];
      data_r_620_sv2v_reg <= data_nn[620];
      data_r_619_sv2v_reg <= data_nn[619];
      data_r_618_sv2v_reg <= data_nn[618];
      data_r_617_sv2v_reg <= data_nn[617];
      data_r_616_sv2v_reg <= data_nn[616];
      data_r_615_sv2v_reg <= data_nn[615];
      data_r_614_sv2v_reg <= data_nn[614];
      data_r_613_sv2v_reg <= data_nn[613];
      data_r_612_sv2v_reg <= data_nn[612];
      data_r_611_sv2v_reg <= data_nn[611];
      data_r_610_sv2v_reg <= data_nn[610];
      data_r_609_sv2v_reg <= data_nn[609];
      data_r_608_sv2v_reg <= data_nn[608];
      data_r_607_sv2v_reg <= data_nn[607];
      data_r_606_sv2v_reg <= data_nn[606];
      data_r_605_sv2v_reg <= data_nn[605];
      data_r_604_sv2v_reg <= data_nn[604];
      data_r_603_sv2v_reg <= data_nn[603];
      data_r_602_sv2v_reg <= data_nn[602];
      data_r_601_sv2v_reg <= data_nn[601];
      data_r_600_sv2v_reg <= data_nn[600];
      data_r_599_sv2v_reg <= data_nn[599];
      data_r_598_sv2v_reg <= data_nn[598];
      data_r_597_sv2v_reg <= data_nn[597];
      data_r_596_sv2v_reg <= data_nn[596];
      data_r_595_sv2v_reg <= data_nn[595];
      data_r_594_sv2v_reg <= data_nn[594];
      data_r_593_sv2v_reg <= data_nn[593];
      data_r_592_sv2v_reg <= data_nn[592];
      data_r_591_sv2v_reg <= data_nn[591];
      data_r_590_sv2v_reg <= data_nn[590];
      data_r_589_sv2v_reg <= data_nn[589];
      data_r_588_sv2v_reg <= data_nn[588];
      data_r_587_sv2v_reg <= data_nn[587];
      data_r_586_sv2v_reg <= data_nn[586];
      data_r_585_sv2v_reg <= data_nn[585];
      data_r_584_sv2v_reg <= data_nn[584];
      data_r_583_sv2v_reg <= data_nn[583];
      data_r_582_sv2v_reg <= data_nn[582];
      data_r_581_sv2v_reg <= data_nn[581];
      data_r_580_sv2v_reg <= data_nn[580];
      data_r_579_sv2v_reg <= data_nn[579];
      data_r_578_sv2v_reg <= data_nn[578];
      data_r_577_sv2v_reg <= data_nn[577];
      data_r_576_sv2v_reg <= data_nn[576];
      data_r_575_sv2v_reg <= data_nn[575];
      data_r_574_sv2v_reg <= data_nn[574];
      data_r_573_sv2v_reg <= data_nn[573];
      data_r_572_sv2v_reg <= data_nn[572];
      data_r_571_sv2v_reg <= data_nn[571];
      data_r_570_sv2v_reg <= data_nn[570];
      data_r_569_sv2v_reg <= data_nn[569];
      data_r_568_sv2v_reg <= data_nn[568];
      data_r_567_sv2v_reg <= data_nn[567];
      data_r_566_sv2v_reg <= data_nn[566];
      data_r_565_sv2v_reg <= data_nn[565];
      data_r_564_sv2v_reg <= data_nn[564];
      data_r_563_sv2v_reg <= data_nn[563];
      data_r_562_sv2v_reg <= data_nn[562];
      data_r_561_sv2v_reg <= data_nn[561];
      data_r_560_sv2v_reg <= data_nn[560];
      data_r_559_sv2v_reg <= data_nn[559];
      data_r_558_sv2v_reg <= data_nn[558];
      data_r_557_sv2v_reg <= data_nn[557];
      data_r_556_sv2v_reg <= data_nn[556];
      data_r_555_sv2v_reg <= data_nn[555];
      data_r_554_sv2v_reg <= data_nn[554];
      data_r_553_sv2v_reg <= data_nn[553];
      data_r_552_sv2v_reg <= data_nn[552];
      data_r_551_sv2v_reg <= data_nn[551];
      data_r_550_sv2v_reg <= data_nn[550];
      data_r_549_sv2v_reg <= data_nn[549];
      data_r_548_sv2v_reg <= data_nn[548];
      data_r_547_sv2v_reg <= data_nn[547];
      data_r_546_sv2v_reg <= data_nn[546];
      data_r_545_sv2v_reg <= data_nn[545];
      data_r_544_sv2v_reg <= data_nn[544];
      data_r_543_sv2v_reg <= data_nn[543];
      data_r_542_sv2v_reg <= data_nn[542];
      data_r_541_sv2v_reg <= data_nn[541];
      data_r_540_sv2v_reg <= data_nn[540];
      data_r_539_sv2v_reg <= data_nn[539];
      data_r_538_sv2v_reg <= data_nn[538];
      data_r_537_sv2v_reg <= data_nn[537];
      data_r_536_sv2v_reg <= data_nn[536];
      data_r_535_sv2v_reg <= data_nn[535];
      data_r_534_sv2v_reg <= data_nn[534];
      data_r_533_sv2v_reg <= data_nn[533];
      data_r_532_sv2v_reg <= data_nn[532];
      data_r_531_sv2v_reg <= data_nn[531];
      data_r_530_sv2v_reg <= data_nn[530];
      data_r_529_sv2v_reg <= data_nn[529];
      data_r_528_sv2v_reg <= data_nn[528];
      data_r_527_sv2v_reg <= data_nn[527];
      data_r_526_sv2v_reg <= data_nn[526];
      data_r_525_sv2v_reg <= data_nn[525];
      data_r_524_sv2v_reg <= data_nn[524];
      data_r_523_sv2v_reg <= data_nn[523];
      data_r_522_sv2v_reg <= data_nn[522];
      data_r_521_sv2v_reg <= data_nn[521];
      data_r_520_sv2v_reg <= data_nn[520];
      data_r_519_sv2v_reg <= data_nn[519];
      data_r_518_sv2v_reg <= data_nn[518];
      data_r_517_sv2v_reg <= data_nn[517];
      data_r_516_sv2v_reg <= data_nn[516];
      data_r_515_sv2v_reg <= data_nn[515];
      data_r_514_sv2v_reg <= data_nn[514];
      data_r_513_sv2v_reg <= data_nn[513];
      data_r_512_sv2v_reg <= data_nn[512];
      data_r_511_sv2v_reg <= data_nn[511];
      data_r_510_sv2v_reg <= data_nn[510];
      data_r_509_sv2v_reg <= data_nn[509];
      data_r_508_sv2v_reg <= data_nn[508];
      data_r_507_sv2v_reg <= data_nn[507];
      data_r_506_sv2v_reg <= data_nn[506];
      data_r_505_sv2v_reg <= data_nn[505];
      data_r_504_sv2v_reg <= data_nn[504];
      data_r_503_sv2v_reg <= data_nn[503];
      data_r_502_sv2v_reg <= data_nn[502];
      data_r_501_sv2v_reg <= data_nn[501];
      data_r_500_sv2v_reg <= data_nn[500];
      data_r_499_sv2v_reg <= data_nn[499];
      data_r_498_sv2v_reg <= data_nn[498];
      data_r_497_sv2v_reg <= data_nn[497];
      data_r_496_sv2v_reg <= data_nn[496];
      data_r_495_sv2v_reg <= data_nn[495];
      data_r_494_sv2v_reg <= data_nn[494];
      data_r_493_sv2v_reg <= data_nn[493];
      data_r_492_sv2v_reg <= data_nn[492];
      data_r_491_sv2v_reg <= data_nn[491];
      data_r_490_sv2v_reg <= data_nn[490];
      data_r_489_sv2v_reg <= data_nn[489];
      data_r_488_sv2v_reg <= data_nn[488];
      data_r_487_sv2v_reg <= data_nn[487];
      data_r_486_sv2v_reg <= data_nn[486];
      data_r_485_sv2v_reg <= data_nn[485];
      data_r_484_sv2v_reg <= data_nn[484];
      data_r_483_sv2v_reg <= data_nn[483];
      data_r_482_sv2v_reg <= data_nn[482];
      data_r_481_sv2v_reg <= data_nn[481];
      data_r_480_sv2v_reg <= data_nn[480];
      data_r_479_sv2v_reg <= data_nn[479];
      data_r_478_sv2v_reg <= data_nn[478];
      data_r_477_sv2v_reg <= data_nn[477];
      data_r_476_sv2v_reg <= data_nn[476];
      data_r_475_sv2v_reg <= data_nn[475];
      data_r_474_sv2v_reg <= data_nn[474];
      data_r_473_sv2v_reg <= data_nn[473];
      data_r_472_sv2v_reg <= data_nn[472];
      data_r_471_sv2v_reg <= data_nn[471];
      data_r_470_sv2v_reg <= data_nn[470];
      data_r_469_sv2v_reg <= data_nn[469];
      data_r_468_sv2v_reg <= data_nn[468];
      data_r_467_sv2v_reg <= data_nn[467];
      data_r_466_sv2v_reg <= data_nn[466];
      data_r_465_sv2v_reg <= data_nn[465];
      data_r_464_sv2v_reg <= data_nn[464];
      data_r_463_sv2v_reg <= data_nn[463];
      data_r_462_sv2v_reg <= data_nn[462];
      data_r_461_sv2v_reg <= data_nn[461];
      data_r_460_sv2v_reg <= data_nn[460];
      data_r_459_sv2v_reg <= data_nn[459];
      data_r_458_sv2v_reg <= data_nn[458];
      data_r_457_sv2v_reg <= data_nn[457];
      data_r_456_sv2v_reg <= data_nn[456];
      data_r_455_sv2v_reg <= data_nn[455];
      data_r_454_sv2v_reg <= data_nn[454];
      data_r_453_sv2v_reg <= data_nn[453];
      data_r_452_sv2v_reg <= data_nn[452];
      data_r_451_sv2v_reg <= data_nn[451];
      data_r_450_sv2v_reg <= data_nn[450];
      data_r_449_sv2v_reg <= data_nn[449];
      data_r_448_sv2v_reg <= data_nn[448];
      data_r_447_sv2v_reg <= data_nn[447];
      data_r_446_sv2v_reg <= data_nn[446];
      data_r_445_sv2v_reg <= data_nn[445];
      data_r_444_sv2v_reg <= data_nn[444];
      data_r_443_sv2v_reg <= data_nn[443];
      data_r_442_sv2v_reg <= data_nn[442];
      data_r_441_sv2v_reg <= data_nn[441];
      data_r_440_sv2v_reg <= data_nn[440];
      data_r_439_sv2v_reg <= data_nn[439];
      data_r_438_sv2v_reg <= data_nn[438];
      data_r_437_sv2v_reg <= data_nn[437];
      data_r_436_sv2v_reg <= data_nn[436];
      data_r_435_sv2v_reg <= data_nn[435];
      data_r_434_sv2v_reg <= data_nn[434];
      data_r_433_sv2v_reg <= data_nn[433];
      data_r_432_sv2v_reg <= data_nn[432];
      data_r_431_sv2v_reg <= data_nn[431];
      data_r_430_sv2v_reg <= data_nn[430];
      data_r_429_sv2v_reg <= data_nn[429];
      data_r_428_sv2v_reg <= data_nn[428];
      data_r_427_sv2v_reg <= data_nn[427];
      data_r_426_sv2v_reg <= data_nn[426];
      data_r_425_sv2v_reg <= data_nn[425];
      data_r_424_sv2v_reg <= data_nn[424];
      data_r_423_sv2v_reg <= data_nn[423];
      data_r_422_sv2v_reg <= data_nn[422];
      data_r_421_sv2v_reg <= data_nn[421];
      data_r_420_sv2v_reg <= data_nn[420];
      data_r_419_sv2v_reg <= data_nn[419];
      data_r_418_sv2v_reg <= data_nn[418];
      data_r_417_sv2v_reg <= data_nn[417];
      data_r_416_sv2v_reg <= data_nn[416];
      data_r_415_sv2v_reg <= data_nn[415];
      data_r_414_sv2v_reg <= data_nn[414];
      data_r_413_sv2v_reg <= data_nn[413];
      data_r_412_sv2v_reg <= data_nn[412];
      data_r_411_sv2v_reg <= data_nn[411];
      data_r_410_sv2v_reg <= data_nn[410];
      data_r_409_sv2v_reg <= data_nn[409];
      data_r_408_sv2v_reg <= data_nn[408];
      data_r_407_sv2v_reg <= data_nn[407];
      data_r_406_sv2v_reg <= data_nn[406];
      data_r_405_sv2v_reg <= data_nn[405];
      data_r_404_sv2v_reg <= data_nn[404];
      data_r_403_sv2v_reg <= data_nn[403];
      data_r_402_sv2v_reg <= data_nn[402];
      data_r_401_sv2v_reg <= data_nn[401];
      data_r_400_sv2v_reg <= data_nn[400];
      data_r_399_sv2v_reg <= data_nn[399];
      data_r_398_sv2v_reg <= data_nn[398];
      data_r_397_sv2v_reg <= data_nn[397];
      data_r_396_sv2v_reg <= data_nn[396];
      data_r_395_sv2v_reg <= data_nn[395];
      data_r_394_sv2v_reg <= data_nn[394];
      data_r_393_sv2v_reg <= data_nn[393];
      data_r_392_sv2v_reg <= data_nn[392];
      data_r_391_sv2v_reg <= data_nn[391];
      data_r_390_sv2v_reg <= data_nn[390];
      data_r_389_sv2v_reg <= data_nn[389];
      data_r_388_sv2v_reg <= data_nn[388];
      data_r_387_sv2v_reg <= data_nn[387];
      data_r_386_sv2v_reg <= data_nn[386];
      data_r_385_sv2v_reg <= data_nn[385];
      data_r_384_sv2v_reg <= data_nn[384];
      data_r_383_sv2v_reg <= data_nn[383];
      data_r_382_sv2v_reg <= data_nn[382];
      data_r_381_sv2v_reg <= data_nn[381];
      data_r_380_sv2v_reg <= data_nn[380];
      data_r_379_sv2v_reg <= data_nn[379];
      data_r_378_sv2v_reg <= data_nn[378];
      data_r_377_sv2v_reg <= data_nn[377];
      data_r_376_sv2v_reg <= data_nn[376];
      data_r_375_sv2v_reg <= data_nn[375];
      data_r_374_sv2v_reg <= data_nn[374];
      data_r_373_sv2v_reg <= data_nn[373];
      data_r_372_sv2v_reg <= data_nn[372];
      data_r_371_sv2v_reg <= data_nn[371];
      data_r_370_sv2v_reg <= data_nn[370];
      data_r_369_sv2v_reg <= data_nn[369];
      data_r_368_sv2v_reg <= data_nn[368];
      data_r_367_sv2v_reg <= data_nn[367];
      data_r_366_sv2v_reg <= data_nn[366];
      data_r_365_sv2v_reg <= data_nn[365];
      data_r_364_sv2v_reg <= data_nn[364];
      data_r_363_sv2v_reg <= data_nn[363];
      data_r_362_sv2v_reg <= data_nn[362];
      data_r_361_sv2v_reg <= data_nn[361];
      data_r_360_sv2v_reg <= data_nn[360];
      data_r_359_sv2v_reg <= data_nn[359];
      data_r_358_sv2v_reg <= data_nn[358];
      data_r_357_sv2v_reg <= data_nn[357];
      data_r_356_sv2v_reg <= data_nn[356];
      data_r_355_sv2v_reg <= data_nn[355];
      data_r_354_sv2v_reg <= data_nn[354];
      data_r_353_sv2v_reg <= data_nn[353];
      data_r_352_sv2v_reg <= data_nn[352];
      data_r_351_sv2v_reg <= data_nn[351];
      data_r_350_sv2v_reg <= data_nn[350];
      data_r_349_sv2v_reg <= data_nn[349];
      data_r_348_sv2v_reg <= data_nn[348];
      data_r_347_sv2v_reg <= data_nn[347];
      data_r_346_sv2v_reg <= data_nn[346];
      data_r_345_sv2v_reg <= data_nn[345];
      data_r_344_sv2v_reg <= data_nn[344];
      data_r_343_sv2v_reg <= data_nn[343];
      data_r_342_sv2v_reg <= data_nn[342];
      data_r_341_sv2v_reg <= data_nn[341];
      data_r_340_sv2v_reg <= data_nn[340];
      data_r_339_sv2v_reg <= data_nn[339];
      data_r_338_sv2v_reg <= data_nn[338];
      data_r_337_sv2v_reg <= data_nn[337];
      data_r_336_sv2v_reg <= data_nn[336];
      data_r_335_sv2v_reg <= data_nn[335];
      data_r_334_sv2v_reg <= data_nn[334];
      data_r_333_sv2v_reg <= data_nn[333];
      data_r_332_sv2v_reg <= data_nn[332];
      data_r_331_sv2v_reg <= data_nn[331];
      data_r_330_sv2v_reg <= data_nn[330];
      data_r_329_sv2v_reg <= data_nn[329];
      data_r_328_sv2v_reg <= data_nn[328];
      data_r_327_sv2v_reg <= data_nn[327];
      data_r_326_sv2v_reg <= data_nn[326];
      data_r_325_sv2v_reg <= data_nn[325];
      data_r_324_sv2v_reg <= data_nn[324];
      data_r_323_sv2v_reg <= data_nn[323];
      data_r_322_sv2v_reg <= data_nn[322];
      data_r_321_sv2v_reg <= data_nn[321];
      data_r_320_sv2v_reg <= data_nn[320];
      data_r_319_sv2v_reg <= data_nn[319];
      data_r_318_sv2v_reg <= data_nn[318];
      data_r_317_sv2v_reg <= data_nn[317];
      data_r_316_sv2v_reg <= data_nn[316];
      data_r_315_sv2v_reg <= data_nn[315];
      data_r_314_sv2v_reg <= data_nn[314];
      data_r_313_sv2v_reg <= data_nn[313];
      data_r_312_sv2v_reg <= data_nn[312];
      data_r_311_sv2v_reg <= data_nn[311];
      data_r_310_sv2v_reg <= data_nn[310];
      data_r_309_sv2v_reg <= data_nn[309];
      data_r_308_sv2v_reg <= data_nn[308];
      data_r_307_sv2v_reg <= data_nn[307];
      data_r_306_sv2v_reg <= data_nn[306];
      data_r_305_sv2v_reg <= data_nn[305];
      data_r_304_sv2v_reg <= data_nn[304];
      data_r_303_sv2v_reg <= data_nn[303];
      data_r_302_sv2v_reg <= data_nn[302];
      data_r_301_sv2v_reg <= data_nn[301];
      data_r_300_sv2v_reg <= data_nn[300];
      data_r_299_sv2v_reg <= data_nn[299];
      data_r_298_sv2v_reg <= data_nn[298];
      data_r_297_sv2v_reg <= data_nn[297];
      data_r_296_sv2v_reg <= data_nn[296];
      data_r_295_sv2v_reg <= data_nn[295];
      data_r_294_sv2v_reg <= data_nn[294];
      data_r_293_sv2v_reg <= data_nn[293];
      data_r_292_sv2v_reg <= data_nn[292];
      data_r_291_sv2v_reg <= data_nn[291];
      data_r_290_sv2v_reg <= data_nn[290];
      data_r_289_sv2v_reg <= data_nn[289];
      data_r_288_sv2v_reg <= data_nn[288];
      data_r_287_sv2v_reg <= data_nn[287];
      data_r_286_sv2v_reg <= data_nn[286];
      data_r_285_sv2v_reg <= data_nn[285];
      data_r_284_sv2v_reg <= data_nn[284];
      data_r_283_sv2v_reg <= data_nn[283];
      data_r_282_sv2v_reg <= data_nn[282];
      data_r_281_sv2v_reg <= data_nn[281];
      data_r_280_sv2v_reg <= data_nn[280];
      data_r_279_sv2v_reg <= data_nn[279];
      data_r_278_sv2v_reg <= data_nn[278];
      data_r_277_sv2v_reg <= data_nn[277];
      data_r_276_sv2v_reg <= data_nn[276];
      data_r_275_sv2v_reg <= data_nn[275];
      data_r_274_sv2v_reg <= data_nn[274];
      data_r_273_sv2v_reg <= data_nn[273];
      data_r_272_sv2v_reg <= data_nn[272];
      data_r_271_sv2v_reg <= data_nn[271];
      data_r_270_sv2v_reg <= data_nn[270];
      data_r_269_sv2v_reg <= data_nn[269];
      data_r_268_sv2v_reg <= data_nn[268];
      data_r_267_sv2v_reg <= data_nn[267];
      data_r_266_sv2v_reg <= data_nn[266];
      data_r_265_sv2v_reg <= data_nn[265];
      data_r_264_sv2v_reg <= data_nn[264];
      data_r_263_sv2v_reg <= data_nn[263];
      data_r_262_sv2v_reg <= data_nn[262];
      data_r_261_sv2v_reg <= data_nn[261];
      data_r_260_sv2v_reg <= data_nn[260];
      data_r_259_sv2v_reg <= data_nn[259];
      data_r_258_sv2v_reg <= data_nn[258];
      data_r_257_sv2v_reg <= data_nn[257];
      data_r_256_sv2v_reg <= data_nn[256];
      data_r_255_sv2v_reg <= data_nn[255];
      data_r_254_sv2v_reg <= data_nn[254];
      data_r_253_sv2v_reg <= data_nn[253];
      data_r_252_sv2v_reg <= data_nn[252];
      data_r_251_sv2v_reg <= data_nn[251];
      data_r_250_sv2v_reg <= data_nn[250];
      data_r_249_sv2v_reg <= data_nn[249];
      data_r_248_sv2v_reg <= data_nn[248];
      data_r_247_sv2v_reg <= data_nn[247];
      data_r_246_sv2v_reg <= data_nn[246];
      data_r_245_sv2v_reg <= data_nn[245];
      data_r_244_sv2v_reg <= data_nn[244];
      data_r_243_sv2v_reg <= data_nn[243];
      data_r_242_sv2v_reg <= data_nn[242];
      data_r_241_sv2v_reg <= data_nn[241];
      data_r_240_sv2v_reg <= data_nn[240];
      data_r_239_sv2v_reg <= data_nn[239];
      data_r_238_sv2v_reg <= data_nn[238];
      data_r_237_sv2v_reg <= data_nn[237];
      data_r_236_sv2v_reg <= data_nn[236];
      data_r_235_sv2v_reg <= data_nn[235];
      data_r_234_sv2v_reg <= data_nn[234];
      data_r_233_sv2v_reg <= data_nn[233];
      data_r_232_sv2v_reg <= data_nn[232];
      data_r_231_sv2v_reg <= data_nn[231];
      data_r_230_sv2v_reg <= data_nn[230];
      data_r_229_sv2v_reg <= data_nn[229];
      data_r_228_sv2v_reg <= data_nn[228];
      data_r_227_sv2v_reg <= data_nn[227];
      data_r_226_sv2v_reg <= data_nn[226];
      data_r_225_sv2v_reg <= data_nn[225];
      data_r_224_sv2v_reg <= data_nn[224];
      data_r_223_sv2v_reg <= data_nn[223];
      data_r_222_sv2v_reg <= data_nn[222];
      data_r_221_sv2v_reg <= data_nn[221];
      data_r_220_sv2v_reg <= data_nn[220];
      data_r_219_sv2v_reg <= data_nn[219];
      data_r_218_sv2v_reg <= data_nn[218];
      data_r_217_sv2v_reg <= data_nn[217];
      data_r_216_sv2v_reg <= data_nn[216];
      data_r_215_sv2v_reg <= data_nn[215];
      data_r_214_sv2v_reg <= data_nn[214];
      data_r_213_sv2v_reg <= data_nn[213];
      data_r_212_sv2v_reg <= data_nn[212];
      data_r_211_sv2v_reg <= data_nn[211];
      data_r_210_sv2v_reg <= data_nn[210];
      data_r_209_sv2v_reg <= data_nn[209];
      data_r_208_sv2v_reg <= data_nn[208];
      data_r_207_sv2v_reg <= data_nn[207];
      data_r_206_sv2v_reg <= data_nn[206];
      data_r_205_sv2v_reg <= data_nn[205];
      data_r_204_sv2v_reg <= data_nn[204];
      data_r_203_sv2v_reg <= data_nn[203];
      data_r_202_sv2v_reg <= data_nn[202];
      data_r_201_sv2v_reg <= data_nn[201];
      data_r_200_sv2v_reg <= data_nn[200];
      data_r_199_sv2v_reg <= data_nn[199];
      data_r_198_sv2v_reg <= data_nn[198];
      data_r_197_sv2v_reg <= data_nn[197];
      data_r_196_sv2v_reg <= data_nn[196];
      data_r_195_sv2v_reg <= data_nn[195];
      data_r_194_sv2v_reg <= data_nn[194];
      data_r_193_sv2v_reg <= data_nn[193];
      data_r_192_sv2v_reg <= data_nn[192];
      data_r_191_sv2v_reg <= data_nn[191];
      data_r_190_sv2v_reg <= data_nn[190];
      data_r_189_sv2v_reg <= data_nn[189];
      data_r_188_sv2v_reg <= data_nn[188];
      data_r_187_sv2v_reg <= data_nn[187];
      data_r_186_sv2v_reg <= data_nn[186];
      data_r_185_sv2v_reg <= data_nn[185];
      data_r_184_sv2v_reg <= data_nn[184];
      data_r_183_sv2v_reg <= data_nn[183];
      data_r_182_sv2v_reg <= data_nn[182];
      data_r_181_sv2v_reg <= data_nn[181];
      data_r_180_sv2v_reg <= data_nn[180];
      data_r_179_sv2v_reg <= data_nn[179];
      data_r_178_sv2v_reg <= data_nn[178];
      data_r_177_sv2v_reg <= data_nn[177];
      data_r_176_sv2v_reg <= data_nn[176];
      data_r_175_sv2v_reg <= data_nn[175];
      data_r_174_sv2v_reg <= data_nn[174];
      data_r_173_sv2v_reg <= data_nn[173];
      data_r_172_sv2v_reg <= data_nn[172];
      data_r_171_sv2v_reg <= data_nn[171];
      data_r_170_sv2v_reg <= data_nn[170];
      data_r_169_sv2v_reg <= data_nn[169];
      data_r_168_sv2v_reg <= data_nn[168];
      data_r_167_sv2v_reg <= data_nn[167];
      data_r_166_sv2v_reg <= data_nn[166];
      data_r_165_sv2v_reg <= data_nn[165];
      data_r_164_sv2v_reg <= data_nn[164];
      data_r_163_sv2v_reg <= data_nn[163];
      data_r_162_sv2v_reg <= data_nn[162];
      data_r_161_sv2v_reg <= data_nn[161];
      data_r_160_sv2v_reg <= data_nn[160];
      data_r_159_sv2v_reg <= data_nn[159];
      data_r_158_sv2v_reg <= data_nn[158];
      data_r_157_sv2v_reg <= data_nn[157];
      data_r_156_sv2v_reg <= data_nn[156];
      data_r_155_sv2v_reg <= data_nn[155];
      data_r_154_sv2v_reg <= data_nn[154];
      data_r_153_sv2v_reg <= data_nn[153];
      data_r_152_sv2v_reg <= data_nn[152];
      data_r_151_sv2v_reg <= data_nn[151];
      data_r_150_sv2v_reg <= data_nn[150];
      data_r_149_sv2v_reg <= data_nn[149];
      data_r_148_sv2v_reg <= data_nn[148];
      data_r_147_sv2v_reg <= data_nn[147];
      data_r_146_sv2v_reg <= data_nn[146];
      data_r_145_sv2v_reg <= data_nn[145];
      data_r_144_sv2v_reg <= data_nn[144];
      data_r_143_sv2v_reg <= data_nn[143];
      data_r_142_sv2v_reg <= data_nn[142];
      data_r_141_sv2v_reg <= data_nn[141];
      data_r_140_sv2v_reg <= data_nn[140];
      data_r_139_sv2v_reg <= data_nn[139];
      data_r_138_sv2v_reg <= data_nn[138];
      data_r_137_sv2v_reg <= data_nn[137];
      data_r_136_sv2v_reg <= data_nn[136];
      data_r_135_sv2v_reg <= data_nn[135];
      data_r_134_sv2v_reg <= data_nn[134];
      data_r_133_sv2v_reg <= data_nn[133];
      data_r_132_sv2v_reg <= data_nn[132];
      data_r_131_sv2v_reg <= data_nn[131];
      data_r_130_sv2v_reg <= data_nn[130];
      data_r_129_sv2v_reg <= data_nn[129];
      data_r_128_sv2v_reg <= data_nn[128];
      data_r_127_sv2v_reg <= data_nn[127];
      data_r_126_sv2v_reg <= data_nn[126];
      data_r_125_sv2v_reg <= data_nn[125];
      data_r_124_sv2v_reg <= data_nn[124];
      data_r_123_sv2v_reg <= data_nn[123];
      data_r_122_sv2v_reg <= data_nn[122];
      data_r_121_sv2v_reg <= data_nn[121];
      data_r_120_sv2v_reg <= data_nn[120];
      data_r_119_sv2v_reg <= data_nn[119];
      data_r_118_sv2v_reg <= data_nn[118];
      data_r_117_sv2v_reg <= data_nn[117];
      data_r_116_sv2v_reg <= data_nn[116];
      data_r_115_sv2v_reg <= data_nn[115];
      data_r_114_sv2v_reg <= data_nn[114];
      data_r_113_sv2v_reg <= data_nn[113];
      data_r_112_sv2v_reg <= data_nn[112];
      data_r_111_sv2v_reg <= data_nn[111];
      data_r_110_sv2v_reg <= data_nn[110];
      data_r_109_sv2v_reg <= data_nn[109];
      data_r_108_sv2v_reg <= data_nn[108];
      data_r_107_sv2v_reg <= data_nn[107];
      data_r_106_sv2v_reg <= data_nn[106];
      data_r_105_sv2v_reg <= data_nn[105];
      data_r_104_sv2v_reg <= data_nn[104];
      data_r_103_sv2v_reg <= data_nn[103];
      data_r_102_sv2v_reg <= data_nn[102];
      data_r_101_sv2v_reg <= data_nn[101];
      data_r_100_sv2v_reg <= data_nn[100];
      data_r_99_sv2v_reg <= data_nn[99];
      data_r_98_sv2v_reg <= data_nn[98];
      data_r_97_sv2v_reg <= data_nn[97];
      data_r_96_sv2v_reg <= data_nn[96];
      data_r_95_sv2v_reg <= data_nn[95];
      data_r_94_sv2v_reg <= data_nn[94];
      data_r_93_sv2v_reg <= data_nn[93];
      data_r_92_sv2v_reg <= data_nn[92];
      data_r_91_sv2v_reg <= data_nn[91];
      data_r_90_sv2v_reg <= data_nn[90];
      data_r_89_sv2v_reg <= data_nn[89];
      data_r_88_sv2v_reg <= data_nn[88];
      data_r_87_sv2v_reg <= data_nn[87];
      data_r_86_sv2v_reg <= data_nn[86];
      data_r_85_sv2v_reg <= data_nn[85];
      data_r_84_sv2v_reg <= data_nn[84];
      data_r_83_sv2v_reg <= data_nn[83];
      data_r_82_sv2v_reg <= data_nn[82];
      data_r_81_sv2v_reg <= data_nn[81];
      data_r_80_sv2v_reg <= data_nn[80];
      data_r_79_sv2v_reg <= data_nn[79];
      data_r_78_sv2v_reg <= data_nn[78];
      data_r_77_sv2v_reg <= data_nn[77];
      data_r_76_sv2v_reg <= data_nn[76];
      data_r_75_sv2v_reg <= data_nn[75];
      data_r_74_sv2v_reg <= data_nn[74];
      data_r_73_sv2v_reg <= data_nn[73];
      data_r_72_sv2v_reg <= data_nn[72];
      data_r_71_sv2v_reg <= data_nn[71];
      data_r_70_sv2v_reg <= data_nn[70];
      data_r_69_sv2v_reg <= data_nn[69];
      data_r_68_sv2v_reg <= data_nn[68];
      data_r_67_sv2v_reg <= data_nn[67];
      data_r_66_sv2v_reg <= data_nn[66];
      data_r_65_sv2v_reg <= data_nn[65];
      data_r_64_sv2v_reg <= data_nn[64];
      data_r_63_sv2v_reg <= data_nn[63];
      data_r_62_sv2v_reg <= data_nn[62];
      data_r_61_sv2v_reg <= data_nn[61];
      data_r_60_sv2v_reg <= data_nn[60];
      data_r_59_sv2v_reg <= data_nn[59];
      data_r_58_sv2v_reg <= data_nn[58];
      data_r_57_sv2v_reg <= data_nn[57];
      data_r_56_sv2v_reg <= data_nn[56];
      data_r_55_sv2v_reg <= data_nn[55];
      data_r_54_sv2v_reg <= data_nn[54];
      data_r_53_sv2v_reg <= data_nn[53];
      data_r_52_sv2v_reg <= data_nn[52];
      data_r_51_sv2v_reg <= data_nn[51];
      data_r_50_sv2v_reg <= data_nn[50];
      data_r_49_sv2v_reg <= data_nn[49];
      data_r_48_sv2v_reg <= data_nn[48];
      data_r_47_sv2v_reg <= data_nn[47];
      data_r_46_sv2v_reg <= data_nn[46];
      data_r_45_sv2v_reg <= data_nn[45];
      data_r_44_sv2v_reg <= data_nn[44];
      data_r_43_sv2v_reg <= data_nn[43];
      data_r_42_sv2v_reg <= data_nn[42];
      data_r_41_sv2v_reg <= data_nn[41];
      data_r_40_sv2v_reg <= data_nn[40];
      data_r_39_sv2v_reg <= data_nn[39];
      data_r_38_sv2v_reg <= data_nn[38];
      data_r_37_sv2v_reg <= data_nn[37];
      data_r_36_sv2v_reg <= data_nn[36];
      data_r_35_sv2v_reg <= data_nn[35];
      data_r_34_sv2v_reg <= data_nn[34];
      data_r_33_sv2v_reg <= data_nn[33];
      data_r_32_sv2v_reg <= data_nn[32];
      data_r_31_sv2v_reg <= data_nn[31];
      data_r_30_sv2v_reg <= data_nn[30];
      data_r_29_sv2v_reg <= data_nn[29];
      data_r_28_sv2v_reg <= data_nn[28];
      data_r_27_sv2v_reg <= data_nn[27];
      data_r_26_sv2v_reg <= data_nn[26];
      data_r_25_sv2v_reg <= data_nn[25];
      data_r_24_sv2v_reg <= data_nn[24];
      data_r_23_sv2v_reg <= data_nn[23];
      data_r_22_sv2v_reg <= data_nn[22];
      data_r_21_sv2v_reg <= data_nn[21];
      data_r_20_sv2v_reg <= data_nn[20];
      data_r_19_sv2v_reg <= data_nn[19];
      data_r_18_sv2v_reg <= data_nn[18];
      data_r_17_sv2v_reg <= data_nn[17];
      data_r_16_sv2v_reg <= data_nn[16];
      data_r_15_sv2v_reg <= data_nn[15];
      data_r_14_sv2v_reg <= data_nn[14];
      data_r_13_sv2v_reg <= data_nn[13];
      data_r_12_sv2v_reg <= data_nn[12];
      data_r_11_sv2v_reg <= data_nn[11];
      data_r_10_sv2v_reg <= data_nn[10];
      data_r_9_sv2v_reg <= data_nn[9];
      data_r_8_sv2v_reg <= data_nn[8];
      data_r_7_sv2v_reg <= data_nn[7];
      data_r_6_sv2v_reg <= data_nn[6];
      data_r_5_sv2v_reg <= data_nn[5];
      data_r_4_sv2v_reg <= data_nn[4];
      data_r_3_sv2v_reg <= data_nn[3];
      data_r_2_sv2v_reg <= data_nn[2];
      data_r_1_sv2v_reg <= data_nn[1];
      data_r_0_sv2v_reg <= data_nn[0];
    end 
  end


endmodule

