

module top
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_i
);

  input [511:0] data_i;
  output [15:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_o;
  output valid_o;

  bsg_parallel_in_serial_out
  wrapper
  (
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .valid_i(valid_i),
    .yumi_i(yumi_i),
    .ready_o(ready_o),
    .valid_o(valid_o)
  );


endmodule



module bsg_parallel_in_serial_out
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_i
);

  input [511:0] data_i;
  output [15:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_o;
  output valid_o;
  wire [15:0] data_o;
  wire ready_o,valid_o,N0,N1,\piso.done_tx_n ,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95;
  wire [4:0] \piso.shift_ctr_r ;
  wire [0:0] \piso.state_n ;
  wire [511:0] \piso.data_r ;
  reg valid_o_sv2v_reg,\piso.data_r_511_sv2v_reg ,\piso.data_r_510_sv2v_reg ,
  \piso.data_r_509_sv2v_reg ,\piso.data_r_508_sv2v_reg ,\piso.data_r_507_sv2v_reg ,
  \piso.data_r_506_sv2v_reg ,\piso.data_r_505_sv2v_reg ,\piso.data_r_504_sv2v_reg ,
  \piso.data_r_503_sv2v_reg ,\piso.data_r_502_sv2v_reg ,\piso.data_r_501_sv2v_reg ,
  \piso.data_r_500_sv2v_reg ,\piso.data_r_499_sv2v_reg ,\piso.data_r_498_sv2v_reg ,
  \piso.data_r_497_sv2v_reg ,\piso.data_r_496_sv2v_reg ,\piso.data_r_495_sv2v_reg ,
  \piso.data_r_494_sv2v_reg ,\piso.data_r_493_sv2v_reg ,\piso.data_r_492_sv2v_reg ,
  \piso.data_r_491_sv2v_reg ,\piso.data_r_490_sv2v_reg ,\piso.data_r_489_sv2v_reg ,
  \piso.data_r_488_sv2v_reg ,\piso.data_r_487_sv2v_reg ,\piso.data_r_486_sv2v_reg ,
  \piso.data_r_485_sv2v_reg ,\piso.data_r_484_sv2v_reg ,\piso.data_r_483_sv2v_reg ,
  \piso.data_r_482_sv2v_reg ,\piso.data_r_481_sv2v_reg ,
  \piso.data_r_480_sv2v_reg ,\piso.data_r_479_sv2v_reg ,\piso.data_r_478_sv2v_reg ,
  \piso.data_r_477_sv2v_reg ,\piso.data_r_476_sv2v_reg ,\piso.data_r_475_sv2v_reg ,
  \piso.data_r_474_sv2v_reg ,\piso.data_r_473_sv2v_reg ,\piso.data_r_472_sv2v_reg ,
  \piso.data_r_471_sv2v_reg ,\piso.data_r_470_sv2v_reg ,\piso.data_r_469_sv2v_reg ,
  \piso.data_r_468_sv2v_reg ,\piso.data_r_467_sv2v_reg ,\piso.data_r_466_sv2v_reg ,
  \piso.data_r_465_sv2v_reg ,\piso.data_r_464_sv2v_reg ,\piso.data_r_463_sv2v_reg ,
  \piso.data_r_462_sv2v_reg ,\piso.data_r_461_sv2v_reg ,\piso.data_r_460_sv2v_reg ,
  \piso.data_r_459_sv2v_reg ,\piso.data_r_458_sv2v_reg ,\piso.data_r_457_sv2v_reg ,
  \piso.data_r_456_sv2v_reg ,\piso.data_r_455_sv2v_reg ,\piso.data_r_454_sv2v_reg ,
  \piso.data_r_453_sv2v_reg ,\piso.data_r_452_sv2v_reg ,\piso.data_r_451_sv2v_reg ,
  \piso.data_r_450_sv2v_reg ,\piso.data_r_449_sv2v_reg ,\piso.data_r_448_sv2v_reg ,
  \piso.data_r_447_sv2v_reg ,\piso.data_r_446_sv2v_reg ,\piso.data_r_445_sv2v_reg ,
  \piso.data_r_444_sv2v_reg ,\piso.data_r_443_sv2v_reg ,\piso.data_r_442_sv2v_reg ,
  \piso.data_r_441_sv2v_reg ,\piso.data_r_440_sv2v_reg ,\piso.data_r_439_sv2v_reg ,
  \piso.data_r_438_sv2v_reg ,\piso.data_r_437_sv2v_reg ,\piso.data_r_436_sv2v_reg ,
  \piso.data_r_435_sv2v_reg ,\piso.data_r_434_sv2v_reg ,\piso.data_r_433_sv2v_reg ,
  \piso.data_r_432_sv2v_reg ,\piso.data_r_431_sv2v_reg ,\piso.data_r_430_sv2v_reg ,
  \piso.data_r_429_sv2v_reg ,\piso.data_r_428_sv2v_reg ,\piso.data_r_427_sv2v_reg ,
  \piso.data_r_426_sv2v_reg ,\piso.data_r_425_sv2v_reg ,\piso.data_r_424_sv2v_reg ,
  \piso.data_r_423_sv2v_reg ,\piso.data_r_422_sv2v_reg ,\piso.data_r_421_sv2v_reg ,
  \piso.data_r_420_sv2v_reg ,\piso.data_r_419_sv2v_reg ,\piso.data_r_418_sv2v_reg ,
  \piso.data_r_417_sv2v_reg ,\piso.data_r_416_sv2v_reg ,\piso.data_r_415_sv2v_reg ,
  \piso.data_r_414_sv2v_reg ,\piso.data_r_413_sv2v_reg ,\piso.data_r_412_sv2v_reg ,
  \piso.data_r_411_sv2v_reg ,\piso.data_r_410_sv2v_reg ,\piso.data_r_409_sv2v_reg ,
  \piso.data_r_408_sv2v_reg ,\piso.data_r_407_sv2v_reg ,\piso.data_r_406_sv2v_reg ,
  \piso.data_r_405_sv2v_reg ,\piso.data_r_404_sv2v_reg ,\piso.data_r_403_sv2v_reg ,
  \piso.data_r_402_sv2v_reg ,\piso.data_r_401_sv2v_reg ,
  \piso.data_r_400_sv2v_reg ,\piso.data_r_399_sv2v_reg ,\piso.data_r_398_sv2v_reg ,
  \piso.data_r_397_sv2v_reg ,\piso.data_r_396_sv2v_reg ,\piso.data_r_395_sv2v_reg ,
  \piso.data_r_394_sv2v_reg ,\piso.data_r_393_sv2v_reg ,\piso.data_r_392_sv2v_reg ,
  \piso.data_r_391_sv2v_reg ,\piso.data_r_390_sv2v_reg ,\piso.data_r_389_sv2v_reg ,
  \piso.data_r_388_sv2v_reg ,\piso.data_r_387_sv2v_reg ,\piso.data_r_386_sv2v_reg ,
  \piso.data_r_385_sv2v_reg ,\piso.data_r_384_sv2v_reg ,\piso.data_r_383_sv2v_reg ,
  \piso.data_r_382_sv2v_reg ,\piso.data_r_381_sv2v_reg ,\piso.data_r_380_sv2v_reg ,
  \piso.data_r_379_sv2v_reg ,\piso.data_r_378_sv2v_reg ,\piso.data_r_377_sv2v_reg ,
  \piso.data_r_376_sv2v_reg ,\piso.data_r_375_sv2v_reg ,\piso.data_r_374_sv2v_reg ,
  \piso.data_r_373_sv2v_reg ,\piso.data_r_372_sv2v_reg ,\piso.data_r_371_sv2v_reg ,
  \piso.data_r_370_sv2v_reg ,\piso.data_r_369_sv2v_reg ,\piso.data_r_368_sv2v_reg ,
  \piso.data_r_367_sv2v_reg ,\piso.data_r_366_sv2v_reg ,\piso.data_r_365_sv2v_reg ,
  \piso.data_r_364_sv2v_reg ,\piso.data_r_363_sv2v_reg ,\piso.data_r_362_sv2v_reg ,
  \piso.data_r_361_sv2v_reg ,\piso.data_r_360_sv2v_reg ,\piso.data_r_359_sv2v_reg ,
  \piso.data_r_358_sv2v_reg ,\piso.data_r_357_sv2v_reg ,\piso.data_r_356_sv2v_reg ,
  \piso.data_r_355_sv2v_reg ,\piso.data_r_354_sv2v_reg ,\piso.data_r_353_sv2v_reg ,
  \piso.data_r_352_sv2v_reg ,\piso.data_r_351_sv2v_reg ,\piso.data_r_350_sv2v_reg ,
  \piso.data_r_349_sv2v_reg ,\piso.data_r_348_sv2v_reg ,\piso.data_r_347_sv2v_reg ,
  \piso.data_r_346_sv2v_reg ,\piso.data_r_345_sv2v_reg ,\piso.data_r_344_sv2v_reg ,
  \piso.data_r_343_sv2v_reg ,\piso.data_r_342_sv2v_reg ,\piso.data_r_341_sv2v_reg ,
  \piso.data_r_340_sv2v_reg ,\piso.data_r_339_sv2v_reg ,\piso.data_r_338_sv2v_reg ,
  \piso.data_r_337_sv2v_reg ,\piso.data_r_336_sv2v_reg ,\piso.data_r_335_sv2v_reg ,
  \piso.data_r_334_sv2v_reg ,\piso.data_r_333_sv2v_reg ,\piso.data_r_332_sv2v_reg ,
  \piso.data_r_331_sv2v_reg ,\piso.data_r_330_sv2v_reg ,\piso.data_r_329_sv2v_reg ,
  \piso.data_r_328_sv2v_reg ,\piso.data_r_327_sv2v_reg ,\piso.data_r_326_sv2v_reg ,
  \piso.data_r_325_sv2v_reg ,\piso.data_r_324_sv2v_reg ,\piso.data_r_323_sv2v_reg ,
  \piso.data_r_322_sv2v_reg ,\piso.data_r_321_sv2v_reg ,
  \piso.data_r_320_sv2v_reg ,\piso.data_r_319_sv2v_reg ,\piso.data_r_318_sv2v_reg ,
  \piso.data_r_317_sv2v_reg ,\piso.data_r_316_sv2v_reg ,\piso.data_r_315_sv2v_reg ,
  \piso.data_r_314_sv2v_reg ,\piso.data_r_313_sv2v_reg ,\piso.data_r_312_sv2v_reg ,
  \piso.data_r_311_sv2v_reg ,\piso.data_r_310_sv2v_reg ,\piso.data_r_309_sv2v_reg ,
  \piso.data_r_308_sv2v_reg ,\piso.data_r_307_sv2v_reg ,\piso.data_r_306_sv2v_reg ,
  \piso.data_r_305_sv2v_reg ,\piso.data_r_304_sv2v_reg ,\piso.data_r_303_sv2v_reg ,
  \piso.data_r_302_sv2v_reg ,\piso.data_r_301_sv2v_reg ,\piso.data_r_300_sv2v_reg ,
  \piso.data_r_299_sv2v_reg ,\piso.data_r_298_sv2v_reg ,\piso.data_r_297_sv2v_reg ,
  \piso.data_r_296_sv2v_reg ,\piso.data_r_295_sv2v_reg ,\piso.data_r_294_sv2v_reg ,
  \piso.data_r_293_sv2v_reg ,\piso.data_r_292_sv2v_reg ,\piso.data_r_291_sv2v_reg ,
  \piso.data_r_290_sv2v_reg ,\piso.data_r_289_sv2v_reg ,\piso.data_r_288_sv2v_reg ,
  \piso.data_r_287_sv2v_reg ,\piso.data_r_286_sv2v_reg ,\piso.data_r_285_sv2v_reg ,
  \piso.data_r_284_sv2v_reg ,\piso.data_r_283_sv2v_reg ,\piso.data_r_282_sv2v_reg ,
  \piso.data_r_281_sv2v_reg ,\piso.data_r_280_sv2v_reg ,\piso.data_r_279_sv2v_reg ,
  \piso.data_r_278_sv2v_reg ,\piso.data_r_277_sv2v_reg ,\piso.data_r_276_sv2v_reg ,
  \piso.data_r_275_sv2v_reg ,\piso.data_r_274_sv2v_reg ,\piso.data_r_273_sv2v_reg ,
  \piso.data_r_272_sv2v_reg ,\piso.data_r_271_sv2v_reg ,\piso.data_r_270_sv2v_reg ,
  \piso.data_r_269_sv2v_reg ,\piso.data_r_268_sv2v_reg ,\piso.data_r_267_sv2v_reg ,
  \piso.data_r_266_sv2v_reg ,\piso.data_r_265_sv2v_reg ,\piso.data_r_264_sv2v_reg ,
  \piso.data_r_263_sv2v_reg ,\piso.data_r_262_sv2v_reg ,\piso.data_r_261_sv2v_reg ,
  \piso.data_r_260_sv2v_reg ,\piso.data_r_259_sv2v_reg ,\piso.data_r_258_sv2v_reg ,
  \piso.data_r_257_sv2v_reg ,\piso.data_r_256_sv2v_reg ,\piso.data_r_255_sv2v_reg ,
  \piso.data_r_254_sv2v_reg ,\piso.data_r_253_sv2v_reg ,\piso.data_r_252_sv2v_reg ,
  \piso.data_r_251_sv2v_reg ,\piso.data_r_250_sv2v_reg ,\piso.data_r_249_sv2v_reg ,
  \piso.data_r_248_sv2v_reg ,\piso.data_r_247_sv2v_reg ,\piso.data_r_246_sv2v_reg ,
  \piso.data_r_245_sv2v_reg ,\piso.data_r_244_sv2v_reg ,\piso.data_r_243_sv2v_reg ,
  \piso.data_r_242_sv2v_reg ,\piso.data_r_241_sv2v_reg ,
  \piso.data_r_240_sv2v_reg ,\piso.data_r_239_sv2v_reg ,\piso.data_r_238_sv2v_reg ,
  \piso.data_r_237_sv2v_reg ,\piso.data_r_236_sv2v_reg ,\piso.data_r_235_sv2v_reg ,
  \piso.data_r_234_sv2v_reg ,\piso.data_r_233_sv2v_reg ,\piso.data_r_232_sv2v_reg ,
  \piso.data_r_231_sv2v_reg ,\piso.data_r_230_sv2v_reg ,\piso.data_r_229_sv2v_reg ,
  \piso.data_r_228_sv2v_reg ,\piso.data_r_227_sv2v_reg ,\piso.data_r_226_sv2v_reg ,
  \piso.data_r_225_sv2v_reg ,\piso.data_r_224_sv2v_reg ,\piso.data_r_223_sv2v_reg ,
  \piso.data_r_222_sv2v_reg ,\piso.data_r_221_sv2v_reg ,\piso.data_r_220_sv2v_reg ,
  \piso.data_r_219_sv2v_reg ,\piso.data_r_218_sv2v_reg ,\piso.data_r_217_sv2v_reg ,
  \piso.data_r_216_sv2v_reg ,\piso.data_r_215_sv2v_reg ,\piso.data_r_214_sv2v_reg ,
  \piso.data_r_213_sv2v_reg ,\piso.data_r_212_sv2v_reg ,\piso.data_r_211_sv2v_reg ,
  \piso.data_r_210_sv2v_reg ,\piso.data_r_209_sv2v_reg ,\piso.data_r_208_sv2v_reg ,
  \piso.data_r_207_sv2v_reg ,\piso.data_r_206_sv2v_reg ,\piso.data_r_205_sv2v_reg ,
  \piso.data_r_204_sv2v_reg ,\piso.data_r_203_sv2v_reg ,\piso.data_r_202_sv2v_reg ,
  \piso.data_r_201_sv2v_reg ,\piso.data_r_200_sv2v_reg ,\piso.data_r_199_sv2v_reg ,
  \piso.data_r_198_sv2v_reg ,\piso.data_r_197_sv2v_reg ,\piso.data_r_196_sv2v_reg ,
  \piso.data_r_195_sv2v_reg ,\piso.data_r_194_sv2v_reg ,\piso.data_r_193_sv2v_reg ,
  \piso.data_r_192_sv2v_reg ,\piso.data_r_191_sv2v_reg ,\piso.data_r_190_sv2v_reg ,
  \piso.data_r_189_sv2v_reg ,\piso.data_r_188_sv2v_reg ,\piso.data_r_187_sv2v_reg ,
  \piso.data_r_186_sv2v_reg ,\piso.data_r_185_sv2v_reg ,\piso.data_r_184_sv2v_reg ,
  \piso.data_r_183_sv2v_reg ,\piso.data_r_182_sv2v_reg ,\piso.data_r_181_sv2v_reg ,
  \piso.data_r_180_sv2v_reg ,\piso.data_r_179_sv2v_reg ,\piso.data_r_178_sv2v_reg ,
  \piso.data_r_177_sv2v_reg ,\piso.data_r_176_sv2v_reg ,\piso.data_r_175_sv2v_reg ,
  \piso.data_r_174_sv2v_reg ,\piso.data_r_173_sv2v_reg ,\piso.data_r_172_sv2v_reg ,
  \piso.data_r_171_sv2v_reg ,\piso.data_r_170_sv2v_reg ,\piso.data_r_169_sv2v_reg ,
  \piso.data_r_168_sv2v_reg ,\piso.data_r_167_sv2v_reg ,\piso.data_r_166_sv2v_reg ,
  \piso.data_r_165_sv2v_reg ,\piso.data_r_164_sv2v_reg ,\piso.data_r_163_sv2v_reg ,
  \piso.data_r_162_sv2v_reg ,\piso.data_r_161_sv2v_reg ,
  \piso.data_r_160_sv2v_reg ,\piso.data_r_159_sv2v_reg ,\piso.data_r_158_sv2v_reg ,
  \piso.data_r_157_sv2v_reg ,\piso.data_r_156_sv2v_reg ,\piso.data_r_155_sv2v_reg ,
  \piso.data_r_154_sv2v_reg ,\piso.data_r_153_sv2v_reg ,\piso.data_r_152_sv2v_reg ,
  \piso.data_r_151_sv2v_reg ,\piso.data_r_150_sv2v_reg ,\piso.data_r_149_sv2v_reg ,
  \piso.data_r_148_sv2v_reg ,\piso.data_r_147_sv2v_reg ,\piso.data_r_146_sv2v_reg ,
  \piso.data_r_145_sv2v_reg ,\piso.data_r_144_sv2v_reg ,\piso.data_r_143_sv2v_reg ,
  \piso.data_r_142_sv2v_reg ,\piso.data_r_141_sv2v_reg ,\piso.data_r_140_sv2v_reg ,
  \piso.data_r_139_sv2v_reg ,\piso.data_r_138_sv2v_reg ,\piso.data_r_137_sv2v_reg ,
  \piso.data_r_136_sv2v_reg ,\piso.data_r_135_sv2v_reg ,\piso.data_r_134_sv2v_reg ,
  \piso.data_r_133_sv2v_reg ,\piso.data_r_132_sv2v_reg ,\piso.data_r_131_sv2v_reg ,
  \piso.data_r_130_sv2v_reg ,\piso.data_r_129_sv2v_reg ,\piso.data_r_128_sv2v_reg ,
  \piso.data_r_127_sv2v_reg ,\piso.data_r_126_sv2v_reg ,\piso.data_r_125_sv2v_reg ,
  \piso.data_r_124_sv2v_reg ,\piso.data_r_123_sv2v_reg ,\piso.data_r_122_sv2v_reg ,
  \piso.data_r_121_sv2v_reg ,\piso.data_r_120_sv2v_reg ,\piso.data_r_119_sv2v_reg ,
  \piso.data_r_118_sv2v_reg ,\piso.data_r_117_sv2v_reg ,\piso.data_r_116_sv2v_reg ,
  \piso.data_r_115_sv2v_reg ,\piso.data_r_114_sv2v_reg ,\piso.data_r_113_sv2v_reg ,
  \piso.data_r_112_sv2v_reg ,\piso.data_r_111_sv2v_reg ,\piso.data_r_110_sv2v_reg ,
  \piso.data_r_109_sv2v_reg ,\piso.data_r_108_sv2v_reg ,\piso.data_r_107_sv2v_reg ,
  \piso.data_r_106_sv2v_reg ,\piso.data_r_105_sv2v_reg ,\piso.data_r_104_sv2v_reg ,
  \piso.data_r_103_sv2v_reg ,\piso.data_r_102_sv2v_reg ,\piso.data_r_101_sv2v_reg ,
  \piso.data_r_100_sv2v_reg ,\piso.data_r_99_sv2v_reg ,\piso.data_r_98_sv2v_reg ,
  \piso.data_r_97_sv2v_reg ,\piso.data_r_96_sv2v_reg ,\piso.data_r_95_sv2v_reg ,
  \piso.data_r_94_sv2v_reg ,\piso.data_r_93_sv2v_reg ,\piso.data_r_92_sv2v_reg ,
  \piso.data_r_91_sv2v_reg ,\piso.data_r_90_sv2v_reg ,\piso.data_r_89_sv2v_reg ,
  \piso.data_r_88_sv2v_reg ,\piso.data_r_87_sv2v_reg ,\piso.data_r_86_sv2v_reg ,
  \piso.data_r_85_sv2v_reg ,\piso.data_r_84_sv2v_reg ,\piso.data_r_83_sv2v_reg ,
  \piso.data_r_82_sv2v_reg ,\piso.data_r_81_sv2v_reg ,\piso.data_r_80_sv2v_reg ,
  \piso.data_r_79_sv2v_reg ,\piso.data_r_78_sv2v_reg ,\piso.data_r_77_sv2v_reg ,
  \piso.data_r_76_sv2v_reg ,\piso.data_r_75_sv2v_reg ,\piso.data_r_74_sv2v_reg ,
  \piso.data_r_73_sv2v_reg ,\piso.data_r_72_sv2v_reg ,\piso.data_r_71_sv2v_reg ,
  \piso.data_r_70_sv2v_reg ,\piso.data_r_69_sv2v_reg ,\piso.data_r_68_sv2v_reg ,\piso.data_r_67_sv2v_reg ,
  \piso.data_r_66_sv2v_reg ,\piso.data_r_65_sv2v_reg ,\piso.data_r_64_sv2v_reg ,
  \piso.data_r_63_sv2v_reg ,\piso.data_r_62_sv2v_reg ,\piso.data_r_61_sv2v_reg ,
  \piso.data_r_60_sv2v_reg ,\piso.data_r_59_sv2v_reg ,\piso.data_r_58_sv2v_reg ,
  \piso.data_r_57_sv2v_reg ,\piso.data_r_56_sv2v_reg ,\piso.data_r_55_sv2v_reg ,
  \piso.data_r_54_sv2v_reg ,\piso.data_r_53_sv2v_reg ,\piso.data_r_52_sv2v_reg ,
  \piso.data_r_51_sv2v_reg ,\piso.data_r_50_sv2v_reg ,\piso.data_r_49_sv2v_reg ,
  \piso.data_r_48_sv2v_reg ,\piso.data_r_47_sv2v_reg ,\piso.data_r_46_sv2v_reg ,
  \piso.data_r_45_sv2v_reg ,\piso.data_r_44_sv2v_reg ,\piso.data_r_43_sv2v_reg ,
  \piso.data_r_42_sv2v_reg ,\piso.data_r_41_sv2v_reg ,\piso.data_r_40_sv2v_reg ,
  \piso.data_r_39_sv2v_reg ,\piso.data_r_38_sv2v_reg ,\piso.data_r_37_sv2v_reg ,
  \piso.data_r_36_sv2v_reg ,\piso.data_r_35_sv2v_reg ,\piso.data_r_34_sv2v_reg ,
  \piso.data_r_33_sv2v_reg ,\piso.data_r_32_sv2v_reg ,\piso.data_r_31_sv2v_reg ,
  \piso.data_r_30_sv2v_reg ,\piso.data_r_29_sv2v_reg ,\piso.data_r_28_sv2v_reg ,\piso.data_r_27_sv2v_reg ,
  \piso.data_r_26_sv2v_reg ,\piso.data_r_25_sv2v_reg ,\piso.data_r_24_sv2v_reg ,
  \piso.data_r_23_sv2v_reg ,\piso.data_r_22_sv2v_reg ,\piso.data_r_21_sv2v_reg ,
  \piso.data_r_20_sv2v_reg ,\piso.data_r_19_sv2v_reg ,\piso.data_r_18_sv2v_reg ,
  \piso.data_r_17_sv2v_reg ,\piso.data_r_16_sv2v_reg ,\piso.data_r_15_sv2v_reg ,
  \piso.data_r_14_sv2v_reg ,\piso.data_r_13_sv2v_reg ,\piso.data_r_12_sv2v_reg ,
  \piso.data_r_11_sv2v_reg ,\piso.data_r_10_sv2v_reg ,\piso.data_r_9_sv2v_reg ,
  \piso.data_r_8_sv2v_reg ,\piso.data_r_7_sv2v_reg ,\piso.data_r_6_sv2v_reg ,
  \piso.data_r_5_sv2v_reg ,\piso.data_r_4_sv2v_reg ,\piso.data_r_3_sv2v_reg ,
  \piso.data_r_2_sv2v_reg ,\piso.data_r_1_sv2v_reg ,\piso.data_r_0_sv2v_reg ,
  \piso.shift_ctr_r_4_sv2v_reg ,\piso.shift_ctr_r_3_sv2v_reg ,\piso.shift_ctr_r_2_sv2v_reg ,
  \piso.shift_ctr_r_1_sv2v_reg ,\piso.shift_ctr_r_0_sv2v_reg ;
  assign valid_o = valid_o_sv2v_reg;
  assign \piso.data_r [511] = \piso.data_r_511_sv2v_reg ;
  assign \piso.data_r [510] = \piso.data_r_510_sv2v_reg ;
  assign \piso.data_r [509] = \piso.data_r_509_sv2v_reg ;
  assign \piso.data_r [508] = \piso.data_r_508_sv2v_reg ;
  assign \piso.data_r [507] = \piso.data_r_507_sv2v_reg ;
  assign \piso.data_r [506] = \piso.data_r_506_sv2v_reg ;
  assign \piso.data_r [505] = \piso.data_r_505_sv2v_reg ;
  assign \piso.data_r [504] = \piso.data_r_504_sv2v_reg ;
  assign \piso.data_r [503] = \piso.data_r_503_sv2v_reg ;
  assign \piso.data_r [502] = \piso.data_r_502_sv2v_reg ;
  assign \piso.data_r [501] = \piso.data_r_501_sv2v_reg ;
  assign \piso.data_r [500] = \piso.data_r_500_sv2v_reg ;
  assign \piso.data_r [499] = \piso.data_r_499_sv2v_reg ;
  assign \piso.data_r [498] = \piso.data_r_498_sv2v_reg ;
  assign \piso.data_r [497] = \piso.data_r_497_sv2v_reg ;
  assign \piso.data_r [496] = \piso.data_r_496_sv2v_reg ;
  assign \piso.data_r [495] = \piso.data_r_495_sv2v_reg ;
  assign \piso.data_r [494] = \piso.data_r_494_sv2v_reg ;
  assign \piso.data_r [493] = \piso.data_r_493_sv2v_reg ;
  assign \piso.data_r [492] = \piso.data_r_492_sv2v_reg ;
  assign \piso.data_r [491] = \piso.data_r_491_sv2v_reg ;
  assign \piso.data_r [490] = \piso.data_r_490_sv2v_reg ;
  assign \piso.data_r [489] = \piso.data_r_489_sv2v_reg ;
  assign \piso.data_r [488] = \piso.data_r_488_sv2v_reg ;
  assign \piso.data_r [487] = \piso.data_r_487_sv2v_reg ;
  assign \piso.data_r [486] = \piso.data_r_486_sv2v_reg ;
  assign \piso.data_r [485] = \piso.data_r_485_sv2v_reg ;
  assign \piso.data_r [484] = \piso.data_r_484_sv2v_reg ;
  assign \piso.data_r [483] = \piso.data_r_483_sv2v_reg ;
  assign \piso.data_r [482] = \piso.data_r_482_sv2v_reg ;
  assign \piso.data_r [481] = \piso.data_r_481_sv2v_reg ;
  assign \piso.data_r [480] = \piso.data_r_480_sv2v_reg ;
  assign \piso.data_r [479] = \piso.data_r_479_sv2v_reg ;
  assign \piso.data_r [478] = \piso.data_r_478_sv2v_reg ;
  assign \piso.data_r [477] = \piso.data_r_477_sv2v_reg ;
  assign \piso.data_r [476] = \piso.data_r_476_sv2v_reg ;
  assign \piso.data_r [475] = \piso.data_r_475_sv2v_reg ;
  assign \piso.data_r [474] = \piso.data_r_474_sv2v_reg ;
  assign \piso.data_r [473] = \piso.data_r_473_sv2v_reg ;
  assign \piso.data_r [472] = \piso.data_r_472_sv2v_reg ;
  assign \piso.data_r [471] = \piso.data_r_471_sv2v_reg ;
  assign \piso.data_r [470] = \piso.data_r_470_sv2v_reg ;
  assign \piso.data_r [469] = \piso.data_r_469_sv2v_reg ;
  assign \piso.data_r [468] = \piso.data_r_468_sv2v_reg ;
  assign \piso.data_r [467] = \piso.data_r_467_sv2v_reg ;
  assign \piso.data_r [466] = \piso.data_r_466_sv2v_reg ;
  assign \piso.data_r [465] = \piso.data_r_465_sv2v_reg ;
  assign \piso.data_r [464] = \piso.data_r_464_sv2v_reg ;
  assign \piso.data_r [463] = \piso.data_r_463_sv2v_reg ;
  assign \piso.data_r [462] = \piso.data_r_462_sv2v_reg ;
  assign \piso.data_r [461] = \piso.data_r_461_sv2v_reg ;
  assign \piso.data_r [460] = \piso.data_r_460_sv2v_reg ;
  assign \piso.data_r [459] = \piso.data_r_459_sv2v_reg ;
  assign \piso.data_r [458] = \piso.data_r_458_sv2v_reg ;
  assign \piso.data_r [457] = \piso.data_r_457_sv2v_reg ;
  assign \piso.data_r [456] = \piso.data_r_456_sv2v_reg ;
  assign \piso.data_r [455] = \piso.data_r_455_sv2v_reg ;
  assign \piso.data_r [454] = \piso.data_r_454_sv2v_reg ;
  assign \piso.data_r [453] = \piso.data_r_453_sv2v_reg ;
  assign \piso.data_r [452] = \piso.data_r_452_sv2v_reg ;
  assign \piso.data_r [451] = \piso.data_r_451_sv2v_reg ;
  assign \piso.data_r [450] = \piso.data_r_450_sv2v_reg ;
  assign \piso.data_r [449] = \piso.data_r_449_sv2v_reg ;
  assign \piso.data_r [448] = \piso.data_r_448_sv2v_reg ;
  assign \piso.data_r [447] = \piso.data_r_447_sv2v_reg ;
  assign \piso.data_r [446] = \piso.data_r_446_sv2v_reg ;
  assign \piso.data_r [445] = \piso.data_r_445_sv2v_reg ;
  assign \piso.data_r [444] = \piso.data_r_444_sv2v_reg ;
  assign \piso.data_r [443] = \piso.data_r_443_sv2v_reg ;
  assign \piso.data_r [442] = \piso.data_r_442_sv2v_reg ;
  assign \piso.data_r [441] = \piso.data_r_441_sv2v_reg ;
  assign \piso.data_r [440] = \piso.data_r_440_sv2v_reg ;
  assign \piso.data_r [439] = \piso.data_r_439_sv2v_reg ;
  assign \piso.data_r [438] = \piso.data_r_438_sv2v_reg ;
  assign \piso.data_r [437] = \piso.data_r_437_sv2v_reg ;
  assign \piso.data_r [436] = \piso.data_r_436_sv2v_reg ;
  assign \piso.data_r [435] = \piso.data_r_435_sv2v_reg ;
  assign \piso.data_r [434] = \piso.data_r_434_sv2v_reg ;
  assign \piso.data_r [433] = \piso.data_r_433_sv2v_reg ;
  assign \piso.data_r [432] = \piso.data_r_432_sv2v_reg ;
  assign \piso.data_r [431] = \piso.data_r_431_sv2v_reg ;
  assign \piso.data_r [430] = \piso.data_r_430_sv2v_reg ;
  assign \piso.data_r [429] = \piso.data_r_429_sv2v_reg ;
  assign \piso.data_r [428] = \piso.data_r_428_sv2v_reg ;
  assign \piso.data_r [427] = \piso.data_r_427_sv2v_reg ;
  assign \piso.data_r [426] = \piso.data_r_426_sv2v_reg ;
  assign \piso.data_r [425] = \piso.data_r_425_sv2v_reg ;
  assign \piso.data_r [424] = \piso.data_r_424_sv2v_reg ;
  assign \piso.data_r [423] = \piso.data_r_423_sv2v_reg ;
  assign \piso.data_r [422] = \piso.data_r_422_sv2v_reg ;
  assign \piso.data_r [421] = \piso.data_r_421_sv2v_reg ;
  assign \piso.data_r [420] = \piso.data_r_420_sv2v_reg ;
  assign \piso.data_r [419] = \piso.data_r_419_sv2v_reg ;
  assign \piso.data_r [418] = \piso.data_r_418_sv2v_reg ;
  assign \piso.data_r [417] = \piso.data_r_417_sv2v_reg ;
  assign \piso.data_r [416] = \piso.data_r_416_sv2v_reg ;
  assign \piso.data_r [415] = \piso.data_r_415_sv2v_reg ;
  assign \piso.data_r [414] = \piso.data_r_414_sv2v_reg ;
  assign \piso.data_r [413] = \piso.data_r_413_sv2v_reg ;
  assign \piso.data_r [412] = \piso.data_r_412_sv2v_reg ;
  assign \piso.data_r [411] = \piso.data_r_411_sv2v_reg ;
  assign \piso.data_r [410] = \piso.data_r_410_sv2v_reg ;
  assign \piso.data_r [409] = \piso.data_r_409_sv2v_reg ;
  assign \piso.data_r [408] = \piso.data_r_408_sv2v_reg ;
  assign \piso.data_r [407] = \piso.data_r_407_sv2v_reg ;
  assign \piso.data_r [406] = \piso.data_r_406_sv2v_reg ;
  assign \piso.data_r [405] = \piso.data_r_405_sv2v_reg ;
  assign \piso.data_r [404] = \piso.data_r_404_sv2v_reg ;
  assign \piso.data_r [403] = \piso.data_r_403_sv2v_reg ;
  assign \piso.data_r [402] = \piso.data_r_402_sv2v_reg ;
  assign \piso.data_r [401] = \piso.data_r_401_sv2v_reg ;
  assign \piso.data_r [400] = \piso.data_r_400_sv2v_reg ;
  assign \piso.data_r [399] = \piso.data_r_399_sv2v_reg ;
  assign \piso.data_r [398] = \piso.data_r_398_sv2v_reg ;
  assign \piso.data_r [397] = \piso.data_r_397_sv2v_reg ;
  assign \piso.data_r [396] = \piso.data_r_396_sv2v_reg ;
  assign \piso.data_r [395] = \piso.data_r_395_sv2v_reg ;
  assign \piso.data_r [394] = \piso.data_r_394_sv2v_reg ;
  assign \piso.data_r [393] = \piso.data_r_393_sv2v_reg ;
  assign \piso.data_r [392] = \piso.data_r_392_sv2v_reg ;
  assign \piso.data_r [391] = \piso.data_r_391_sv2v_reg ;
  assign \piso.data_r [390] = \piso.data_r_390_sv2v_reg ;
  assign \piso.data_r [389] = \piso.data_r_389_sv2v_reg ;
  assign \piso.data_r [388] = \piso.data_r_388_sv2v_reg ;
  assign \piso.data_r [387] = \piso.data_r_387_sv2v_reg ;
  assign \piso.data_r [386] = \piso.data_r_386_sv2v_reg ;
  assign \piso.data_r [385] = \piso.data_r_385_sv2v_reg ;
  assign \piso.data_r [384] = \piso.data_r_384_sv2v_reg ;
  assign \piso.data_r [383] = \piso.data_r_383_sv2v_reg ;
  assign \piso.data_r [382] = \piso.data_r_382_sv2v_reg ;
  assign \piso.data_r [381] = \piso.data_r_381_sv2v_reg ;
  assign \piso.data_r [380] = \piso.data_r_380_sv2v_reg ;
  assign \piso.data_r [379] = \piso.data_r_379_sv2v_reg ;
  assign \piso.data_r [378] = \piso.data_r_378_sv2v_reg ;
  assign \piso.data_r [377] = \piso.data_r_377_sv2v_reg ;
  assign \piso.data_r [376] = \piso.data_r_376_sv2v_reg ;
  assign \piso.data_r [375] = \piso.data_r_375_sv2v_reg ;
  assign \piso.data_r [374] = \piso.data_r_374_sv2v_reg ;
  assign \piso.data_r [373] = \piso.data_r_373_sv2v_reg ;
  assign \piso.data_r [372] = \piso.data_r_372_sv2v_reg ;
  assign \piso.data_r [371] = \piso.data_r_371_sv2v_reg ;
  assign \piso.data_r [370] = \piso.data_r_370_sv2v_reg ;
  assign \piso.data_r [369] = \piso.data_r_369_sv2v_reg ;
  assign \piso.data_r [368] = \piso.data_r_368_sv2v_reg ;
  assign \piso.data_r [367] = \piso.data_r_367_sv2v_reg ;
  assign \piso.data_r [366] = \piso.data_r_366_sv2v_reg ;
  assign \piso.data_r [365] = \piso.data_r_365_sv2v_reg ;
  assign \piso.data_r [364] = \piso.data_r_364_sv2v_reg ;
  assign \piso.data_r [363] = \piso.data_r_363_sv2v_reg ;
  assign \piso.data_r [362] = \piso.data_r_362_sv2v_reg ;
  assign \piso.data_r [361] = \piso.data_r_361_sv2v_reg ;
  assign \piso.data_r [360] = \piso.data_r_360_sv2v_reg ;
  assign \piso.data_r [359] = \piso.data_r_359_sv2v_reg ;
  assign \piso.data_r [358] = \piso.data_r_358_sv2v_reg ;
  assign \piso.data_r [357] = \piso.data_r_357_sv2v_reg ;
  assign \piso.data_r [356] = \piso.data_r_356_sv2v_reg ;
  assign \piso.data_r [355] = \piso.data_r_355_sv2v_reg ;
  assign \piso.data_r [354] = \piso.data_r_354_sv2v_reg ;
  assign \piso.data_r [353] = \piso.data_r_353_sv2v_reg ;
  assign \piso.data_r [352] = \piso.data_r_352_sv2v_reg ;
  assign \piso.data_r [351] = \piso.data_r_351_sv2v_reg ;
  assign \piso.data_r [350] = \piso.data_r_350_sv2v_reg ;
  assign \piso.data_r [349] = \piso.data_r_349_sv2v_reg ;
  assign \piso.data_r [348] = \piso.data_r_348_sv2v_reg ;
  assign \piso.data_r [347] = \piso.data_r_347_sv2v_reg ;
  assign \piso.data_r [346] = \piso.data_r_346_sv2v_reg ;
  assign \piso.data_r [345] = \piso.data_r_345_sv2v_reg ;
  assign \piso.data_r [344] = \piso.data_r_344_sv2v_reg ;
  assign \piso.data_r [343] = \piso.data_r_343_sv2v_reg ;
  assign \piso.data_r [342] = \piso.data_r_342_sv2v_reg ;
  assign \piso.data_r [341] = \piso.data_r_341_sv2v_reg ;
  assign \piso.data_r [340] = \piso.data_r_340_sv2v_reg ;
  assign \piso.data_r [339] = \piso.data_r_339_sv2v_reg ;
  assign \piso.data_r [338] = \piso.data_r_338_sv2v_reg ;
  assign \piso.data_r [337] = \piso.data_r_337_sv2v_reg ;
  assign \piso.data_r [336] = \piso.data_r_336_sv2v_reg ;
  assign \piso.data_r [335] = \piso.data_r_335_sv2v_reg ;
  assign \piso.data_r [334] = \piso.data_r_334_sv2v_reg ;
  assign \piso.data_r [333] = \piso.data_r_333_sv2v_reg ;
  assign \piso.data_r [332] = \piso.data_r_332_sv2v_reg ;
  assign \piso.data_r [331] = \piso.data_r_331_sv2v_reg ;
  assign \piso.data_r [330] = \piso.data_r_330_sv2v_reg ;
  assign \piso.data_r [329] = \piso.data_r_329_sv2v_reg ;
  assign \piso.data_r [328] = \piso.data_r_328_sv2v_reg ;
  assign \piso.data_r [327] = \piso.data_r_327_sv2v_reg ;
  assign \piso.data_r [326] = \piso.data_r_326_sv2v_reg ;
  assign \piso.data_r [325] = \piso.data_r_325_sv2v_reg ;
  assign \piso.data_r [324] = \piso.data_r_324_sv2v_reg ;
  assign \piso.data_r [323] = \piso.data_r_323_sv2v_reg ;
  assign \piso.data_r [322] = \piso.data_r_322_sv2v_reg ;
  assign \piso.data_r [321] = \piso.data_r_321_sv2v_reg ;
  assign \piso.data_r [320] = \piso.data_r_320_sv2v_reg ;
  assign \piso.data_r [319] = \piso.data_r_319_sv2v_reg ;
  assign \piso.data_r [318] = \piso.data_r_318_sv2v_reg ;
  assign \piso.data_r [317] = \piso.data_r_317_sv2v_reg ;
  assign \piso.data_r [316] = \piso.data_r_316_sv2v_reg ;
  assign \piso.data_r [315] = \piso.data_r_315_sv2v_reg ;
  assign \piso.data_r [314] = \piso.data_r_314_sv2v_reg ;
  assign \piso.data_r [313] = \piso.data_r_313_sv2v_reg ;
  assign \piso.data_r [312] = \piso.data_r_312_sv2v_reg ;
  assign \piso.data_r [311] = \piso.data_r_311_sv2v_reg ;
  assign \piso.data_r [310] = \piso.data_r_310_sv2v_reg ;
  assign \piso.data_r [309] = \piso.data_r_309_sv2v_reg ;
  assign \piso.data_r [308] = \piso.data_r_308_sv2v_reg ;
  assign \piso.data_r [307] = \piso.data_r_307_sv2v_reg ;
  assign \piso.data_r [306] = \piso.data_r_306_sv2v_reg ;
  assign \piso.data_r [305] = \piso.data_r_305_sv2v_reg ;
  assign \piso.data_r [304] = \piso.data_r_304_sv2v_reg ;
  assign \piso.data_r [303] = \piso.data_r_303_sv2v_reg ;
  assign \piso.data_r [302] = \piso.data_r_302_sv2v_reg ;
  assign \piso.data_r [301] = \piso.data_r_301_sv2v_reg ;
  assign \piso.data_r [300] = \piso.data_r_300_sv2v_reg ;
  assign \piso.data_r [299] = \piso.data_r_299_sv2v_reg ;
  assign \piso.data_r [298] = \piso.data_r_298_sv2v_reg ;
  assign \piso.data_r [297] = \piso.data_r_297_sv2v_reg ;
  assign \piso.data_r [296] = \piso.data_r_296_sv2v_reg ;
  assign \piso.data_r [295] = \piso.data_r_295_sv2v_reg ;
  assign \piso.data_r [294] = \piso.data_r_294_sv2v_reg ;
  assign \piso.data_r [293] = \piso.data_r_293_sv2v_reg ;
  assign \piso.data_r [292] = \piso.data_r_292_sv2v_reg ;
  assign \piso.data_r [291] = \piso.data_r_291_sv2v_reg ;
  assign \piso.data_r [290] = \piso.data_r_290_sv2v_reg ;
  assign \piso.data_r [289] = \piso.data_r_289_sv2v_reg ;
  assign \piso.data_r [288] = \piso.data_r_288_sv2v_reg ;
  assign \piso.data_r [287] = \piso.data_r_287_sv2v_reg ;
  assign \piso.data_r [286] = \piso.data_r_286_sv2v_reg ;
  assign \piso.data_r [285] = \piso.data_r_285_sv2v_reg ;
  assign \piso.data_r [284] = \piso.data_r_284_sv2v_reg ;
  assign \piso.data_r [283] = \piso.data_r_283_sv2v_reg ;
  assign \piso.data_r [282] = \piso.data_r_282_sv2v_reg ;
  assign \piso.data_r [281] = \piso.data_r_281_sv2v_reg ;
  assign \piso.data_r [280] = \piso.data_r_280_sv2v_reg ;
  assign \piso.data_r [279] = \piso.data_r_279_sv2v_reg ;
  assign \piso.data_r [278] = \piso.data_r_278_sv2v_reg ;
  assign \piso.data_r [277] = \piso.data_r_277_sv2v_reg ;
  assign \piso.data_r [276] = \piso.data_r_276_sv2v_reg ;
  assign \piso.data_r [275] = \piso.data_r_275_sv2v_reg ;
  assign \piso.data_r [274] = \piso.data_r_274_sv2v_reg ;
  assign \piso.data_r [273] = \piso.data_r_273_sv2v_reg ;
  assign \piso.data_r [272] = \piso.data_r_272_sv2v_reg ;
  assign \piso.data_r [271] = \piso.data_r_271_sv2v_reg ;
  assign \piso.data_r [270] = \piso.data_r_270_sv2v_reg ;
  assign \piso.data_r [269] = \piso.data_r_269_sv2v_reg ;
  assign \piso.data_r [268] = \piso.data_r_268_sv2v_reg ;
  assign \piso.data_r [267] = \piso.data_r_267_sv2v_reg ;
  assign \piso.data_r [266] = \piso.data_r_266_sv2v_reg ;
  assign \piso.data_r [265] = \piso.data_r_265_sv2v_reg ;
  assign \piso.data_r [264] = \piso.data_r_264_sv2v_reg ;
  assign \piso.data_r [263] = \piso.data_r_263_sv2v_reg ;
  assign \piso.data_r [262] = \piso.data_r_262_sv2v_reg ;
  assign \piso.data_r [261] = \piso.data_r_261_sv2v_reg ;
  assign \piso.data_r [260] = \piso.data_r_260_sv2v_reg ;
  assign \piso.data_r [259] = \piso.data_r_259_sv2v_reg ;
  assign \piso.data_r [258] = \piso.data_r_258_sv2v_reg ;
  assign \piso.data_r [257] = \piso.data_r_257_sv2v_reg ;
  assign \piso.data_r [256] = \piso.data_r_256_sv2v_reg ;
  assign \piso.data_r [255] = \piso.data_r_255_sv2v_reg ;
  assign \piso.data_r [254] = \piso.data_r_254_sv2v_reg ;
  assign \piso.data_r [253] = \piso.data_r_253_sv2v_reg ;
  assign \piso.data_r [252] = \piso.data_r_252_sv2v_reg ;
  assign \piso.data_r [251] = \piso.data_r_251_sv2v_reg ;
  assign \piso.data_r [250] = \piso.data_r_250_sv2v_reg ;
  assign \piso.data_r [249] = \piso.data_r_249_sv2v_reg ;
  assign \piso.data_r [248] = \piso.data_r_248_sv2v_reg ;
  assign \piso.data_r [247] = \piso.data_r_247_sv2v_reg ;
  assign \piso.data_r [246] = \piso.data_r_246_sv2v_reg ;
  assign \piso.data_r [245] = \piso.data_r_245_sv2v_reg ;
  assign \piso.data_r [244] = \piso.data_r_244_sv2v_reg ;
  assign \piso.data_r [243] = \piso.data_r_243_sv2v_reg ;
  assign \piso.data_r [242] = \piso.data_r_242_sv2v_reg ;
  assign \piso.data_r [241] = \piso.data_r_241_sv2v_reg ;
  assign \piso.data_r [240] = \piso.data_r_240_sv2v_reg ;
  assign \piso.data_r [239] = \piso.data_r_239_sv2v_reg ;
  assign \piso.data_r [238] = \piso.data_r_238_sv2v_reg ;
  assign \piso.data_r [237] = \piso.data_r_237_sv2v_reg ;
  assign \piso.data_r [236] = \piso.data_r_236_sv2v_reg ;
  assign \piso.data_r [235] = \piso.data_r_235_sv2v_reg ;
  assign \piso.data_r [234] = \piso.data_r_234_sv2v_reg ;
  assign \piso.data_r [233] = \piso.data_r_233_sv2v_reg ;
  assign \piso.data_r [232] = \piso.data_r_232_sv2v_reg ;
  assign \piso.data_r [231] = \piso.data_r_231_sv2v_reg ;
  assign \piso.data_r [230] = \piso.data_r_230_sv2v_reg ;
  assign \piso.data_r [229] = \piso.data_r_229_sv2v_reg ;
  assign \piso.data_r [228] = \piso.data_r_228_sv2v_reg ;
  assign \piso.data_r [227] = \piso.data_r_227_sv2v_reg ;
  assign \piso.data_r [226] = \piso.data_r_226_sv2v_reg ;
  assign \piso.data_r [225] = \piso.data_r_225_sv2v_reg ;
  assign \piso.data_r [224] = \piso.data_r_224_sv2v_reg ;
  assign \piso.data_r [223] = \piso.data_r_223_sv2v_reg ;
  assign \piso.data_r [222] = \piso.data_r_222_sv2v_reg ;
  assign \piso.data_r [221] = \piso.data_r_221_sv2v_reg ;
  assign \piso.data_r [220] = \piso.data_r_220_sv2v_reg ;
  assign \piso.data_r [219] = \piso.data_r_219_sv2v_reg ;
  assign \piso.data_r [218] = \piso.data_r_218_sv2v_reg ;
  assign \piso.data_r [217] = \piso.data_r_217_sv2v_reg ;
  assign \piso.data_r [216] = \piso.data_r_216_sv2v_reg ;
  assign \piso.data_r [215] = \piso.data_r_215_sv2v_reg ;
  assign \piso.data_r [214] = \piso.data_r_214_sv2v_reg ;
  assign \piso.data_r [213] = \piso.data_r_213_sv2v_reg ;
  assign \piso.data_r [212] = \piso.data_r_212_sv2v_reg ;
  assign \piso.data_r [211] = \piso.data_r_211_sv2v_reg ;
  assign \piso.data_r [210] = \piso.data_r_210_sv2v_reg ;
  assign \piso.data_r [209] = \piso.data_r_209_sv2v_reg ;
  assign \piso.data_r [208] = \piso.data_r_208_sv2v_reg ;
  assign \piso.data_r [207] = \piso.data_r_207_sv2v_reg ;
  assign \piso.data_r [206] = \piso.data_r_206_sv2v_reg ;
  assign \piso.data_r [205] = \piso.data_r_205_sv2v_reg ;
  assign \piso.data_r [204] = \piso.data_r_204_sv2v_reg ;
  assign \piso.data_r [203] = \piso.data_r_203_sv2v_reg ;
  assign \piso.data_r [202] = \piso.data_r_202_sv2v_reg ;
  assign \piso.data_r [201] = \piso.data_r_201_sv2v_reg ;
  assign \piso.data_r [200] = \piso.data_r_200_sv2v_reg ;
  assign \piso.data_r [199] = \piso.data_r_199_sv2v_reg ;
  assign \piso.data_r [198] = \piso.data_r_198_sv2v_reg ;
  assign \piso.data_r [197] = \piso.data_r_197_sv2v_reg ;
  assign \piso.data_r [196] = \piso.data_r_196_sv2v_reg ;
  assign \piso.data_r [195] = \piso.data_r_195_sv2v_reg ;
  assign \piso.data_r [194] = \piso.data_r_194_sv2v_reg ;
  assign \piso.data_r [193] = \piso.data_r_193_sv2v_reg ;
  assign \piso.data_r [192] = \piso.data_r_192_sv2v_reg ;
  assign \piso.data_r [191] = \piso.data_r_191_sv2v_reg ;
  assign \piso.data_r [190] = \piso.data_r_190_sv2v_reg ;
  assign \piso.data_r [189] = \piso.data_r_189_sv2v_reg ;
  assign \piso.data_r [188] = \piso.data_r_188_sv2v_reg ;
  assign \piso.data_r [187] = \piso.data_r_187_sv2v_reg ;
  assign \piso.data_r [186] = \piso.data_r_186_sv2v_reg ;
  assign \piso.data_r [185] = \piso.data_r_185_sv2v_reg ;
  assign \piso.data_r [184] = \piso.data_r_184_sv2v_reg ;
  assign \piso.data_r [183] = \piso.data_r_183_sv2v_reg ;
  assign \piso.data_r [182] = \piso.data_r_182_sv2v_reg ;
  assign \piso.data_r [181] = \piso.data_r_181_sv2v_reg ;
  assign \piso.data_r [180] = \piso.data_r_180_sv2v_reg ;
  assign \piso.data_r [179] = \piso.data_r_179_sv2v_reg ;
  assign \piso.data_r [178] = \piso.data_r_178_sv2v_reg ;
  assign \piso.data_r [177] = \piso.data_r_177_sv2v_reg ;
  assign \piso.data_r [176] = \piso.data_r_176_sv2v_reg ;
  assign \piso.data_r [175] = \piso.data_r_175_sv2v_reg ;
  assign \piso.data_r [174] = \piso.data_r_174_sv2v_reg ;
  assign \piso.data_r [173] = \piso.data_r_173_sv2v_reg ;
  assign \piso.data_r [172] = \piso.data_r_172_sv2v_reg ;
  assign \piso.data_r [171] = \piso.data_r_171_sv2v_reg ;
  assign \piso.data_r [170] = \piso.data_r_170_sv2v_reg ;
  assign \piso.data_r [169] = \piso.data_r_169_sv2v_reg ;
  assign \piso.data_r [168] = \piso.data_r_168_sv2v_reg ;
  assign \piso.data_r [167] = \piso.data_r_167_sv2v_reg ;
  assign \piso.data_r [166] = \piso.data_r_166_sv2v_reg ;
  assign \piso.data_r [165] = \piso.data_r_165_sv2v_reg ;
  assign \piso.data_r [164] = \piso.data_r_164_sv2v_reg ;
  assign \piso.data_r [163] = \piso.data_r_163_sv2v_reg ;
  assign \piso.data_r [162] = \piso.data_r_162_sv2v_reg ;
  assign \piso.data_r [161] = \piso.data_r_161_sv2v_reg ;
  assign \piso.data_r [160] = \piso.data_r_160_sv2v_reg ;
  assign \piso.data_r [159] = \piso.data_r_159_sv2v_reg ;
  assign \piso.data_r [158] = \piso.data_r_158_sv2v_reg ;
  assign \piso.data_r [157] = \piso.data_r_157_sv2v_reg ;
  assign \piso.data_r [156] = \piso.data_r_156_sv2v_reg ;
  assign \piso.data_r [155] = \piso.data_r_155_sv2v_reg ;
  assign \piso.data_r [154] = \piso.data_r_154_sv2v_reg ;
  assign \piso.data_r [153] = \piso.data_r_153_sv2v_reg ;
  assign \piso.data_r [152] = \piso.data_r_152_sv2v_reg ;
  assign \piso.data_r [151] = \piso.data_r_151_sv2v_reg ;
  assign \piso.data_r [150] = \piso.data_r_150_sv2v_reg ;
  assign \piso.data_r [149] = \piso.data_r_149_sv2v_reg ;
  assign \piso.data_r [148] = \piso.data_r_148_sv2v_reg ;
  assign \piso.data_r [147] = \piso.data_r_147_sv2v_reg ;
  assign \piso.data_r [146] = \piso.data_r_146_sv2v_reg ;
  assign \piso.data_r [145] = \piso.data_r_145_sv2v_reg ;
  assign \piso.data_r [144] = \piso.data_r_144_sv2v_reg ;
  assign \piso.data_r [143] = \piso.data_r_143_sv2v_reg ;
  assign \piso.data_r [142] = \piso.data_r_142_sv2v_reg ;
  assign \piso.data_r [141] = \piso.data_r_141_sv2v_reg ;
  assign \piso.data_r [140] = \piso.data_r_140_sv2v_reg ;
  assign \piso.data_r [139] = \piso.data_r_139_sv2v_reg ;
  assign \piso.data_r [138] = \piso.data_r_138_sv2v_reg ;
  assign \piso.data_r [137] = \piso.data_r_137_sv2v_reg ;
  assign \piso.data_r [136] = \piso.data_r_136_sv2v_reg ;
  assign \piso.data_r [135] = \piso.data_r_135_sv2v_reg ;
  assign \piso.data_r [134] = \piso.data_r_134_sv2v_reg ;
  assign \piso.data_r [133] = \piso.data_r_133_sv2v_reg ;
  assign \piso.data_r [132] = \piso.data_r_132_sv2v_reg ;
  assign \piso.data_r [131] = \piso.data_r_131_sv2v_reg ;
  assign \piso.data_r [130] = \piso.data_r_130_sv2v_reg ;
  assign \piso.data_r [129] = \piso.data_r_129_sv2v_reg ;
  assign \piso.data_r [128] = \piso.data_r_128_sv2v_reg ;
  assign \piso.data_r [127] = \piso.data_r_127_sv2v_reg ;
  assign \piso.data_r [126] = \piso.data_r_126_sv2v_reg ;
  assign \piso.data_r [125] = \piso.data_r_125_sv2v_reg ;
  assign \piso.data_r [124] = \piso.data_r_124_sv2v_reg ;
  assign \piso.data_r [123] = \piso.data_r_123_sv2v_reg ;
  assign \piso.data_r [122] = \piso.data_r_122_sv2v_reg ;
  assign \piso.data_r [121] = \piso.data_r_121_sv2v_reg ;
  assign \piso.data_r [120] = \piso.data_r_120_sv2v_reg ;
  assign \piso.data_r [119] = \piso.data_r_119_sv2v_reg ;
  assign \piso.data_r [118] = \piso.data_r_118_sv2v_reg ;
  assign \piso.data_r [117] = \piso.data_r_117_sv2v_reg ;
  assign \piso.data_r [116] = \piso.data_r_116_sv2v_reg ;
  assign \piso.data_r [115] = \piso.data_r_115_sv2v_reg ;
  assign \piso.data_r [114] = \piso.data_r_114_sv2v_reg ;
  assign \piso.data_r [113] = \piso.data_r_113_sv2v_reg ;
  assign \piso.data_r [112] = \piso.data_r_112_sv2v_reg ;
  assign \piso.data_r [111] = \piso.data_r_111_sv2v_reg ;
  assign \piso.data_r [110] = \piso.data_r_110_sv2v_reg ;
  assign \piso.data_r [109] = \piso.data_r_109_sv2v_reg ;
  assign \piso.data_r [108] = \piso.data_r_108_sv2v_reg ;
  assign \piso.data_r [107] = \piso.data_r_107_sv2v_reg ;
  assign \piso.data_r [106] = \piso.data_r_106_sv2v_reg ;
  assign \piso.data_r [105] = \piso.data_r_105_sv2v_reg ;
  assign \piso.data_r [104] = \piso.data_r_104_sv2v_reg ;
  assign \piso.data_r [103] = \piso.data_r_103_sv2v_reg ;
  assign \piso.data_r [102] = \piso.data_r_102_sv2v_reg ;
  assign \piso.data_r [101] = \piso.data_r_101_sv2v_reg ;
  assign \piso.data_r [100] = \piso.data_r_100_sv2v_reg ;
  assign \piso.data_r [99] = \piso.data_r_99_sv2v_reg ;
  assign \piso.data_r [98] = \piso.data_r_98_sv2v_reg ;
  assign \piso.data_r [97] = \piso.data_r_97_sv2v_reg ;
  assign \piso.data_r [96] = \piso.data_r_96_sv2v_reg ;
  assign \piso.data_r [95] = \piso.data_r_95_sv2v_reg ;
  assign \piso.data_r [94] = \piso.data_r_94_sv2v_reg ;
  assign \piso.data_r [93] = \piso.data_r_93_sv2v_reg ;
  assign \piso.data_r [92] = \piso.data_r_92_sv2v_reg ;
  assign \piso.data_r [91] = \piso.data_r_91_sv2v_reg ;
  assign \piso.data_r [90] = \piso.data_r_90_sv2v_reg ;
  assign \piso.data_r [89] = \piso.data_r_89_sv2v_reg ;
  assign \piso.data_r [88] = \piso.data_r_88_sv2v_reg ;
  assign \piso.data_r [87] = \piso.data_r_87_sv2v_reg ;
  assign \piso.data_r [86] = \piso.data_r_86_sv2v_reg ;
  assign \piso.data_r [85] = \piso.data_r_85_sv2v_reg ;
  assign \piso.data_r [84] = \piso.data_r_84_sv2v_reg ;
  assign \piso.data_r [83] = \piso.data_r_83_sv2v_reg ;
  assign \piso.data_r [82] = \piso.data_r_82_sv2v_reg ;
  assign \piso.data_r [81] = \piso.data_r_81_sv2v_reg ;
  assign \piso.data_r [80] = \piso.data_r_80_sv2v_reg ;
  assign \piso.data_r [79] = \piso.data_r_79_sv2v_reg ;
  assign \piso.data_r [78] = \piso.data_r_78_sv2v_reg ;
  assign \piso.data_r [77] = \piso.data_r_77_sv2v_reg ;
  assign \piso.data_r [76] = \piso.data_r_76_sv2v_reg ;
  assign \piso.data_r [75] = \piso.data_r_75_sv2v_reg ;
  assign \piso.data_r [74] = \piso.data_r_74_sv2v_reg ;
  assign \piso.data_r [73] = \piso.data_r_73_sv2v_reg ;
  assign \piso.data_r [72] = \piso.data_r_72_sv2v_reg ;
  assign \piso.data_r [71] = \piso.data_r_71_sv2v_reg ;
  assign \piso.data_r [70] = \piso.data_r_70_sv2v_reg ;
  assign \piso.data_r [69] = \piso.data_r_69_sv2v_reg ;
  assign \piso.data_r [68] = \piso.data_r_68_sv2v_reg ;
  assign \piso.data_r [67] = \piso.data_r_67_sv2v_reg ;
  assign \piso.data_r [66] = \piso.data_r_66_sv2v_reg ;
  assign \piso.data_r [65] = \piso.data_r_65_sv2v_reg ;
  assign \piso.data_r [64] = \piso.data_r_64_sv2v_reg ;
  assign \piso.data_r [63] = \piso.data_r_63_sv2v_reg ;
  assign \piso.data_r [62] = \piso.data_r_62_sv2v_reg ;
  assign \piso.data_r [61] = \piso.data_r_61_sv2v_reg ;
  assign \piso.data_r [60] = \piso.data_r_60_sv2v_reg ;
  assign \piso.data_r [59] = \piso.data_r_59_sv2v_reg ;
  assign \piso.data_r [58] = \piso.data_r_58_sv2v_reg ;
  assign \piso.data_r [57] = \piso.data_r_57_sv2v_reg ;
  assign \piso.data_r [56] = \piso.data_r_56_sv2v_reg ;
  assign \piso.data_r [55] = \piso.data_r_55_sv2v_reg ;
  assign \piso.data_r [54] = \piso.data_r_54_sv2v_reg ;
  assign \piso.data_r [53] = \piso.data_r_53_sv2v_reg ;
  assign \piso.data_r [52] = \piso.data_r_52_sv2v_reg ;
  assign \piso.data_r [51] = \piso.data_r_51_sv2v_reg ;
  assign \piso.data_r [50] = \piso.data_r_50_sv2v_reg ;
  assign \piso.data_r [49] = \piso.data_r_49_sv2v_reg ;
  assign \piso.data_r [48] = \piso.data_r_48_sv2v_reg ;
  assign \piso.data_r [47] = \piso.data_r_47_sv2v_reg ;
  assign \piso.data_r [46] = \piso.data_r_46_sv2v_reg ;
  assign \piso.data_r [45] = \piso.data_r_45_sv2v_reg ;
  assign \piso.data_r [44] = \piso.data_r_44_sv2v_reg ;
  assign \piso.data_r [43] = \piso.data_r_43_sv2v_reg ;
  assign \piso.data_r [42] = \piso.data_r_42_sv2v_reg ;
  assign \piso.data_r [41] = \piso.data_r_41_sv2v_reg ;
  assign \piso.data_r [40] = \piso.data_r_40_sv2v_reg ;
  assign \piso.data_r [39] = \piso.data_r_39_sv2v_reg ;
  assign \piso.data_r [38] = \piso.data_r_38_sv2v_reg ;
  assign \piso.data_r [37] = \piso.data_r_37_sv2v_reg ;
  assign \piso.data_r [36] = \piso.data_r_36_sv2v_reg ;
  assign \piso.data_r [35] = \piso.data_r_35_sv2v_reg ;
  assign \piso.data_r [34] = \piso.data_r_34_sv2v_reg ;
  assign \piso.data_r [33] = \piso.data_r_33_sv2v_reg ;
  assign \piso.data_r [32] = \piso.data_r_32_sv2v_reg ;
  assign \piso.data_r [31] = \piso.data_r_31_sv2v_reg ;
  assign \piso.data_r [30] = \piso.data_r_30_sv2v_reg ;
  assign \piso.data_r [29] = \piso.data_r_29_sv2v_reg ;
  assign \piso.data_r [28] = \piso.data_r_28_sv2v_reg ;
  assign \piso.data_r [27] = \piso.data_r_27_sv2v_reg ;
  assign \piso.data_r [26] = \piso.data_r_26_sv2v_reg ;
  assign \piso.data_r [25] = \piso.data_r_25_sv2v_reg ;
  assign \piso.data_r [24] = \piso.data_r_24_sv2v_reg ;
  assign \piso.data_r [23] = \piso.data_r_23_sv2v_reg ;
  assign \piso.data_r [22] = \piso.data_r_22_sv2v_reg ;
  assign \piso.data_r [21] = \piso.data_r_21_sv2v_reg ;
  assign \piso.data_r [20] = \piso.data_r_20_sv2v_reg ;
  assign \piso.data_r [19] = \piso.data_r_19_sv2v_reg ;
  assign \piso.data_r [18] = \piso.data_r_18_sv2v_reg ;
  assign \piso.data_r [17] = \piso.data_r_17_sv2v_reg ;
  assign \piso.data_r [16] = \piso.data_r_16_sv2v_reg ;
  assign \piso.data_r [15] = \piso.data_r_15_sv2v_reg ;
  assign \piso.data_r [14] = \piso.data_r_14_sv2v_reg ;
  assign \piso.data_r [13] = \piso.data_r_13_sv2v_reg ;
  assign \piso.data_r [12] = \piso.data_r_12_sv2v_reg ;
  assign \piso.data_r [11] = \piso.data_r_11_sv2v_reg ;
  assign \piso.data_r [10] = \piso.data_r_10_sv2v_reg ;
  assign \piso.data_r [9] = \piso.data_r_9_sv2v_reg ;
  assign \piso.data_r [8] = \piso.data_r_8_sv2v_reg ;
  assign \piso.data_r [7] = \piso.data_r_7_sv2v_reg ;
  assign \piso.data_r [6] = \piso.data_r_6_sv2v_reg ;
  assign \piso.data_r [5] = \piso.data_r_5_sv2v_reg ;
  assign \piso.data_r [4] = \piso.data_r_4_sv2v_reg ;
  assign \piso.data_r [3] = \piso.data_r_3_sv2v_reg ;
  assign \piso.data_r [2] = \piso.data_r_2_sv2v_reg ;
  assign \piso.data_r [1] = \piso.data_r_1_sv2v_reg ;
  assign \piso.data_r [0] = \piso.data_r_0_sv2v_reg ;
  assign \piso.shift_ctr_r [4] = \piso.shift_ctr_r_4_sv2v_reg ;
  assign \piso.shift_ctr_r [3] = \piso.shift_ctr_r_3_sv2v_reg ;
  assign \piso.shift_ctr_r [2] = \piso.shift_ctr_r_2_sv2v_reg ;
  assign \piso.shift_ctr_r [1] = \piso.shift_ctr_r_1_sv2v_reg ;
  assign \piso.shift_ctr_r [0] = \piso.shift_ctr_r_0_sv2v_reg ;
  assign data_o[15] = (N54)? \piso.data_r [15] : 
                      (N56)? \piso.data_r [31] : 
                      (N58)? \piso.data_r [47] : 
                      (N60)? \piso.data_r [63] : 
                      (N62)? \piso.data_r [79] : 
                      (N64)? \piso.data_r [95] : 
                      (N66)? \piso.data_r [111] : 
                      (N68)? \piso.data_r [127] : 
                      (N70)? \piso.data_r [143] : 
                      (N72)? \piso.data_r [159] : 
                      (N74)? \piso.data_r [175] : 
                      (N76)? \piso.data_r [191] : 
                      (N78)? \piso.data_r [207] : 
                      (N80)? \piso.data_r [223] : 
                      (N82)? \piso.data_r [239] : 
                      (N84)? \piso.data_r [255] : 
                      (N55)? \piso.data_r [271] : 
                      (N57)? \piso.data_r [287] : 
                      (N59)? \piso.data_r [303] : 
                      (N61)? \piso.data_r [319] : 
                      (N63)? \piso.data_r [335] : 
                      (N65)? \piso.data_r [351] : 
                      (N67)? \piso.data_r [367] : 
                      (N69)? \piso.data_r [383] : 
                      (N71)? \piso.data_r [399] : 
                      (N73)? \piso.data_r [415] : 
                      (N75)? \piso.data_r [431] : 
                      (N77)? \piso.data_r [447] : 
                      (N79)? \piso.data_r [463] : 
                      (N81)? \piso.data_r [479] : 
                      (N83)? \piso.data_r [495] : 
                      (N85)? \piso.data_r [511] : 1'b0;
  assign data_o[14] = (N54)? \piso.data_r [14] : 
                      (N56)? \piso.data_r [30] : 
                      (N58)? \piso.data_r [46] : 
                      (N60)? \piso.data_r [62] : 
                      (N62)? \piso.data_r [78] : 
                      (N64)? \piso.data_r [94] : 
                      (N66)? \piso.data_r [110] : 
                      (N68)? \piso.data_r [126] : 
                      (N70)? \piso.data_r [142] : 
                      (N72)? \piso.data_r [158] : 
                      (N74)? \piso.data_r [174] : 
                      (N76)? \piso.data_r [190] : 
                      (N78)? \piso.data_r [206] : 
                      (N80)? \piso.data_r [222] : 
                      (N82)? \piso.data_r [238] : 
                      (N84)? \piso.data_r [254] : 
                      (N55)? \piso.data_r [270] : 
                      (N57)? \piso.data_r [286] : 
                      (N59)? \piso.data_r [302] : 
                      (N61)? \piso.data_r [318] : 
                      (N63)? \piso.data_r [334] : 
                      (N65)? \piso.data_r [350] : 
                      (N67)? \piso.data_r [366] : 
                      (N69)? \piso.data_r [382] : 
                      (N71)? \piso.data_r [398] : 
                      (N73)? \piso.data_r [414] : 
                      (N75)? \piso.data_r [430] : 
                      (N77)? \piso.data_r [446] : 
                      (N79)? \piso.data_r [462] : 
                      (N81)? \piso.data_r [478] : 
                      (N83)? \piso.data_r [494] : 
                      (N85)? \piso.data_r [510] : 1'b0;
  assign data_o[13] = (N54)? \piso.data_r [13] : 
                      (N56)? \piso.data_r [29] : 
                      (N58)? \piso.data_r [45] : 
                      (N60)? \piso.data_r [61] : 
                      (N62)? \piso.data_r [77] : 
                      (N64)? \piso.data_r [93] : 
                      (N66)? \piso.data_r [109] : 
                      (N68)? \piso.data_r [125] : 
                      (N70)? \piso.data_r [141] : 
                      (N72)? \piso.data_r [157] : 
                      (N74)? \piso.data_r [173] : 
                      (N76)? \piso.data_r [189] : 
                      (N78)? \piso.data_r [205] : 
                      (N80)? \piso.data_r [221] : 
                      (N82)? \piso.data_r [237] : 
                      (N84)? \piso.data_r [253] : 
                      (N55)? \piso.data_r [269] : 
                      (N57)? \piso.data_r [285] : 
                      (N59)? \piso.data_r [301] : 
                      (N61)? \piso.data_r [317] : 
                      (N63)? \piso.data_r [333] : 
                      (N65)? \piso.data_r [349] : 
                      (N67)? \piso.data_r [365] : 
                      (N69)? \piso.data_r [381] : 
                      (N71)? \piso.data_r [397] : 
                      (N73)? \piso.data_r [413] : 
                      (N75)? \piso.data_r [429] : 
                      (N77)? \piso.data_r [445] : 
                      (N79)? \piso.data_r [461] : 
                      (N81)? \piso.data_r [477] : 
                      (N83)? \piso.data_r [493] : 
                      (N85)? \piso.data_r [509] : 1'b0;
  assign data_o[12] = (N54)? \piso.data_r [12] : 
                      (N56)? \piso.data_r [28] : 
                      (N58)? \piso.data_r [44] : 
                      (N60)? \piso.data_r [60] : 
                      (N62)? \piso.data_r [76] : 
                      (N64)? \piso.data_r [92] : 
                      (N66)? \piso.data_r [108] : 
                      (N68)? \piso.data_r [124] : 
                      (N70)? \piso.data_r [140] : 
                      (N72)? \piso.data_r [156] : 
                      (N74)? \piso.data_r [172] : 
                      (N76)? \piso.data_r [188] : 
                      (N78)? \piso.data_r [204] : 
                      (N80)? \piso.data_r [220] : 
                      (N82)? \piso.data_r [236] : 
                      (N84)? \piso.data_r [252] : 
                      (N55)? \piso.data_r [268] : 
                      (N57)? \piso.data_r [284] : 
                      (N59)? \piso.data_r [300] : 
                      (N61)? \piso.data_r [316] : 
                      (N63)? \piso.data_r [332] : 
                      (N65)? \piso.data_r [348] : 
                      (N67)? \piso.data_r [364] : 
                      (N69)? \piso.data_r [380] : 
                      (N71)? \piso.data_r [396] : 
                      (N73)? \piso.data_r [412] : 
                      (N75)? \piso.data_r [428] : 
                      (N77)? \piso.data_r [444] : 
                      (N79)? \piso.data_r [460] : 
                      (N81)? \piso.data_r [476] : 
                      (N83)? \piso.data_r [492] : 
                      (N85)? \piso.data_r [508] : 1'b0;
  assign data_o[11] = (N54)? \piso.data_r [11] : 
                      (N56)? \piso.data_r [27] : 
                      (N58)? \piso.data_r [43] : 
                      (N60)? \piso.data_r [59] : 
                      (N62)? \piso.data_r [75] : 
                      (N64)? \piso.data_r [91] : 
                      (N66)? \piso.data_r [107] : 
                      (N68)? \piso.data_r [123] : 
                      (N70)? \piso.data_r [139] : 
                      (N72)? \piso.data_r [155] : 
                      (N74)? \piso.data_r [171] : 
                      (N76)? \piso.data_r [187] : 
                      (N78)? \piso.data_r [203] : 
                      (N80)? \piso.data_r [219] : 
                      (N82)? \piso.data_r [235] : 
                      (N84)? \piso.data_r [251] : 
                      (N55)? \piso.data_r [267] : 
                      (N57)? \piso.data_r [283] : 
                      (N59)? \piso.data_r [299] : 
                      (N61)? \piso.data_r [315] : 
                      (N63)? \piso.data_r [331] : 
                      (N65)? \piso.data_r [347] : 
                      (N67)? \piso.data_r [363] : 
                      (N69)? \piso.data_r [379] : 
                      (N71)? \piso.data_r [395] : 
                      (N73)? \piso.data_r [411] : 
                      (N75)? \piso.data_r [427] : 
                      (N77)? \piso.data_r [443] : 
                      (N79)? \piso.data_r [459] : 
                      (N81)? \piso.data_r [475] : 
                      (N83)? \piso.data_r [491] : 
                      (N85)? \piso.data_r [507] : 1'b0;
  assign data_o[10] = (N54)? \piso.data_r [10] : 
                      (N56)? \piso.data_r [26] : 
                      (N58)? \piso.data_r [42] : 
                      (N60)? \piso.data_r [58] : 
                      (N62)? \piso.data_r [74] : 
                      (N64)? \piso.data_r [90] : 
                      (N66)? \piso.data_r [106] : 
                      (N68)? \piso.data_r [122] : 
                      (N70)? \piso.data_r [138] : 
                      (N72)? \piso.data_r [154] : 
                      (N74)? \piso.data_r [170] : 
                      (N76)? \piso.data_r [186] : 
                      (N78)? \piso.data_r [202] : 
                      (N80)? \piso.data_r [218] : 
                      (N82)? \piso.data_r [234] : 
                      (N84)? \piso.data_r [250] : 
                      (N55)? \piso.data_r [266] : 
                      (N57)? \piso.data_r [282] : 
                      (N59)? \piso.data_r [298] : 
                      (N61)? \piso.data_r [314] : 
                      (N63)? \piso.data_r [330] : 
                      (N65)? \piso.data_r [346] : 
                      (N67)? \piso.data_r [362] : 
                      (N69)? \piso.data_r [378] : 
                      (N71)? \piso.data_r [394] : 
                      (N73)? \piso.data_r [410] : 
                      (N75)? \piso.data_r [426] : 
                      (N77)? \piso.data_r [442] : 
                      (N79)? \piso.data_r [458] : 
                      (N81)? \piso.data_r [474] : 
                      (N83)? \piso.data_r [490] : 
                      (N85)? \piso.data_r [506] : 1'b0;
  assign data_o[9] = (N54)? \piso.data_r [9] : 
                     (N56)? \piso.data_r [25] : 
                     (N58)? \piso.data_r [41] : 
                     (N60)? \piso.data_r [57] : 
                     (N62)? \piso.data_r [73] : 
                     (N64)? \piso.data_r [89] : 
                     (N66)? \piso.data_r [105] : 
                     (N68)? \piso.data_r [121] : 
                     (N70)? \piso.data_r [137] : 
                     (N72)? \piso.data_r [153] : 
                     (N74)? \piso.data_r [169] : 
                     (N76)? \piso.data_r [185] : 
                     (N78)? \piso.data_r [201] : 
                     (N80)? \piso.data_r [217] : 
                     (N82)? \piso.data_r [233] : 
                     (N84)? \piso.data_r [249] : 
                     (N55)? \piso.data_r [265] : 
                     (N57)? \piso.data_r [281] : 
                     (N59)? \piso.data_r [297] : 
                     (N61)? \piso.data_r [313] : 
                     (N63)? \piso.data_r [329] : 
                     (N65)? \piso.data_r [345] : 
                     (N67)? \piso.data_r [361] : 
                     (N69)? \piso.data_r [377] : 
                     (N71)? \piso.data_r [393] : 
                     (N73)? \piso.data_r [409] : 
                     (N75)? \piso.data_r [425] : 
                     (N77)? \piso.data_r [441] : 
                     (N79)? \piso.data_r [457] : 
                     (N81)? \piso.data_r [473] : 
                     (N83)? \piso.data_r [489] : 
                     (N85)? \piso.data_r [505] : 1'b0;
  assign data_o[8] = (N54)? \piso.data_r [8] : 
                     (N56)? \piso.data_r [24] : 
                     (N58)? \piso.data_r [40] : 
                     (N60)? \piso.data_r [56] : 
                     (N62)? \piso.data_r [72] : 
                     (N64)? \piso.data_r [88] : 
                     (N66)? \piso.data_r [104] : 
                     (N68)? \piso.data_r [120] : 
                     (N70)? \piso.data_r [136] : 
                     (N72)? \piso.data_r [152] : 
                     (N74)? \piso.data_r [168] : 
                     (N76)? \piso.data_r [184] : 
                     (N78)? \piso.data_r [200] : 
                     (N80)? \piso.data_r [216] : 
                     (N82)? \piso.data_r [232] : 
                     (N84)? \piso.data_r [248] : 
                     (N55)? \piso.data_r [264] : 
                     (N57)? \piso.data_r [280] : 
                     (N59)? \piso.data_r [296] : 
                     (N61)? \piso.data_r [312] : 
                     (N63)? \piso.data_r [328] : 
                     (N65)? \piso.data_r [344] : 
                     (N67)? \piso.data_r [360] : 
                     (N69)? \piso.data_r [376] : 
                     (N71)? \piso.data_r [392] : 
                     (N73)? \piso.data_r [408] : 
                     (N75)? \piso.data_r [424] : 
                     (N77)? \piso.data_r [440] : 
                     (N79)? \piso.data_r [456] : 
                     (N81)? \piso.data_r [472] : 
                     (N83)? \piso.data_r [488] : 
                     (N85)? \piso.data_r [504] : 1'b0;
  assign data_o[7] = (N54)? \piso.data_r [7] : 
                     (N56)? \piso.data_r [23] : 
                     (N58)? \piso.data_r [39] : 
                     (N60)? \piso.data_r [55] : 
                     (N62)? \piso.data_r [71] : 
                     (N64)? \piso.data_r [87] : 
                     (N66)? \piso.data_r [103] : 
                     (N68)? \piso.data_r [119] : 
                     (N70)? \piso.data_r [135] : 
                     (N72)? \piso.data_r [151] : 
                     (N74)? \piso.data_r [167] : 
                     (N76)? \piso.data_r [183] : 
                     (N78)? \piso.data_r [199] : 
                     (N80)? \piso.data_r [215] : 
                     (N82)? \piso.data_r [231] : 
                     (N84)? \piso.data_r [247] : 
                     (N55)? \piso.data_r [263] : 
                     (N57)? \piso.data_r [279] : 
                     (N59)? \piso.data_r [295] : 
                     (N61)? \piso.data_r [311] : 
                     (N63)? \piso.data_r [327] : 
                     (N65)? \piso.data_r [343] : 
                     (N67)? \piso.data_r [359] : 
                     (N69)? \piso.data_r [375] : 
                     (N71)? \piso.data_r [391] : 
                     (N73)? \piso.data_r [407] : 
                     (N75)? \piso.data_r [423] : 
                     (N77)? \piso.data_r [439] : 
                     (N79)? \piso.data_r [455] : 
                     (N81)? \piso.data_r [471] : 
                     (N83)? \piso.data_r [487] : 
                     (N85)? \piso.data_r [503] : 1'b0;
  assign data_o[6] = (N54)? \piso.data_r [6] : 
                     (N56)? \piso.data_r [22] : 
                     (N58)? \piso.data_r [38] : 
                     (N60)? \piso.data_r [54] : 
                     (N62)? \piso.data_r [70] : 
                     (N64)? \piso.data_r [86] : 
                     (N66)? \piso.data_r [102] : 
                     (N68)? \piso.data_r [118] : 
                     (N70)? \piso.data_r [134] : 
                     (N72)? \piso.data_r [150] : 
                     (N74)? \piso.data_r [166] : 
                     (N76)? \piso.data_r [182] : 
                     (N78)? \piso.data_r [198] : 
                     (N80)? \piso.data_r [214] : 
                     (N82)? \piso.data_r [230] : 
                     (N84)? \piso.data_r [246] : 
                     (N55)? \piso.data_r [262] : 
                     (N57)? \piso.data_r [278] : 
                     (N59)? \piso.data_r [294] : 
                     (N61)? \piso.data_r [310] : 
                     (N63)? \piso.data_r [326] : 
                     (N65)? \piso.data_r [342] : 
                     (N67)? \piso.data_r [358] : 
                     (N69)? \piso.data_r [374] : 
                     (N71)? \piso.data_r [390] : 
                     (N73)? \piso.data_r [406] : 
                     (N75)? \piso.data_r [422] : 
                     (N77)? \piso.data_r [438] : 
                     (N79)? \piso.data_r [454] : 
                     (N81)? \piso.data_r [470] : 
                     (N83)? \piso.data_r [486] : 
                     (N85)? \piso.data_r [502] : 1'b0;
  assign data_o[5] = (N54)? \piso.data_r [5] : 
                     (N56)? \piso.data_r [21] : 
                     (N58)? \piso.data_r [37] : 
                     (N60)? \piso.data_r [53] : 
                     (N62)? \piso.data_r [69] : 
                     (N64)? \piso.data_r [85] : 
                     (N66)? \piso.data_r [101] : 
                     (N68)? \piso.data_r [117] : 
                     (N70)? \piso.data_r [133] : 
                     (N72)? \piso.data_r [149] : 
                     (N74)? \piso.data_r [165] : 
                     (N76)? \piso.data_r [181] : 
                     (N78)? \piso.data_r [197] : 
                     (N80)? \piso.data_r [213] : 
                     (N82)? \piso.data_r [229] : 
                     (N84)? \piso.data_r [245] : 
                     (N55)? \piso.data_r [261] : 
                     (N57)? \piso.data_r [277] : 
                     (N59)? \piso.data_r [293] : 
                     (N61)? \piso.data_r [309] : 
                     (N63)? \piso.data_r [325] : 
                     (N65)? \piso.data_r [341] : 
                     (N67)? \piso.data_r [357] : 
                     (N69)? \piso.data_r [373] : 
                     (N71)? \piso.data_r [389] : 
                     (N73)? \piso.data_r [405] : 
                     (N75)? \piso.data_r [421] : 
                     (N77)? \piso.data_r [437] : 
                     (N79)? \piso.data_r [453] : 
                     (N81)? \piso.data_r [469] : 
                     (N83)? \piso.data_r [485] : 
                     (N85)? \piso.data_r [501] : 1'b0;
  assign data_o[4] = (N54)? \piso.data_r [4] : 
                     (N56)? \piso.data_r [20] : 
                     (N58)? \piso.data_r [36] : 
                     (N60)? \piso.data_r [52] : 
                     (N62)? \piso.data_r [68] : 
                     (N64)? \piso.data_r [84] : 
                     (N66)? \piso.data_r [100] : 
                     (N68)? \piso.data_r [116] : 
                     (N70)? \piso.data_r [132] : 
                     (N72)? \piso.data_r [148] : 
                     (N74)? \piso.data_r [164] : 
                     (N76)? \piso.data_r [180] : 
                     (N78)? \piso.data_r [196] : 
                     (N80)? \piso.data_r [212] : 
                     (N82)? \piso.data_r [228] : 
                     (N84)? \piso.data_r [244] : 
                     (N55)? \piso.data_r [260] : 
                     (N57)? \piso.data_r [276] : 
                     (N59)? \piso.data_r [292] : 
                     (N61)? \piso.data_r [308] : 
                     (N63)? \piso.data_r [324] : 
                     (N65)? \piso.data_r [340] : 
                     (N67)? \piso.data_r [356] : 
                     (N69)? \piso.data_r [372] : 
                     (N71)? \piso.data_r [388] : 
                     (N73)? \piso.data_r [404] : 
                     (N75)? \piso.data_r [420] : 
                     (N77)? \piso.data_r [436] : 
                     (N79)? \piso.data_r [452] : 
                     (N81)? \piso.data_r [468] : 
                     (N83)? \piso.data_r [484] : 
                     (N85)? \piso.data_r [500] : 1'b0;
  assign data_o[3] = (N54)? \piso.data_r [3] : 
                     (N56)? \piso.data_r [19] : 
                     (N58)? \piso.data_r [35] : 
                     (N60)? \piso.data_r [51] : 
                     (N62)? \piso.data_r [67] : 
                     (N64)? \piso.data_r [83] : 
                     (N66)? \piso.data_r [99] : 
                     (N68)? \piso.data_r [115] : 
                     (N70)? \piso.data_r [131] : 
                     (N72)? \piso.data_r [147] : 
                     (N74)? \piso.data_r [163] : 
                     (N76)? \piso.data_r [179] : 
                     (N78)? \piso.data_r [195] : 
                     (N80)? \piso.data_r [211] : 
                     (N82)? \piso.data_r [227] : 
                     (N84)? \piso.data_r [243] : 
                     (N55)? \piso.data_r [259] : 
                     (N57)? \piso.data_r [275] : 
                     (N59)? \piso.data_r [291] : 
                     (N61)? \piso.data_r [307] : 
                     (N63)? \piso.data_r [323] : 
                     (N65)? \piso.data_r [339] : 
                     (N67)? \piso.data_r [355] : 
                     (N69)? \piso.data_r [371] : 
                     (N71)? \piso.data_r [387] : 
                     (N73)? \piso.data_r [403] : 
                     (N75)? \piso.data_r [419] : 
                     (N77)? \piso.data_r [435] : 
                     (N79)? \piso.data_r [451] : 
                     (N81)? \piso.data_r [467] : 
                     (N83)? \piso.data_r [483] : 
                     (N85)? \piso.data_r [499] : 1'b0;
  assign data_o[2] = (N54)? \piso.data_r [2] : 
                     (N56)? \piso.data_r [18] : 
                     (N58)? \piso.data_r [34] : 
                     (N60)? \piso.data_r [50] : 
                     (N62)? \piso.data_r [66] : 
                     (N64)? \piso.data_r [82] : 
                     (N66)? \piso.data_r [98] : 
                     (N68)? \piso.data_r [114] : 
                     (N70)? \piso.data_r [130] : 
                     (N72)? \piso.data_r [146] : 
                     (N74)? \piso.data_r [162] : 
                     (N76)? \piso.data_r [178] : 
                     (N78)? \piso.data_r [194] : 
                     (N80)? \piso.data_r [210] : 
                     (N82)? \piso.data_r [226] : 
                     (N84)? \piso.data_r [242] : 
                     (N55)? \piso.data_r [258] : 
                     (N57)? \piso.data_r [274] : 
                     (N59)? \piso.data_r [290] : 
                     (N61)? \piso.data_r [306] : 
                     (N63)? \piso.data_r [322] : 
                     (N65)? \piso.data_r [338] : 
                     (N67)? \piso.data_r [354] : 
                     (N69)? \piso.data_r [370] : 
                     (N71)? \piso.data_r [386] : 
                     (N73)? \piso.data_r [402] : 
                     (N75)? \piso.data_r [418] : 
                     (N77)? \piso.data_r [434] : 
                     (N79)? \piso.data_r [450] : 
                     (N81)? \piso.data_r [466] : 
                     (N83)? \piso.data_r [482] : 
                     (N85)? \piso.data_r [498] : 1'b0;
  assign data_o[1] = (N54)? \piso.data_r [1] : 
                     (N56)? \piso.data_r [17] : 
                     (N58)? \piso.data_r [33] : 
                     (N60)? \piso.data_r [49] : 
                     (N62)? \piso.data_r [65] : 
                     (N64)? \piso.data_r [81] : 
                     (N66)? \piso.data_r [97] : 
                     (N68)? \piso.data_r [113] : 
                     (N70)? \piso.data_r [129] : 
                     (N72)? \piso.data_r [145] : 
                     (N74)? \piso.data_r [161] : 
                     (N76)? \piso.data_r [177] : 
                     (N78)? \piso.data_r [193] : 
                     (N80)? \piso.data_r [209] : 
                     (N82)? \piso.data_r [225] : 
                     (N84)? \piso.data_r [241] : 
                     (N55)? \piso.data_r [257] : 
                     (N57)? \piso.data_r [273] : 
                     (N59)? \piso.data_r [289] : 
                     (N61)? \piso.data_r [305] : 
                     (N63)? \piso.data_r [321] : 
                     (N65)? \piso.data_r [337] : 
                     (N67)? \piso.data_r [353] : 
                     (N69)? \piso.data_r [369] : 
                     (N71)? \piso.data_r [385] : 
                     (N73)? \piso.data_r [401] : 
                     (N75)? \piso.data_r [417] : 
                     (N77)? \piso.data_r [433] : 
                     (N79)? \piso.data_r [449] : 
                     (N81)? \piso.data_r [465] : 
                     (N83)? \piso.data_r [481] : 
                     (N85)? \piso.data_r [497] : 1'b0;
  assign data_o[0] = (N54)? \piso.data_r [0] : 
                     (N56)? \piso.data_r [16] : 
                     (N58)? \piso.data_r [32] : 
                     (N60)? \piso.data_r [48] : 
                     (N62)? \piso.data_r [64] : 
                     (N64)? \piso.data_r [80] : 
                     (N66)? \piso.data_r [96] : 
                     (N68)? \piso.data_r [112] : 
                     (N70)? \piso.data_r [128] : 
                     (N72)? \piso.data_r [144] : 
                     (N74)? \piso.data_r [160] : 
                     (N76)? \piso.data_r [176] : 
                     (N78)? \piso.data_r [192] : 
                     (N80)? \piso.data_r [208] : 
                     (N82)? \piso.data_r [224] : 
                     (N84)? \piso.data_r [240] : 
                     (N55)? \piso.data_r [256] : 
                     (N57)? \piso.data_r [272] : 
                     (N59)? \piso.data_r [288] : 
                     (N61)? \piso.data_r [304] : 
                     (N63)? \piso.data_r [320] : 
                     (N65)? \piso.data_r [336] : 
                     (N67)? \piso.data_r [352] : 
                     (N69)? \piso.data_r [368] : 
                     (N71)? \piso.data_r [384] : 
                     (N73)? \piso.data_r [400] : 
                     (N75)? \piso.data_r [416] : 
                     (N77)? \piso.data_r [432] : 
                     (N79)? \piso.data_r [448] : 
                     (N81)? \piso.data_r [464] : 
                     (N83)? \piso.data_r [480] : 
                     (N85)? \piso.data_r [496] : 1'b0;
  assign N88 = ~valid_o;
  assign N89 = \piso.shift_ctr_r [3] & \piso.shift_ctr_r [4];
  assign N90 = \piso.shift_ctr_r [2] & N89;
  assign N91 = \piso.shift_ctr_r [1] & N90;
  assign N92 = \piso.shift_ctr_r [0] & N91;
  assign { N20, N19, N18, N17, N16 } = \piso.shift_ctr_r  + 1'b1;
  assign \piso.state_n [0] = (N0)? 1'b1 : 
                             (N5)? 1'b0 : 1'b0;
  assign N0 = N2;
  assign { N13, N12, N11, N10, N9 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N8)? { N20, N19, N18, N17, N16 } : 1'b0;
  assign N1 = N7;
  assign \piso.done_tx_n  = N93 & yumi_i;
  assign N93 = valid_o & N92;
  assign ready_o = N88 | \piso.done_tx_n ;
  assign N2 = ready_o & valid_i;
  assign N3 = \piso.done_tx_n  | N2;
  assign N4 = ~N2;
  assign N5 = \piso.done_tx_n  & N4;
  assign N6 = ready_o & valid_i;
  assign N7 = ready_o & valid_i;
  assign N8 = ~N7;
  assign N14 = N94 & N95;
  assign N94 = valid_o & yumi_i;
  assign N95 = ~\piso.done_tx_n ;
  assign N15 = ~N14;
  assign N21 = ~\piso.shift_ctr_r [0];
  assign N22 = ~\piso.shift_ctr_r [1];
  assign N23 = N21 & N22;
  assign N24 = N21 & \piso.shift_ctr_r [1];
  assign N25 = \piso.shift_ctr_r [0] & N22;
  assign N26 = \piso.shift_ctr_r [0] & \piso.shift_ctr_r [1];
  assign N27 = ~\piso.shift_ctr_r [2];
  assign N28 = N23 & N27;
  assign N29 = N23 & \piso.shift_ctr_r [2];
  assign N30 = N25 & N27;
  assign N31 = N25 & \piso.shift_ctr_r [2];
  assign N32 = N24 & N27;
  assign N33 = N24 & \piso.shift_ctr_r [2];
  assign N34 = N26 & N27;
  assign N35 = N26 & \piso.shift_ctr_r [2];
  assign N36 = ~\piso.shift_ctr_r [3];
  assign N37 = N28 & N36;
  assign N38 = N28 & \piso.shift_ctr_r [3];
  assign N39 = N30 & N36;
  assign N40 = N30 & \piso.shift_ctr_r [3];
  assign N41 = N32 & N36;
  assign N42 = N32 & \piso.shift_ctr_r [3];
  assign N43 = N34 & N36;
  assign N44 = N34 & \piso.shift_ctr_r [3];
  assign N45 = N29 & N36;
  assign N46 = N29 & \piso.shift_ctr_r [3];
  assign N47 = N31 & N36;
  assign N48 = N31 & \piso.shift_ctr_r [3];
  assign N49 = N33 & N36;
  assign N50 = N33 & \piso.shift_ctr_r [3];
  assign N51 = N35 & N36;
  assign N52 = N35 & \piso.shift_ctr_r [3];
  assign N53 = ~\piso.shift_ctr_r [4];
  assign N54 = N37 & N53;
  assign N55 = N37 & \piso.shift_ctr_r [4];
  assign N56 = N39 & N53;
  assign N57 = N39 & \piso.shift_ctr_r [4];
  assign N58 = N41 & N53;
  assign N59 = N41 & \piso.shift_ctr_r [4];
  assign N60 = N43 & N53;
  assign N61 = N43 & \piso.shift_ctr_r [4];
  assign N62 = N45 & N53;
  assign N63 = N45 & \piso.shift_ctr_r [4];
  assign N64 = N47 & N53;
  assign N65 = N47 & \piso.shift_ctr_r [4];
  assign N66 = N49 & N53;
  assign N67 = N49 & \piso.shift_ctr_r [4];
  assign N68 = N51 & N53;
  assign N69 = N51 & \piso.shift_ctr_r [4];
  assign N70 = N38 & N53;
  assign N71 = N38 & \piso.shift_ctr_r [4];
  assign N72 = N40 & N53;
  assign N73 = N40 & \piso.shift_ctr_r [4];
  assign N74 = N42 & N53;
  assign N75 = N42 & \piso.shift_ctr_r [4];
  assign N76 = N44 & N53;
  assign N77 = N44 & \piso.shift_ctr_r [4];
  assign N78 = N46 & N53;
  assign N79 = N46 & \piso.shift_ctr_r [4];
  assign N80 = N48 & N53;
  assign N81 = N48 & \piso.shift_ctr_r [4];
  assign N82 = N50 & N53;
  assign N83 = N50 & \piso.shift_ctr_r [4];
  assign N84 = N52 & N53;
  assign N85 = N52 & \piso.shift_ctr_r [4];
  assign N86 = N15 & N8;
  assign N87 = ~N86;

  always @(posedge clk_i) begin
    if(reset_i) begin
      valid_o_sv2v_reg <= 1'b0;
    end else if(N3) begin
      valid_o_sv2v_reg <= \piso.state_n [0];
    end 
    if(reset_i) begin
      \piso.data_r_511_sv2v_reg  <= 1'b0;
      \piso.data_r_510_sv2v_reg  <= 1'b0;
      \piso.data_r_509_sv2v_reg  <= 1'b0;
      \piso.data_r_508_sv2v_reg  <= 1'b0;
      \piso.data_r_507_sv2v_reg  <= 1'b0;
      \piso.data_r_506_sv2v_reg  <= 1'b0;
      \piso.data_r_505_sv2v_reg  <= 1'b0;
      \piso.data_r_504_sv2v_reg  <= 1'b0;
      \piso.data_r_503_sv2v_reg  <= 1'b0;
      \piso.data_r_502_sv2v_reg  <= 1'b0;
      \piso.data_r_501_sv2v_reg  <= 1'b0;
      \piso.data_r_500_sv2v_reg  <= 1'b0;
      \piso.data_r_499_sv2v_reg  <= 1'b0;
      \piso.data_r_498_sv2v_reg  <= 1'b0;
      \piso.data_r_497_sv2v_reg  <= 1'b0;
      \piso.data_r_496_sv2v_reg  <= 1'b0;
      \piso.data_r_495_sv2v_reg  <= 1'b0;
      \piso.data_r_494_sv2v_reg  <= 1'b0;
      \piso.data_r_493_sv2v_reg  <= 1'b0;
      \piso.data_r_492_sv2v_reg  <= 1'b0;
      \piso.data_r_491_sv2v_reg  <= 1'b0;
      \piso.data_r_490_sv2v_reg  <= 1'b0;
      \piso.data_r_489_sv2v_reg  <= 1'b0;
      \piso.data_r_488_sv2v_reg  <= 1'b0;
      \piso.data_r_487_sv2v_reg  <= 1'b0;
      \piso.data_r_486_sv2v_reg  <= 1'b0;
      \piso.data_r_485_sv2v_reg  <= 1'b0;
      \piso.data_r_484_sv2v_reg  <= 1'b0;
      \piso.data_r_483_sv2v_reg  <= 1'b0;
      \piso.data_r_482_sv2v_reg  <= 1'b0;
      \piso.data_r_481_sv2v_reg  <= 1'b0;
      \piso.data_r_480_sv2v_reg  <= 1'b0;
      \piso.data_r_479_sv2v_reg  <= 1'b0;
      \piso.data_r_478_sv2v_reg  <= 1'b0;
      \piso.data_r_477_sv2v_reg  <= 1'b0;
      \piso.data_r_476_sv2v_reg  <= 1'b0;
      \piso.data_r_475_sv2v_reg  <= 1'b0;
      \piso.data_r_474_sv2v_reg  <= 1'b0;
      \piso.data_r_473_sv2v_reg  <= 1'b0;
      \piso.data_r_472_sv2v_reg  <= 1'b0;
      \piso.data_r_471_sv2v_reg  <= 1'b0;
      \piso.data_r_470_sv2v_reg  <= 1'b0;
      \piso.data_r_469_sv2v_reg  <= 1'b0;
      \piso.data_r_468_sv2v_reg  <= 1'b0;
      \piso.data_r_467_sv2v_reg  <= 1'b0;
      \piso.data_r_466_sv2v_reg  <= 1'b0;
      \piso.data_r_465_sv2v_reg  <= 1'b0;
      \piso.data_r_464_sv2v_reg  <= 1'b0;
      \piso.data_r_463_sv2v_reg  <= 1'b0;
      \piso.data_r_462_sv2v_reg  <= 1'b0;
      \piso.data_r_461_sv2v_reg  <= 1'b0;
      \piso.data_r_460_sv2v_reg  <= 1'b0;
      \piso.data_r_459_sv2v_reg  <= 1'b0;
      \piso.data_r_458_sv2v_reg  <= 1'b0;
      \piso.data_r_457_sv2v_reg  <= 1'b0;
      \piso.data_r_456_sv2v_reg  <= 1'b0;
      \piso.data_r_455_sv2v_reg  <= 1'b0;
      \piso.data_r_454_sv2v_reg  <= 1'b0;
      \piso.data_r_453_sv2v_reg  <= 1'b0;
      \piso.data_r_452_sv2v_reg  <= 1'b0;
      \piso.data_r_451_sv2v_reg  <= 1'b0;
      \piso.data_r_450_sv2v_reg  <= 1'b0;
      \piso.data_r_449_sv2v_reg  <= 1'b0;
      \piso.data_r_448_sv2v_reg  <= 1'b0;
      \piso.data_r_447_sv2v_reg  <= 1'b0;
      \piso.data_r_446_sv2v_reg  <= 1'b0;
      \piso.data_r_445_sv2v_reg  <= 1'b0;
      \piso.data_r_444_sv2v_reg  <= 1'b0;
      \piso.data_r_443_sv2v_reg  <= 1'b0;
      \piso.data_r_442_sv2v_reg  <= 1'b0;
      \piso.data_r_441_sv2v_reg  <= 1'b0;
      \piso.data_r_440_sv2v_reg  <= 1'b0;
      \piso.data_r_439_sv2v_reg  <= 1'b0;
      \piso.data_r_438_sv2v_reg  <= 1'b0;
      \piso.data_r_437_sv2v_reg  <= 1'b0;
      \piso.data_r_436_sv2v_reg  <= 1'b0;
      \piso.data_r_435_sv2v_reg  <= 1'b0;
      \piso.data_r_434_sv2v_reg  <= 1'b0;
      \piso.data_r_433_sv2v_reg  <= 1'b0;
      \piso.data_r_432_sv2v_reg  <= 1'b0;
      \piso.data_r_431_sv2v_reg  <= 1'b0;
      \piso.data_r_430_sv2v_reg  <= 1'b0;
      \piso.data_r_429_sv2v_reg  <= 1'b0;
      \piso.data_r_428_sv2v_reg  <= 1'b0;
      \piso.data_r_427_sv2v_reg  <= 1'b0;
      \piso.data_r_426_sv2v_reg  <= 1'b0;
      \piso.data_r_425_sv2v_reg  <= 1'b0;
      \piso.data_r_424_sv2v_reg  <= 1'b0;
      \piso.data_r_423_sv2v_reg  <= 1'b0;
      \piso.data_r_422_sv2v_reg  <= 1'b0;
      \piso.data_r_421_sv2v_reg  <= 1'b0;
      \piso.data_r_420_sv2v_reg  <= 1'b0;
      \piso.data_r_419_sv2v_reg  <= 1'b0;
      \piso.data_r_418_sv2v_reg  <= 1'b0;
      \piso.data_r_417_sv2v_reg  <= 1'b0;
      \piso.data_r_416_sv2v_reg  <= 1'b0;
      \piso.data_r_415_sv2v_reg  <= 1'b0;
      \piso.data_r_414_sv2v_reg  <= 1'b0;
      \piso.data_r_413_sv2v_reg  <= 1'b0;
      \piso.data_r_412_sv2v_reg  <= 1'b0;
      \piso.data_r_411_sv2v_reg  <= 1'b0;
      \piso.data_r_410_sv2v_reg  <= 1'b0;
      \piso.data_r_409_sv2v_reg  <= 1'b0;
      \piso.data_r_408_sv2v_reg  <= 1'b0;
      \piso.data_r_407_sv2v_reg  <= 1'b0;
      \piso.data_r_406_sv2v_reg  <= 1'b0;
      \piso.data_r_405_sv2v_reg  <= 1'b0;
      \piso.data_r_404_sv2v_reg  <= 1'b0;
      \piso.data_r_403_sv2v_reg  <= 1'b0;
      \piso.data_r_402_sv2v_reg  <= 1'b0;
      \piso.data_r_401_sv2v_reg  <= 1'b0;
      \piso.data_r_400_sv2v_reg  <= 1'b0;
      \piso.data_r_399_sv2v_reg  <= 1'b0;
      \piso.data_r_398_sv2v_reg  <= 1'b0;
      \piso.data_r_397_sv2v_reg  <= 1'b0;
      \piso.data_r_396_sv2v_reg  <= 1'b0;
      \piso.data_r_395_sv2v_reg  <= 1'b0;
      \piso.data_r_394_sv2v_reg  <= 1'b0;
      \piso.data_r_393_sv2v_reg  <= 1'b0;
      \piso.data_r_392_sv2v_reg  <= 1'b0;
      \piso.data_r_391_sv2v_reg  <= 1'b0;
      \piso.data_r_390_sv2v_reg  <= 1'b0;
      \piso.data_r_389_sv2v_reg  <= 1'b0;
      \piso.data_r_388_sv2v_reg  <= 1'b0;
      \piso.data_r_387_sv2v_reg  <= 1'b0;
      \piso.data_r_386_sv2v_reg  <= 1'b0;
      \piso.data_r_385_sv2v_reg  <= 1'b0;
      \piso.data_r_384_sv2v_reg  <= 1'b0;
      \piso.data_r_383_sv2v_reg  <= 1'b0;
      \piso.data_r_382_sv2v_reg  <= 1'b0;
      \piso.data_r_381_sv2v_reg  <= 1'b0;
      \piso.data_r_380_sv2v_reg  <= 1'b0;
      \piso.data_r_379_sv2v_reg  <= 1'b0;
      \piso.data_r_378_sv2v_reg  <= 1'b0;
      \piso.data_r_377_sv2v_reg  <= 1'b0;
      \piso.data_r_376_sv2v_reg  <= 1'b0;
      \piso.data_r_375_sv2v_reg  <= 1'b0;
      \piso.data_r_374_sv2v_reg  <= 1'b0;
      \piso.data_r_373_sv2v_reg  <= 1'b0;
      \piso.data_r_372_sv2v_reg  <= 1'b0;
      \piso.data_r_371_sv2v_reg  <= 1'b0;
      \piso.data_r_370_sv2v_reg  <= 1'b0;
      \piso.data_r_369_sv2v_reg  <= 1'b0;
      \piso.data_r_368_sv2v_reg  <= 1'b0;
      \piso.data_r_367_sv2v_reg  <= 1'b0;
      \piso.data_r_366_sv2v_reg  <= 1'b0;
      \piso.data_r_365_sv2v_reg  <= 1'b0;
      \piso.data_r_364_sv2v_reg  <= 1'b0;
      \piso.data_r_363_sv2v_reg  <= 1'b0;
      \piso.data_r_362_sv2v_reg  <= 1'b0;
      \piso.data_r_361_sv2v_reg  <= 1'b0;
      \piso.data_r_360_sv2v_reg  <= 1'b0;
      \piso.data_r_359_sv2v_reg  <= 1'b0;
      \piso.data_r_358_sv2v_reg  <= 1'b0;
      \piso.data_r_357_sv2v_reg  <= 1'b0;
      \piso.data_r_356_sv2v_reg  <= 1'b0;
      \piso.data_r_355_sv2v_reg  <= 1'b0;
      \piso.data_r_354_sv2v_reg  <= 1'b0;
      \piso.data_r_353_sv2v_reg  <= 1'b0;
      \piso.data_r_352_sv2v_reg  <= 1'b0;
      \piso.data_r_351_sv2v_reg  <= 1'b0;
      \piso.data_r_350_sv2v_reg  <= 1'b0;
      \piso.data_r_349_sv2v_reg  <= 1'b0;
      \piso.data_r_348_sv2v_reg  <= 1'b0;
      \piso.data_r_347_sv2v_reg  <= 1'b0;
      \piso.data_r_346_sv2v_reg  <= 1'b0;
      \piso.data_r_345_sv2v_reg  <= 1'b0;
      \piso.data_r_344_sv2v_reg  <= 1'b0;
      \piso.data_r_343_sv2v_reg  <= 1'b0;
      \piso.data_r_342_sv2v_reg  <= 1'b0;
      \piso.data_r_341_sv2v_reg  <= 1'b0;
      \piso.data_r_340_sv2v_reg  <= 1'b0;
      \piso.data_r_339_sv2v_reg  <= 1'b0;
      \piso.data_r_338_sv2v_reg  <= 1'b0;
      \piso.data_r_337_sv2v_reg  <= 1'b0;
      \piso.data_r_336_sv2v_reg  <= 1'b0;
      \piso.data_r_335_sv2v_reg  <= 1'b0;
      \piso.data_r_334_sv2v_reg  <= 1'b0;
      \piso.data_r_333_sv2v_reg  <= 1'b0;
      \piso.data_r_332_sv2v_reg  <= 1'b0;
      \piso.data_r_331_sv2v_reg  <= 1'b0;
      \piso.data_r_330_sv2v_reg  <= 1'b0;
      \piso.data_r_329_sv2v_reg  <= 1'b0;
      \piso.data_r_328_sv2v_reg  <= 1'b0;
      \piso.data_r_327_sv2v_reg  <= 1'b0;
      \piso.data_r_326_sv2v_reg  <= 1'b0;
      \piso.data_r_325_sv2v_reg  <= 1'b0;
      \piso.data_r_324_sv2v_reg  <= 1'b0;
      \piso.data_r_323_sv2v_reg  <= 1'b0;
      \piso.data_r_322_sv2v_reg  <= 1'b0;
      \piso.data_r_321_sv2v_reg  <= 1'b0;
      \piso.data_r_320_sv2v_reg  <= 1'b0;
      \piso.data_r_319_sv2v_reg  <= 1'b0;
      \piso.data_r_318_sv2v_reg  <= 1'b0;
      \piso.data_r_317_sv2v_reg  <= 1'b0;
      \piso.data_r_316_sv2v_reg  <= 1'b0;
      \piso.data_r_315_sv2v_reg  <= 1'b0;
      \piso.data_r_314_sv2v_reg  <= 1'b0;
      \piso.data_r_313_sv2v_reg  <= 1'b0;
      \piso.data_r_312_sv2v_reg  <= 1'b0;
      \piso.data_r_311_sv2v_reg  <= 1'b0;
      \piso.data_r_310_sv2v_reg  <= 1'b0;
      \piso.data_r_309_sv2v_reg  <= 1'b0;
      \piso.data_r_308_sv2v_reg  <= 1'b0;
      \piso.data_r_307_sv2v_reg  <= 1'b0;
      \piso.data_r_306_sv2v_reg  <= 1'b0;
      \piso.data_r_305_sv2v_reg  <= 1'b0;
      \piso.data_r_304_sv2v_reg  <= 1'b0;
      \piso.data_r_303_sv2v_reg  <= 1'b0;
      \piso.data_r_302_sv2v_reg  <= 1'b0;
      \piso.data_r_301_sv2v_reg  <= 1'b0;
      \piso.data_r_300_sv2v_reg  <= 1'b0;
      \piso.data_r_299_sv2v_reg  <= 1'b0;
      \piso.data_r_298_sv2v_reg  <= 1'b0;
      \piso.data_r_297_sv2v_reg  <= 1'b0;
      \piso.data_r_296_sv2v_reg  <= 1'b0;
      \piso.data_r_295_sv2v_reg  <= 1'b0;
      \piso.data_r_294_sv2v_reg  <= 1'b0;
      \piso.data_r_293_sv2v_reg  <= 1'b0;
      \piso.data_r_292_sv2v_reg  <= 1'b0;
      \piso.data_r_291_sv2v_reg  <= 1'b0;
      \piso.data_r_290_sv2v_reg  <= 1'b0;
      \piso.data_r_289_sv2v_reg  <= 1'b0;
      \piso.data_r_288_sv2v_reg  <= 1'b0;
      \piso.data_r_287_sv2v_reg  <= 1'b0;
      \piso.data_r_286_sv2v_reg  <= 1'b0;
      \piso.data_r_285_sv2v_reg  <= 1'b0;
      \piso.data_r_284_sv2v_reg  <= 1'b0;
      \piso.data_r_283_sv2v_reg  <= 1'b0;
      \piso.data_r_282_sv2v_reg  <= 1'b0;
      \piso.data_r_281_sv2v_reg  <= 1'b0;
      \piso.data_r_280_sv2v_reg  <= 1'b0;
      \piso.data_r_279_sv2v_reg  <= 1'b0;
      \piso.data_r_278_sv2v_reg  <= 1'b0;
      \piso.data_r_277_sv2v_reg  <= 1'b0;
      \piso.data_r_276_sv2v_reg  <= 1'b0;
      \piso.data_r_275_sv2v_reg  <= 1'b0;
      \piso.data_r_274_sv2v_reg  <= 1'b0;
      \piso.data_r_273_sv2v_reg  <= 1'b0;
      \piso.data_r_272_sv2v_reg  <= 1'b0;
      \piso.data_r_271_sv2v_reg  <= 1'b0;
      \piso.data_r_270_sv2v_reg  <= 1'b0;
      \piso.data_r_269_sv2v_reg  <= 1'b0;
      \piso.data_r_268_sv2v_reg  <= 1'b0;
      \piso.data_r_267_sv2v_reg  <= 1'b0;
      \piso.data_r_266_sv2v_reg  <= 1'b0;
      \piso.data_r_265_sv2v_reg  <= 1'b0;
      \piso.data_r_264_sv2v_reg  <= 1'b0;
      \piso.data_r_263_sv2v_reg  <= 1'b0;
      \piso.data_r_262_sv2v_reg  <= 1'b0;
      \piso.data_r_261_sv2v_reg  <= 1'b0;
      \piso.data_r_260_sv2v_reg  <= 1'b0;
      \piso.data_r_259_sv2v_reg  <= 1'b0;
      \piso.data_r_258_sv2v_reg  <= 1'b0;
      \piso.data_r_257_sv2v_reg  <= 1'b0;
      \piso.data_r_256_sv2v_reg  <= 1'b0;
      \piso.data_r_255_sv2v_reg  <= 1'b0;
      \piso.data_r_254_sv2v_reg  <= 1'b0;
      \piso.data_r_253_sv2v_reg  <= 1'b0;
      \piso.data_r_252_sv2v_reg  <= 1'b0;
      \piso.data_r_251_sv2v_reg  <= 1'b0;
      \piso.data_r_250_sv2v_reg  <= 1'b0;
      \piso.data_r_249_sv2v_reg  <= 1'b0;
      \piso.data_r_248_sv2v_reg  <= 1'b0;
      \piso.data_r_247_sv2v_reg  <= 1'b0;
      \piso.data_r_246_sv2v_reg  <= 1'b0;
      \piso.data_r_245_sv2v_reg  <= 1'b0;
      \piso.data_r_244_sv2v_reg  <= 1'b0;
      \piso.data_r_243_sv2v_reg  <= 1'b0;
      \piso.data_r_242_sv2v_reg  <= 1'b0;
      \piso.data_r_241_sv2v_reg  <= 1'b0;
      \piso.data_r_240_sv2v_reg  <= 1'b0;
      \piso.data_r_239_sv2v_reg  <= 1'b0;
      \piso.data_r_238_sv2v_reg  <= 1'b0;
      \piso.data_r_237_sv2v_reg  <= 1'b0;
      \piso.data_r_236_sv2v_reg  <= 1'b0;
      \piso.data_r_235_sv2v_reg  <= 1'b0;
      \piso.data_r_234_sv2v_reg  <= 1'b0;
      \piso.data_r_233_sv2v_reg  <= 1'b0;
      \piso.data_r_232_sv2v_reg  <= 1'b0;
      \piso.data_r_231_sv2v_reg  <= 1'b0;
      \piso.data_r_230_sv2v_reg  <= 1'b0;
      \piso.data_r_229_sv2v_reg  <= 1'b0;
      \piso.data_r_228_sv2v_reg  <= 1'b0;
      \piso.data_r_227_sv2v_reg  <= 1'b0;
      \piso.data_r_226_sv2v_reg  <= 1'b0;
      \piso.data_r_225_sv2v_reg  <= 1'b0;
      \piso.data_r_224_sv2v_reg  <= 1'b0;
      \piso.data_r_223_sv2v_reg  <= 1'b0;
      \piso.data_r_222_sv2v_reg  <= 1'b0;
      \piso.data_r_221_sv2v_reg  <= 1'b0;
      \piso.data_r_220_sv2v_reg  <= 1'b0;
      \piso.data_r_219_sv2v_reg  <= 1'b0;
      \piso.data_r_218_sv2v_reg  <= 1'b0;
      \piso.data_r_217_sv2v_reg  <= 1'b0;
      \piso.data_r_216_sv2v_reg  <= 1'b0;
      \piso.data_r_215_sv2v_reg  <= 1'b0;
      \piso.data_r_214_sv2v_reg  <= 1'b0;
      \piso.data_r_213_sv2v_reg  <= 1'b0;
      \piso.data_r_212_sv2v_reg  <= 1'b0;
      \piso.data_r_211_sv2v_reg  <= 1'b0;
      \piso.data_r_210_sv2v_reg  <= 1'b0;
      \piso.data_r_209_sv2v_reg  <= 1'b0;
      \piso.data_r_208_sv2v_reg  <= 1'b0;
      \piso.data_r_207_sv2v_reg  <= 1'b0;
      \piso.data_r_206_sv2v_reg  <= 1'b0;
      \piso.data_r_205_sv2v_reg  <= 1'b0;
      \piso.data_r_204_sv2v_reg  <= 1'b0;
      \piso.data_r_203_sv2v_reg  <= 1'b0;
      \piso.data_r_202_sv2v_reg  <= 1'b0;
      \piso.data_r_201_sv2v_reg  <= 1'b0;
      \piso.data_r_200_sv2v_reg  <= 1'b0;
      \piso.data_r_199_sv2v_reg  <= 1'b0;
      \piso.data_r_198_sv2v_reg  <= 1'b0;
      \piso.data_r_197_sv2v_reg  <= 1'b0;
      \piso.data_r_196_sv2v_reg  <= 1'b0;
      \piso.data_r_195_sv2v_reg  <= 1'b0;
      \piso.data_r_194_sv2v_reg  <= 1'b0;
      \piso.data_r_193_sv2v_reg  <= 1'b0;
      \piso.data_r_192_sv2v_reg  <= 1'b0;
      \piso.data_r_191_sv2v_reg  <= 1'b0;
      \piso.data_r_190_sv2v_reg  <= 1'b0;
      \piso.data_r_189_sv2v_reg  <= 1'b0;
      \piso.data_r_188_sv2v_reg  <= 1'b0;
      \piso.data_r_187_sv2v_reg  <= 1'b0;
      \piso.data_r_186_sv2v_reg  <= 1'b0;
      \piso.data_r_185_sv2v_reg  <= 1'b0;
      \piso.data_r_184_sv2v_reg  <= 1'b0;
      \piso.data_r_183_sv2v_reg  <= 1'b0;
      \piso.data_r_182_sv2v_reg  <= 1'b0;
      \piso.data_r_181_sv2v_reg  <= 1'b0;
      \piso.data_r_180_sv2v_reg  <= 1'b0;
      \piso.data_r_179_sv2v_reg  <= 1'b0;
      \piso.data_r_178_sv2v_reg  <= 1'b0;
      \piso.data_r_177_sv2v_reg  <= 1'b0;
      \piso.data_r_176_sv2v_reg  <= 1'b0;
      \piso.data_r_175_sv2v_reg  <= 1'b0;
      \piso.data_r_174_sv2v_reg  <= 1'b0;
      \piso.data_r_173_sv2v_reg  <= 1'b0;
      \piso.data_r_172_sv2v_reg  <= 1'b0;
      \piso.data_r_171_sv2v_reg  <= 1'b0;
      \piso.data_r_170_sv2v_reg  <= 1'b0;
      \piso.data_r_169_sv2v_reg  <= 1'b0;
      \piso.data_r_168_sv2v_reg  <= 1'b0;
      \piso.data_r_167_sv2v_reg  <= 1'b0;
      \piso.data_r_166_sv2v_reg  <= 1'b0;
      \piso.data_r_165_sv2v_reg  <= 1'b0;
      \piso.data_r_164_sv2v_reg  <= 1'b0;
      \piso.data_r_163_sv2v_reg  <= 1'b0;
      \piso.data_r_162_sv2v_reg  <= 1'b0;
      \piso.data_r_161_sv2v_reg  <= 1'b0;
      \piso.data_r_160_sv2v_reg  <= 1'b0;
      \piso.data_r_159_sv2v_reg  <= 1'b0;
      \piso.data_r_158_sv2v_reg  <= 1'b0;
      \piso.data_r_157_sv2v_reg  <= 1'b0;
      \piso.data_r_156_sv2v_reg  <= 1'b0;
      \piso.data_r_155_sv2v_reg  <= 1'b0;
      \piso.data_r_154_sv2v_reg  <= 1'b0;
      \piso.data_r_153_sv2v_reg  <= 1'b0;
      \piso.data_r_152_sv2v_reg  <= 1'b0;
      \piso.data_r_151_sv2v_reg  <= 1'b0;
      \piso.data_r_150_sv2v_reg  <= 1'b0;
      \piso.data_r_149_sv2v_reg  <= 1'b0;
      \piso.data_r_148_sv2v_reg  <= 1'b0;
      \piso.data_r_147_sv2v_reg  <= 1'b0;
      \piso.data_r_146_sv2v_reg  <= 1'b0;
      \piso.data_r_145_sv2v_reg  <= 1'b0;
      \piso.data_r_144_sv2v_reg  <= 1'b0;
      \piso.data_r_143_sv2v_reg  <= 1'b0;
      \piso.data_r_142_sv2v_reg  <= 1'b0;
      \piso.data_r_141_sv2v_reg  <= 1'b0;
      \piso.data_r_140_sv2v_reg  <= 1'b0;
      \piso.data_r_139_sv2v_reg  <= 1'b0;
      \piso.data_r_138_sv2v_reg  <= 1'b0;
      \piso.data_r_137_sv2v_reg  <= 1'b0;
      \piso.data_r_136_sv2v_reg  <= 1'b0;
      \piso.data_r_135_sv2v_reg  <= 1'b0;
      \piso.data_r_134_sv2v_reg  <= 1'b0;
      \piso.data_r_133_sv2v_reg  <= 1'b0;
      \piso.data_r_132_sv2v_reg  <= 1'b0;
      \piso.data_r_131_sv2v_reg  <= 1'b0;
      \piso.data_r_130_sv2v_reg  <= 1'b0;
      \piso.data_r_129_sv2v_reg  <= 1'b0;
      \piso.data_r_128_sv2v_reg  <= 1'b0;
      \piso.data_r_127_sv2v_reg  <= 1'b0;
      \piso.data_r_126_sv2v_reg  <= 1'b0;
      \piso.data_r_125_sv2v_reg  <= 1'b0;
      \piso.data_r_124_sv2v_reg  <= 1'b0;
      \piso.data_r_123_sv2v_reg  <= 1'b0;
      \piso.data_r_122_sv2v_reg  <= 1'b0;
      \piso.data_r_121_sv2v_reg  <= 1'b0;
      \piso.data_r_120_sv2v_reg  <= 1'b0;
      \piso.data_r_119_sv2v_reg  <= 1'b0;
      \piso.data_r_118_sv2v_reg  <= 1'b0;
      \piso.data_r_117_sv2v_reg  <= 1'b0;
      \piso.data_r_116_sv2v_reg  <= 1'b0;
      \piso.data_r_115_sv2v_reg  <= 1'b0;
      \piso.data_r_114_sv2v_reg  <= 1'b0;
      \piso.data_r_113_sv2v_reg  <= 1'b0;
      \piso.data_r_112_sv2v_reg  <= 1'b0;
      \piso.data_r_111_sv2v_reg  <= 1'b0;
      \piso.data_r_110_sv2v_reg  <= 1'b0;
      \piso.data_r_109_sv2v_reg  <= 1'b0;
      \piso.data_r_108_sv2v_reg  <= 1'b0;
      \piso.data_r_107_sv2v_reg  <= 1'b0;
      \piso.data_r_106_sv2v_reg  <= 1'b0;
      \piso.data_r_105_sv2v_reg  <= 1'b0;
      \piso.data_r_104_sv2v_reg  <= 1'b0;
      \piso.data_r_103_sv2v_reg  <= 1'b0;
      \piso.data_r_102_sv2v_reg  <= 1'b0;
      \piso.data_r_101_sv2v_reg  <= 1'b0;
      \piso.data_r_100_sv2v_reg  <= 1'b0;
      \piso.data_r_99_sv2v_reg  <= 1'b0;
      \piso.data_r_98_sv2v_reg  <= 1'b0;
      \piso.data_r_97_sv2v_reg  <= 1'b0;
      \piso.data_r_96_sv2v_reg  <= 1'b0;
      \piso.data_r_95_sv2v_reg  <= 1'b0;
      \piso.data_r_94_sv2v_reg  <= 1'b0;
      \piso.data_r_93_sv2v_reg  <= 1'b0;
      \piso.data_r_92_sv2v_reg  <= 1'b0;
      \piso.data_r_91_sv2v_reg  <= 1'b0;
      \piso.data_r_90_sv2v_reg  <= 1'b0;
      \piso.data_r_89_sv2v_reg  <= 1'b0;
      \piso.data_r_88_sv2v_reg  <= 1'b0;
      \piso.data_r_87_sv2v_reg  <= 1'b0;
      \piso.data_r_86_sv2v_reg  <= 1'b0;
      \piso.data_r_85_sv2v_reg  <= 1'b0;
      \piso.data_r_84_sv2v_reg  <= 1'b0;
      \piso.data_r_83_sv2v_reg  <= 1'b0;
      \piso.data_r_82_sv2v_reg  <= 1'b0;
      \piso.data_r_81_sv2v_reg  <= 1'b0;
      \piso.data_r_80_sv2v_reg  <= 1'b0;
      \piso.data_r_79_sv2v_reg  <= 1'b0;
      \piso.data_r_78_sv2v_reg  <= 1'b0;
      \piso.data_r_77_sv2v_reg  <= 1'b0;
      \piso.data_r_76_sv2v_reg  <= 1'b0;
      \piso.data_r_75_sv2v_reg  <= 1'b0;
      \piso.data_r_74_sv2v_reg  <= 1'b0;
      \piso.data_r_73_sv2v_reg  <= 1'b0;
      \piso.data_r_72_sv2v_reg  <= 1'b0;
      \piso.data_r_71_sv2v_reg  <= 1'b0;
      \piso.data_r_70_sv2v_reg  <= 1'b0;
      \piso.data_r_69_sv2v_reg  <= 1'b0;
      \piso.data_r_68_sv2v_reg  <= 1'b0;
      \piso.data_r_67_sv2v_reg  <= 1'b0;
      \piso.data_r_66_sv2v_reg  <= 1'b0;
      \piso.data_r_65_sv2v_reg  <= 1'b0;
      \piso.data_r_64_sv2v_reg  <= 1'b0;
      \piso.data_r_63_sv2v_reg  <= 1'b0;
      \piso.data_r_62_sv2v_reg  <= 1'b0;
      \piso.data_r_61_sv2v_reg  <= 1'b0;
      \piso.data_r_60_sv2v_reg  <= 1'b0;
      \piso.data_r_59_sv2v_reg  <= 1'b0;
      \piso.data_r_58_sv2v_reg  <= 1'b0;
      \piso.data_r_57_sv2v_reg  <= 1'b0;
      \piso.data_r_56_sv2v_reg  <= 1'b0;
      \piso.data_r_55_sv2v_reg  <= 1'b0;
      \piso.data_r_54_sv2v_reg  <= 1'b0;
      \piso.data_r_53_sv2v_reg  <= 1'b0;
      \piso.data_r_52_sv2v_reg  <= 1'b0;
      \piso.data_r_51_sv2v_reg  <= 1'b0;
      \piso.data_r_50_sv2v_reg  <= 1'b0;
      \piso.data_r_49_sv2v_reg  <= 1'b0;
      \piso.data_r_48_sv2v_reg  <= 1'b0;
      \piso.data_r_47_sv2v_reg  <= 1'b0;
      \piso.data_r_46_sv2v_reg  <= 1'b0;
      \piso.data_r_45_sv2v_reg  <= 1'b0;
      \piso.data_r_44_sv2v_reg  <= 1'b0;
      \piso.data_r_43_sv2v_reg  <= 1'b0;
      \piso.data_r_42_sv2v_reg  <= 1'b0;
      \piso.data_r_41_sv2v_reg  <= 1'b0;
      \piso.data_r_40_sv2v_reg  <= 1'b0;
      \piso.data_r_39_sv2v_reg  <= 1'b0;
      \piso.data_r_38_sv2v_reg  <= 1'b0;
      \piso.data_r_37_sv2v_reg  <= 1'b0;
      \piso.data_r_36_sv2v_reg  <= 1'b0;
      \piso.data_r_35_sv2v_reg  <= 1'b0;
      \piso.data_r_34_sv2v_reg  <= 1'b0;
      \piso.data_r_33_sv2v_reg  <= 1'b0;
      \piso.data_r_32_sv2v_reg  <= 1'b0;
      \piso.data_r_31_sv2v_reg  <= 1'b0;
      \piso.data_r_30_sv2v_reg  <= 1'b0;
      \piso.data_r_29_sv2v_reg  <= 1'b0;
      \piso.data_r_28_sv2v_reg  <= 1'b0;
      \piso.data_r_27_sv2v_reg  <= 1'b0;
      \piso.data_r_26_sv2v_reg  <= 1'b0;
      \piso.data_r_25_sv2v_reg  <= 1'b0;
      \piso.data_r_24_sv2v_reg  <= 1'b0;
      \piso.data_r_23_sv2v_reg  <= 1'b0;
      \piso.data_r_22_sv2v_reg  <= 1'b0;
      \piso.data_r_21_sv2v_reg  <= 1'b0;
      \piso.data_r_20_sv2v_reg  <= 1'b0;
      \piso.data_r_19_sv2v_reg  <= 1'b0;
      \piso.data_r_18_sv2v_reg  <= 1'b0;
      \piso.data_r_17_sv2v_reg  <= 1'b0;
      \piso.data_r_16_sv2v_reg  <= 1'b0;
      \piso.data_r_15_sv2v_reg  <= 1'b0;
      \piso.data_r_14_sv2v_reg  <= 1'b0;
      \piso.data_r_13_sv2v_reg  <= 1'b0;
      \piso.data_r_12_sv2v_reg  <= 1'b0;
      \piso.data_r_11_sv2v_reg  <= 1'b0;
      \piso.data_r_10_sv2v_reg  <= 1'b0;
      \piso.data_r_9_sv2v_reg  <= 1'b0;
      \piso.data_r_8_sv2v_reg  <= 1'b0;
      \piso.data_r_7_sv2v_reg  <= 1'b0;
      \piso.data_r_6_sv2v_reg  <= 1'b0;
      \piso.data_r_5_sv2v_reg  <= 1'b0;
      \piso.data_r_4_sv2v_reg  <= 1'b0;
      \piso.data_r_3_sv2v_reg  <= 1'b0;
      \piso.data_r_2_sv2v_reg  <= 1'b0;
      \piso.data_r_1_sv2v_reg  <= 1'b0;
      \piso.data_r_0_sv2v_reg  <= 1'b0;
    end else if(N6) begin
      \piso.data_r_511_sv2v_reg  <= data_i[511];
      \piso.data_r_510_sv2v_reg  <= data_i[510];
      \piso.data_r_509_sv2v_reg  <= data_i[509];
      \piso.data_r_508_sv2v_reg  <= data_i[508];
      \piso.data_r_507_sv2v_reg  <= data_i[507];
      \piso.data_r_506_sv2v_reg  <= data_i[506];
      \piso.data_r_505_sv2v_reg  <= data_i[505];
      \piso.data_r_504_sv2v_reg  <= data_i[504];
      \piso.data_r_503_sv2v_reg  <= data_i[503];
      \piso.data_r_502_sv2v_reg  <= data_i[502];
      \piso.data_r_501_sv2v_reg  <= data_i[501];
      \piso.data_r_500_sv2v_reg  <= data_i[500];
      \piso.data_r_499_sv2v_reg  <= data_i[499];
      \piso.data_r_498_sv2v_reg  <= data_i[498];
      \piso.data_r_497_sv2v_reg  <= data_i[497];
      \piso.data_r_496_sv2v_reg  <= data_i[496];
      \piso.data_r_495_sv2v_reg  <= data_i[495];
      \piso.data_r_494_sv2v_reg  <= data_i[494];
      \piso.data_r_493_sv2v_reg  <= data_i[493];
      \piso.data_r_492_sv2v_reg  <= data_i[492];
      \piso.data_r_491_sv2v_reg  <= data_i[491];
      \piso.data_r_490_sv2v_reg  <= data_i[490];
      \piso.data_r_489_sv2v_reg  <= data_i[489];
      \piso.data_r_488_sv2v_reg  <= data_i[488];
      \piso.data_r_487_sv2v_reg  <= data_i[487];
      \piso.data_r_486_sv2v_reg  <= data_i[486];
      \piso.data_r_485_sv2v_reg  <= data_i[485];
      \piso.data_r_484_sv2v_reg  <= data_i[484];
      \piso.data_r_483_sv2v_reg  <= data_i[483];
      \piso.data_r_482_sv2v_reg  <= data_i[482];
      \piso.data_r_481_sv2v_reg  <= data_i[481];
      \piso.data_r_480_sv2v_reg  <= data_i[480];
      \piso.data_r_479_sv2v_reg  <= data_i[479];
      \piso.data_r_478_sv2v_reg  <= data_i[478];
      \piso.data_r_477_sv2v_reg  <= data_i[477];
      \piso.data_r_476_sv2v_reg  <= data_i[476];
      \piso.data_r_475_sv2v_reg  <= data_i[475];
      \piso.data_r_474_sv2v_reg  <= data_i[474];
      \piso.data_r_473_sv2v_reg  <= data_i[473];
      \piso.data_r_472_sv2v_reg  <= data_i[472];
      \piso.data_r_471_sv2v_reg  <= data_i[471];
      \piso.data_r_470_sv2v_reg  <= data_i[470];
      \piso.data_r_469_sv2v_reg  <= data_i[469];
      \piso.data_r_468_sv2v_reg  <= data_i[468];
      \piso.data_r_467_sv2v_reg  <= data_i[467];
      \piso.data_r_466_sv2v_reg  <= data_i[466];
      \piso.data_r_465_sv2v_reg  <= data_i[465];
      \piso.data_r_464_sv2v_reg  <= data_i[464];
      \piso.data_r_463_sv2v_reg  <= data_i[463];
      \piso.data_r_462_sv2v_reg  <= data_i[462];
      \piso.data_r_461_sv2v_reg  <= data_i[461];
      \piso.data_r_460_sv2v_reg  <= data_i[460];
      \piso.data_r_459_sv2v_reg  <= data_i[459];
      \piso.data_r_458_sv2v_reg  <= data_i[458];
      \piso.data_r_457_sv2v_reg  <= data_i[457];
      \piso.data_r_456_sv2v_reg  <= data_i[456];
      \piso.data_r_455_sv2v_reg  <= data_i[455];
      \piso.data_r_454_sv2v_reg  <= data_i[454];
      \piso.data_r_453_sv2v_reg  <= data_i[453];
      \piso.data_r_452_sv2v_reg  <= data_i[452];
      \piso.data_r_451_sv2v_reg  <= data_i[451];
      \piso.data_r_450_sv2v_reg  <= data_i[450];
      \piso.data_r_449_sv2v_reg  <= data_i[449];
      \piso.data_r_448_sv2v_reg  <= data_i[448];
      \piso.data_r_447_sv2v_reg  <= data_i[447];
      \piso.data_r_446_sv2v_reg  <= data_i[446];
      \piso.data_r_445_sv2v_reg  <= data_i[445];
      \piso.data_r_444_sv2v_reg  <= data_i[444];
      \piso.data_r_443_sv2v_reg  <= data_i[443];
      \piso.data_r_442_sv2v_reg  <= data_i[442];
      \piso.data_r_441_sv2v_reg  <= data_i[441];
      \piso.data_r_440_sv2v_reg  <= data_i[440];
      \piso.data_r_439_sv2v_reg  <= data_i[439];
      \piso.data_r_438_sv2v_reg  <= data_i[438];
      \piso.data_r_437_sv2v_reg  <= data_i[437];
      \piso.data_r_436_sv2v_reg  <= data_i[436];
      \piso.data_r_435_sv2v_reg  <= data_i[435];
      \piso.data_r_434_sv2v_reg  <= data_i[434];
      \piso.data_r_433_sv2v_reg  <= data_i[433];
      \piso.data_r_432_sv2v_reg  <= data_i[432];
      \piso.data_r_431_sv2v_reg  <= data_i[431];
      \piso.data_r_430_sv2v_reg  <= data_i[430];
      \piso.data_r_429_sv2v_reg  <= data_i[429];
      \piso.data_r_428_sv2v_reg  <= data_i[428];
      \piso.data_r_427_sv2v_reg  <= data_i[427];
      \piso.data_r_426_sv2v_reg  <= data_i[426];
      \piso.data_r_425_sv2v_reg  <= data_i[425];
      \piso.data_r_424_sv2v_reg  <= data_i[424];
      \piso.data_r_423_sv2v_reg  <= data_i[423];
      \piso.data_r_422_sv2v_reg  <= data_i[422];
      \piso.data_r_421_sv2v_reg  <= data_i[421];
      \piso.data_r_420_sv2v_reg  <= data_i[420];
      \piso.data_r_419_sv2v_reg  <= data_i[419];
      \piso.data_r_418_sv2v_reg  <= data_i[418];
      \piso.data_r_417_sv2v_reg  <= data_i[417];
      \piso.data_r_416_sv2v_reg  <= data_i[416];
      \piso.data_r_415_sv2v_reg  <= data_i[415];
      \piso.data_r_414_sv2v_reg  <= data_i[414];
      \piso.data_r_413_sv2v_reg  <= data_i[413];
      \piso.data_r_412_sv2v_reg  <= data_i[412];
      \piso.data_r_411_sv2v_reg  <= data_i[411];
      \piso.data_r_410_sv2v_reg  <= data_i[410];
      \piso.data_r_409_sv2v_reg  <= data_i[409];
      \piso.data_r_408_sv2v_reg  <= data_i[408];
      \piso.data_r_407_sv2v_reg  <= data_i[407];
      \piso.data_r_406_sv2v_reg  <= data_i[406];
      \piso.data_r_405_sv2v_reg  <= data_i[405];
      \piso.data_r_404_sv2v_reg  <= data_i[404];
      \piso.data_r_403_sv2v_reg  <= data_i[403];
      \piso.data_r_402_sv2v_reg  <= data_i[402];
      \piso.data_r_401_sv2v_reg  <= data_i[401];
      \piso.data_r_400_sv2v_reg  <= data_i[400];
      \piso.data_r_399_sv2v_reg  <= data_i[399];
      \piso.data_r_398_sv2v_reg  <= data_i[398];
      \piso.data_r_397_sv2v_reg  <= data_i[397];
      \piso.data_r_396_sv2v_reg  <= data_i[396];
      \piso.data_r_395_sv2v_reg  <= data_i[395];
      \piso.data_r_394_sv2v_reg  <= data_i[394];
      \piso.data_r_393_sv2v_reg  <= data_i[393];
      \piso.data_r_392_sv2v_reg  <= data_i[392];
      \piso.data_r_391_sv2v_reg  <= data_i[391];
      \piso.data_r_390_sv2v_reg  <= data_i[390];
      \piso.data_r_389_sv2v_reg  <= data_i[389];
      \piso.data_r_388_sv2v_reg  <= data_i[388];
      \piso.data_r_387_sv2v_reg  <= data_i[387];
      \piso.data_r_386_sv2v_reg  <= data_i[386];
      \piso.data_r_385_sv2v_reg  <= data_i[385];
      \piso.data_r_384_sv2v_reg  <= data_i[384];
      \piso.data_r_383_sv2v_reg  <= data_i[383];
      \piso.data_r_382_sv2v_reg  <= data_i[382];
      \piso.data_r_381_sv2v_reg  <= data_i[381];
      \piso.data_r_380_sv2v_reg  <= data_i[380];
      \piso.data_r_379_sv2v_reg  <= data_i[379];
      \piso.data_r_378_sv2v_reg  <= data_i[378];
      \piso.data_r_377_sv2v_reg  <= data_i[377];
      \piso.data_r_376_sv2v_reg  <= data_i[376];
      \piso.data_r_375_sv2v_reg  <= data_i[375];
      \piso.data_r_374_sv2v_reg  <= data_i[374];
      \piso.data_r_373_sv2v_reg  <= data_i[373];
      \piso.data_r_372_sv2v_reg  <= data_i[372];
      \piso.data_r_371_sv2v_reg  <= data_i[371];
      \piso.data_r_370_sv2v_reg  <= data_i[370];
      \piso.data_r_369_sv2v_reg  <= data_i[369];
      \piso.data_r_368_sv2v_reg  <= data_i[368];
      \piso.data_r_367_sv2v_reg  <= data_i[367];
      \piso.data_r_366_sv2v_reg  <= data_i[366];
      \piso.data_r_365_sv2v_reg  <= data_i[365];
      \piso.data_r_364_sv2v_reg  <= data_i[364];
      \piso.data_r_363_sv2v_reg  <= data_i[363];
      \piso.data_r_362_sv2v_reg  <= data_i[362];
      \piso.data_r_361_sv2v_reg  <= data_i[361];
      \piso.data_r_360_sv2v_reg  <= data_i[360];
      \piso.data_r_359_sv2v_reg  <= data_i[359];
      \piso.data_r_358_sv2v_reg  <= data_i[358];
      \piso.data_r_357_sv2v_reg  <= data_i[357];
      \piso.data_r_356_sv2v_reg  <= data_i[356];
      \piso.data_r_355_sv2v_reg  <= data_i[355];
      \piso.data_r_354_sv2v_reg  <= data_i[354];
      \piso.data_r_353_sv2v_reg  <= data_i[353];
      \piso.data_r_352_sv2v_reg  <= data_i[352];
      \piso.data_r_351_sv2v_reg  <= data_i[351];
      \piso.data_r_350_sv2v_reg  <= data_i[350];
      \piso.data_r_349_sv2v_reg  <= data_i[349];
      \piso.data_r_348_sv2v_reg  <= data_i[348];
      \piso.data_r_347_sv2v_reg  <= data_i[347];
      \piso.data_r_346_sv2v_reg  <= data_i[346];
      \piso.data_r_345_sv2v_reg  <= data_i[345];
      \piso.data_r_344_sv2v_reg  <= data_i[344];
      \piso.data_r_343_sv2v_reg  <= data_i[343];
      \piso.data_r_342_sv2v_reg  <= data_i[342];
      \piso.data_r_341_sv2v_reg  <= data_i[341];
      \piso.data_r_340_sv2v_reg  <= data_i[340];
      \piso.data_r_339_sv2v_reg  <= data_i[339];
      \piso.data_r_338_sv2v_reg  <= data_i[338];
      \piso.data_r_337_sv2v_reg  <= data_i[337];
      \piso.data_r_336_sv2v_reg  <= data_i[336];
      \piso.data_r_335_sv2v_reg  <= data_i[335];
      \piso.data_r_334_sv2v_reg  <= data_i[334];
      \piso.data_r_333_sv2v_reg  <= data_i[333];
      \piso.data_r_332_sv2v_reg  <= data_i[332];
      \piso.data_r_331_sv2v_reg  <= data_i[331];
      \piso.data_r_330_sv2v_reg  <= data_i[330];
      \piso.data_r_329_sv2v_reg  <= data_i[329];
      \piso.data_r_328_sv2v_reg  <= data_i[328];
      \piso.data_r_327_sv2v_reg  <= data_i[327];
      \piso.data_r_326_sv2v_reg  <= data_i[326];
      \piso.data_r_325_sv2v_reg  <= data_i[325];
      \piso.data_r_324_sv2v_reg  <= data_i[324];
      \piso.data_r_323_sv2v_reg  <= data_i[323];
      \piso.data_r_322_sv2v_reg  <= data_i[322];
      \piso.data_r_321_sv2v_reg  <= data_i[321];
      \piso.data_r_320_sv2v_reg  <= data_i[320];
      \piso.data_r_319_sv2v_reg  <= data_i[319];
      \piso.data_r_318_sv2v_reg  <= data_i[318];
      \piso.data_r_317_sv2v_reg  <= data_i[317];
      \piso.data_r_316_sv2v_reg  <= data_i[316];
      \piso.data_r_315_sv2v_reg  <= data_i[315];
      \piso.data_r_314_sv2v_reg  <= data_i[314];
      \piso.data_r_313_sv2v_reg  <= data_i[313];
      \piso.data_r_312_sv2v_reg  <= data_i[312];
      \piso.data_r_311_sv2v_reg  <= data_i[311];
      \piso.data_r_310_sv2v_reg  <= data_i[310];
      \piso.data_r_309_sv2v_reg  <= data_i[309];
      \piso.data_r_308_sv2v_reg  <= data_i[308];
      \piso.data_r_307_sv2v_reg  <= data_i[307];
      \piso.data_r_306_sv2v_reg  <= data_i[306];
      \piso.data_r_305_sv2v_reg  <= data_i[305];
      \piso.data_r_304_sv2v_reg  <= data_i[304];
      \piso.data_r_303_sv2v_reg  <= data_i[303];
      \piso.data_r_302_sv2v_reg  <= data_i[302];
      \piso.data_r_301_sv2v_reg  <= data_i[301];
      \piso.data_r_300_sv2v_reg  <= data_i[300];
      \piso.data_r_299_sv2v_reg  <= data_i[299];
      \piso.data_r_298_sv2v_reg  <= data_i[298];
      \piso.data_r_297_sv2v_reg  <= data_i[297];
      \piso.data_r_296_sv2v_reg  <= data_i[296];
      \piso.data_r_295_sv2v_reg  <= data_i[295];
      \piso.data_r_294_sv2v_reg  <= data_i[294];
      \piso.data_r_293_sv2v_reg  <= data_i[293];
      \piso.data_r_292_sv2v_reg  <= data_i[292];
      \piso.data_r_291_sv2v_reg  <= data_i[291];
      \piso.data_r_290_sv2v_reg  <= data_i[290];
      \piso.data_r_289_sv2v_reg  <= data_i[289];
      \piso.data_r_288_sv2v_reg  <= data_i[288];
      \piso.data_r_287_sv2v_reg  <= data_i[287];
      \piso.data_r_286_sv2v_reg  <= data_i[286];
      \piso.data_r_285_sv2v_reg  <= data_i[285];
      \piso.data_r_284_sv2v_reg  <= data_i[284];
      \piso.data_r_283_sv2v_reg  <= data_i[283];
      \piso.data_r_282_sv2v_reg  <= data_i[282];
      \piso.data_r_281_sv2v_reg  <= data_i[281];
      \piso.data_r_280_sv2v_reg  <= data_i[280];
      \piso.data_r_279_sv2v_reg  <= data_i[279];
      \piso.data_r_278_sv2v_reg  <= data_i[278];
      \piso.data_r_277_sv2v_reg  <= data_i[277];
      \piso.data_r_276_sv2v_reg  <= data_i[276];
      \piso.data_r_275_sv2v_reg  <= data_i[275];
      \piso.data_r_274_sv2v_reg  <= data_i[274];
      \piso.data_r_273_sv2v_reg  <= data_i[273];
      \piso.data_r_272_sv2v_reg  <= data_i[272];
      \piso.data_r_271_sv2v_reg  <= data_i[271];
      \piso.data_r_270_sv2v_reg  <= data_i[270];
      \piso.data_r_269_sv2v_reg  <= data_i[269];
      \piso.data_r_268_sv2v_reg  <= data_i[268];
      \piso.data_r_267_sv2v_reg  <= data_i[267];
      \piso.data_r_266_sv2v_reg  <= data_i[266];
      \piso.data_r_265_sv2v_reg  <= data_i[265];
      \piso.data_r_264_sv2v_reg  <= data_i[264];
      \piso.data_r_263_sv2v_reg  <= data_i[263];
      \piso.data_r_262_sv2v_reg  <= data_i[262];
      \piso.data_r_261_sv2v_reg  <= data_i[261];
      \piso.data_r_260_sv2v_reg  <= data_i[260];
      \piso.data_r_259_sv2v_reg  <= data_i[259];
      \piso.data_r_258_sv2v_reg  <= data_i[258];
      \piso.data_r_257_sv2v_reg  <= data_i[257];
      \piso.data_r_256_sv2v_reg  <= data_i[256];
      \piso.data_r_255_sv2v_reg  <= data_i[255];
      \piso.data_r_254_sv2v_reg  <= data_i[254];
      \piso.data_r_253_sv2v_reg  <= data_i[253];
      \piso.data_r_252_sv2v_reg  <= data_i[252];
      \piso.data_r_251_sv2v_reg  <= data_i[251];
      \piso.data_r_250_sv2v_reg  <= data_i[250];
      \piso.data_r_249_sv2v_reg  <= data_i[249];
      \piso.data_r_248_sv2v_reg  <= data_i[248];
      \piso.data_r_247_sv2v_reg  <= data_i[247];
      \piso.data_r_246_sv2v_reg  <= data_i[246];
      \piso.data_r_245_sv2v_reg  <= data_i[245];
      \piso.data_r_244_sv2v_reg  <= data_i[244];
      \piso.data_r_243_sv2v_reg  <= data_i[243];
      \piso.data_r_242_sv2v_reg  <= data_i[242];
      \piso.data_r_241_sv2v_reg  <= data_i[241];
      \piso.data_r_240_sv2v_reg  <= data_i[240];
      \piso.data_r_239_sv2v_reg  <= data_i[239];
      \piso.data_r_238_sv2v_reg  <= data_i[238];
      \piso.data_r_237_sv2v_reg  <= data_i[237];
      \piso.data_r_236_sv2v_reg  <= data_i[236];
      \piso.data_r_235_sv2v_reg  <= data_i[235];
      \piso.data_r_234_sv2v_reg  <= data_i[234];
      \piso.data_r_233_sv2v_reg  <= data_i[233];
      \piso.data_r_232_sv2v_reg  <= data_i[232];
      \piso.data_r_231_sv2v_reg  <= data_i[231];
      \piso.data_r_230_sv2v_reg  <= data_i[230];
      \piso.data_r_229_sv2v_reg  <= data_i[229];
      \piso.data_r_228_sv2v_reg  <= data_i[228];
      \piso.data_r_227_sv2v_reg  <= data_i[227];
      \piso.data_r_226_sv2v_reg  <= data_i[226];
      \piso.data_r_225_sv2v_reg  <= data_i[225];
      \piso.data_r_224_sv2v_reg  <= data_i[224];
      \piso.data_r_223_sv2v_reg  <= data_i[223];
      \piso.data_r_222_sv2v_reg  <= data_i[222];
      \piso.data_r_221_sv2v_reg  <= data_i[221];
      \piso.data_r_220_sv2v_reg  <= data_i[220];
      \piso.data_r_219_sv2v_reg  <= data_i[219];
      \piso.data_r_218_sv2v_reg  <= data_i[218];
      \piso.data_r_217_sv2v_reg  <= data_i[217];
      \piso.data_r_216_sv2v_reg  <= data_i[216];
      \piso.data_r_215_sv2v_reg  <= data_i[215];
      \piso.data_r_214_sv2v_reg  <= data_i[214];
      \piso.data_r_213_sv2v_reg  <= data_i[213];
      \piso.data_r_212_sv2v_reg  <= data_i[212];
      \piso.data_r_211_sv2v_reg  <= data_i[211];
      \piso.data_r_210_sv2v_reg  <= data_i[210];
      \piso.data_r_209_sv2v_reg  <= data_i[209];
      \piso.data_r_208_sv2v_reg  <= data_i[208];
      \piso.data_r_207_sv2v_reg  <= data_i[207];
      \piso.data_r_206_sv2v_reg  <= data_i[206];
      \piso.data_r_205_sv2v_reg  <= data_i[205];
      \piso.data_r_204_sv2v_reg  <= data_i[204];
      \piso.data_r_203_sv2v_reg  <= data_i[203];
      \piso.data_r_202_sv2v_reg  <= data_i[202];
      \piso.data_r_201_sv2v_reg  <= data_i[201];
      \piso.data_r_200_sv2v_reg  <= data_i[200];
      \piso.data_r_199_sv2v_reg  <= data_i[199];
      \piso.data_r_198_sv2v_reg  <= data_i[198];
      \piso.data_r_197_sv2v_reg  <= data_i[197];
      \piso.data_r_196_sv2v_reg  <= data_i[196];
      \piso.data_r_195_sv2v_reg  <= data_i[195];
      \piso.data_r_194_sv2v_reg  <= data_i[194];
      \piso.data_r_193_sv2v_reg  <= data_i[193];
      \piso.data_r_192_sv2v_reg  <= data_i[192];
      \piso.data_r_191_sv2v_reg  <= data_i[191];
      \piso.data_r_190_sv2v_reg  <= data_i[190];
      \piso.data_r_189_sv2v_reg  <= data_i[189];
      \piso.data_r_188_sv2v_reg  <= data_i[188];
      \piso.data_r_187_sv2v_reg  <= data_i[187];
      \piso.data_r_186_sv2v_reg  <= data_i[186];
      \piso.data_r_185_sv2v_reg  <= data_i[185];
      \piso.data_r_184_sv2v_reg  <= data_i[184];
      \piso.data_r_183_sv2v_reg  <= data_i[183];
      \piso.data_r_182_sv2v_reg  <= data_i[182];
      \piso.data_r_181_sv2v_reg  <= data_i[181];
      \piso.data_r_180_sv2v_reg  <= data_i[180];
      \piso.data_r_179_sv2v_reg  <= data_i[179];
      \piso.data_r_178_sv2v_reg  <= data_i[178];
      \piso.data_r_177_sv2v_reg  <= data_i[177];
      \piso.data_r_176_sv2v_reg  <= data_i[176];
      \piso.data_r_175_sv2v_reg  <= data_i[175];
      \piso.data_r_174_sv2v_reg  <= data_i[174];
      \piso.data_r_173_sv2v_reg  <= data_i[173];
      \piso.data_r_172_sv2v_reg  <= data_i[172];
      \piso.data_r_171_sv2v_reg  <= data_i[171];
      \piso.data_r_170_sv2v_reg  <= data_i[170];
      \piso.data_r_169_sv2v_reg  <= data_i[169];
      \piso.data_r_168_sv2v_reg  <= data_i[168];
      \piso.data_r_167_sv2v_reg  <= data_i[167];
      \piso.data_r_166_sv2v_reg  <= data_i[166];
      \piso.data_r_165_sv2v_reg  <= data_i[165];
      \piso.data_r_164_sv2v_reg  <= data_i[164];
      \piso.data_r_163_sv2v_reg  <= data_i[163];
      \piso.data_r_162_sv2v_reg  <= data_i[162];
      \piso.data_r_161_sv2v_reg  <= data_i[161];
      \piso.data_r_160_sv2v_reg  <= data_i[160];
      \piso.data_r_159_sv2v_reg  <= data_i[159];
      \piso.data_r_158_sv2v_reg  <= data_i[158];
      \piso.data_r_157_sv2v_reg  <= data_i[157];
      \piso.data_r_156_sv2v_reg  <= data_i[156];
      \piso.data_r_155_sv2v_reg  <= data_i[155];
      \piso.data_r_154_sv2v_reg  <= data_i[154];
      \piso.data_r_153_sv2v_reg  <= data_i[153];
      \piso.data_r_152_sv2v_reg  <= data_i[152];
      \piso.data_r_151_sv2v_reg  <= data_i[151];
      \piso.data_r_150_sv2v_reg  <= data_i[150];
      \piso.data_r_149_sv2v_reg  <= data_i[149];
      \piso.data_r_148_sv2v_reg  <= data_i[148];
      \piso.data_r_147_sv2v_reg  <= data_i[147];
      \piso.data_r_146_sv2v_reg  <= data_i[146];
      \piso.data_r_145_sv2v_reg  <= data_i[145];
      \piso.data_r_144_sv2v_reg  <= data_i[144];
      \piso.data_r_143_sv2v_reg  <= data_i[143];
      \piso.data_r_142_sv2v_reg  <= data_i[142];
      \piso.data_r_141_sv2v_reg  <= data_i[141];
      \piso.data_r_140_sv2v_reg  <= data_i[140];
      \piso.data_r_139_sv2v_reg  <= data_i[139];
      \piso.data_r_138_sv2v_reg  <= data_i[138];
      \piso.data_r_137_sv2v_reg  <= data_i[137];
      \piso.data_r_136_sv2v_reg  <= data_i[136];
      \piso.data_r_135_sv2v_reg  <= data_i[135];
      \piso.data_r_134_sv2v_reg  <= data_i[134];
      \piso.data_r_133_sv2v_reg  <= data_i[133];
      \piso.data_r_132_sv2v_reg  <= data_i[132];
      \piso.data_r_131_sv2v_reg  <= data_i[131];
      \piso.data_r_130_sv2v_reg  <= data_i[130];
      \piso.data_r_129_sv2v_reg  <= data_i[129];
      \piso.data_r_128_sv2v_reg  <= data_i[128];
      \piso.data_r_127_sv2v_reg  <= data_i[127];
      \piso.data_r_126_sv2v_reg  <= data_i[126];
      \piso.data_r_125_sv2v_reg  <= data_i[125];
      \piso.data_r_124_sv2v_reg  <= data_i[124];
      \piso.data_r_123_sv2v_reg  <= data_i[123];
      \piso.data_r_122_sv2v_reg  <= data_i[122];
      \piso.data_r_121_sv2v_reg  <= data_i[121];
      \piso.data_r_120_sv2v_reg  <= data_i[120];
      \piso.data_r_119_sv2v_reg  <= data_i[119];
      \piso.data_r_118_sv2v_reg  <= data_i[118];
      \piso.data_r_117_sv2v_reg  <= data_i[117];
      \piso.data_r_116_sv2v_reg  <= data_i[116];
      \piso.data_r_115_sv2v_reg  <= data_i[115];
      \piso.data_r_114_sv2v_reg  <= data_i[114];
      \piso.data_r_113_sv2v_reg  <= data_i[113];
      \piso.data_r_112_sv2v_reg  <= data_i[112];
      \piso.data_r_111_sv2v_reg  <= data_i[111];
      \piso.data_r_110_sv2v_reg  <= data_i[110];
      \piso.data_r_109_sv2v_reg  <= data_i[109];
      \piso.data_r_108_sv2v_reg  <= data_i[108];
      \piso.data_r_107_sv2v_reg  <= data_i[107];
      \piso.data_r_106_sv2v_reg  <= data_i[106];
      \piso.data_r_105_sv2v_reg  <= data_i[105];
      \piso.data_r_104_sv2v_reg  <= data_i[104];
      \piso.data_r_103_sv2v_reg  <= data_i[103];
      \piso.data_r_102_sv2v_reg  <= data_i[102];
      \piso.data_r_101_sv2v_reg  <= data_i[101];
      \piso.data_r_100_sv2v_reg  <= data_i[100];
      \piso.data_r_99_sv2v_reg  <= data_i[99];
      \piso.data_r_98_sv2v_reg  <= data_i[98];
      \piso.data_r_97_sv2v_reg  <= data_i[97];
      \piso.data_r_96_sv2v_reg  <= data_i[96];
      \piso.data_r_95_sv2v_reg  <= data_i[95];
      \piso.data_r_94_sv2v_reg  <= data_i[94];
      \piso.data_r_93_sv2v_reg  <= data_i[93];
      \piso.data_r_92_sv2v_reg  <= data_i[92];
      \piso.data_r_91_sv2v_reg  <= data_i[91];
      \piso.data_r_90_sv2v_reg  <= data_i[90];
      \piso.data_r_89_sv2v_reg  <= data_i[89];
      \piso.data_r_88_sv2v_reg  <= data_i[88];
      \piso.data_r_87_sv2v_reg  <= data_i[87];
      \piso.data_r_86_sv2v_reg  <= data_i[86];
      \piso.data_r_85_sv2v_reg  <= data_i[85];
      \piso.data_r_84_sv2v_reg  <= data_i[84];
      \piso.data_r_83_sv2v_reg  <= data_i[83];
      \piso.data_r_82_sv2v_reg  <= data_i[82];
      \piso.data_r_81_sv2v_reg  <= data_i[81];
      \piso.data_r_80_sv2v_reg  <= data_i[80];
      \piso.data_r_79_sv2v_reg  <= data_i[79];
      \piso.data_r_78_sv2v_reg  <= data_i[78];
      \piso.data_r_77_sv2v_reg  <= data_i[77];
      \piso.data_r_76_sv2v_reg  <= data_i[76];
      \piso.data_r_75_sv2v_reg  <= data_i[75];
      \piso.data_r_74_sv2v_reg  <= data_i[74];
      \piso.data_r_73_sv2v_reg  <= data_i[73];
      \piso.data_r_72_sv2v_reg  <= data_i[72];
      \piso.data_r_71_sv2v_reg  <= data_i[71];
      \piso.data_r_70_sv2v_reg  <= data_i[70];
      \piso.data_r_69_sv2v_reg  <= data_i[69];
      \piso.data_r_68_sv2v_reg  <= data_i[68];
      \piso.data_r_67_sv2v_reg  <= data_i[67];
      \piso.data_r_66_sv2v_reg  <= data_i[66];
      \piso.data_r_65_sv2v_reg  <= data_i[65];
      \piso.data_r_64_sv2v_reg  <= data_i[64];
      \piso.data_r_63_sv2v_reg  <= data_i[63];
      \piso.data_r_62_sv2v_reg  <= data_i[62];
      \piso.data_r_61_sv2v_reg  <= data_i[61];
      \piso.data_r_60_sv2v_reg  <= data_i[60];
      \piso.data_r_59_sv2v_reg  <= data_i[59];
      \piso.data_r_58_sv2v_reg  <= data_i[58];
      \piso.data_r_57_sv2v_reg  <= data_i[57];
      \piso.data_r_56_sv2v_reg  <= data_i[56];
      \piso.data_r_55_sv2v_reg  <= data_i[55];
      \piso.data_r_54_sv2v_reg  <= data_i[54];
      \piso.data_r_53_sv2v_reg  <= data_i[53];
      \piso.data_r_52_sv2v_reg  <= data_i[52];
      \piso.data_r_51_sv2v_reg  <= data_i[51];
      \piso.data_r_50_sv2v_reg  <= data_i[50];
      \piso.data_r_49_sv2v_reg  <= data_i[49];
      \piso.data_r_48_sv2v_reg  <= data_i[48];
      \piso.data_r_47_sv2v_reg  <= data_i[47];
      \piso.data_r_46_sv2v_reg  <= data_i[46];
      \piso.data_r_45_sv2v_reg  <= data_i[45];
      \piso.data_r_44_sv2v_reg  <= data_i[44];
      \piso.data_r_43_sv2v_reg  <= data_i[43];
      \piso.data_r_42_sv2v_reg  <= data_i[42];
      \piso.data_r_41_sv2v_reg  <= data_i[41];
      \piso.data_r_40_sv2v_reg  <= data_i[40];
      \piso.data_r_39_sv2v_reg  <= data_i[39];
      \piso.data_r_38_sv2v_reg  <= data_i[38];
      \piso.data_r_37_sv2v_reg  <= data_i[37];
      \piso.data_r_36_sv2v_reg  <= data_i[36];
      \piso.data_r_35_sv2v_reg  <= data_i[35];
      \piso.data_r_34_sv2v_reg  <= data_i[34];
      \piso.data_r_33_sv2v_reg  <= data_i[33];
      \piso.data_r_32_sv2v_reg  <= data_i[32];
      \piso.data_r_31_sv2v_reg  <= data_i[31];
      \piso.data_r_30_sv2v_reg  <= data_i[30];
      \piso.data_r_29_sv2v_reg  <= data_i[29];
      \piso.data_r_28_sv2v_reg  <= data_i[28];
      \piso.data_r_27_sv2v_reg  <= data_i[27];
      \piso.data_r_26_sv2v_reg  <= data_i[26];
      \piso.data_r_25_sv2v_reg  <= data_i[25];
      \piso.data_r_24_sv2v_reg  <= data_i[24];
      \piso.data_r_23_sv2v_reg  <= data_i[23];
      \piso.data_r_22_sv2v_reg  <= data_i[22];
      \piso.data_r_21_sv2v_reg  <= data_i[21];
      \piso.data_r_20_sv2v_reg  <= data_i[20];
      \piso.data_r_19_sv2v_reg  <= data_i[19];
      \piso.data_r_18_sv2v_reg  <= data_i[18];
      \piso.data_r_17_sv2v_reg  <= data_i[17];
      \piso.data_r_16_sv2v_reg  <= data_i[16];
      \piso.data_r_15_sv2v_reg  <= data_i[15];
      \piso.data_r_14_sv2v_reg  <= data_i[14];
      \piso.data_r_13_sv2v_reg  <= data_i[13];
      \piso.data_r_12_sv2v_reg  <= data_i[12];
      \piso.data_r_11_sv2v_reg  <= data_i[11];
      \piso.data_r_10_sv2v_reg  <= data_i[10];
      \piso.data_r_9_sv2v_reg  <= data_i[9];
      \piso.data_r_8_sv2v_reg  <= data_i[8];
      \piso.data_r_7_sv2v_reg  <= data_i[7];
      \piso.data_r_6_sv2v_reg  <= data_i[6];
      \piso.data_r_5_sv2v_reg  <= data_i[5];
      \piso.data_r_4_sv2v_reg  <= data_i[4];
      \piso.data_r_3_sv2v_reg  <= data_i[3];
      \piso.data_r_2_sv2v_reg  <= data_i[2];
      \piso.data_r_1_sv2v_reg  <= data_i[1];
      \piso.data_r_0_sv2v_reg  <= data_i[0];
    end 
    if(reset_i) begin
      \piso.shift_ctr_r_4_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_3_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_2_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_1_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_0_sv2v_reg  <= 1'b0;
    end else if(N87) begin
      \piso.shift_ctr_r_4_sv2v_reg  <= N13;
      \piso.shift_ctr_r_3_sv2v_reg  <= N12;
      \piso.shift_ctr_r_2_sv2v_reg  <= N11;
      \piso.shift_ctr_r_1_sv2v_reg  <= N10;
      \piso.shift_ctr_r_0_sv2v_reg  <= N9;
    end 
  end


endmodule

