

module top
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_i
);

  input [4095:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_o;
  output valid_o;

  bsg_parallel_in_serial_out
  wrapper
  (
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .valid_i(valid_i),
    .yumi_i(yumi_i),
    .ready_o(ready_o),
    .valid_o(valid_o)
  );


endmodule



module bsg_array_reverse_width_p32_els_p128
(
  i,
  o
);

  input [4095:0] i;
  output [4095:0] o;
  wire [4095:0] o;
  assign o[4095] = i[31];
  assign o[4094] = i[30];
  assign o[4093] = i[29];
  assign o[4092] = i[28];
  assign o[4091] = i[27];
  assign o[4090] = i[26];
  assign o[4089] = i[25];
  assign o[4088] = i[24];
  assign o[4087] = i[23];
  assign o[4086] = i[22];
  assign o[4085] = i[21];
  assign o[4084] = i[20];
  assign o[4083] = i[19];
  assign o[4082] = i[18];
  assign o[4081] = i[17];
  assign o[4080] = i[16];
  assign o[4079] = i[15];
  assign o[4078] = i[14];
  assign o[4077] = i[13];
  assign o[4076] = i[12];
  assign o[4075] = i[11];
  assign o[4074] = i[10];
  assign o[4073] = i[9];
  assign o[4072] = i[8];
  assign o[4071] = i[7];
  assign o[4070] = i[6];
  assign o[4069] = i[5];
  assign o[4068] = i[4];
  assign o[4067] = i[3];
  assign o[4066] = i[2];
  assign o[4065] = i[1];
  assign o[4064] = i[0];
  assign o[4063] = i[63];
  assign o[4062] = i[62];
  assign o[4061] = i[61];
  assign o[4060] = i[60];
  assign o[4059] = i[59];
  assign o[4058] = i[58];
  assign o[4057] = i[57];
  assign o[4056] = i[56];
  assign o[4055] = i[55];
  assign o[4054] = i[54];
  assign o[4053] = i[53];
  assign o[4052] = i[52];
  assign o[4051] = i[51];
  assign o[4050] = i[50];
  assign o[4049] = i[49];
  assign o[4048] = i[48];
  assign o[4047] = i[47];
  assign o[4046] = i[46];
  assign o[4045] = i[45];
  assign o[4044] = i[44];
  assign o[4043] = i[43];
  assign o[4042] = i[42];
  assign o[4041] = i[41];
  assign o[4040] = i[40];
  assign o[4039] = i[39];
  assign o[4038] = i[38];
  assign o[4037] = i[37];
  assign o[4036] = i[36];
  assign o[4035] = i[35];
  assign o[4034] = i[34];
  assign o[4033] = i[33];
  assign o[4032] = i[32];
  assign o[4031] = i[95];
  assign o[4030] = i[94];
  assign o[4029] = i[93];
  assign o[4028] = i[92];
  assign o[4027] = i[91];
  assign o[4026] = i[90];
  assign o[4025] = i[89];
  assign o[4024] = i[88];
  assign o[4023] = i[87];
  assign o[4022] = i[86];
  assign o[4021] = i[85];
  assign o[4020] = i[84];
  assign o[4019] = i[83];
  assign o[4018] = i[82];
  assign o[4017] = i[81];
  assign o[4016] = i[80];
  assign o[4015] = i[79];
  assign o[4014] = i[78];
  assign o[4013] = i[77];
  assign o[4012] = i[76];
  assign o[4011] = i[75];
  assign o[4010] = i[74];
  assign o[4009] = i[73];
  assign o[4008] = i[72];
  assign o[4007] = i[71];
  assign o[4006] = i[70];
  assign o[4005] = i[69];
  assign o[4004] = i[68];
  assign o[4003] = i[67];
  assign o[4002] = i[66];
  assign o[4001] = i[65];
  assign o[4000] = i[64];
  assign o[3999] = i[127];
  assign o[3998] = i[126];
  assign o[3997] = i[125];
  assign o[3996] = i[124];
  assign o[3995] = i[123];
  assign o[3994] = i[122];
  assign o[3993] = i[121];
  assign o[3992] = i[120];
  assign o[3991] = i[119];
  assign o[3990] = i[118];
  assign o[3989] = i[117];
  assign o[3988] = i[116];
  assign o[3987] = i[115];
  assign o[3986] = i[114];
  assign o[3985] = i[113];
  assign o[3984] = i[112];
  assign o[3983] = i[111];
  assign o[3982] = i[110];
  assign o[3981] = i[109];
  assign o[3980] = i[108];
  assign o[3979] = i[107];
  assign o[3978] = i[106];
  assign o[3977] = i[105];
  assign o[3976] = i[104];
  assign o[3975] = i[103];
  assign o[3974] = i[102];
  assign o[3973] = i[101];
  assign o[3972] = i[100];
  assign o[3971] = i[99];
  assign o[3970] = i[98];
  assign o[3969] = i[97];
  assign o[3968] = i[96];
  assign o[3967] = i[159];
  assign o[3966] = i[158];
  assign o[3965] = i[157];
  assign o[3964] = i[156];
  assign o[3963] = i[155];
  assign o[3962] = i[154];
  assign o[3961] = i[153];
  assign o[3960] = i[152];
  assign o[3959] = i[151];
  assign o[3958] = i[150];
  assign o[3957] = i[149];
  assign o[3956] = i[148];
  assign o[3955] = i[147];
  assign o[3954] = i[146];
  assign o[3953] = i[145];
  assign o[3952] = i[144];
  assign o[3951] = i[143];
  assign o[3950] = i[142];
  assign o[3949] = i[141];
  assign o[3948] = i[140];
  assign o[3947] = i[139];
  assign o[3946] = i[138];
  assign o[3945] = i[137];
  assign o[3944] = i[136];
  assign o[3943] = i[135];
  assign o[3942] = i[134];
  assign o[3941] = i[133];
  assign o[3940] = i[132];
  assign o[3939] = i[131];
  assign o[3938] = i[130];
  assign o[3937] = i[129];
  assign o[3936] = i[128];
  assign o[3935] = i[191];
  assign o[3934] = i[190];
  assign o[3933] = i[189];
  assign o[3932] = i[188];
  assign o[3931] = i[187];
  assign o[3930] = i[186];
  assign o[3929] = i[185];
  assign o[3928] = i[184];
  assign o[3927] = i[183];
  assign o[3926] = i[182];
  assign o[3925] = i[181];
  assign o[3924] = i[180];
  assign o[3923] = i[179];
  assign o[3922] = i[178];
  assign o[3921] = i[177];
  assign o[3920] = i[176];
  assign o[3919] = i[175];
  assign o[3918] = i[174];
  assign o[3917] = i[173];
  assign o[3916] = i[172];
  assign o[3915] = i[171];
  assign o[3914] = i[170];
  assign o[3913] = i[169];
  assign o[3912] = i[168];
  assign o[3911] = i[167];
  assign o[3910] = i[166];
  assign o[3909] = i[165];
  assign o[3908] = i[164];
  assign o[3907] = i[163];
  assign o[3906] = i[162];
  assign o[3905] = i[161];
  assign o[3904] = i[160];
  assign o[3903] = i[223];
  assign o[3902] = i[222];
  assign o[3901] = i[221];
  assign o[3900] = i[220];
  assign o[3899] = i[219];
  assign o[3898] = i[218];
  assign o[3897] = i[217];
  assign o[3896] = i[216];
  assign o[3895] = i[215];
  assign o[3894] = i[214];
  assign o[3893] = i[213];
  assign o[3892] = i[212];
  assign o[3891] = i[211];
  assign o[3890] = i[210];
  assign o[3889] = i[209];
  assign o[3888] = i[208];
  assign o[3887] = i[207];
  assign o[3886] = i[206];
  assign o[3885] = i[205];
  assign o[3884] = i[204];
  assign o[3883] = i[203];
  assign o[3882] = i[202];
  assign o[3881] = i[201];
  assign o[3880] = i[200];
  assign o[3879] = i[199];
  assign o[3878] = i[198];
  assign o[3877] = i[197];
  assign o[3876] = i[196];
  assign o[3875] = i[195];
  assign o[3874] = i[194];
  assign o[3873] = i[193];
  assign o[3872] = i[192];
  assign o[3871] = i[255];
  assign o[3870] = i[254];
  assign o[3869] = i[253];
  assign o[3868] = i[252];
  assign o[3867] = i[251];
  assign o[3866] = i[250];
  assign o[3865] = i[249];
  assign o[3864] = i[248];
  assign o[3863] = i[247];
  assign o[3862] = i[246];
  assign o[3861] = i[245];
  assign o[3860] = i[244];
  assign o[3859] = i[243];
  assign o[3858] = i[242];
  assign o[3857] = i[241];
  assign o[3856] = i[240];
  assign o[3855] = i[239];
  assign o[3854] = i[238];
  assign o[3853] = i[237];
  assign o[3852] = i[236];
  assign o[3851] = i[235];
  assign o[3850] = i[234];
  assign o[3849] = i[233];
  assign o[3848] = i[232];
  assign o[3847] = i[231];
  assign o[3846] = i[230];
  assign o[3845] = i[229];
  assign o[3844] = i[228];
  assign o[3843] = i[227];
  assign o[3842] = i[226];
  assign o[3841] = i[225];
  assign o[3840] = i[224];
  assign o[3839] = i[287];
  assign o[3838] = i[286];
  assign o[3837] = i[285];
  assign o[3836] = i[284];
  assign o[3835] = i[283];
  assign o[3834] = i[282];
  assign o[3833] = i[281];
  assign o[3832] = i[280];
  assign o[3831] = i[279];
  assign o[3830] = i[278];
  assign o[3829] = i[277];
  assign o[3828] = i[276];
  assign o[3827] = i[275];
  assign o[3826] = i[274];
  assign o[3825] = i[273];
  assign o[3824] = i[272];
  assign o[3823] = i[271];
  assign o[3822] = i[270];
  assign o[3821] = i[269];
  assign o[3820] = i[268];
  assign o[3819] = i[267];
  assign o[3818] = i[266];
  assign o[3817] = i[265];
  assign o[3816] = i[264];
  assign o[3815] = i[263];
  assign o[3814] = i[262];
  assign o[3813] = i[261];
  assign o[3812] = i[260];
  assign o[3811] = i[259];
  assign o[3810] = i[258];
  assign o[3809] = i[257];
  assign o[3808] = i[256];
  assign o[3807] = i[319];
  assign o[3806] = i[318];
  assign o[3805] = i[317];
  assign o[3804] = i[316];
  assign o[3803] = i[315];
  assign o[3802] = i[314];
  assign o[3801] = i[313];
  assign o[3800] = i[312];
  assign o[3799] = i[311];
  assign o[3798] = i[310];
  assign o[3797] = i[309];
  assign o[3796] = i[308];
  assign o[3795] = i[307];
  assign o[3794] = i[306];
  assign o[3793] = i[305];
  assign o[3792] = i[304];
  assign o[3791] = i[303];
  assign o[3790] = i[302];
  assign o[3789] = i[301];
  assign o[3788] = i[300];
  assign o[3787] = i[299];
  assign o[3786] = i[298];
  assign o[3785] = i[297];
  assign o[3784] = i[296];
  assign o[3783] = i[295];
  assign o[3782] = i[294];
  assign o[3781] = i[293];
  assign o[3780] = i[292];
  assign o[3779] = i[291];
  assign o[3778] = i[290];
  assign o[3777] = i[289];
  assign o[3776] = i[288];
  assign o[3775] = i[351];
  assign o[3774] = i[350];
  assign o[3773] = i[349];
  assign o[3772] = i[348];
  assign o[3771] = i[347];
  assign o[3770] = i[346];
  assign o[3769] = i[345];
  assign o[3768] = i[344];
  assign o[3767] = i[343];
  assign o[3766] = i[342];
  assign o[3765] = i[341];
  assign o[3764] = i[340];
  assign o[3763] = i[339];
  assign o[3762] = i[338];
  assign o[3761] = i[337];
  assign o[3760] = i[336];
  assign o[3759] = i[335];
  assign o[3758] = i[334];
  assign o[3757] = i[333];
  assign o[3756] = i[332];
  assign o[3755] = i[331];
  assign o[3754] = i[330];
  assign o[3753] = i[329];
  assign o[3752] = i[328];
  assign o[3751] = i[327];
  assign o[3750] = i[326];
  assign o[3749] = i[325];
  assign o[3748] = i[324];
  assign o[3747] = i[323];
  assign o[3746] = i[322];
  assign o[3745] = i[321];
  assign o[3744] = i[320];
  assign o[3743] = i[383];
  assign o[3742] = i[382];
  assign o[3741] = i[381];
  assign o[3740] = i[380];
  assign o[3739] = i[379];
  assign o[3738] = i[378];
  assign o[3737] = i[377];
  assign o[3736] = i[376];
  assign o[3735] = i[375];
  assign o[3734] = i[374];
  assign o[3733] = i[373];
  assign o[3732] = i[372];
  assign o[3731] = i[371];
  assign o[3730] = i[370];
  assign o[3729] = i[369];
  assign o[3728] = i[368];
  assign o[3727] = i[367];
  assign o[3726] = i[366];
  assign o[3725] = i[365];
  assign o[3724] = i[364];
  assign o[3723] = i[363];
  assign o[3722] = i[362];
  assign o[3721] = i[361];
  assign o[3720] = i[360];
  assign o[3719] = i[359];
  assign o[3718] = i[358];
  assign o[3717] = i[357];
  assign o[3716] = i[356];
  assign o[3715] = i[355];
  assign o[3714] = i[354];
  assign o[3713] = i[353];
  assign o[3712] = i[352];
  assign o[3711] = i[415];
  assign o[3710] = i[414];
  assign o[3709] = i[413];
  assign o[3708] = i[412];
  assign o[3707] = i[411];
  assign o[3706] = i[410];
  assign o[3705] = i[409];
  assign o[3704] = i[408];
  assign o[3703] = i[407];
  assign o[3702] = i[406];
  assign o[3701] = i[405];
  assign o[3700] = i[404];
  assign o[3699] = i[403];
  assign o[3698] = i[402];
  assign o[3697] = i[401];
  assign o[3696] = i[400];
  assign o[3695] = i[399];
  assign o[3694] = i[398];
  assign o[3693] = i[397];
  assign o[3692] = i[396];
  assign o[3691] = i[395];
  assign o[3690] = i[394];
  assign o[3689] = i[393];
  assign o[3688] = i[392];
  assign o[3687] = i[391];
  assign o[3686] = i[390];
  assign o[3685] = i[389];
  assign o[3684] = i[388];
  assign o[3683] = i[387];
  assign o[3682] = i[386];
  assign o[3681] = i[385];
  assign o[3680] = i[384];
  assign o[3679] = i[447];
  assign o[3678] = i[446];
  assign o[3677] = i[445];
  assign o[3676] = i[444];
  assign o[3675] = i[443];
  assign o[3674] = i[442];
  assign o[3673] = i[441];
  assign o[3672] = i[440];
  assign o[3671] = i[439];
  assign o[3670] = i[438];
  assign o[3669] = i[437];
  assign o[3668] = i[436];
  assign o[3667] = i[435];
  assign o[3666] = i[434];
  assign o[3665] = i[433];
  assign o[3664] = i[432];
  assign o[3663] = i[431];
  assign o[3662] = i[430];
  assign o[3661] = i[429];
  assign o[3660] = i[428];
  assign o[3659] = i[427];
  assign o[3658] = i[426];
  assign o[3657] = i[425];
  assign o[3656] = i[424];
  assign o[3655] = i[423];
  assign o[3654] = i[422];
  assign o[3653] = i[421];
  assign o[3652] = i[420];
  assign o[3651] = i[419];
  assign o[3650] = i[418];
  assign o[3649] = i[417];
  assign o[3648] = i[416];
  assign o[3647] = i[479];
  assign o[3646] = i[478];
  assign o[3645] = i[477];
  assign o[3644] = i[476];
  assign o[3643] = i[475];
  assign o[3642] = i[474];
  assign o[3641] = i[473];
  assign o[3640] = i[472];
  assign o[3639] = i[471];
  assign o[3638] = i[470];
  assign o[3637] = i[469];
  assign o[3636] = i[468];
  assign o[3635] = i[467];
  assign o[3634] = i[466];
  assign o[3633] = i[465];
  assign o[3632] = i[464];
  assign o[3631] = i[463];
  assign o[3630] = i[462];
  assign o[3629] = i[461];
  assign o[3628] = i[460];
  assign o[3627] = i[459];
  assign o[3626] = i[458];
  assign o[3625] = i[457];
  assign o[3624] = i[456];
  assign o[3623] = i[455];
  assign o[3622] = i[454];
  assign o[3621] = i[453];
  assign o[3620] = i[452];
  assign o[3619] = i[451];
  assign o[3618] = i[450];
  assign o[3617] = i[449];
  assign o[3616] = i[448];
  assign o[3615] = i[511];
  assign o[3614] = i[510];
  assign o[3613] = i[509];
  assign o[3612] = i[508];
  assign o[3611] = i[507];
  assign o[3610] = i[506];
  assign o[3609] = i[505];
  assign o[3608] = i[504];
  assign o[3607] = i[503];
  assign o[3606] = i[502];
  assign o[3605] = i[501];
  assign o[3604] = i[500];
  assign o[3603] = i[499];
  assign o[3602] = i[498];
  assign o[3601] = i[497];
  assign o[3600] = i[496];
  assign o[3599] = i[495];
  assign o[3598] = i[494];
  assign o[3597] = i[493];
  assign o[3596] = i[492];
  assign o[3595] = i[491];
  assign o[3594] = i[490];
  assign o[3593] = i[489];
  assign o[3592] = i[488];
  assign o[3591] = i[487];
  assign o[3590] = i[486];
  assign o[3589] = i[485];
  assign o[3588] = i[484];
  assign o[3587] = i[483];
  assign o[3586] = i[482];
  assign o[3585] = i[481];
  assign o[3584] = i[480];
  assign o[3583] = i[543];
  assign o[3582] = i[542];
  assign o[3581] = i[541];
  assign o[3580] = i[540];
  assign o[3579] = i[539];
  assign o[3578] = i[538];
  assign o[3577] = i[537];
  assign o[3576] = i[536];
  assign o[3575] = i[535];
  assign o[3574] = i[534];
  assign o[3573] = i[533];
  assign o[3572] = i[532];
  assign o[3571] = i[531];
  assign o[3570] = i[530];
  assign o[3569] = i[529];
  assign o[3568] = i[528];
  assign o[3567] = i[527];
  assign o[3566] = i[526];
  assign o[3565] = i[525];
  assign o[3564] = i[524];
  assign o[3563] = i[523];
  assign o[3562] = i[522];
  assign o[3561] = i[521];
  assign o[3560] = i[520];
  assign o[3559] = i[519];
  assign o[3558] = i[518];
  assign o[3557] = i[517];
  assign o[3556] = i[516];
  assign o[3555] = i[515];
  assign o[3554] = i[514];
  assign o[3553] = i[513];
  assign o[3552] = i[512];
  assign o[3551] = i[575];
  assign o[3550] = i[574];
  assign o[3549] = i[573];
  assign o[3548] = i[572];
  assign o[3547] = i[571];
  assign o[3546] = i[570];
  assign o[3545] = i[569];
  assign o[3544] = i[568];
  assign o[3543] = i[567];
  assign o[3542] = i[566];
  assign o[3541] = i[565];
  assign o[3540] = i[564];
  assign o[3539] = i[563];
  assign o[3538] = i[562];
  assign o[3537] = i[561];
  assign o[3536] = i[560];
  assign o[3535] = i[559];
  assign o[3534] = i[558];
  assign o[3533] = i[557];
  assign o[3532] = i[556];
  assign o[3531] = i[555];
  assign o[3530] = i[554];
  assign o[3529] = i[553];
  assign o[3528] = i[552];
  assign o[3527] = i[551];
  assign o[3526] = i[550];
  assign o[3525] = i[549];
  assign o[3524] = i[548];
  assign o[3523] = i[547];
  assign o[3522] = i[546];
  assign o[3521] = i[545];
  assign o[3520] = i[544];
  assign o[3519] = i[607];
  assign o[3518] = i[606];
  assign o[3517] = i[605];
  assign o[3516] = i[604];
  assign o[3515] = i[603];
  assign o[3514] = i[602];
  assign o[3513] = i[601];
  assign o[3512] = i[600];
  assign o[3511] = i[599];
  assign o[3510] = i[598];
  assign o[3509] = i[597];
  assign o[3508] = i[596];
  assign o[3507] = i[595];
  assign o[3506] = i[594];
  assign o[3505] = i[593];
  assign o[3504] = i[592];
  assign o[3503] = i[591];
  assign o[3502] = i[590];
  assign o[3501] = i[589];
  assign o[3500] = i[588];
  assign o[3499] = i[587];
  assign o[3498] = i[586];
  assign o[3497] = i[585];
  assign o[3496] = i[584];
  assign o[3495] = i[583];
  assign o[3494] = i[582];
  assign o[3493] = i[581];
  assign o[3492] = i[580];
  assign o[3491] = i[579];
  assign o[3490] = i[578];
  assign o[3489] = i[577];
  assign o[3488] = i[576];
  assign o[3487] = i[639];
  assign o[3486] = i[638];
  assign o[3485] = i[637];
  assign o[3484] = i[636];
  assign o[3483] = i[635];
  assign o[3482] = i[634];
  assign o[3481] = i[633];
  assign o[3480] = i[632];
  assign o[3479] = i[631];
  assign o[3478] = i[630];
  assign o[3477] = i[629];
  assign o[3476] = i[628];
  assign o[3475] = i[627];
  assign o[3474] = i[626];
  assign o[3473] = i[625];
  assign o[3472] = i[624];
  assign o[3471] = i[623];
  assign o[3470] = i[622];
  assign o[3469] = i[621];
  assign o[3468] = i[620];
  assign o[3467] = i[619];
  assign o[3466] = i[618];
  assign o[3465] = i[617];
  assign o[3464] = i[616];
  assign o[3463] = i[615];
  assign o[3462] = i[614];
  assign o[3461] = i[613];
  assign o[3460] = i[612];
  assign o[3459] = i[611];
  assign o[3458] = i[610];
  assign o[3457] = i[609];
  assign o[3456] = i[608];
  assign o[3455] = i[671];
  assign o[3454] = i[670];
  assign o[3453] = i[669];
  assign o[3452] = i[668];
  assign o[3451] = i[667];
  assign o[3450] = i[666];
  assign o[3449] = i[665];
  assign o[3448] = i[664];
  assign o[3447] = i[663];
  assign o[3446] = i[662];
  assign o[3445] = i[661];
  assign o[3444] = i[660];
  assign o[3443] = i[659];
  assign o[3442] = i[658];
  assign o[3441] = i[657];
  assign o[3440] = i[656];
  assign o[3439] = i[655];
  assign o[3438] = i[654];
  assign o[3437] = i[653];
  assign o[3436] = i[652];
  assign o[3435] = i[651];
  assign o[3434] = i[650];
  assign o[3433] = i[649];
  assign o[3432] = i[648];
  assign o[3431] = i[647];
  assign o[3430] = i[646];
  assign o[3429] = i[645];
  assign o[3428] = i[644];
  assign o[3427] = i[643];
  assign o[3426] = i[642];
  assign o[3425] = i[641];
  assign o[3424] = i[640];
  assign o[3423] = i[703];
  assign o[3422] = i[702];
  assign o[3421] = i[701];
  assign o[3420] = i[700];
  assign o[3419] = i[699];
  assign o[3418] = i[698];
  assign o[3417] = i[697];
  assign o[3416] = i[696];
  assign o[3415] = i[695];
  assign o[3414] = i[694];
  assign o[3413] = i[693];
  assign o[3412] = i[692];
  assign o[3411] = i[691];
  assign o[3410] = i[690];
  assign o[3409] = i[689];
  assign o[3408] = i[688];
  assign o[3407] = i[687];
  assign o[3406] = i[686];
  assign o[3405] = i[685];
  assign o[3404] = i[684];
  assign o[3403] = i[683];
  assign o[3402] = i[682];
  assign o[3401] = i[681];
  assign o[3400] = i[680];
  assign o[3399] = i[679];
  assign o[3398] = i[678];
  assign o[3397] = i[677];
  assign o[3396] = i[676];
  assign o[3395] = i[675];
  assign o[3394] = i[674];
  assign o[3393] = i[673];
  assign o[3392] = i[672];
  assign o[3391] = i[735];
  assign o[3390] = i[734];
  assign o[3389] = i[733];
  assign o[3388] = i[732];
  assign o[3387] = i[731];
  assign o[3386] = i[730];
  assign o[3385] = i[729];
  assign o[3384] = i[728];
  assign o[3383] = i[727];
  assign o[3382] = i[726];
  assign o[3381] = i[725];
  assign o[3380] = i[724];
  assign o[3379] = i[723];
  assign o[3378] = i[722];
  assign o[3377] = i[721];
  assign o[3376] = i[720];
  assign o[3375] = i[719];
  assign o[3374] = i[718];
  assign o[3373] = i[717];
  assign o[3372] = i[716];
  assign o[3371] = i[715];
  assign o[3370] = i[714];
  assign o[3369] = i[713];
  assign o[3368] = i[712];
  assign o[3367] = i[711];
  assign o[3366] = i[710];
  assign o[3365] = i[709];
  assign o[3364] = i[708];
  assign o[3363] = i[707];
  assign o[3362] = i[706];
  assign o[3361] = i[705];
  assign o[3360] = i[704];
  assign o[3359] = i[767];
  assign o[3358] = i[766];
  assign o[3357] = i[765];
  assign o[3356] = i[764];
  assign o[3355] = i[763];
  assign o[3354] = i[762];
  assign o[3353] = i[761];
  assign o[3352] = i[760];
  assign o[3351] = i[759];
  assign o[3350] = i[758];
  assign o[3349] = i[757];
  assign o[3348] = i[756];
  assign o[3347] = i[755];
  assign o[3346] = i[754];
  assign o[3345] = i[753];
  assign o[3344] = i[752];
  assign o[3343] = i[751];
  assign o[3342] = i[750];
  assign o[3341] = i[749];
  assign o[3340] = i[748];
  assign o[3339] = i[747];
  assign o[3338] = i[746];
  assign o[3337] = i[745];
  assign o[3336] = i[744];
  assign o[3335] = i[743];
  assign o[3334] = i[742];
  assign o[3333] = i[741];
  assign o[3332] = i[740];
  assign o[3331] = i[739];
  assign o[3330] = i[738];
  assign o[3329] = i[737];
  assign o[3328] = i[736];
  assign o[3327] = i[799];
  assign o[3326] = i[798];
  assign o[3325] = i[797];
  assign o[3324] = i[796];
  assign o[3323] = i[795];
  assign o[3322] = i[794];
  assign o[3321] = i[793];
  assign o[3320] = i[792];
  assign o[3319] = i[791];
  assign o[3318] = i[790];
  assign o[3317] = i[789];
  assign o[3316] = i[788];
  assign o[3315] = i[787];
  assign o[3314] = i[786];
  assign o[3313] = i[785];
  assign o[3312] = i[784];
  assign o[3311] = i[783];
  assign o[3310] = i[782];
  assign o[3309] = i[781];
  assign o[3308] = i[780];
  assign o[3307] = i[779];
  assign o[3306] = i[778];
  assign o[3305] = i[777];
  assign o[3304] = i[776];
  assign o[3303] = i[775];
  assign o[3302] = i[774];
  assign o[3301] = i[773];
  assign o[3300] = i[772];
  assign o[3299] = i[771];
  assign o[3298] = i[770];
  assign o[3297] = i[769];
  assign o[3296] = i[768];
  assign o[3295] = i[831];
  assign o[3294] = i[830];
  assign o[3293] = i[829];
  assign o[3292] = i[828];
  assign o[3291] = i[827];
  assign o[3290] = i[826];
  assign o[3289] = i[825];
  assign o[3288] = i[824];
  assign o[3287] = i[823];
  assign o[3286] = i[822];
  assign o[3285] = i[821];
  assign o[3284] = i[820];
  assign o[3283] = i[819];
  assign o[3282] = i[818];
  assign o[3281] = i[817];
  assign o[3280] = i[816];
  assign o[3279] = i[815];
  assign o[3278] = i[814];
  assign o[3277] = i[813];
  assign o[3276] = i[812];
  assign o[3275] = i[811];
  assign o[3274] = i[810];
  assign o[3273] = i[809];
  assign o[3272] = i[808];
  assign o[3271] = i[807];
  assign o[3270] = i[806];
  assign o[3269] = i[805];
  assign o[3268] = i[804];
  assign o[3267] = i[803];
  assign o[3266] = i[802];
  assign o[3265] = i[801];
  assign o[3264] = i[800];
  assign o[3263] = i[863];
  assign o[3262] = i[862];
  assign o[3261] = i[861];
  assign o[3260] = i[860];
  assign o[3259] = i[859];
  assign o[3258] = i[858];
  assign o[3257] = i[857];
  assign o[3256] = i[856];
  assign o[3255] = i[855];
  assign o[3254] = i[854];
  assign o[3253] = i[853];
  assign o[3252] = i[852];
  assign o[3251] = i[851];
  assign o[3250] = i[850];
  assign o[3249] = i[849];
  assign o[3248] = i[848];
  assign o[3247] = i[847];
  assign o[3246] = i[846];
  assign o[3245] = i[845];
  assign o[3244] = i[844];
  assign o[3243] = i[843];
  assign o[3242] = i[842];
  assign o[3241] = i[841];
  assign o[3240] = i[840];
  assign o[3239] = i[839];
  assign o[3238] = i[838];
  assign o[3237] = i[837];
  assign o[3236] = i[836];
  assign o[3235] = i[835];
  assign o[3234] = i[834];
  assign o[3233] = i[833];
  assign o[3232] = i[832];
  assign o[3231] = i[895];
  assign o[3230] = i[894];
  assign o[3229] = i[893];
  assign o[3228] = i[892];
  assign o[3227] = i[891];
  assign o[3226] = i[890];
  assign o[3225] = i[889];
  assign o[3224] = i[888];
  assign o[3223] = i[887];
  assign o[3222] = i[886];
  assign o[3221] = i[885];
  assign o[3220] = i[884];
  assign o[3219] = i[883];
  assign o[3218] = i[882];
  assign o[3217] = i[881];
  assign o[3216] = i[880];
  assign o[3215] = i[879];
  assign o[3214] = i[878];
  assign o[3213] = i[877];
  assign o[3212] = i[876];
  assign o[3211] = i[875];
  assign o[3210] = i[874];
  assign o[3209] = i[873];
  assign o[3208] = i[872];
  assign o[3207] = i[871];
  assign o[3206] = i[870];
  assign o[3205] = i[869];
  assign o[3204] = i[868];
  assign o[3203] = i[867];
  assign o[3202] = i[866];
  assign o[3201] = i[865];
  assign o[3200] = i[864];
  assign o[3199] = i[927];
  assign o[3198] = i[926];
  assign o[3197] = i[925];
  assign o[3196] = i[924];
  assign o[3195] = i[923];
  assign o[3194] = i[922];
  assign o[3193] = i[921];
  assign o[3192] = i[920];
  assign o[3191] = i[919];
  assign o[3190] = i[918];
  assign o[3189] = i[917];
  assign o[3188] = i[916];
  assign o[3187] = i[915];
  assign o[3186] = i[914];
  assign o[3185] = i[913];
  assign o[3184] = i[912];
  assign o[3183] = i[911];
  assign o[3182] = i[910];
  assign o[3181] = i[909];
  assign o[3180] = i[908];
  assign o[3179] = i[907];
  assign o[3178] = i[906];
  assign o[3177] = i[905];
  assign o[3176] = i[904];
  assign o[3175] = i[903];
  assign o[3174] = i[902];
  assign o[3173] = i[901];
  assign o[3172] = i[900];
  assign o[3171] = i[899];
  assign o[3170] = i[898];
  assign o[3169] = i[897];
  assign o[3168] = i[896];
  assign o[3167] = i[959];
  assign o[3166] = i[958];
  assign o[3165] = i[957];
  assign o[3164] = i[956];
  assign o[3163] = i[955];
  assign o[3162] = i[954];
  assign o[3161] = i[953];
  assign o[3160] = i[952];
  assign o[3159] = i[951];
  assign o[3158] = i[950];
  assign o[3157] = i[949];
  assign o[3156] = i[948];
  assign o[3155] = i[947];
  assign o[3154] = i[946];
  assign o[3153] = i[945];
  assign o[3152] = i[944];
  assign o[3151] = i[943];
  assign o[3150] = i[942];
  assign o[3149] = i[941];
  assign o[3148] = i[940];
  assign o[3147] = i[939];
  assign o[3146] = i[938];
  assign o[3145] = i[937];
  assign o[3144] = i[936];
  assign o[3143] = i[935];
  assign o[3142] = i[934];
  assign o[3141] = i[933];
  assign o[3140] = i[932];
  assign o[3139] = i[931];
  assign o[3138] = i[930];
  assign o[3137] = i[929];
  assign o[3136] = i[928];
  assign o[3135] = i[991];
  assign o[3134] = i[990];
  assign o[3133] = i[989];
  assign o[3132] = i[988];
  assign o[3131] = i[987];
  assign o[3130] = i[986];
  assign o[3129] = i[985];
  assign o[3128] = i[984];
  assign o[3127] = i[983];
  assign o[3126] = i[982];
  assign o[3125] = i[981];
  assign o[3124] = i[980];
  assign o[3123] = i[979];
  assign o[3122] = i[978];
  assign o[3121] = i[977];
  assign o[3120] = i[976];
  assign o[3119] = i[975];
  assign o[3118] = i[974];
  assign o[3117] = i[973];
  assign o[3116] = i[972];
  assign o[3115] = i[971];
  assign o[3114] = i[970];
  assign o[3113] = i[969];
  assign o[3112] = i[968];
  assign o[3111] = i[967];
  assign o[3110] = i[966];
  assign o[3109] = i[965];
  assign o[3108] = i[964];
  assign o[3107] = i[963];
  assign o[3106] = i[962];
  assign o[3105] = i[961];
  assign o[3104] = i[960];
  assign o[3103] = i[1023];
  assign o[3102] = i[1022];
  assign o[3101] = i[1021];
  assign o[3100] = i[1020];
  assign o[3099] = i[1019];
  assign o[3098] = i[1018];
  assign o[3097] = i[1017];
  assign o[3096] = i[1016];
  assign o[3095] = i[1015];
  assign o[3094] = i[1014];
  assign o[3093] = i[1013];
  assign o[3092] = i[1012];
  assign o[3091] = i[1011];
  assign o[3090] = i[1010];
  assign o[3089] = i[1009];
  assign o[3088] = i[1008];
  assign o[3087] = i[1007];
  assign o[3086] = i[1006];
  assign o[3085] = i[1005];
  assign o[3084] = i[1004];
  assign o[3083] = i[1003];
  assign o[3082] = i[1002];
  assign o[3081] = i[1001];
  assign o[3080] = i[1000];
  assign o[3079] = i[999];
  assign o[3078] = i[998];
  assign o[3077] = i[997];
  assign o[3076] = i[996];
  assign o[3075] = i[995];
  assign o[3074] = i[994];
  assign o[3073] = i[993];
  assign o[3072] = i[992];
  assign o[3071] = i[1055];
  assign o[3070] = i[1054];
  assign o[3069] = i[1053];
  assign o[3068] = i[1052];
  assign o[3067] = i[1051];
  assign o[3066] = i[1050];
  assign o[3065] = i[1049];
  assign o[3064] = i[1048];
  assign o[3063] = i[1047];
  assign o[3062] = i[1046];
  assign o[3061] = i[1045];
  assign o[3060] = i[1044];
  assign o[3059] = i[1043];
  assign o[3058] = i[1042];
  assign o[3057] = i[1041];
  assign o[3056] = i[1040];
  assign o[3055] = i[1039];
  assign o[3054] = i[1038];
  assign o[3053] = i[1037];
  assign o[3052] = i[1036];
  assign o[3051] = i[1035];
  assign o[3050] = i[1034];
  assign o[3049] = i[1033];
  assign o[3048] = i[1032];
  assign o[3047] = i[1031];
  assign o[3046] = i[1030];
  assign o[3045] = i[1029];
  assign o[3044] = i[1028];
  assign o[3043] = i[1027];
  assign o[3042] = i[1026];
  assign o[3041] = i[1025];
  assign o[3040] = i[1024];
  assign o[3039] = i[1087];
  assign o[3038] = i[1086];
  assign o[3037] = i[1085];
  assign o[3036] = i[1084];
  assign o[3035] = i[1083];
  assign o[3034] = i[1082];
  assign o[3033] = i[1081];
  assign o[3032] = i[1080];
  assign o[3031] = i[1079];
  assign o[3030] = i[1078];
  assign o[3029] = i[1077];
  assign o[3028] = i[1076];
  assign o[3027] = i[1075];
  assign o[3026] = i[1074];
  assign o[3025] = i[1073];
  assign o[3024] = i[1072];
  assign o[3023] = i[1071];
  assign o[3022] = i[1070];
  assign o[3021] = i[1069];
  assign o[3020] = i[1068];
  assign o[3019] = i[1067];
  assign o[3018] = i[1066];
  assign o[3017] = i[1065];
  assign o[3016] = i[1064];
  assign o[3015] = i[1063];
  assign o[3014] = i[1062];
  assign o[3013] = i[1061];
  assign o[3012] = i[1060];
  assign o[3011] = i[1059];
  assign o[3010] = i[1058];
  assign o[3009] = i[1057];
  assign o[3008] = i[1056];
  assign o[3007] = i[1119];
  assign o[3006] = i[1118];
  assign o[3005] = i[1117];
  assign o[3004] = i[1116];
  assign o[3003] = i[1115];
  assign o[3002] = i[1114];
  assign o[3001] = i[1113];
  assign o[3000] = i[1112];
  assign o[2999] = i[1111];
  assign o[2998] = i[1110];
  assign o[2997] = i[1109];
  assign o[2996] = i[1108];
  assign o[2995] = i[1107];
  assign o[2994] = i[1106];
  assign o[2993] = i[1105];
  assign o[2992] = i[1104];
  assign o[2991] = i[1103];
  assign o[2990] = i[1102];
  assign o[2989] = i[1101];
  assign o[2988] = i[1100];
  assign o[2987] = i[1099];
  assign o[2986] = i[1098];
  assign o[2985] = i[1097];
  assign o[2984] = i[1096];
  assign o[2983] = i[1095];
  assign o[2982] = i[1094];
  assign o[2981] = i[1093];
  assign o[2980] = i[1092];
  assign o[2979] = i[1091];
  assign o[2978] = i[1090];
  assign o[2977] = i[1089];
  assign o[2976] = i[1088];
  assign o[2975] = i[1151];
  assign o[2974] = i[1150];
  assign o[2973] = i[1149];
  assign o[2972] = i[1148];
  assign o[2971] = i[1147];
  assign o[2970] = i[1146];
  assign o[2969] = i[1145];
  assign o[2968] = i[1144];
  assign o[2967] = i[1143];
  assign o[2966] = i[1142];
  assign o[2965] = i[1141];
  assign o[2964] = i[1140];
  assign o[2963] = i[1139];
  assign o[2962] = i[1138];
  assign o[2961] = i[1137];
  assign o[2960] = i[1136];
  assign o[2959] = i[1135];
  assign o[2958] = i[1134];
  assign o[2957] = i[1133];
  assign o[2956] = i[1132];
  assign o[2955] = i[1131];
  assign o[2954] = i[1130];
  assign o[2953] = i[1129];
  assign o[2952] = i[1128];
  assign o[2951] = i[1127];
  assign o[2950] = i[1126];
  assign o[2949] = i[1125];
  assign o[2948] = i[1124];
  assign o[2947] = i[1123];
  assign o[2946] = i[1122];
  assign o[2945] = i[1121];
  assign o[2944] = i[1120];
  assign o[2943] = i[1183];
  assign o[2942] = i[1182];
  assign o[2941] = i[1181];
  assign o[2940] = i[1180];
  assign o[2939] = i[1179];
  assign o[2938] = i[1178];
  assign o[2937] = i[1177];
  assign o[2936] = i[1176];
  assign o[2935] = i[1175];
  assign o[2934] = i[1174];
  assign o[2933] = i[1173];
  assign o[2932] = i[1172];
  assign o[2931] = i[1171];
  assign o[2930] = i[1170];
  assign o[2929] = i[1169];
  assign o[2928] = i[1168];
  assign o[2927] = i[1167];
  assign o[2926] = i[1166];
  assign o[2925] = i[1165];
  assign o[2924] = i[1164];
  assign o[2923] = i[1163];
  assign o[2922] = i[1162];
  assign o[2921] = i[1161];
  assign o[2920] = i[1160];
  assign o[2919] = i[1159];
  assign o[2918] = i[1158];
  assign o[2917] = i[1157];
  assign o[2916] = i[1156];
  assign o[2915] = i[1155];
  assign o[2914] = i[1154];
  assign o[2913] = i[1153];
  assign o[2912] = i[1152];
  assign o[2911] = i[1215];
  assign o[2910] = i[1214];
  assign o[2909] = i[1213];
  assign o[2908] = i[1212];
  assign o[2907] = i[1211];
  assign o[2906] = i[1210];
  assign o[2905] = i[1209];
  assign o[2904] = i[1208];
  assign o[2903] = i[1207];
  assign o[2902] = i[1206];
  assign o[2901] = i[1205];
  assign o[2900] = i[1204];
  assign o[2899] = i[1203];
  assign o[2898] = i[1202];
  assign o[2897] = i[1201];
  assign o[2896] = i[1200];
  assign o[2895] = i[1199];
  assign o[2894] = i[1198];
  assign o[2893] = i[1197];
  assign o[2892] = i[1196];
  assign o[2891] = i[1195];
  assign o[2890] = i[1194];
  assign o[2889] = i[1193];
  assign o[2888] = i[1192];
  assign o[2887] = i[1191];
  assign o[2886] = i[1190];
  assign o[2885] = i[1189];
  assign o[2884] = i[1188];
  assign o[2883] = i[1187];
  assign o[2882] = i[1186];
  assign o[2881] = i[1185];
  assign o[2880] = i[1184];
  assign o[2879] = i[1247];
  assign o[2878] = i[1246];
  assign o[2877] = i[1245];
  assign o[2876] = i[1244];
  assign o[2875] = i[1243];
  assign o[2874] = i[1242];
  assign o[2873] = i[1241];
  assign o[2872] = i[1240];
  assign o[2871] = i[1239];
  assign o[2870] = i[1238];
  assign o[2869] = i[1237];
  assign o[2868] = i[1236];
  assign o[2867] = i[1235];
  assign o[2866] = i[1234];
  assign o[2865] = i[1233];
  assign o[2864] = i[1232];
  assign o[2863] = i[1231];
  assign o[2862] = i[1230];
  assign o[2861] = i[1229];
  assign o[2860] = i[1228];
  assign o[2859] = i[1227];
  assign o[2858] = i[1226];
  assign o[2857] = i[1225];
  assign o[2856] = i[1224];
  assign o[2855] = i[1223];
  assign o[2854] = i[1222];
  assign o[2853] = i[1221];
  assign o[2852] = i[1220];
  assign o[2851] = i[1219];
  assign o[2850] = i[1218];
  assign o[2849] = i[1217];
  assign o[2848] = i[1216];
  assign o[2847] = i[1279];
  assign o[2846] = i[1278];
  assign o[2845] = i[1277];
  assign o[2844] = i[1276];
  assign o[2843] = i[1275];
  assign o[2842] = i[1274];
  assign o[2841] = i[1273];
  assign o[2840] = i[1272];
  assign o[2839] = i[1271];
  assign o[2838] = i[1270];
  assign o[2837] = i[1269];
  assign o[2836] = i[1268];
  assign o[2835] = i[1267];
  assign o[2834] = i[1266];
  assign o[2833] = i[1265];
  assign o[2832] = i[1264];
  assign o[2831] = i[1263];
  assign o[2830] = i[1262];
  assign o[2829] = i[1261];
  assign o[2828] = i[1260];
  assign o[2827] = i[1259];
  assign o[2826] = i[1258];
  assign o[2825] = i[1257];
  assign o[2824] = i[1256];
  assign o[2823] = i[1255];
  assign o[2822] = i[1254];
  assign o[2821] = i[1253];
  assign o[2820] = i[1252];
  assign o[2819] = i[1251];
  assign o[2818] = i[1250];
  assign o[2817] = i[1249];
  assign o[2816] = i[1248];
  assign o[2815] = i[1311];
  assign o[2814] = i[1310];
  assign o[2813] = i[1309];
  assign o[2812] = i[1308];
  assign o[2811] = i[1307];
  assign o[2810] = i[1306];
  assign o[2809] = i[1305];
  assign o[2808] = i[1304];
  assign o[2807] = i[1303];
  assign o[2806] = i[1302];
  assign o[2805] = i[1301];
  assign o[2804] = i[1300];
  assign o[2803] = i[1299];
  assign o[2802] = i[1298];
  assign o[2801] = i[1297];
  assign o[2800] = i[1296];
  assign o[2799] = i[1295];
  assign o[2798] = i[1294];
  assign o[2797] = i[1293];
  assign o[2796] = i[1292];
  assign o[2795] = i[1291];
  assign o[2794] = i[1290];
  assign o[2793] = i[1289];
  assign o[2792] = i[1288];
  assign o[2791] = i[1287];
  assign o[2790] = i[1286];
  assign o[2789] = i[1285];
  assign o[2788] = i[1284];
  assign o[2787] = i[1283];
  assign o[2786] = i[1282];
  assign o[2785] = i[1281];
  assign o[2784] = i[1280];
  assign o[2783] = i[1343];
  assign o[2782] = i[1342];
  assign o[2781] = i[1341];
  assign o[2780] = i[1340];
  assign o[2779] = i[1339];
  assign o[2778] = i[1338];
  assign o[2777] = i[1337];
  assign o[2776] = i[1336];
  assign o[2775] = i[1335];
  assign o[2774] = i[1334];
  assign o[2773] = i[1333];
  assign o[2772] = i[1332];
  assign o[2771] = i[1331];
  assign o[2770] = i[1330];
  assign o[2769] = i[1329];
  assign o[2768] = i[1328];
  assign o[2767] = i[1327];
  assign o[2766] = i[1326];
  assign o[2765] = i[1325];
  assign o[2764] = i[1324];
  assign o[2763] = i[1323];
  assign o[2762] = i[1322];
  assign o[2761] = i[1321];
  assign o[2760] = i[1320];
  assign o[2759] = i[1319];
  assign o[2758] = i[1318];
  assign o[2757] = i[1317];
  assign o[2756] = i[1316];
  assign o[2755] = i[1315];
  assign o[2754] = i[1314];
  assign o[2753] = i[1313];
  assign o[2752] = i[1312];
  assign o[2751] = i[1375];
  assign o[2750] = i[1374];
  assign o[2749] = i[1373];
  assign o[2748] = i[1372];
  assign o[2747] = i[1371];
  assign o[2746] = i[1370];
  assign o[2745] = i[1369];
  assign o[2744] = i[1368];
  assign o[2743] = i[1367];
  assign o[2742] = i[1366];
  assign o[2741] = i[1365];
  assign o[2740] = i[1364];
  assign o[2739] = i[1363];
  assign o[2738] = i[1362];
  assign o[2737] = i[1361];
  assign o[2736] = i[1360];
  assign o[2735] = i[1359];
  assign o[2734] = i[1358];
  assign o[2733] = i[1357];
  assign o[2732] = i[1356];
  assign o[2731] = i[1355];
  assign o[2730] = i[1354];
  assign o[2729] = i[1353];
  assign o[2728] = i[1352];
  assign o[2727] = i[1351];
  assign o[2726] = i[1350];
  assign o[2725] = i[1349];
  assign o[2724] = i[1348];
  assign o[2723] = i[1347];
  assign o[2722] = i[1346];
  assign o[2721] = i[1345];
  assign o[2720] = i[1344];
  assign o[2719] = i[1407];
  assign o[2718] = i[1406];
  assign o[2717] = i[1405];
  assign o[2716] = i[1404];
  assign o[2715] = i[1403];
  assign o[2714] = i[1402];
  assign o[2713] = i[1401];
  assign o[2712] = i[1400];
  assign o[2711] = i[1399];
  assign o[2710] = i[1398];
  assign o[2709] = i[1397];
  assign o[2708] = i[1396];
  assign o[2707] = i[1395];
  assign o[2706] = i[1394];
  assign o[2705] = i[1393];
  assign o[2704] = i[1392];
  assign o[2703] = i[1391];
  assign o[2702] = i[1390];
  assign o[2701] = i[1389];
  assign o[2700] = i[1388];
  assign o[2699] = i[1387];
  assign o[2698] = i[1386];
  assign o[2697] = i[1385];
  assign o[2696] = i[1384];
  assign o[2695] = i[1383];
  assign o[2694] = i[1382];
  assign o[2693] = i[1381];
  assign o[2692] = i[1380];
  assign o[2691] = i[1379];
  assign o[2690] = i[1378];
  assign o[2689] = i[1377];
  assign o[2688] = i[1376];
  assign o[2687] = i[1439];
  assign o[2686] = i[1438];
  assign o[2685] = i[1437];
  assign o[2684] = i[1436];
  assign o[2683] = i[1435];
  assign o[2682] = i[1434];
  assign o[2681] = i[1433];
  assign o[2680] = i[1432];
  assign o[2679] = i[1431];
  assign o[2678] = i[1430];
  assign o[2677] = i[1429];
  assign o[2676] = i[1428];
  assign o[2675] = i[1427];
  assign o[2674] = i[1426];
  assign o[2673] = i[1425];
  assign o[2672] = i[1424];
  assign o[2671] = i[1423];
  assign o[2670] = i[1422];
  assign o[2669] = i[1421];
  assign o[2668] = i[1420];
  assign o[2667] = i[1419];
  assign o[2666] = i[1418];
  assign o[2665] = i[1417];
  assign o[2664] = i[1416];
  assign o[2663] = i[1415];
  assign o[2662] = i[1414];
  assign o[2661] = i[1413];
  assign o[2660] = i[1412];
  assign o[2659] = i[1411];
  assign o[2658] = i[1410];
  assign o[2657] = i[1409];
  assign o[2656] = i[1408];
  assign o[2655] = i[1471];
  assign o[2654] = i[1470];
  assign o[2653] = i[1469];
  assign o[2652] = i[1468];
  assign o[2651] = i[1467];
  assign o[2650] = i[1466];
  assign o[2649] = i[1465];
  assign o[2648] = i[1464];
  assign o[2647] = i[1463];
  assign o[2646] = i[1462];
  assign o[2645] = i[1461];
  assign o[2644] = i[1460];
  assign o[2643] = i[1459];
  assign o[2642] = i[1458];
  assign o[2641] = i[1457];
  assign o[2640] = i[1456];
  assign o[2639] = i[1455];
  assign o[2638] = i[1454];
  assign o[2637] = i[1453];
  assign o[2636] = i[1452];
  assign o[2635] = i[1451];
  assign o[2634] = i[1450];
  assign o[2633] = i[1449];
  assign o[2632] = i[1448];
  assign o[2631] = i[1447];
  assign o[2630] = i[1446];
  assign o[2629] = i[1445];
  assign o[2628] = i[1444];
  assign o[2627] = i[1443];
  assign o[2626] = i[1442];
  assign o[2625] = i[1441];
  assign o[2624] = i[1440];
  assign o[2623] = i[1503];
  assign o[2622] = i[1502];
  assign o[2621] = i[1501];
  assign o[2620] = i[1500];
  assign o[2619] = i[1499];
  assign o[2618] = i[1498];
  assign o[2617] = i[1497];
  assign o[2616] = i[1496];
  assign o[2615] = i[1495];
  assign o[2614] = i[1494];
  assign o[2613] = i[1493];
  assign o[2612] = i[1492];
  assign o[2611] = i[1491];
  assign o[2610] = i[1490];
  assign o[2609] = i[1489];
  assign o[2608] = i[1488];
  assign o[2607] = i[1487];
  assign o[2606] = i[1486];
  assign o[2605] = i[1485];
  assign o[2604] = i[1484];
  assign o[2603] = i[1483];
  assign o[2602] = i[1482];
  assign o[2601] = i[1481];
  assign o[2600] = i[1480];
  assign o[2599] = i[1479];
  assign o[2598] = i[1478];
  assign o[2597] = i[1477];
  assign o[2596] = i[1476];
  assign o[2595] = i[1475];
  assign o[2594] = i[1474];
  assign o[2593] = i[1473];
  assign o[2592] = i[1472];
  assign o[2591] = i[1535];
  assign o[2590] = i[1534];
  assign o[2589] = i[1533];
  assign o[2588] = i[1532];
  assign o[2587] = i[1531];
  assign o[2586] = i[1530];
  assign o[2585] = i[1529];
  assign o[2584] = i[1528];
  assign o[2583] = i[1527];
  assign o[2582] = i[1526];
  assign o[2581] = i[1525];
  assign o[2580] = i[1524];
  assign o[2579] = i[1523];
  assign o[2578] = i[1522];
  assign o[2577] = i[1521];
  assign o[2576] = i[1520];
  assign o[2575] = i[1519];
  assign o[2574] = i[1518];
  assign o[2573] = i[1517];
  assign o[2572] = i[1516];
  assign o[2571] = i[1515];
  assign o[2570] = i[1514];
  assign o[2569] = i[1513];
  assign o[2568] = i[1512];
  assign o[2567] = i[1511];
  assign o[2566] = i[1510];
  assign o[2565] = i[1509];
  assign o[2564] = i[1508];
  assign o[2563] = i[1507];
  assign o[2562] = i[1506];
  assign o[2561] = i[1505];
  assign o[2560] = i[1504];
  assign o[2559] = i[1567];
  assign o[2558] = i[1566];
  assign o[2557] = i[1565];
  assign o[2556] = i[1564];
  assign o[2555] = i[1563];
  assign o[2554] = i[1562];
  assign o[2553] = i[1561];
  assign o[2552] = i[1560];
  assign o[2551] = i[1559];
  assign o[2550] = i[1558];
  assign o[2549] = i[1557];
  assign o[2548] = i[1556];
  assign o[2547] = i[1555];
  assign o[2546] = i[1554];
  assign o[2545] = i[1553];
  assign o[2544] = i[1552];
  assign o[2543] = i[1551];
  assign o[2542] = i[1550];
  assign o[2541] = i[1549];
  assign o[2540] = i[1548];
  assign o[2539] = i[1547];
  assign o[2538] = i[1546];
  assign o[2537] = i[1545];
  assign o[2536] = i[1544];
  assign o[2535] = i[1543];
  assign o[2534] = i[1542];
  assign o[2533] = i[1541];
  assign o[2532] = i[1540];
  assign o[2531] = i[1539];
  assign o[2530] = i[1538];
  assign o[2529] = i[1537];
  assign o[2528] = i[1536];
  assign o[2527] = i[1599];
  assign o[2526] = i[1598];
  assign o[2525] = i[1597];
  assign o[2524] = i[1596];
  assign o[2523] = i[1595];
  assign o[2522] = i[1594];
  assign o[2521] = i[1593];
  assign o[2520] = i[1592];
  assign o[2519] = i[1591];
  assign o[2518] = i[1590];
  assign o[2517] = i[1589];
  assign o[2516] = i[1588];
  assign o[2515] = i[1587];
  assign o[2514] = i[1586];
  assign o[2513] = i[1585];
  assign o[2512] = i[1584];
  assign o[2511] = i[1583];
  assign o[2510] = i[1582];
  assign o[2509] = i[1581];
  assign o[2508] = i[1580];
  assign o[2507] = i[1579];
  assign o[2506] = i[1578];
  assign o[2505] = i[1577];
  assign o[2504] = i[1576];
  assign o[2503] = i[1575];
  assign o[2502] = i[1574];
  assign o[2501] = i[1573];
  assign o[2500] = i[1572];
  assign o[2499] = i[1571];
  assign o[2498] = i[1570];
  assign o[2497] = i[1569];
  assign o[2496] = i[1568];
  assign o[2495] = i[1631];
  assign o[2494] = i[1630];
  assign o[2493] = i[1629];
  assign o[2492] = i[1628];
  assign o[2491] = i[1627];
  assign o[2490] = i[1626];
  assign o[2489] = i[1625];
  assign o[2488] = i[1624];
  assign o[2487] = i[1623];
  assign o[2486] = i[1622];
  assign o[2485] = i[1621];
  assign o[2484] = i[1620];
  assign o[2483] = i[1619];
  assign o[2482] = i[1618];
  assign o[2481] = i[1617];
  assign o[2480] = i[1616];
  assign o[2479] = i[1615];
  assign o[2478] = i[1614];
  assign o[2477] = i[1613];
  assign o[2476] = i[1612];
  assign o[2475] = i[1611];
  assign o[2474] = i[1610];
  assign o[2473] = i[1609];
  assign o[2472] = i[1608];
  assign o[2471] = i[1607];
  assign o[2470] = i[1606];
  assign o[2469] = i[1605];
  assign o[2468] = i[1604];
  assign o[2467] = i[1603];
  assign o[2466] = i[1602];
  assign o[2465] = i[1601];
  assign o[2464] = i[1600];
  assign o[2463] = i[1663];
  assign o[2462] = i[1662];
  assign o[2461] = i[1661];
  assign o[2460] = i[1660];
  assign o[2459] = i[1659];
  assign o[2458] = i[1658];
  assign o[2457] = i[1657];
  assign o[2456] = i[1656];
  assign o[2455] = i[1655];
  assign o[2454] = i[1654];
  assign o[2453] = i[1653];
  assign o[2452] = i[1652];
  assign o[2451] = i[1651];
  assign o[2450] = i[1650];
  assign o[2449] = i[1649];
  assign o[2448] = i[1648];
  assign o[2447] = i[1647];
  assign o[2446] = i[1646];
  assign o[2445] = i[1645];
  assign o[2444] = i[1644];
  assign o[2443] = i[1643];
  assign o[2442] = i[1642];
  assign o[2441] = i[1641];
  assign o[2440] = i[1640];
  assign o[2439] = i[1639];
  assign o[2438] = i[1638];
  assign o[2437] = i[1637];
  assign o[2436] = i[1636];
  assign o[2435] = i[1635];
  assign o[2434] = i[1634];
  assign o[2433] = i[1633];
  assign o[2432] = i[1632];
  assign o[2431] = i[1695];
  assign o[2430] = i[1694];
  assign o[2429] = i[1693];
  assign o[2428] = i[1692];
  assign o[2427] = i[1691];
  assign o[2426] = i[1690];
  assign o[2425] = i[1689];
  assign o[2424] = i[1688];
  assign o[2423] = i[1687];
  assign o[2422] = i[1686];
  assign o[2421] = i[1685];
  assign o[2420] = i[1684];
  assign o[2419] = i[1683];
  assign o[2418] = i[1682];
  assign o[2417] = i[1681];
  assign o[2416] = i[1680];
  assign o[2415] = i[1679];
  assign o[2414] = i[1678];
  assign o[2413] = i[1677];
  assign o[2412] = i[1676];
  assign o[2411] = i[1675];
  assign o[2410] = i[1674];
  assign o[2409] = i[1673];
  assign o[2408] = i[1672];
  assign o[2407] = i[1671];
  assign o[2406] = i[1670];
  assign o[2405] = i[1669];
  assign o[2404] = i[1668];
  assign o[2403] = i[1667];
  assign o[2402] = i[1666];
  assign o[2401] = i[1665];
  assign o[2400] = i[1664];
  assign o[2399] = i[1727];
  assign o[2398] = i[1726];
  assign o[2397] = i[1725];
  assign o[2396] = i[1724];
  assign o[2395] = i[1723];
  assign o[2394] = i[1722];
  assign o[2393] = i[1721];
  assign o[2392] = i[1720];
  assign o[2391] = i[1719];
  assign o[2390] = i[1718];
  assign o[2389] = i[1717];
  assign o[2388] = i[1716];
  assign o[2387] = i[1715];
  assign o[2386] = i[1714];
  assign o[2385] = i[1713];
  assign o[2384] = i[1712];
  assign o[2383] = i[1711];
  assign o[2382] = i[1710];
  assign o[2381] = i[1709];
  assign o[2380] = i[1708];
  assign o[2379] = i[1707];
  assign o[2378] = i[1706];
  assign o[2377] = i[1705];
  assign o[2376] = i[1704];
  assign o[2375] = i[1703];
  assign o[2374] = i[1702];
  assign o[2373] = i[1701];
  assign o[2372] = i[1700];
  assign o[2371] = i[1699];
  assign o[2370] = i[1698];
  assign o[2369] = i[1697];
  assign o[2368] = i[1696];
  assign o[2367] = i[1759];
  assign o[2366] = i[1758];
  assign o[2365] = i[1757];
  assign o[2364] = i[1756];
  assign o[2363] = i[1755];
  assign o[2362] = i[1754];
  assign o[2361] = i[1753];
  assign o[2360] = i[1752];
  assign o[2359] = i[1751];
  assign o[2358] = i[1750];
  assign o[2357] = i[1749];
  assign o[2356] = i[1748];
  assign o[2355] = i[1747];
  assign o[2354] = i[1746];
  assign o[2353] = i[1745];
  assign o[2352] = i[1744];
  assign o[2351] = i[1743];
  assign o[2350] = i[1742];
  assign o[2349] = i[1741];
  assign o[2348] = i[1740];
  assign o[2347] = i[1739];
  assign o[2346] = i[1738];
  assign o[2345] = i[1737];
  assign o[2344] = i[1736];
  assign o[2343] = i[1735];
  assign o[2342] = i[1734];
  assign o[2341] = i[1733];
  assign o[2340] = i[1732];
  assign o[2339] = i[1731];
  assign o[2338] = i[1730];
  assign o[2337] = i[1729];
  assign o[2336] = i[1728];
  assign o[2335] = i[1791];
  assign o[2334] = i[1790];
  assign o[2333] = i[1789];
  assign o[2332] = i[1788];
  assign o[2331] = i[1787];
  assign o[2330] = i[1786];
  assign o[2329] = i[1785];
  assign o[2328] = i[1784];
  assign o[2327] = i[1783];
  assign o[2326] = i[1782];
  assign o[2325] = i[1781];
  assign o[2324] = i[1780];
  assign o[2323] = i[1779];
  assign o[2322] = i[1778];
  assign o[2321] = i[1777];
  assign o[2320] = i[1776];
  assign o[2319] = i[1775];
  assign o[2318] = i[1774];
  assign o[2317] = i[1773];
  assign o[2316] = i[1772];
  assign o[2315] = i[1771];
  assign o[2314] = i[1770];
  assign o[2313] = i[1769];
  assign o[2312] = i[1768];
  assign o[2311] = i[1767];
  assign o[2310] = i[1766];
  assign o[2309] = i[1765];
  assign o[2308] = i[1764];
  assign o[2307] = i[1763];
  assign o[2306] = i[1762];
  assign o[2305] = i[1761];
  assign o[2304] = i[1760];
  assign o[2303] = i[1823];
  assign o[2302] = i[1822];
  assign o[2301] = i[1821];
  assign o[2300] = i[1820];
  assign o[2299] = i[1819];
  assign o[2298] = i[1818];
  assign o[2297] = i[1817];
  assign o[2296] = i[1816];
  assign o[2295] = i[1815];
  assign o[2294] = i[1814];
  assign o[2293] = i[1813];
  assign o[2292] = i[1812];
  assign o[2291] = i[1811];
  assign o[2290] = i[1810];
  assign o[2289] = i[1809];
  assign o[2288] = i[1808];
  assign o[2287] = i[1807];
  assign o[2286] = i[1806];
  assign o[2285] = i[1805];
  assign o[2284] = i[1804];
  assign o[2283] = i[1803];
  assign o[2282] = i[1802];
  assign o[2281] = i[1801];
  assign o[2280] = i[1800];
  assign o[2279] = i[1799];
  assign o[2278] = i[1798];
  assign o[2277] = i[1797];
  assign o[2276] = i[1796];
  assign o[2275] = i[1795];
  assign o[2274] = i[1794];
  assign o[2273] = i[1793];
  assign o[2272] = i[1792];
  assign o[2271] = i[1855];
  assign o[2270] = i[1854];
  assign o[2269] = i[1853];
  assign o[2268] = i[1852];
  assign o[2267] = i[1851];
  assign o[2266] = i[1850];
  assign o[2265] = i[1849];
  assign o[2264] = i[1848];
  assign o[2263] = i[1847];
  assign o[2262] = i[1846];
  assign o[2261] = i[1845];
  assign o[2260] = i[1844];
  assign o[2259] = i[1843];
  assign o[2258] = i[1842];
  assign o[2257] = i[1841];
  assign o[2256] = i[1840];
  assign o[2255] = i[1839];
  assign o[2254] = i[1838];
  assign o[2253] = i[1837];
  assign o[2252] = i[1836];
  assign o[2251] = i[1835];
  assign o[2250] = i[1834];
  assign o[2249] = i[1833];
  assign o[2248] = i[1832];
  assign o[2247] = i[1831];
  assign o[2246] = i[1830];
  assign o[2245] = i[1829];
  assign o[2244] = i[1828];
  assign o[2243] = i[1827];
  assign o[2242] = i[1826];
  assign o[2241] = i[1825];
  assign o[2240] = i[1824];
  assign o[2239] = i[1887];
  assign o[2238] = i[1886];
  assign o[2237] = i[1885];
  assign o[2236] = i[1884];
  assign o[2235] = i[1883];
  assign o[2234] = i[1882];
  assign o[2233] = i[1881];
  assign o[2232] = i[1880];
  assign o[2231] = i[1879];
  assign o[2230] = i[1878];
  assign o[2229] = i[1877];
  assign o[2228] = i[1876];
  assign o[2227] = i[1875];
  assign o[2226] = i[1874];
  assign o[2225] = i[1873];
  assign o[2224] = i[1872];
  assign o[2223] = i[1871];
  assign o[2222] = i[1870];
  assign o[2221] = i[1869];
  assign o[2220] = i[1868];
  assign o[2219] = i[1867];
  assign o[2218] = i[1866];
  assign o[2217] = i[1865];
  assign o[2216] = i[1864];
  assign o[2215] = i[1863];
  assign o[2214] = i[1862];
  assign o[2213] = i[1861];
  assign o[2212] = i[1860];
  assign o[2211] = i[1859];
  assign o[2210] = i[1858];
  assign o[2209] = i[1857];
  assign o[2208] = i[1856];
  assign o[2207] = i[1919];
  assign o[2206] = i[1918];
  assign o[2205] = i[1917];
  assign o[2204] = i[1916];
  assign o[2203] = i[1915];
  assign o[2202] = i[1914];
  assign o[2201] = i[1913];
  assign o[2200] = i[1912];
  assign o[2199] = i[1911];
  assign o[2198] = i[1910];
  assign o[2197] = i[1909];
  assign o[2196] = i[1908];
  assign o[2195] = i[1907];
  assign o[2194] = i[1906];
  assign o[2193] = i[1905];
  assign o[2192] = i[1904];
  assign o[2191] = i[1903];
  assign o[2190] = i[1902];
  assign o[2189] = i[1901];
  assign o[2188] = i[1900];
  assign o[2187] = i[1899];
  assign o[2186] = i[1898];
  assign o[2185] = i[1897];
  assign o[2184] = i[1896];
  assign o[2183] = i[1895];
  assign o[2182] = i[1894];
  assign o[2181] = i[1893];
  assign o[2180] = i[1892];
  assign o[2179] = i[1891];
  assign o[2178] = i[1890];
  assign o[2177] = i[1889];
  assign o[2176] = i[1888];
  assign o[2175] = i[1951];
  assign o[2174] = i[1950];
  assign o[2173] = i[1949];
  assign o[2172] = i[1948];
  assign o[2171] = i[1947];
  assign o[2170] = i[1946];
  assign o[2169] = i[1945];
  assign o[2168] = i[1944];
  assign o[2167] = i[1943];
  assign o[2166] = i[1942];
  assign o[2165] = i[1941];
  assign o[2164] = i[1940];
  assign o[2163] = i[1939];
  assign o[2162] = i[1938];
  assign o[2161] = i[1937];
  assign o[2160] = i[1936];
  assign o[2159] = i[1935];
  assign o[2158] = i[1934];
  assign o[2157] = i[1933];
  assign o[2156] = i[1932];
  assign o[2155] = i[1931];
  assign o[2154] = i[1930];
  assign o[2153] = i[1929];
  assign o[2152] = i[1928];
  assign o[2151] = i[1927];
  assign o[2150] = i[1926];
  assign o[2149] = i[1925];
  assign o[2148] = i[1924];
  assign o[2147] = i[1923];
  assign o[2146] = i[1922];
  assign o[2145] = i[1921];
  assign o[2144] = i[1920];
  assign o[2143] = i[1983];
  assign o[2142] = i[1982];
  assign o[2141] = i[1981];
  assign o[2140] = i[1980];
  assign o[2139] = i[1979];
  assign o[2138] = i[1978];
  assign o[2137] = i[1977];
  assign o[2136] = i[1976];
  assign o[2135] = i[1975];
  assign o[2134] = i[1974];
  assign o[2133] = i[1973];
  assign o[2132] = i[1972];
  assign o[2131] = i[1971];
  assign o[2130] = i[1970];
  assign o[2129] = i[1969];
  assign o[2128] = i[1968];
  assign o[2127] = i[1967];
  assign o[2126] = i[1966];
  assign o[2125] = i[1965];
  assign o[2124] = i[1964];
  assign o[2123] = i[1963];
  assign o[2122] = i[1962];
  assign o[2121] = i[1961];
  assign o[2120] = i[1960];
  assign o[2119] = i[1959];
  assign o[2118] = i[1958];
  assign o[2117] = i[1957];
  assign o[2116] = i[1956];
  assign o[2115] = i[1955];
  assign o[2114] = i[1954];
  assign o[2113] = i[1953];
  assign o[2112] = i[1952];
  assign o[2111] = i[2015];
  assign o[2110] = i[2014];
  assign o[2109] = i[2013];
  assign o[2108] = i[2012];
  assign o[2107] = i[2011];
  assign o[2106] = i[2010];
  assign o[2105] = i[2009];
  assign o[2104] = i[2008];
  assign o[2103] = i[2007];
  assign o[2102] = i[2006];
  assign o[2101] = i[2005];
  assign o[2100] = i[2004];
  assign o[2099] = i[2003];
  assign o[2098] = i[2002];
  assign o[2097] = i[2001];
  assign o[2096] = i[2000];
  assign o[2095] = i[1999];
  assign o[2094] = i[1998];
  assign o[2093] = i[1997];
  assign o[2092] = i[1996];
  assign o[2091] = i[1995];
  assign o[2090] = i[1994];
  assign o[2089] = i[1993];
  assign o[2088] = i[1992];
  assign o[2087] = i[1991];
  assign o[2086] = i[1990];
  assign o[2085] = i[1989];
  assign o[2084] = i[1988];
  assign o[2083] = i[1987];
  assign o[2082] = i[1986];
  assign o[2081] = i[1985];
  assign o[2080] = i[1984];
  assign o[2079] = i[2047];
  assign o[2078] = i[2046];
  assign o[2077] = i[2045];
  assign o[2076] = i[2044];
  assign o[2075] = i[2043];
  assign o[2074] = i[2042];
  assign o[2073] = i[2041];
  assign o[2072] = i[2040];
  assign o[2071] = i[2039];
  assign o[2070] = i[2038];
  assign o[2069] = i[2037];
  assign o[2068] = i[2036];
  assign o[2067] = i[2035];
  assign o[2066] = i[2034];
  assign o[2065] = i[2033];
  assign o[2064] = i[2032];
  assign o[2063] = i[2031];
  assign o[2062] = i[2030];
  assign o[2061] = i[2029];
  assign o[2060] = i[2028];
  assign o[2059] = i[2027];
  assign o[2058] = i[2026];
  assign o[2057] = i[2025];
  assign o[2056] = i[2024];
  assign o[2055] = i[2023];
  assign o[2054] = i[2022];
  assign o[2053] = i[2021];
  assign o[2052] = i[2020];
  assign o[2051] = i[2019];
  assign o[2050] = i[2018];
  assign o[2049] = i[2017];
  assign o[2048] = i[2016];
  assign o[2047] = i[2079];
  assign o[2046] = i[2078];
  assign o[2045] = i[2077];
  assign o[2044] = i[2076];
  assign o[2043] = i[2075];
  assign o[2042] = i[2074];
  assign o[2041] = i[2073];
  assign o[2040] = i[2072];
  assign o[2039] = i[2071];
  assign o[2038] = i[2070];
  assign o[2037] = i[2069];
  assign o[2036] = i[2068];
  assign o[2035] = i[2067];
  assign o[2034] = i[2066];
  assign o[2033] = i[2065];
  assign o[2032] = i[2064];
  assign o[2031] = i[2063];
  assign o[2030] = i[2062];
  assign o[2029] = i[2061];
  assign o[2028] = i[2060];
  assign o[2027] = i[2059];
  assign o[2026] = i[2058];
  assign o[2025] = i[2057];
  assign o[2024] = i[2056];
  assign o[2023] = i[2055];
  assign o[2022] = i[2054];
  assign o[2021] = i[2053];
  assign o[2020] = i[2052];
  assign o[2019] = i[2051];
  assign o[2018] = i[2050];
  assign o[2017] = i[2049];
  assign o[2016] = i[2048];
  assign o[2015] = i[2111];
  assign o[2014] = i[2110];
  assign o[2013] = i[2109];
  assign o[2012] = i[2108];
  assign o[2011] = i[2107];
  assign o[2010] = i[2106];
  assign o[2009] = i[2105];
  assign o[2008] = i[2104];
  assign o[2007] = i[2103];
  assign o[2006] = i[2102];
  assign o[2005] = i[2101];
  assign o[2004] = i[2100];
  assign o[2003] = i[2099];
  assign o[2002] = i[2098];
  assign o[2001] = i[2097];
  assign o[2000] = i[2096];
  assign o[1999] = i[2095];
  assign o[1998] = i[2094];
  assign o[1997] = i[2093];
  assign o[1996] = i[2092];
  assign o[1995] = i[2091];
  assign o[1994] = i[2090];
  assign o[1993] = i[2089];
  assign o[1992] = i[2088];
  assign o[1991] = i[2087];
  assign o[1990] = i[2086];
  assign o[1989] = i[2085];
  assign o[1988] = i[2084];
  assign o[1987] = i[2083];
  assign o[1986] = i[2082];
  assign o[1985] = i[2081];
  assign o[1984] = i[2080];
  assign o[1983] = i[2143];
  assign o[1982] = i[2142];
  assign o[1981] = i[2141];
  assign o[1980] = i[2140];
  assign o[1979] = i[2139];
  assign o[1978] = i[2138];
  assign o[1977] = i[2137];
  assign o[1976] = i[2136];
  assign o[1975] = i[2135];
  assign o[1974] = i[2134];
  assign o[1973] = i[2133];
  assign o[1972] = i[2132];
  assign o[1971] = i[2131];
  assign o[1970] = i[2130];
  assign o[1969] = i[2129];
  assign o[1968] = i[2128];
  assign o[1967] = i[2127];
  assign o[1966] = i[2126];
  assign o[1965] = i[2125];
  assign o[1964] = i[2124];
  assign o[1963] = i[2123];
  assign o[1962] = i[2122];
  assign o[1961] = i[2121];
  assign o[1960] = i[2120];
  assign o[1959] = i[2119];
  assign o[1958] = i[2118];
  assign o[1957] = i[2117];
  assign o[1956] = i[2116];
  assign o[1955] = i[2115];
  assign o[1954] = i[2114];
  assign o[1953] = i[2113];
  assign o[1952] = i[2112];
  assign o[1951] = i[2175];
  assign o[1950] = i[2174];
  assign o[1949] = i[2173];
  assign o[1948] = i[2172];
  assign o[1947] = i[2171];
  assign o[1946] = i[2170];
  assign o[1945] = i[2169];
  assign o[1944] = i[2168];
  assign o[1943] = i[2167];
  assign o[1942] = i[2166];
  assign o[1941] = i[2165];
  assign o[1940] = i[2164];
  assign o[1939] = i[2163];
  assign o[1938] = i[2162];
  assign o[1937] = i[2161];
  assign o[1936] = i[2160];
  assign o[1935] = i[2159];
  assign o[1934] = i[2158];
  assign o[1933] = i[2157];
  assign o[1932] = i[2156];
  assign o[1931] = i[2155];
  assign o[1930] = i[2154];
  assign o[1929] = i[2153];
  assign o[1928] = i[2152];
  assign o[1927] = i[2151];
  assign o[1926] = i[2150];
  assign o[1925] = i[2149];
  assign o[1924] = i[2148];
  assign o[1923] = i[2147];
  assign o[1922] = i[2146];
  assign o[1921] = i[2145];
  assign o[1920] = i[2144];
  assign o[1919] = i[2207];
  assign o[1918] = i[2206];
  assign o[1917] = i[2205];
  assign o[1916] = i[2204];
  assign o[1915] = i[2203];
  assign o[1914] = i[2202];
  assign o[1913] = i[2201];
  assign o[1912] = i[2200];
  assign o[1911] = i[2199];
  assign o[1910] = i[2198];
  assign o[1909] = i[2197];
  assign o[1908] = i[2196];
  assign o[1907] = i[2195];
  assign o[1906] = i[2194];
  assign o[1905] = i[2193];
  assign o[1904] = i[2192];
  assign o[1903] = i[2191];
  assign o[1902] = i[2190];
  assign o[1901] = i[2189];
  assign o[1900] = i[2188];
  assign o[1899] = i[2187];
  assign o[1898] = i[2186];
  assign o[1897] = i[2185];
  assign o[1896] = i[2184];
  assign o[1895] = i[2183];
  assign o[1894] = i[2182];
  assign o[1893] = i[2181];
  assign o[1892] = i[2180];
  assign o[1891] = i[2179];
  assign o[1890] = i[2178];
  assign o[1889] = i[2177];
  assign o[1888] = i[2176];
  assign o[1887] = i[2239];
  assign o[1886] = i[2238];
  assign o[1885] = i[2237];
  assign o[1884] = i[2236];
  assign o[1883] = i[2235];
  assign o[1882] = i[2234];
  assign o[1881] = i[2233];
  assign o[1880] = i[2232];
  assign o[1879] = i[2231];
  assign o[1878] = i[2230];
  assign o[1877] = i[2229];
  assign o[1876] = i[2228];
  assign o[1875] = i[2227];
  assign o[1874] = i[2226];
  assign o[1873] = i[2225];
  assign o[1872] = i[2224];
  assign o[1871] = i[2223];
  assign o[1870] = i[2222];
  assign o[1869] = i[2221];
  assign o[1868] = i[2220];
  assign o[1867] = i[2219];
  assign o[1866] = i[2218];
  assign o[1865] = i[2217];
  assign o[1864] = i[2216];
  assign o[1863] = i[2215];
  assign o[1862] = i[2214];
  assign o[1861] = i[2213];
  assign o[1860] = i[2212];
  assign o[1859] = i[2211];
  assign o[1858] = i[2210];
  assign o[1857] = i[2209];
  assign o[1856] = i[2208];
  assign o[1855] = i[2271];
  assign o[1854] = i[2270];
  assign o[1853] = i[2269];
  assign o[1852] = i[2268];
  assign o[1851] = i[2267];
  assign o[1850] = i[2266];
  assign o[1849] = i[2265];
  assign o[1848] = i[2264];
  assign o[1847] = i[2263];
  assign o[1846] = i[2262];
  assign o[1845] = i[2261];
  assign o[1844] = i[2260];
  assign o[1843] = i[2259];
  assign o[1842] = i[2258];
  assign o[1841] = i[2257];
  assign o[1840] = i[2256];
  assign o[1839] = i[2255];
  assign o[1838] = i[2254];
  assign o[1837] = i[2253];
  assign o[1836] = i[2252];
  assign o[1835] = i[2251];
  assign o[1834] = i[2250];
  assign o[1833] = i[2249];
  assign o[1832] = i[2248];
  assign o[1831] = i[2247];
  assign o[1830] = i[2246];
  assign o[1829] = i[2245];
  assign o[1828] = i[2244];
  assign o[1827] = i[2243];
  assign o[1826] = i[2242];
  assign o[1825] = i[2241];
  assign o[1824] = i[2240];
  assign o[1823] = i[2303];
  assign o[1822] = i[2302];
  assign o[1821] = i[2301];
  assign o[1820] = i[2300];
  assign o[1819] = i[2299];
  assign o[1818] = i[2298];
  assign o[1817] = i[2297];
  assign o[1816] = i[2296];
  assign o[1815] = i[2295];
  assign o[1814] = i[2294];
  assign o[1813] = i[2293];
  assign o[1812] = i[2292];
  assign o[1811] = i[2291];
  assign o[1810] = i[2290];
  assign o[1809] = i[2289];
  assign o[1808] = i[2288];
  assign o[1807] = i[2287];
  assign o[1806] = i[2286];
  assign o[1805] = i[2285];
  assign o[1804] = i[2284];
  assign o[1803] = i[2283];
  assign o[1802] = i[2282];
  assign o[1801] = i[2281];
  assign o[1800] = i[2280];
  assign o[1799] = i[2279];
  assign o[1798] = i[2278];
  assign o[1797] = i[2277];
  assign o[1796] = i[2276];
  assign o[1795] = i[2275];
  assign o[1794] = i[2274];
  assign o[1793] = i[2273];
  assign o[1792] = i[2272];
  assign o[1791] = i[2335];
  assign o[1790] = i[2334];
  assign o[1789] = i[2333];
  assign o[1788] = i[2332];
  assign o[1787] = i[2331];
  assign o[1786] = i[2330];
  assign o[1785] = i[2329];
  assign o[1784] = i[2328];
  assign o[1783] = i[2327];
  assign o[1782] = i[2326];
  assign o[1781] = i[2325];
  assign o[1780] = i[2324];
  assign o[1779] = i[2323];
  assign o[1778] = i[2322];
  assign o[1777] = i[2321];
  assign o[1776] = i[2320];
  assign o[1775] = i[2319];
  assign o[1774] = i[2318];
  assign o[1773] = i[2317];
  assign o[1772] = i[2316];
  assign o[1771] = i[2315];
  assign o[1770] = i[2314];
  assign o[1769] = i[2313];
  assign o[1768] = i[2312];
  assign o[1767] = i[2311];
  assign o[1766] = i[2310];
  assign o[1765] = i[2309];
  assign o[1764] = i[2308];
  assign o[1763] = i[2307];
  assign o[1762] = i[2306];
  assign o[1761] = i[2305];
  assign o[1760] = i[2304];
  assign o[1759] = i[2367];
  assign o[1758] = i[2366];
  assign o[1757] = i[2365];
  assign o[1756] = i[2364];
  assign o[1755] = i[2363];
  assign o[1754] = i[2362];
  assign o[1753] = i[2361];
  assign o[1752] = i[2360];
  assign o[1751] = i[2359];
  assign o[1750] = i[2358];
  assign o[1749] = i[2357];
  assign o[1748] = i[2356];
  assign o[1747] = i[2355];
  assign o[1746] = i[2354];
  assign o[1745] = i[2353];
  assign o[1744] = i[2352];
  assign o[1743] = i[2351];
  assign o[1742] = i[2350];
  assign o[1741] = i[2349];
  assign o[1740] = i[2348];
  assign o[1739] = i[2347];
  assign o[1738] = i[2346];
  assign o[1737] = i[2345];
  assign o[1736] = i[2344];
  assign o[1735] = i[2343];
  assign o[1734] = i[2342];
  assign o[1733] = i[2341];
  assign o[1732] = i[2340];
  assign o[1731] = i[2339];
  assign o[1730] = i[2338];
  assign o[1729] = i[2337];
  assign o[1728] = i[2336];
  assign o[1727] = i[2399];
  assign o[1726] = i[2398];
  assign o[1725] = i[2397];
  assign o[1724] = i[2396];
  assign o[1723] = i[2395];
  assign o[1722] = i[2394];
  assign o[1721] = i[2393];
  assign o[1720] = i[2392];
  assign o[1719] = i[2391];
  assign o[1718] = i[2390];
  assign o[1717] = i[2389];
  assign o[1716] = i[2388];
  assign o[1715] = i[2387];
  assign o[1714] = i[2386];
  assign o[1713] = i[2385];
  assign o[1712] = i[2384];
  assign o[1711] = i[2383];
  assign o[1710] = i[2382];
  assign o[1709] = i[2381];
  assign o[1708] = i[2380];
  assign o[1707] = i[2379];
  assign o[1706] = i[2378];
  assign o[1705] = i[2377];
  assign o[1704] = i[2376];
  assign o[1703] = i[2375];
  assign o[1702] = i[2374];
  assign o[1701] = i[2373];
  assign o[1700] = i[2372];
  assign o[1699] = i[2371];
  assign o[1698] = i[2370];
  assign o[1697] = i[2369];
  assign o[1696] = i[2368];
  assign o[1695] = i[2431];
  assign o[1694] = i[2430];
  assign o[1693] = i[2429];
  assign o[1692] = i[2428];
  assign o[1691] = i[2427];
  assign o[1690] = i[2426];
  assign o[1689] = i[2425];
  assign o[1688] = i[2424];
  assign o[1687] = i[2423];
  assign o[1686] = i[2422];
  assign o[1685] = i[2421];
  assign o[1684] = i[2420];
  assign o[1683] = i[2419];
  assign o[1682] = i[2418];
  assign o[1681] = i[2417];
  assign o[1680] = i[2416];
  assign o[1679] = i[2415];
  assign o[1678] = i[2414];
  assign o[1677] = i[2413];
  assign o[1676] = i[2412];
  assign o[1675] = i[2411];
  assign o[1674] = i[2410];
  assign o[1673] = i[2409];
  assign o[1672] = i[2408];
  assign o[1671] = i[2407];
  assign o[1670] = i[2406];
  assign o[1669] = i[2405];
  assign o[1668] = i[2404];
  assign o[1667] = i[2403];
  assign o[1666] = i[2402];
  assign o[1665] = i[2401];
  assign o[1664] = i[2400];
  assign o[1663] = i[2463];
  assign o[1662] = i[2462];
  assign o[1661] = i[2461];
  assign o[1660] = i[2460];
  assign o[1659] = i[2459];
  assign o[1658] = i[2458];
  assign o[1657] = i[2457];
  assign o[1656] = i[2456];
  assign o[1655] = i[2455];
  assign o[1654] = i[2454];
  assign o[1653] = i[2453];
  assign o[1652] = i[2452];
  assign o[1651] = i[2451];
  assign o[1650] = i[2450];
  assign o[1649] = i[2449];
  assign o[1648] = i[2448];
  assign o[1647] = i[2447];
  assign o[1646] = i[2446];
  assign o[1645] = i[2445];
  assign o[1644] = i[2444];
  assign o[1643] = i[2443];
  assign o[1642] = i[2442];
  assign o[1641] = i[2441];
  assign o[1640] = i[2440];
  assign o[1639] = i[2439];
  assign o[1638] = i[2438];
  assign o[1637] = i[2437];
  assign o[1636] = i[2436];
  assign o[1635] = i[2435];
  assign o[1634] = i[2434];
  assign o[1633] = i[2433];
  assign o[1632] = i[2432];
  assign o[1631] = i[2495];
  assign o[1630] = i[2494];
  assign o[1629] = i[2493];
  assign o[1628] = i[2492];
  assign o[1627] = i[2491];
  assign o[1626] = i[2490];
  assign o[1625] = i[2489];
  assign o[1624] = i[2488];
  assign o[1623] = i[2487];
  assign o[1622] = i[2486];
  assign o[1621] = i[2485];
  assign o[1620] = i[2484];
  assign o[1619] = i[2483];
  assign o[1618] = i[2482];
  assign o[1617] = i[2481];
  assign o[1616] = i[2480];
  assign o[1615] = i[2479];
  assign o[1614] = i[2478];
  assign o[1613] = i[2477];
  assign o[1612] = i[2476];
  assign o[1611] = i[2475];
  assign o[1610] = i[2474];
  assign o[1609] = i[2473];
  assign o[1608] = i[2472];
  assign o[1607] = i[2471];
  assign o[1606] = i[2470];
  assign o[1605] = i[2469];
  assign o[1604] = i[2468];
  assign o[1603] = i[2467];
  assign o[1602] = i[2466];
  assign o[1601] = i[2465];
  assign o[1600] = i[2464];
  assign o[1599] = i[2527];
  assign o[1598] = i[2526];
  assign o[1597] = i[2525];
  assign o[1596] = i[2524];
  assign o[1595] = i[2523];
  assign o[1594] = i[2522];
  assign o[1593] = i[2521];
  assign o[1592] = i[2520];
  assign o[1591] = i[2519];
  assign o[1590] = i[2518];
  assign o[1589] = i[2517];
  assign o[1588] = i[2516];
  assign o[1587] = i[2515];
  assign o[1586] = i[2514];
  assign o[1585] = i[2513];
  assign o[1584] = i[2512];
  assign o[1583] = i[2511];
  assign o[1582] = i[2510];
  assign o[1581] = i[2509];
  assign o[1580] = i[2508];
  assign o[1579] = i[2507];
  assign o[1578] = i[2506];
  assign o[1577] = i[2505];
  assign o[1576] = i[2504];
  assign o[1575] = i[2503];
  assign o[1574] = i[2502];
  assign o[1573] = i[2501];
  assign o[1572] = i[2500];
  assign o[1571] = i[2499];
  assign o[1570] = i[2498];
  assign o[1569] = i[2497];
  assign o[1568] = i[2496];
  assign o[1567] = i[2559];
  assign o[1566] = i[2558];
  assign o[1565] = i[2557];
  assign o[1564] = i[2556];
  assign o[1563] = i[2555];
  assign o[1562] = i[2554];
  assign o[1561] = i[2553];
  assign o[1560] = i[2552];
  assign o[1559] = i[2551];
  assign o[1558] = i[2550];
  assign o[1557] = i[2549];
  assign o[1556] = i[2548];
  assign o[1555] = i[2547];
  assign o[1554] = i[2546];
  assign o[1553] = i[2545];
  assign o[1552] = i[2544];
  assign o[1551] = i[2543];
  assign o[1550] = i[2542];
  assign o[1549] = i[2541];
  assign o[1548] = i[2540];
  assign o[1547] = i[2539];
  assign o[1546] = i[2538];
  assign o[1545] = i[2537];
  assign o[1544] = i[2536];
  assign o[1543] = i[2535];
  assign o[1542] = i[2534];
  assign o[1541] = i[2533];
  assign o[1540] = i[2532];
  assign o[1539] = i[2531];
  assign o[1538] = i[2530];
  assign o[1537] = i[2529];
  assign o[1536] = i[2528];
  assign o[1535] = i[2591];
  assign o[1534] = i[2590];
  assign o[1533] = i[2589];
  assign o[1532] = i[2588];
  assign o[1531] = i[2587];
  assign o[1530] = i[2586];
  assign o[1529] = i[2585];
  assign o[1528] = i[2584];
  assign o[1527] = i[2583];
  assign o[1526] = i[2582];
  assign o[1525] = i[2581];
  assign o[1524] = i[2580];
  assign o[1523] = i[2579];
  assign o[1522] = i[2578];
  assign o[1521] = i[2577];
  assign o[1520] = i[2576];
  assign o[1519] = i[2575];
  assign o[1518] = i[2574];
  assign o[1517] = i[2573];
  assign o[1516] = i[2572];
  assign o[1515] = i[2571];
  assign o[1514] = i[2570];
  assign o[1513] = i[2569];
  assign o[1512] = i[2568];
  assign o[1511] = i[2567];
  assign o[1510] = i[2566];
  assign o[1509] = i[2565];
  assign o[1508] = i[2564];
  assign o[1507] = i[2563];
  assign o[1506] = i[2562];
  assign o[1505] = i[2561];
  assign o[1504] = i[2560];
  assign o[1503] = i[2623];
  assign o[1502] = i[2622];
  assign o[1501] = i[2621];
  assign o[1500] = i[2620];
  assign o[1499] = i[2619];
  assign o[1498] = i[2618];
  assign o[1497] = i[2617];
  assign o[1496] = i[2616];
  assign o[1495] = i[2615];
  assign o[1494] = i[2614];
  assign o[1493] = i[2613];
  assign o[1492] = i[2612];
  assign o[1491] = i[2611];
  assign o[1490] = i[2610];
  assign o[1489] = i[2609];
  assign o[1488] = i[2608];
  assign o[1487] = i[2607];
  assign o[1486] = i[2606];
  assign o[1485] = i[2605];
  assign o[1484] = i[2604];
  assign o[1483] = i[2603];
  assign o[1482] = i[2602];
  assign o[1481] = i[2601];
  assign o[1480] = i[2600];
  assign o[1479] = i[2599];
  assign o[1478] = i[2598];
  assign o[1477] = i[2597];
  assign o[1476] = i[2596];
  assign o[1475] = i[2595];
  assign o[1474] = i[2594];
  assign o[1473] = i[2593];
  assign o[1472] = i[2592];
  assign o[1471] = i[2655];
  assign o[1470] = i[2654];
  assign o[1469] = i[2653];
  assign o[1468] = i[2652];
  assign o[1467] = i[2651];
  assign o[1466] = i[2650];
  assign o[1465] = i[2649];
  assign o[1464] = i[2648];
  assign o[1463] = i[2647];
  assign o[1462] = i[2646];
  assign o[1461] = i[2645];
  assign o[1460] = i[2644];
  assign o[1459] = i[2643];
  assign o[1458] = i[2642];
  assign o[1457] = i[2641];
  assign o[1456] = i[2640];
  assign o[1455] = i[2639];
  assign o[1454] = i[2638];
  assign o[1453] = i[2637];
  assign o[1452] = i[2636];
  assign o[1451] = i[2635];
  assign o[1450] = i[2634];
  assign o[1449] = i[2633];
  assign o[1448] = i[2632];
  assign o[1447] = i[2631];
  assign o[1446] = i[2630];
  assign o[1445] = i[2629];
  assign o[1444] = i[2628];
  assign o[1443] = i[2627];
  assign o[1442] = i[2626];
  assign o[1441] = i[2625];
  assign o[1440] = i[2624];
  assign o[1439] = i[2687];
  assign o[1438] = i[2686];
  assign o[1437] = i[2685];
  assign o[1436] = i[2684];
  assign o[1435] = i[2683];
  assign o[1434] = i[2682];
  assign o[1433] = i[2681];
  assign o[1432] = i[2680];
  assign o[1431] = i[2679];
  assign o[1430] = i[2678];
  assign o[1429] = i[2677];
  assign o[1428] = i[2676];
  assign o[1427] = i[2675];
  assign o[1426] = i[2674];
  assign o[1425] = i[2673];
  assign o[1424] = i[2672];
  assign o[1423] = i[2671];
  assign o[1422] = i[2670];
  assign o[1421] = i[2669];
  assign o[1420] = i[2668];
  assign o[1419] = i[2667];
  assign o[1418] = i[2666];
  assign o[1417] = i[2665];
  assign o[1416] = i[2664];
  assign o[1415] = i[2663];
  assign o[1414] = i[2662];
  assign o[1413] = i[2661];
  assign o[1412] = i[2660];
  assign o[1411] = i[2659];
  assign o[1410] = i[2658];
  assign o[1409] = i[2657];
  assign o[1408] = i[2656];
  assign o[1407] = i[2719];
  assign o[1406] = i[2718];
  assign o[1405] = i[2717];
  assign o[1404] = i[2716];
  assign o[1403] = i[2715];
  assign o[1402] = i[2714];
  assign o[1401] = i[2713];
  assign o[1400] = i[2712];
  assign o[1399] = i[2711];
  assign o[1398] = i[2710];
  assign o[1397] = i[2709];
  assign o[1396] = i[2708];
  assign o[1395] = i[2707];
  assign o[1394] = i[2706];
  assign o[1393] = i[2705];
  assign o[1392] = i[2704];
  assign o[1391] = i[2703];
  assign o[1390] = i[2702];
  assign o[1389] = i[2701];
  assign o[1388] = i[2700];
  assign o[1387] = i[2699];
  assign o[1386] = i[2698];
  assign o[1385] = i[2697];
  assign o[1384] = i[2696];
  assign o[1383] = i[2695];
  assign o[1382] = i[2694];
  assign o[1381] = i[2693];
  assign o[1380] = i[2692];
  assign o[1379] = i[2691];
  assign o[1378] = i[2690];
  assign o[1377] = i[2689];
  assign o[1376] = i[2688];
  assign o[1375] = i[2751];
  assign o[1374] = i[2750];
  assign o[1373] = i[2749];
  assign o[1372] = i[2748];
  assign o[1371] = i[2747];
  assign o[1370] = i[2746];
  assign o[1369] = i[2745];
  assign o[1368] = i[2744];
  assign o[1367] = i[2743];
  assign o[1366] = i[2742];
  assign o[1365] = i[2741];
  assign o[1364] = i[2740];
  assign o[1363] = i[2739];
  assign o[1362] = i[2738];
  assign o[1361] = i[2737];
  assign o[1360] = i[2736];
  assign o[1359] = i[2735];
  assign o[1358] = i[2734];
  assign o[1357] = i[2733];
  assign o[1356] = i[2732];
  assign o[1355] = i[2731];
  assign o[1354] = i[2730];
  assign o[1353] = i[2729];
  assign o[1352] = i[2728];
  assign o[1351] = i[2727];
  assign o[1350] = i[2726];
  assign o[1349] = i[2725];
  assign o[1348] = i[2724];
  assign o[1347] = i[2723];
  assign o[1346] = i[2722];
  assign o[1345] = i[2721];
  assign o[1344] = i[2720];
  assign o[1343] = i[2783];
  assign o[1342] = i[2782];
  assign o[1341] = i[2781];
  assign o[1340] = i[2780];
  assign o[1339] = i[2779];
  assign o[1338] = i[2778];
  assign o[1337] = i[2777];
  assign o[1336] = i[2776];
  assign o[1335] = i[2775];
  assign o[1334] = i[2774];
  assign o[1333] = i[2773];
  assign o[1332] = i[2772];
  assign o[1331] = i[2771];
  assign o[1330] = i[2770];
  assign o[1329] = i[2769];
  assign o[1328] = i[2768];
  assign o[1327] = i[2767];
  assign o[1326] = i[2766];
  assign o[1325] = i[2765];
  assign o[1324] = i[2764];
  assign o[1323] = i[2763];
  assign o[1322] = i[2762];
  assign o[1321] = i[2761];
  assign o[1320] = i[2760];
  assign o[1319] = i[2759];
  assign o[1318] = i[2758];
  assign o[1317] = i[2757];
  assign o[1316] = i[2756];
  assign o[1315] = i[2755];
  assign o[1314] = i[2754];
  assign o[1313] = i[2753];
  assign o[1312] = i[2752];
  assign o[1311] = i[2815];
  assign o[1310] = i[2814];
  assign o[1309] = i[2813];
  assign o[1308] = i[2812];
  assign o[1307] = i[2811];
  assign o[1306] = i[2810];
  assign o[1305] = i[2809];
  assign o[1304] = i[2808];
  assign o[1303] = i[2807];
  assign o[1302] = i[2806];
  assign o[1301] = i[2805];
  assign o[1300] = i[2804];
  assign o[1299] = i[2803];
  assign o[1298] = i[2802];
  assign o[1297] = i[2801];
  assign o[1296] = i[2800];
  assign o[1295] = i[2799];
  assign o[1294] = i[2798];
  assign o[1293] = i[2797];
  assign o[1292] = i[2796];
  assign o[1291] = i[2795];
  assign o[1290] = i[2794];
  assign o[1289] = i[2793];
  assign o[1288] = i[2792];
  assign o[1287] = i[2791];
  assign o[1286] = i[2790];
  assign o[1285] = i[2789];
  assign o[1284] = i[2788];
  assign o[1283] = i[2787];
  assign o[1282] = i[2786];
  assign o[1281] = i[2785];
  assign o[1280] = i[2784];
  assign o[1279] = i[2847];
  assign o[1278] = i[2846];
  assign o[1277] = i[2845];
  assign o[1276] = i[2844];
  assign o[1275] = i[2843];
  assign o[1274] = i[2842];
  assign o[1273] = i[2841];
  assign o[1272] = i[2840];
  assign o[1271] = i[2839];
  assign o[1270] = i[2838];
  assign o[1269] = i[2837];
  assign o[1268] = i[2836];
  assign o[1267] = i[2835];
  assign o[1266] = i[2834];
  assign o[1265] = i[2833];
  assign o[1264] = i[2832];
  assign o[1263] = i[2831];
  assign o[1262] = i[2830];
  assign o[1261] = i[2829];
  assign o[1260] = i[2828];
  assign o[1259] = i[2827];
  assign o[1258] = i[2826];
  assign o[1257] = i[2825];
  assign o[1256] = i[2824];
  assign o[1255] = i[2823];
  assign o[1254] = i[2822];
  assign o[1253] = i[2821];
  assign o[1252] = i[2820];
  assign o[1251] = i[2819];
  assign o[1250] = i[2818];
  assign o[1249] = i[2817];
  assign o[1248] = i[2816];
  assign o[1247] = i[2879];
  assign o[1246] = i[2878];
  assign o[1245] = i[2877];
  assign o[1244] = i[2876];
  assign o[1243] = i[2875];
  assign o[1242] = i[2874];
  assign o[1241] = i[2873];
  assign o[1240] = i[2872];
  assign o[1239] = i[2871];
  assign o[1238] = i[2870];
  assign o[1237] = i[2869];
  assign o[1236] = i[2868];
  assign o[1235] = i[2867];
  assign o[1234] = i[2866];
  assign o[1233] = i[2865];
  assign o[1232] = i[2864];
  assign o[1231] = i[2863];
  assign o[1230] = i[2862];
  assign o[1229] = i[2861];
  assign o[1228] = i[2860];
  assign o[1227] = i[2859];
  assign o[1226] = i[2858];
  assign o[1225] = i[2857];
  assign o[1224] = i[2856];
  assign o[1223] = i[2855];
  assign o[1222] = i[2854];
  assign o[1221] = i[2853];
  assign o[1220] = i[2852];
  assign o[1219] = i[2851];
  assign o[1218] = i[2850];
  assign o[1217] = i[2849];
  assign o[1216] = i[2848];
  assign o[1215] = i[2911];
  assign o[1214] = i[2910];
  assign o[1213] = i[2909];
  assign o[1212] = i[2908];
  assign o[1211] = i[2907];
  assign o[1210] = i[2906];
  assign o[1209] = i[2905];
  assign o[1208] = i[2904];
  assign o[1207] = i[2903];
  assign o[1206] = i[2902];
  assign o[1205] = i[2901];
  assign o[1204] = i[2900];
  assign o[1203] = i[2899];
  assign o[1202] = i[2898];
  assign o[1201] = i[2897];
  assign o[1200] = i[2896];
  assign o[1199] = i[2895];
  assign o[1198] = i[2894];
  assign o[1197] = i[2893];
  assign o[1196] = i[2892];
  assign o[1195] = i[2891];
  assign o[1194] = i[2890];
  assign o[1193] = i[2889];
  assign o[1192] = i[2888];
  assign o[1191] = i[2887];
  assign o[1190] = i[2886];
  assign o[1189] = i[2885];
  assign o[1188] = i[2884];
  assign o[1187] = i[2883];
  assign o[1186] = i[2882];
  assign o[1185] = i[2881];
  assign o[1184] = i[2880];
  assign o[1183] = i[2943];
  assign o[1182] = i[2942];
  assign o[1181] = i[2941];
  assign o[1180] = i[2940];
  assign o[1179] = i[2939];
  assign o[1178] = i[2938];
  assign o[1177] = i[2937];
  assign o[1176] = i[2936];
  assign o[1175] = i[2935];
  assign o[1174] = i[2934];
  assign o[1173] = i[2933];
  assign o[1172] = i[2932];
  assign o[1171] = i[2931];
  assign o[1170] = i[2930];
  assign o[1169] = i[2929];
  assign o[1168] = i[2928];
  assign o[1167] = i[2927];
  assign o[1166] = i[2926];
  assign o[1165] = i[2925];
  assign o[1164] = i[2924];
  assign o[1163] = i[2923];
  assign o[1162] = i[2922];
  assign o[1161] = i[2921];
  assign o[1160] = i[2920];
  assign o[1159] = i[2919];
  assign o[1158] = i[2918];
  assign o[1157] = i[2917];
  assign o[1156] = i[2916];
  assign o[1155] = i[2915];
  assign o[1154] = i[2914];
  assign o[1153] = i[2913];
  assign o[1152] = i[2912];
  assign o[1151] = i[2975];
  assign o[1150] = i[2974];
  assign o[1149] = i[2973];
  assign o[1148] = i[2972];
  assign o[1147] = i[2971];
  assign o[1146] = i[2970];
  assign o[1145] = i[2969];
  assign o[1144] = i[2968];
  assign o[1143] = i[2967];
  assign o[1142] = i[2966];
  assign o[1141] = i[2965];
  assign o[1140] = i[2964];
  assign o[1139] = i[2963];
  assign o[1138] = i[2962];
  assign o[1137] = i[2961];
  assign o[1136] = i[2960];
  assign o[1135] = i[2959];
  assign o[1134] = i[2958];
  assign o[1133] = i[2957];
  assign o[1132] = i[2956];
  assign o[1131] = i[2955];
  assign o[1130] = i[2954];
  assign o[1129] = i[2953];
  assign o[1128] = i[2952];
  assign o[1127] = i[2951];
  assign o[1126] = i[2950];
  assign o[1125] = i[2949];
  assign o[1124] = i[2948];
  assign o[1123] = i[2947];
  assign o[1122] = i[2946];
  assign o[1121] = i[2945];
  assign o[1120] = i[2944];
  assign o[1119] = i[3007];
  assign o[1118] = i[3006];
  assign o[1117] = i[3005];
  assign o[1116] = i[3004];
  assign o[1115] = i[3003];
  assign o[1114] = i[3002];
  assign o[1113] = i[3001];
  assign o[1112] = i[3000];
  assign o[1111] = i[2999];
  assign o[1110] = i[2998];
  assign o[1109] = i[2997];
  assign o[1108] = i[2996];
  assign o[1107] = i[2995];
  assign o[1106] = i[2994];
  assign o[1105] = i[2993];
  assign o[1104] = i[2992];
  assign o[1103] = i[2991];
  assign o[1102] = i[2990];
  assign o[1101] = i[2989];
  assign o[1100] = i[2988];
  assign o[1099] = i[2987];
  assign o[1098] = i[2986];
  assign o[1097] = i[2985];
  assign o[1096] = i[2984];
  assign o[1095] = i[2983];
  assign o[1094] = i[2982];
  assign o[1093] = i[2981];
  assign o[1092] = i[2980];
  assign o[1091] = i[2979];
  assign o[1090] = i[2978];
  assign o[1089] = i[2977];
  assign o[1088] = i[2976];
  assign o[1087] = i[3039];
  assign o[1086] = i[3038];
  assign o[1085] = i[3037];
  assign o[1084] = i[3036];
  assign o[1083] = i[3035];
  assign o[1082] = i[3034];
  assign o[1081] = i[3033];
  assign o[1080] = i[3032];
  assign o[1079] = i[3031];
  assign o[1078] = i[3030];
  assign o[1077] = i[3029];
  assign o[1076] = i[3028];
  assign o[1075] = i[3027];
  assign o[1074] = i[3026];
  assign o[1073] = i[3025];
  assign o[1072] = i[3024];
  assign o[1071] = i[3023];
  assign o[1070] = i[3022];
  assign o[1069] = i[3021];
  assign o[1068] = i[3020];
  assign o[1067] = i[3019];
  assign o[1066] = i[3018];
  assign o[1065] = i[3017];
  assign o[1064] = i[3016];
  assign o[1063] = i[3015];
  assign o[1062] = i[3014];
  assign o[1061] = i[3013];
  assign o[1060] = i[3012];
  assign o[1059] = i[3011];
  assign o[1058] = i[3010];
  assign o[1057] = i[3009];
  assign o[1056] = i[3008];
  assign o[1055] = i[3071];
  assign o[1054] = i[3070];
  assign o[1053] = i[3069];
  assign o[1052] = i[3068];
  assign o[1051] = i[3067];
  assign o[1050] = i[3066];
  assign o[1049] = i[3065];
  assign o[1048] = i[3064];
  assign o[1047] = i[3063];
  assign o[1046] = i[3062];
  assign o[1045] = i[3061];
  assign o[1044] = i[3060];
  assign o[1043] = i[3059];
  assign o[1042] = i[3058];
  assign o[1041] = i[3057];
  assign o[1040] = i[3056];
  assign o[1039] = i[3055];
  assign o[1038] = i[3054];
  assign o[1037] = i[3053];
  assign o[1036] = i[3052];
  assign o[1035] = i[3051];
  assign o[1034] = i[3050];
  assign o[1033] = i[3049];
  assign o[1032] = i[3048];
  assign o[1031] = i[3047];
  assign o[1030] = i[3046];
  assign o[1029] = i[3045];
  assign o[1028] = i[3044];
  assign o[1027] = i[3043];
  assign o[1026] = i[3042];
  assign o[1025] = i[3041];
  assign o[1024] = i[3040];
  assign o[1023] = i[3103];
  assign o[1022] = i[3102];
  assign o[1021] = i[3101];
  assign o[1020] = i[3100];
  assign o[1019] = i[3099];
  assign o[1018] = i[3098];
  assign o[1017] = i[3097];
  assign o[1016] = i[3096];
  assign o[1015] = i[3095];
  assign o[1014] = i[3094];
  assign o[1013] = i[3093];
  assign o[1012] = i[3092];
  assign o[1011] = i[3091];
  assign o[1010] = i[3090];
  assign o[1009] = i[3089];
  assign o[1008] = i[3088];
  assign o[1007] = i[3087];
  assign o[1006] = i[3086];
  assign o[1005] = i[3085];
  assign o[1004] = i[3084];
  assign o[1003] = i[3083];
  assign o[1002] = i[3082];
  assign o[1001] = i[3081];
  assign o[1000] = i[3080];
  assign o[999] = i[3079];
  assign o[998] = i[3078];
  assign o[997] = i[3077];
  assign o[996] = i[3076];
  assign o[995] = i[3075];
  assign o[994] = i[3074];
  assign o[993] = i[3073];
  assign o[992] = i[3072];
  assign o[991] = i[3135];
  assign o[990] = i[3134];
  assign o[989] = i[3133];
  assign o[988] = i[3132];
  assign o[987] = i[3131];
  assign o[986] = i[3130];
  assign o[985] = i[3129];
  assign o[984] = i[3128];
  assign o[983] = i[3127];
  assign o[982] = i[3126];
  assign o[981] = i[3125];
  assign o[980] = i[3124];
  assign o[979] = i[3123];
  assign o[978] = i[3122];
  assign o[977] = i[3121];
  assign o[976] = i[3120];
  assign o[975] = i[3119];
  assign o[974] = i[3118];
  assign o[973] = i[3117];
  assign o[972] = i[3116];
  assign o[971] = i[3115];
  assign o[970] = i[3114];
  assign o[969] = i[3113];
  assign o[968] = i[3112];
  assign o[967] = i[3111];
  assign o[966] = i[3110];
  assign o[965] = i[3109];
  assign o[964] = i[3108];
  assign o[963] = i[3107];
  assign o[962] = i[3106];
  assign o[961] = i[3105];
  assign o[960] = i[3104];
  assign o[959] = i[3167];
  assign o[958] = i[3166];
  assign o[957] = i[3165];
  assign o[956] = i[3164];
  assign o[955] = i[3163];
  assign o[954] = i[3162];
  assign o[953] = i[3161];
  assign o[952] = i[3160];
  assign o[951] = i[3159];
  assign o[950] = i[3158];
  assign o[949] = i[3157];
  assign o[948] = i[3156];
  assign o[947] = i[3155];
  assign o[946] = i[3154];
  assign o[945] = i[3153];
  assign o[944] = i[3152];
  assign o[943] = i[3151];
  assign o[942] = i[3150];
  assign o[941] = i[3149];
  assign o[940] = i[3148];
  assign o[939] = i[3147];
  assign o[938] = i[3146];
  assign o[937] = i[3145];
  assign o[936] = i[3144];
  assign o[935] = i[3143];
  assign o[934] = i[3142];
  assign o[933] = i[3141];
  assign o[932] = i[3140];
  assign o[931] = i[3139];
  assign o[930] = i[3138];
  assign o[929] = i[3137];
  assign o[928] = i[3136];
  assign o[927] = i[3199];
  assign o[926] = i[3198];
  assign o[925] = i[3197];
  assign o[924] = i[3196];
  assign o[923] = i[3195];
  assign o[922] = i[3194];
  assign o[921] = i[3193];
  assign o[920] = i[3192];
  assign o[919] = i[3191];
  assign o[918] = i[3190];
  assign o[917] = i[3189];
  assign o[916] = i[3188];
  assign o[915] = i[3187];
  assign o[914] = i[3186];
  assign o[913] = i[3185];
  assign o[912] = i[3184];
  assign o[911] = i[3183];
  assign o[910] = i[3182];
  assign o[909] = i[3181];
  assign o[908] = i[3180];
  assign o[907] = i[3179];
  assign o[906] = i[3178];
  assign o[905] = i[3177];
  assign o[904] = i[3176];
  assign o[903] = i[3175];
  assign o[902] = i[3174];
  assign o[901] = i[3173];
  assign o[900] = i[3172];
  assign o[899] = i[3171];
  assign o[898] = i[3170];
  assign o[897] = i[3169];
  assign o[896] = i[3168];
  assign o[895] = i[3231];
  assign o[894] = i[3230];
  assign o[893] = i[3229];
  assign o[892] = i[3228];
  assign o[891] = i[3227];
  assign o[890] = i[3226];
  assign o[889] = i[3225];
  assign o[888] = i[3224];
  assign o[887] = i[3223];
  assign o[886] = i[3222];
  assign o[885] = i[3221];
  assign o[884] = i[3220];
  assign o[883] = i[3219];
  assign o[882] = i[3218];
  assign o[881] = i[3217];
  assign o[880] = i[3216];
  assign o[879] = i[3215];
  assign o[878] = i[3214];
  assign o[877] = i[3213];
  assign o[876] = i[3212];
  assign o[875] = i[3211];
  assign o[874] = i[3210];
  assign o[873] = i[3209];
  assign o[872] = i[3208];
  assign o[871] = i[3207];
  assign o[870] = i[3206];
  assign o[869] = i[3205];
  assign o[868] = i[3204];
  assign o[867] = i[3203];
  assign o[866] = i[3202];
  assign o[865] = i[3201];
  assign o[864] = i[3200];
  assign o[863] = i[3263];
  assign o[862] = i[3262];
  assign o[861] = i[3261];
  assign o[860] = i[3260];
  assign o[859] = i[3259];
  assign o[858] = i[3258];
  assign o[857] = i[3257];
  assign o[856] = i[3256];
  assign o[855] = i[3255];
  assign o[854] = i[3254];
  assign o[853] = i[3253];
  assign o[852] = i[3252];
  assign o[851] = i[3251];
  assign o[850] = i[3250];
  assign o[849] = i[3249];
  assign o[848] = i[3248];
  assign o[847] = i[3247];
  assign o[846] = i[3246];
  assign o[845] = i[3245];
  assign o[844] = i[3244];
  assign o[843] = i[3243];
  assign o[842] = i[3242];
  assign o[841] = i[3241];
  assign o[840] = i[3240];
  assign o[839] = i[3239];
  assign o[838] = i[3238];
  assign o[837] = i[3237];
  assign o[836] = i[3236];
  assign o[835] = i[3235];
  assign o[834] = i[3234];
  assign o[833] = i[3233];
  assign o[832] = i[3232];
  assign o[831] = i[3295];
  assign o[830] = i[3294];
  assign o[829] = i[3293];
  assign o[828] = i[3292];
  assign o[827] = i[3291];
  assign o[826] = i[3290];
  assign o[825] = i[3289];
  assign o[824] = i[3288];
  assign o[823] = i[3287];
  assign o[822] = i[3286];
  assign o[821] = i[3285];
  assign o[820] = i[3284];
  assign o[819] = i[3283];
  assign o[818] = i[3282];
  assign o[817] = i[3281];
  assign o[816] = i[3280];
  assign o[815] = i[3279];
  assign o[814] = i[3278];
  assign o[813] = i[3277];
  assign o[812] = i[3276];
  assign o[811] = i[3275];
  assign o[810] = i[3274];
  assign o[809] = i[3273];
  assign o[808] = i[3272];
  assign o[807] = i[3271];
  assign o[806] = i[3270];
  assign o[805] = i[3269];
  assign o[804] = i[3268];
  assign o[803] = i[3267];
  assign o[802] = i[3266];
  assign o[801] = i[3265];
  assign o[800] = i[3264];
  assign o[799] = i[3327];
  assign o[798] = i[3326];
  assign o[797] = i[3325];
  assign o[796] = i[3324];
  assign o[795] = i[3323];
  assign o[794] = i[3322];
  assign o[793] = i[3321];
  assign o[792] = i[3320];
  assign o[791] = i[3319];
  assign o[790] = i[3318];
  assign o[789] = i[3317];
  assign o[788] = i[3316];
  assign o[787] = i[3315];
  assign o[786] = i[3314];
  assign o[785] = i[3313];
  assign o[784] = i[3312];
  assign o[783] = i[3311];
  assign o[782] = i[3310];
  assign o[781] = i[3309];
  assign o[780] = i[3308];
  assign o[779] = i[3307];
  assign o[778] = i[3306];
  assign o[777] = i[3305];
  assign o[776] = i[3304];
  assign o[775] = i[3303];
  assign o[774] = i[3302];
  assign o[773] = i[3301];
  assign o[772] = i[3300];
  assign o[771] = i[3299];
  assign o[770] = i[3298];
  assign o[769] = i[3297];
  assign o[768] = i[3296];
  assign o[767] = i[3359];
  assign o[766] = i[3358];
  assign o[765] = i[3357];
  assign o[764] = i[3356];
  assign o[763] = i[3355];
  assign o[762] = i[3354];
  assign o[761] = i[3353];
  assign o[760] = i[3352];
  assign o[759] = i[3351];
  assign o[758] = i[3350];
  assign o[757] = i[3349];
  assign o[756] = i[3348];
  assign o[755] = i[3347];
  assign o[754] = i[3346];
  assign o[753] = i[3345];
  assign o[752] = i[3344];
  assign o[751] = i[3343];
  assign o[750] = i[3342];
  assign o[749] = i[3341];
  assign o[748] = i[3340];
  assign o[747] = i[3339];
  assign o[746] = i[3338];
  assign o[745] = i[3337];
  assign o[744] = i[3336];
  assign o[743] = i[3335];
  assign o[742] = i[3334];
  assign o[741] = i[3333];
  assign o[740] = i[3332];
  assign o[739] = i[3331];
  assign o[738] = i[3330];
  assign o[737] = i[3329];
  assign o[736] = i[3328];
  assign o[735] = i[3391];
  assign o[734] = i[3390];
  assign o[733] = i[3389];
  assign o[732] = i[3388];
  assign o[731] = i[3387];
  assign o[730] = i[3386];
  assign o[729] = i[3385];
  assign o[728] = i[3384];
  assign o[727] = i[3383];
  assign o[726] = i[3382];
  assign o[725] = i[3381];
  assign o[724] = i[3380];
  assign o[723] = i[3379];
  assign o[722] = i[3378];
  assign o[721] = i[3377];
  assign o[720] = i[3376];
  assign o[719] = i[3375];
  assign o[718] = i[3374];
  assign o[717] = i[3373];
  assign o[716] = i[3372];
  assign o[715] = i[3371];
  assign o[714] = i[3370];
  assign o[713] = i[3369];
  assign o[712] = i[3368];
  assign o[711] = i[3367];
  assign o[710] = i[3366];
  assign o[709] = i[3365];
  assign o[708] = i[3364];
  assign o[707] = i[3363];
  assign o[706] = i[3362];
  assign o[705] = i[3361];
  assign o[704] = i[3360];
  assign o[703] = i[3423];
  assign o[702] = i[3422];
  assign o[701] = i[3421];
  assign o[700] = i[3420];
  assign o[699] = i[3419];
  assign o[698] = i[3418];
  assign o[697] = i[3417];
  assign o[696] = i[3416];
  assign o[695] = i[3415];
  assign o[694] = i[3414];
  assign o[693] = i[3413];
  assign o[692] = i[3412];
  assign o[691] = i[3411];
  assign o[690] = i[3410];
  assign o[689] = i[3409];
  assign o[688] = i[3408];
  assign o[687] = i[3407];
  assign o[686] = i[3406];
  assign o[685] = i[3405];
  assign o[684] = i[3404];
  assign o[683] = i[3403];
  assign o[682] = i[3402];
  assign o[681] = i[3401];
  assign o[680] = i[3400];
  assign o[679] = i[3399];
  assign o[678] = i[3398];
  assign o[677] = i[3397];
  assign o[676] = i[3396];
  assign o[675] = i[3395];
  assign o[674] = i[3394];
  assign o[673] = i[3393];
  assign o[672] = i[3392];
  assign o[671] = i[3455];
  assign o[670] = i[3454];
  assign o[669] = i[3453];
  assign o[668] = i[3452];
  assign o[667] = i[3451];
  assign o[666] = i[3450];
  assign o[665] = i[3449];
  assign o[664] = i[3448];
  assign o[663] = i[3447];
  assign o[662] = i[3446];
  assign o[661] = i[3445];
  assign o[660] = i[3444];
  assign o[659] = i[3443];
  assign o[658] = i[3442];
  assign o[657] = i[3441];
  assign o[656] = i[3440];
  assign o[655] = i[3439];
  assign o[654] = i[3438];
  assign o[653] = i[3437];
  assign o[652] = i[3436];
  assign o[651] = i[3435];
  assign o[650] = i[3434];
  assign o[649] = i[3433];
  assign o[648] = i[3432];
  assign o[647] = i[3431];
  assign o[646] = i[3430];
  assign o[645] = i[3429];
  assign o[644] = i[3428];
  assign o[643] = i[3427];
  assign o[642] = i[3426];
  assign o[641] = i[3425];
  assign o[640] = i[3424];
  assign o[639] = i[3487];
  assign o[638] = i[3486];
  assign o[637] = i[3485];
  assign o[636] = i[3484];
  assign o[635] = i[3483];
  assign o[634] = i[3482];
  assign o[633] = i[3481];
  assign o[632] = i[3480];
  assign o[631] = i[3479];
  assign o[630] = i[3478];
  assign o[629] = i[3477];
  assign o[628] = i[3476];
  assign o[627] = i[3475];
  assign o[626] = i[3474];
  assign o[625] = i[3473];
  assign o[624] = i[3472];
  assign o[623] = i[3471];
  assign o[622] = i[3470];
  assign o[621] = i[3469];
  assign o[620] = i[3468];
  assign o[619] = i[3467];
  assign o[618] = i[3466];
  assign o[617] = i[3465];
  assign o[616] = i[3464];
  assign o[615] = i[3463];
  assign o[614] = i[3462];
  assign o[613] = i[3461];
  assign o[612] = i[3460];
  assign o[611] = i[3459];
  assign o[610] = i[3458];
  assign o[609] = i[3457];
  assign o[608] = i[3456];
  assign o[607] = i[3519];
  assign o[606] = i[3518];
  assign o[605] = i[3517];
  assign o[604] = i[3516];
  assign o[603] = i[3515];
  assign o[602] = i[3514];
  assign o[601] = i[3513];
  assign o[600] = i[3512];
  assign o[599] = i[3511];
  assign o[598] = i[3510];
  assign o[597] = i[3509];
  assign o[596] = i[3508];
  assign o[595] = i[3507];
  assign o[594] = i[3506];
  assign o[593] = i[3505];
  assign o[592] = i[3504];
  assign o[591] = i[3503];
  assign o[590] = i[3502];
  assign o[589] = i[3501];
  assign o[588] = i[3500];
  assign o[587] = i[3499];
  assign o[586] = i[3498];
  assign o[585] = i[3497];
  assign o[584] = i[3496];
  assign o[583] = i[3495];
  assign o[582] = i[3494];
  assign o[581] = i[3493];
  assign o[580] = i[3492];
  assign o[579] = i[3491];
  assign o[578] = i[3490];
  assign o[577] = i[3489];
  assign o[576] = i[3488];
  assign o[575] = i[3551];
  assign o[574] = i[3550];
  assign o[573] = i[3549];
  assign o[572] = i[3548];
  assign o[571] = i[3547];
  assign o[570] = i[3546];
  assign o[569] = i[3545];
  assign o[568] = i[3544];
  assign o[567] = i[3543];
  assign o[566] = i[3542];
  assign o[565] = i[3541];
  assign o[564] = i[3540];
  assign o[563] = i[3539];
  assign o[562] = i[3538];
  assign o[561] = i[3537];
  assign o[560] = i[3536];
  assign o[559] = i[3535];
  assign o[558] = i[3534];
  assign o[557] = i[3533];
  assign o[556] = i[3532];
  assign o[555] = i[3531];
  assign o[554] = i[3530];
  assign o[553] = i[3529];
  assign o[552] = i[3528];
  assign o[551] = i[3527];
  assign o[550] = i[3526];
  assign o[549] = i[3525];
  assign o[548] = i[3524];
  assign o[547] = i[3523];
  assign o[546] = i[3522];
  assign o[545] = i[3521];
  assign o[544] = i[3520];
  assign o[543] = i[3583];
  assign o[542] = i[3582];
  assign o[541] = i[3581];
  assign o[540] = i[3580];
  assign o[539] = i[3579];
  assign o[538] = i[3578];
  assign o[537] = i[3577];
  assign o[536] = i[3576];
  assign o[535] = i[3575];
  assign o[534] = i[3574];
  assign o[533] = i[3573];
  assign o[532] = i[3572];
  assign o[531] = i[3571];
  assign o[530] = i[3570];
  assign o[529] = i[3569];
  assign o[528] = i[3568];
  assign o[527] = i[3567];
  assign o[526] = i[3566];
  assign o[525] = i[3565];
  assign o[524] = i[3564];
  assign o[523] = i[3563];
  assign o[522] = i[3562];
  assign o[521] = i[3561];
  assign o[520] = i[3560];
  assign o[519] = i[3559];
  assign o[518] = i[3558];
  assign o[517] = i[3557];
  assign o[516] = i[3556];
  assign o[515] = i[3555];
  assign o[514] = i[3554];
  assign o[513] = i[3553];
  assign o[512] = i[3552];
  assign o[511] = i[3615];
  assign o[510] = i[3614];
  assign o[509] = i[3613];
  assign o[508] = i[3612];
  assign o[507] = i[3611];
  assign o[506] = i[3610];
  assign o[505] = i[3609];
  assign o[504] = i[3608];
  assign o[503] = i[3607];
  assign o[502] = i[3606];
  assign o[501] = i[3605];
  assign o[500] = i[3604];
  assign o[499] = i[3603];
  assign o[498] = i[3602];
  assign o[497] = i[3601];
  assign o[496] = i[3600];
  assign o[495] = i[3599];
  assign o[494] = i[3598];
  assign o[493] = i[3597];
  assign o[492] = i[3596];
  assign o[491] = i[3595];
  assign o[490] = i[3594];
  assign o[489] = i[3593];
  assign o[488] = i[3592];
  assign o[487] = i[3591];
  assign o[486] = i[3590];
  assign o[485] = i[3589];
  assign o[484] = i[3588];
  assign o[483] = i[3587];
  assign o[482] = i[3586];
  assign o[481] = i[3585];
  assign o[480] = i[3584];
  assign o[479] = i[3647];
  assign o[478] = i[3646];
  assign o[477] = i[3645];
  assign o[476] = i[3644];
  assign o[475] = i[3643];
  assign o[474] = i[3642];
  assign o[473] = i[3641];
  assign o[472] = i[3640];
  assign o[471] = i[3639];
  assign o[470] = i[3638];
  assign o[469] = i[3637];
  assign o[468] = i[3636];
  assign o[467] = i[3635];
  assign o[466] = i[3634];
  assign o[465] = i[3633];
  assign o[464] = i[3632];
  assign o[463] = i[3631];
  assign o[462] = i[3630];
  assign o[461] = i[3629];
  assign o[460] = i[3628];
  assign o[459] = i[3627];
  assign o[458] = i[3626];
  assign o[457] = i[3625];
  assign o[456] = i[3624];
  assign o[455] = i[3623];
  assign o[454] = i[3622];
  assign o[453] = i[3621];
  assign o[452] = i[3620];
  assign o[451] = i[3619];
  assign o[450] = i[3618];
  assign o[449] = i[3617];
  assign o[448] = i[3616];
  assign o[447] = i[3679];
  assign o[446] = i[3678];
  assign o[445] = i[3677];
  assign o[444] = i[3676];
  assign o[443] = i[3675];
  assign o[442] = i[3674];
  assign o[441] = i[3673];
  assign o[440] = i[3672];
  assign o[439] = i[3671];
  assign o[438] = i[3670];
  assign o[437] = i[3669];
  assign o[436] = i[3668];
  assign o[435] = i[3667];
  assign o[434] = i[3666];
  assign o[433] = i[3665];
  assign o[432] = i[3664];
  assign o[431] = i[3663];
  assign o[430] = i[3662];
  assign o[429] = i[3661];
  assign o[428] = i[3660];
  assign o[427] = i[3659];
  assign o[426] = i[3658];
  assign o[425] = i[3657];
  assign o[424] = i[3656];
  assign o[423] = i[3655];
  assign o[422] = i[3654];
  assign o[421] = i[3653];
  assign o[420] = i[3652];
  assign o[419] = i[3651];
  assign o[418] = i[3650];
  assign o[417] = i[3649];
  assign o[416] = i[3648];
  assign o[415] = i[3711];
  assign o[414] = i[3710];
  assign o[413] = i[3709];
  assign o[412] = i[3708];
  assign o[411] = i[3707];
  assign o[410] = i[3706];
  assign o[409] = i[3705];
  assign o[408] = i[3704];
  assign o[407] = i[3703];
  assign o[406] = i[3702];
  assign o[405] = i[3701];
  assign o[404] = i[3700];
  assign o[403] = i[3699];
  assign o[402] = i[3698];
  assign o[401] = i[3697];
  assign o[400] = i[3696];
  assign o[399] = i[3695];
  assign o[398] = i[3694];
  assign o[397] = i[3693];
  assign o[396] = i[3692];
  assign o[395] = i[3691];
  assign o[394] = i[3690];
  assign o[393] = i[3689];
  assign o[392] = i[3688];
  assign o[391] = i[3687];
  assign o[390] = i[3686];
  assign o[389] = i[3685];
  assign o[388] = i[3684];
  assign o[387] = i[3683];
  assign o[386] = i[3682];
  assign o[385] = i[3681];
  assign o[384] = i[3680];
  assign o[383] = i[3743];
  assign o[382] = i[3742];
  assign o[381] = i[3741];
  assign o[380] = i[3740];
  assign o[379] = i[3739];
  assign o[378] = i[3738];
  assign o[377] = i[3737];
  assign o[376] = i[3736];
  assign o[375] = i[3735];
  assign o[374] = i[3734];
  assign o[373] = i[3733];
  assign o[372] = i[3732];
  assign o[371] = i[3731];
  assign o[370] = i[3730];
  assign o[369] = i[3729];
  assign o[368] = i[3728];
  assign o[367] = i[3727];
  assign o[366] = i[3726];
  assign o[365] = i[3725];
  assign o[364] = i[3724];
  assign o[363] = i[3723];
  assign o[362] = i[3722];
  assign o[361] = i[3721];
  assign o[360] = i[3720];
  assign o[359] = i[3719];
  assign o[358] = i[3718];
  assign o[357] = i[3717];
  assign o[356] = i[3716];
  assign o[355] = i[3715];
  assign o[354] = i[3714];
  assign o[353] = i[3713];
  assign o[352] = i[3712];
  assign o[351] = i[3775];
  assign o[350] = i[3774];
  assign o[349] = i[3773];
  assign o[348] = i[3772];
  assign o[347] = i[3771];
  assign o[346] = i[3770];
  assign o[345] = i[3769];
  assign o[344] = i[3768];
  assign o[343] = i[3767];
  assign o[342] = i[3766];
  assign o[341] = i[3765];
  assign o[340] = i[3764];
  assign o[339] = i[3763];
  assign o[338] = i[3762];
  assign o[337] = i[3761];
  assign o[336] = i[3760];
  assign o[335] = i[3759];
  assign o[334] = i[3758];
  assign o[333] = i[3757];
  assign o[332] = i[3756];
  assign o[331] = i[3755];
  assign o[330] = i[3754];
  assign o[329] = i[3753];
  assign o[328] = i[3752];
  assign o[327] = i[3751];
  assign o[326] = i[3750];
  assign o[325] = i[3749];
  assign o[324] = i[3748];
  assign o[323] = i[3747];
  assign o[322] = i[3746];
  assign o[321] = i[3745];
  assign o[320] = i[3744];
  assign o[319] = i[3807];
  assign o[318] = i[3806];
  assign o[317] = i[3805];
  assign o[316] = i[3804];
  assign o[315] = i[3803];
  assign o[314] = i[3802];
  assign o[313] = i[3801];
  assign o[312] = i[3800];
  assign o[311] = i[3799];
  assign o[310] = i[3798];
  assign o[309] = i[3797];
  assign o[308] = i[3796];
  assign o[307] = i[3795];
  assign o[306] = i[3794];
  assign o[305] = i[3793];
  assign o[304] = i[3792];
  assign o[303] = i[3791];
  assign o[302] = i[3790];
  assign o[301] = i[3789];
  assign o[300] = i[3788];
  assign o[299] = i[3787];
  assign o[298] = i[3786];
  assign o[297] = i[3785];
  assign o[296] = i[3784];
  assign o[295] = i[3783];
  assign o[294] = i[3782];
  assign o[293] = i[3781];
  assign o[292] = i[3780];
  assign o[291] = i[3779];
  assign o[290] = i[3778];
  assign o[289] = i[3777];
  assign o[288] = i[3776];
  assign o[287] = i[3839];
  assign o[286] = i[3838];
  assign o[285] = i[3837];
  assign o[284] = i[3836];
  assign o[283] = i[3835];
  assign o[282] = i[3834];
  assign o[281] = i[3833];
  assign o[280] = i[3832];
  assign o[279] = i[3831];
  assign o[278] = i[3830];
  assign o[277] = i[3829];
  assign o[276] = i[3828];
  assign o[275] = i[3827];
  assign o[274] = i[3826];
  assign o[273] = i[3825];
  assign o[272] = i[3824];
  assign o[271] = i[3823];
  assign o[270] = i[3822];
  assign o[269] = i[3821];
  assign o[268] = i[3820];
  assign o[267] = i[3819];
  assign o[266] = i[3818];
  assign o[265] = i[3817];
  assign o[264] = i[3816];
  assign o[263] = i[3815];
  assign o[262] = i[3814];
  assign o[261] = i[3813];
  assign o[260] = i[3812];
  assign o[259] = i[3811];
  assign o[258] = i[3810];
  assign o[257] = i[3809];
  assign o[256] = i[3808];
  assign o[255] = i[3871];
  assign o[254] = i[3870];
  assign o[253] = i[3869];
  assign o[252] = i[3868];
  assign o[251] = i[3867];
  assign o[250] = i[3866];
  assign o[249] = i[3865];
  assign o[248] = i[3864];
  assign o[247] = i[3863];
  assign o[246] = i[3862];
  assign o[245] = i[3861];
  assign o[244] = i[3860];
  assign o[243] = i[3859];
  assign o[242] = i[3858];
  assign o[241] = i[3857];
  assign o[240] = i[3856];
  assign o[239] = i[3855];
  assign o[238] = i[3854];
  assign o[237] = i[3853];
  assign o[236] = i[3852];
  assign o[235] = i[3851];
  assign o[234] = i[3850];
  assign o[233] = i[3849];
  assign o[232] = i[3848];
  assign o[231] = i[3847];
  assign o[230] = i[3846];
  assign o[229] = i[3845];
  assign o[228] = i[3844];
  assign o[227] = i[3843];
  assign o[226] = i[3842];
  assign o[225] = i[3841];
  assign o[224] = i[3840];
  assign o[223] = i[3903];
  assign o[222] = i[3902];
  assign o[221] = i[3901];
  assign o[220] = i[3900];
  assign o[219] = i[3899];
  assign o[218] = i[3898];
  assign o[217] = i[3897];
  assign o[216] = i[3896];
  assign o[215] = i[3895];
  assign o[214] = i[3894];
  assign o[213] = i[3893];
  assign o[212] = i[3892];
  assign o[211] = i[3891];
  assign o[210] = i[3890];
  assign o[209] = i[3889];
  assign o[208] = i[3888];
  assign o[207] = i[3887];
  assign o[206] = i[3886];
  assign o[205] = i[3885];
  assign o[204] = i[3884];
  assign o[203] = i[3883];
  assign o[202] = i[3882];
  assign o[201] = i[3881];
  assign o[200] = i[3880];
  assign o[199] = i[3879];
  assign o[198] = i[3878];
  assign o[197] = i[3877];
  assign o[196] = i[3876];
  assign o[195] = i[3875];
  assign o[194] = i[3874];
  assign o[193] = i[3873];
  assign o[192] = i[3872];
  assign o[191] = i[3935];
  assign o[190] = i[3934];
  assign o[189] = i[3933];
  assign o[188] = i[3932];
  assign o[187] = i[3931];
  assign o[186] = i[3930];
  assign o[185] = i[3929];
  assign o[184] = i[3928];
  assign o[183] = i[3927];
  assign o[182] = i[3926];
  assign o[181] = i[3925];
  assign o[180] = i[3924];
  assign o[179] = i[3923];
  assign o[178] = i[3922];
  assign o[177] = i[3921];
  assign o[176] = i[3920];
  assign o[175] = i[3919];
  assign o[174] = i[3918];
  assign o[173] = i[3917];
  assign o[172] = i[3916];
  assign o[171] = i[3915];
  assign o[170] = i[3914];
  assign o[169] = i[3913];
  assign o[168] = i[3912];
  assign o[167] = i[3911];
  assign o[166] = i[3910];
  assign o[165] = i[3909];
  assign o[164] = i[3908];
  assign o[163] = i[3907];
  assign o[162] = i[3906];
  assign o[161] = i[3905];
  assign o[160] = i[3904];
  assign o[159] = i[3967];
  assign o[158] = i[3966];
  assign o[157] = i[3965];
  assign o[156] = i[3964];
  assign o[155] = i[3963];
  assign o[154] = i[3962];
  assign o[153] = i[3961];
  assign o[152] = i[3960];
  assign o[151] = i[3959];
  assign o[150] = i[3958];
  assign o[149] = i[3957];
  assign o[148] = i[3956];
  assign o[147] = i[3955];
  assign o[146] = i[3954];
  assign o[145] = i[3953];
  assign o[144] = i[3952];
  assign o[143] = i[3951];
  assign o[142] = i[3950];
  assign o[141] = i[3949];
  assign o[140] = i[3948];
  assign o[139] = i[3947];
  assign o[138] = i[3946];
  assign o[137] = i[3945];
  assign o[136] = i[3944];
  assign o[135] = i[3943];
  assign o[134] = i[3942];
  assign o[133] = i[3941];
  assign o[132] = i[3940];
  assign o[131] = i[3939];
  assign o[130] = i[3938];
  assign o[129] = i[3937];
  assign o[128] = i[3936];
  assign o[127] = i[3999];
  assign o[126] = i[3998];
  assign o[125] = i[3997];
  assign o[124] = i[3996];
  assign o[123] = i[3995];
  assign o[122] = i[3994];
  assign o[121] = i[3993];
  assign o[120] = i[3992];
  assign o[119] = i[3991];
  assign o[118] = i[3990];
  assign o[117] = i[3989];
  assign o[116] = i[3988];
  assign o[115] = i[3987];
  assign o[114] = i[3986];
  assign o[113] = i[3985];
  assign o[112] = i[3984];
  assign o[111] = i[3983];
  assign o[110] = i[3982];
  assign o[109] = i[3981];
  assign o[108] = i[3980];
  assign o[107] = i[3979];
  assign o[106] = i[3978];
  assign o[105] = i[3977];
  assign o[104] = i[3976];
  assign o[103] = i[3975];
  assign o[102] = i[3974];
  assign o[101] = i[3973];
  assign o[100] = i[3972];
  assign o[99] = i[3971];
  assign o[98] = i[3970];
  assign o[97] = i[3969];
  assign o[96] = i[3968];
  assign o[95] = i[4031];
  assign o[94] = i[4030];
  assign o[93] = i[4029];
  assign o[92] = i[4028];
  assign o[91] = i[4027];
  assign o[90] = i[4026];
  assign o[89] = i[4025];
  assign o[88] = i[4024];
  assign o[87] = i[4023];
  assign o[86] = i[4022];
  assign o[85] = i[4021];
  assign o[84] = i[4020];
  assign o[83] = i[4019];
  assign o[82] = i[4018];
  assign o[81] = i[4017];
  assign o[80] = i[4016];
  assign o[79] = i[4015];
  assign o[78] = i[4014];
  assign o[77] = i[4013];
  assign o[76] = i[4012];
  assign o[75] = i[4011];
  assign o[74] = i[4010];
  assign o[73] = i[4009];
  assign o[72] = i[4008];
  assign o[71] = i[4007];
  assign o[70] = i[4006];
  assign o[69] = i[4005];
  assign o[68] = i[4004];
  assign o[67] = i[4003];
  assign o[66] = i[4002];
  assign o[65] = i[4001];
  assign o[64] = i[4000];
  assign o[63] = i[4063];
  assign o[62] = i[4062];
  assign o[61] = i[4061];
  assign o[60] = i[4060];
  assign o[59] = i[4059];
  assign o[58] = i[4058];
  assign o[57] = i[4057];
  assign o[56] = i[4056];
  assign o[55] = i[4055];
  assign o[54] = i[4054];
  assign o[53] = i[4053];
  assign o[52] = i[4052];
  assign o[51] = i[4051];
  assign o[50] = i[4050];
  assign o[49] = i[4049];
  assign o[48] = i[4048];
  assign o[47] = i[4047];
  assign o[46] = i[4046];
  assign o[45] = i[4045];
  assign o[44] = i[4044];
  assign o[43] = i[4043];
  assign o[42] = i[4042];
  assign o[41] = i[4041];
  assign o[40] = i[4040];
  assign o[39] = i[4039];
  assign o[38] = i[4038];
  assign o[37] = i[4037];
  assign o[36] = i[4036];
  assign o[35] = i[4035];
  assign o[34] = i[4034];
  assign o[33] = i[4033];
  assign o[32] = i[4032];
  assign o[31] = i[4095];
  assign o[30] = i[4094];
  assign o[29] = i[4093];
  assign o[28] = i[4092];
  assign o[27] = i[4091];
  assign o[26] = i[4090];
  assign o[25] = i[4089];
  assign o[24] = i[4088];
  assign o[23] = i[4087];
  assign o[22] = i[4086];
  assign o[21] = i[4085];
  assign o[20] = i[4084];
  assign o[19] = i[4083];
  assign o[18] = i[4082];
  assign o[17] = i[4081];
  assign o[16] = i[4080];
  assign o[15] = i[4079];
  assign o[14] = i[4078];
  assign o[13] = i[4077];
  assign o[12] = i[4076];
  assign o[11] = i[4075];
  assign o[10] = i[4074];
  assign o[9] = i[4073];
  assign o[8] = i[4072];
  assign o[7] = i[4071];
  assign o[6] = i[4070];
  assign o[5] = i[4069];
  assign o[4] = i[4068];
  assign o[3] = i[4067];
  assign o[2] = i[4066];
  assign o[1] = i[4065];
  assign o[0] = i[4064];

endmodule



module bsg_parallel_in_serial_out
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_i
);

  input [4095:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_o;
  output valid_o;
  wire [31:0] data_o;
  wire ready_o,valid_o,N0,N1,\piso.done_tx_n ,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,
  N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295;
  wire [6:0] \piso.shift_ctr_r ;
  wire [0:0] \piso.state_n ;
  wire [4095:0] \piso.data_li ,\piso.data_r ;
  reg valid_o_sv2v_reg,\piso.data_r_4095_sv2v_reg ,\piso.data_r_4094_sv2v_reg ,
  \piso.data_r_4093_sv2v_reg ,\piso.data_r_4092_sv2v_reg ,\piso.data_r_4091_sv2v_reg ,
  \piso.data_r_4090_sv2v_reg ,\piso.data_r_4089_sv2v_reg ,
  \piso.data_r_4088_sv2v_reg ,\piso.data_r_4087_sv2v_reg ,\piso.data_r_4086_sv2v_reg ,
  \piso.data_r_4085_sv2v_reg ,\piso.data_r_4084_sv2v_reg ,\piso.data_r_4083_sv2v_reg ,
  \piso.data_r_4082_sv2v_reg ,\piso.data_r_4081_sv2v_reg ,\piso.data_r_4080_sv2v_reg ,
  \piso.data_r_4079_sv2v_reg ,\piso.data_r_4078_sv2v_reg ,\piso.data_r_4077_sv2v_reg ,
  \piso.data_r_4076_sv2v_reg ,\piso.data_r_4075_sv2v_reg ,\piso.data_r_4074_sv2v_reg ,
  \piso.data_r_4073_sv2v_reg ,\piso.data_r_4072_sv2v_reg ,\piso.data_r_4071_sv2v_reg ,
  \piso.data_r_4070_sv2v_reg ,\piso.data_r_4069_sv2v_reg ,
  \piso.data_r_4068_sv2v_reg ,\piso.data_r_4067_sv2v_reg ,\piso.data_r_4066_sv2v_reg ,
  \piso.data_r_4065_sv2v_reg ,\piso.data_r_4064_sv2v_reg ,\piso.data_r_4063_sv2v_reg ,
  \piso.data_r_4062_sv2v_reg ,\piso.data_r_4061_sv2v_reg ,\piso.data_r_4060_sv2v_reg ,
  \piso.data_r_4059_sv2v_reg ,\piso.data_r_4058_sv2v_reg ,\piso.data_r_4057_sv2v_reg ,
  \piso.data_r_4056_sv2v_reg ,\piso.data_r_4055_sv2v_reg ,\piso.data_r_4054_sv2v_reg ,
  \piso.data_r_4053_sv2v_reg ,\piso.data_r_4052_sv2v_reg ,\piso.data_r_4051_sv2v_reg ,
  \piso.data_r_4050_sv2v_reg ,\piso.data_r_4049_sv2v_reg ,
  \piso.data_r_4048_sv2v_reg ,\piso.data_r_4047_sv2v_reg ,\piso.data_r_4046_sv2v_reg ,
  \piso.data_r_4045_sv2v_reg ,\piso.data_r_4044_sv2v_reg ,\piso.data_r_4043_sv2v_reg ,
  \piso.data_r_4042_sv2v_reg ,\piso.data_r_4041_sv2v_reg ,\piso.data_r_4040_sv2v_reg ,
  \piso.data_r_4039_sv2v_reg ,\piso.data_r_4038_sv2v_reg ,\piso.data_r_4037_sv2v_reg ,
  \piso.data_r_4036_sv2v_reg ,\piso.data_r_4035_sv2v_reg ,\piso.data_r_4034_sv2v_reg ,
  \piso.data_r_4033_sv2v_reg ,\piso.data_r_4032_sv2v_reg ,\piso.data_r_4031_sv2v_reg ,
  \piso.data_r_4030_sv2v_reg ,\piso.data_r_4029_sv2v_reg ,
  \piso.data_r_4028_sv2v_reg ,\piso.data_r_4027_sv2v_reg ,\piso.data_r_4026_sv2v_reg ,
  \piso.data_r_4025_sv2v_reg ,\piso.data_r_4024_sv2v_reg ,\piso.data_r_4023_sv2v_reg ,
  \piso.data_r_4022_sv2v_reg ,\piso.data_r_4021_sv2v_reg ,\piso.data_r_4020_sv2v_reg ,
  \piso.data_r_4019_sv2v_reg ,\piso.data_r_4018_sv2v_reg ,\piso.data_r_4017_sv2v_reg ,
  \piso.data_r_4016_sv2v_reg ,\piso.data_r_4015_sv2v_reg ,\piso.data_r_4014_sv2v_reg ,
  \piso.data_r_4013_sv2v_reg ,\piso.data_r_4012_sv2v_reg ,\piso.data_r_4011_sv2v_reg ,
  \piso.data_r_4010_sv2v_reg ,\piso.data_r_4009_sv2v_reg ,
  \piso.data_r_4008_sv2v_reg ,\piso.data_r_4007_sv2v_reg ,\piso.data_r_4006_sv2v_reg ,
  \piso.data_r_4005_sv2v_reg ,\piso.data_r_4004_sv2v_reg ,\piso.data_r_4003_sv2v_reg ,
  \piso.data_r_4002_sv2v_reg ,\piso.data_r_4001_sv2v_reg ,\piso.data_r_4000_sv2v_reg ,
  \piso.data_r_3999_sv2v_reg ,\piso.data_r_3998_sv2v_reg ,\piso.data_r_3997_sv2v_reg ,
  \piso.data_r_3996_sv2v_reg ,\piso.data_r_3995_sv2v_reg ,\piso.data_r_3994_sv2v_reg ,
  \piso.data_r_3993_sv2v_reg ,\piso.data_r_3992_sv2v_reg ,\piso.data_r_3991_sv2v_reg ,
  \piso.data_r_3990_sv2v_reg ,\piso.data_r_3989_sv2v_reg ,
  \piso.data_r_3988_sv2v_reg ,\piso.data_r_3987_sv2v_reg ,\piso.data_r_3986_sv2v_reg ,
  \piso.data_r_3985_sv2v_reg ,\piso.data_r_3984_sv2v_reg ,\piso.data_r_3983_sv2v_reg ,
  \piso.data_r_3982_sv2v_reg ,\piso.data_r_3981_sv2v_reg ,\piso.data_r_3980_sv2v_reg ,
  \piso.data_r_3979_sv2v_reg ,\piso.data_r_3978_sv2v_reg ,\piso.data_r_3977_sv2v_reg ,
  \piso.data_r_3976_sv2v_reg ,\piso.data_r_3975_sv2v_reg ,\piso.data_r_3974_sv2v_reg ,
  \piso.data_r_3973_sv2v_reg ,\piso.data_r_3972_sv2v_reg ,\piso.data_r_3971_sv2v_reg ,
  \piso.data_r_3970_sv2v_reg ,\piso.data_r_3969_sv2v_reg ,
  \piso.data_r_3968_sv2v_reg ,\piso.data_r_3967_sv2v_reg ,\piso.data_r_3966_sv2v_reg ,
  \piso.data_r_3965_sv2v_reg ,\piso.data_r_3964_sv2v_reg ,\piso.data_r_3963_sv2v_reg ,
  \piso.data_r_3962_sv2v_reg ,\piso.data_r_3961_sv2v_reg ,\piso.data_r_3960_sv2v_reg ,
  \piso.data_r_3959_sv2v_reg ,\piso.data_r_3958_sv2v_reg ,\piso.data_r_3957_sv2v_reg ,
  \piso.data_r_3956_sv2v_reg ,\piso.data_r_3955_sv2v_reg ,\piso.data_r_3954_sv2v_reg ,
  \piso.data_r_3953_sv2v_reg ,\piso.data_r_3952_sv2v_reg ,\piso.data_r_3951_sv2v_reg ,
  \piso.data_r_3950_sv2v_reg ,\piso.data_r_3949_sv2v_reg ,
  \piso.data_r_3948_sv2v_reg ,\piso.data_r_3947_sv2v_reg ,\piso.data_r_3946_sv2v_reg ,
  \piso.data_r_3945_sv2v_reg ,\piso.data_r_3944_sv2v_reg ,\piso.data_r_3943_sv2v_reg ,
  \piso.data_r_3942_sv2v_reg ,\piso.data_r_3941_sv2v_reg ,\piso.data_r_3940_sv2v_reg ,
  \piso.data_r_3939_sv2v_reg ,\piso.data_r_3938_sv2v_reg ,\piso.data_r_3937_sv2v_reg ,
  \piso.data_r_3936_sv2v_reg ,\piso.data_r_3935_sv2v_reg ,\piso.data_r_3934_sv2v_reg ,
  \piso.data_r_3933_sv2v_reg ,\piso.data_r_3932_sv2v_reg ,\piso.data_r_3931_sv2v_reg ,
  \piso.data_r_3930_sv2v_reg ,\piso.data_r_3929_sv2v_reg ,
  \piso.data_r_3928_sv2v_reg ,\piso.data_r_3927_sv2v_reg ,\piso.data_r_3926_sv2v_reg ,
  \piso.data_r_3925_sv2v_reg ,\piso.data_r_3924_sv2v_reg ,\piso.data_r_3923_sv2v_reg ,
  \piso.data_r_3922_sv2v_reg ,\piso.data_r_3921_sv2v_reg ,\piso.data_r_3920_sv2v_reg ,
  \piso.data_r_3919_sv2v_reg ,\piso.data_r_3918_sv2v_reg ,\piso.data_r_3917_sv2v_reg ,
  \piso.data_r_3916_sv2v_reg ,\piso.data_r_3915_sv2v_reg ,\piso.data_r_3914_sv2v_reg ,
  \piso.data_r_3913_sv2v_reg ,\piso.data_r_3912_sv2v_reg ,\piso.data_r_3911_sv2v_reg ,
  \piso.data_r_3910_sv2v_reg ,\piso.data_r_3909_sv2v_reg ,
  \piso.data_r_3908_sv2v_reg ,\piso.data_r_3907_sv2v_reg ,\piso.data_r_3906_sv2v_reg ,
  \piso.data_r_3905_sv2v_reg ,\piso.data_r_3904_sv2v_reg ,\piso.data_r_3903_sv2v_reg ,
  \piso.data_r_3902_sv2v_reg ,\piso.data_r_3901_sv2v_reg ,\piso.data_r_3900_sv2v_reg ,
  \piso.data_r_3899_sv2v_reg ,\piso.data_r_3898_sv2v_reg ,\piso.data_r_3897_sv2v_reg ,
  \piso.data_r_3896_sv2v_reg ,\piso.data_r_3895_sv2v_reg ,\piso.data_r_3894_sv2v_reg ,
  \piso.data_r_3893_sv2v_reg ,\piso.data_r_3892_sv2v_reg ,\piso.data_r_3891_sv2v_reg ,
  \piso.data_r_3890_sv2v_reg ,\piso.data_r_3889_sv2v_reg ,
  \piso.data_r_3888_sv2v_reg ,\piso.data_r_3887_sv2v_reg ,\piso.data_r_3886_sv2v_reg ,
  \piso.data_r_3885_sv2v_reg ,\piso.data_r_3884_sv2v_reg ,\piso.data_r_3883_sv2v_reg ,
  \piso.data_r_3882_sv2v_reg ,\piso.data_r_3881_sv2v_reg ,\piso.data_r_3880_sv2v_reg ,
  \piso.data_r_3879_sv2v_reg ,\piso.data_r_3878_sv2v_reg ,\piso.data_r_3877_sv2v_reg ,
  \piso.data_r_3876_sv2v_reg ,\piso.data_r_3875_sv2v_reg ,\piso.data_r_3874_sv2v_reg ,
  \piso.data_r_3873_sv2v_reg ,\piso.data_r_3872_sv2v_reg ,\piso.data_r_3871_sv2v_reg ,
  \piso.data_r_3870_sv2v_reg ,\piso.data_r_3869_sv2v_reg ,
  \piso.data_r_3868_sv2v_reg ,\piso.data_r_3867_sv2v_reg ,\piso.data_r_3866_sv2v_reg ,
  \piso.data_r_3865_sv2v_reg ,\piso.data_r_3864_sv2v_reg ,\piso.data_r_3863_sv2v_reg ,
  \piso.data_r_3862_sv2v_reg ,\piso.data_r_3861_sv2v_reg ,\piso.data_r_3860_sv2v_reg ,
  \piso.data_r_3859_sv2v_reg ,\piso.data_r_3858_sv2v_reg ,\piso.data_r_3857_sv2v_reg ,
  \piso.data_r_3856_sv2v_reg ,\piso.data_r_3855_sv2v_reg ,\piso.data_r_3854_sv2v_reg ,
  \piso.data_r_3853_sv2v_reg ,\piso.data_r_3852_sv2v_reg ,\piso.data_r_3851_sv2v_reg ,
  \piso.data_r_3850_sv2v_reg ,\piso.data_r_3849_sv2v_reg ,
  \piso.data_r_3848_sv2v_reg ,\piso.data_r_3847_sv2v_reg ,\piso.data_r_3846_sv2v_reg ,
  \piso.data_r_3845_sv2v_reg ,\piso.data_r_3844_sv2v_reg ,\piso.data_r_3843_sv2v_reg ,
  \piso.data_r_3842_sv2v_reg ,\piso.data_r_3841_sv2v_reg ,\piso.data_r_3840_sv2v_reg ,
  \piso.data_r_3839_sv2v_reg ,\piso.data_r_3838_sv2v_reg ,\piso.data_r_3837_sv2v_reg ,
  \piso.data_r_3836_sv2v_reg ,\piso.data_r_3835_sv2v_reg ,\piso.data_r_3834_sv2v_reg ,
  \piso.data_r_3833_sv2v_reg ,\piso.data_r_3832_sv2v_reg ,\piso.data_r_3831_sv2v_reg ,
  \piso.data_r_3830_sv2v_reg ,\piso.data_r_3829_sv2v_reg ,
  \piso.data_r_3828_sv2v_reg ,\piso.data_r_3827_sv2v_reg ,\piso.data_r_3826_sv2v_reg ,
  \piso.data_r_3825_sv2v_reg ,\piso.data_r_3824_sv2v_reg ,\piso.data_r_3823_sv2v_reg ,
  \piso.data_r_3822_sv2v_reg ,\piso.data_r_3821_sv2v_reg ,\piso.data_r_3820_sv2v_reg ,
  \piso.data_r_3819_sv2v_reg ,\piso.data_r_3818_sv2v_reg ,\piso.data_r_3817_sv2v_reg ,
  \piso.data_r_3816_sv2v_reg ,\piso.data_r_3815_sv2v_reg ,\piso.data_r_3814_sv2v_reg ,
  \piso.data_r_3813_sv2v_reg ,\piso.data_r_3812_sv2v_reg ,\piso.data_r_3811_sv2v_reg ,
  \piso.data_r_3810_sv2v_reg ,\piso.data_r_3809_sv2v_reg ,
  \piso.data_r_3808_sv2v_reg ,\piso.data_r_3807_sv2v_reg ,\piso.data_r_3806_sv2v_reg ,
  \piso.data_r_3805_sv2v_reg ,\piso.data_r_3804_sv2v_reg ,\piso.data_r_3803_sv2v_reg ,
  \piso.data_r_3802_sv2v_reg ,\piso.data_r_3801_sv2v_reg ,\piso.data_r_3800_sv2v_reg ,
  \piso.data_r_3799_sv2v_reg ,\piso.data_r_3798_sv2v_reg ,\piso.data_r_3797_sv2v_reg ,
  \piso.data_r_3796_sv2v_reg ,\piso.data_r_3795_sv2v_reg ,\piso.data_r_3794_sv2v_reg ,
  \piso.data_r_3793_sv2v_reg ,\piso.data_r_3792_sv2v_reg ,\piso.data_r_3791_sv2v_reg ,
  \piso.data_r_3790_sv2v_reg ,\piso.data_r_3789_sv2v_reg ,
  \piso.data_r_3788_sv2v_reg ,\piso.data_r_3787_sv2v_reg ,\piso.data_r_3786_sv2v_reg ,
  \piso.data_r_3785_sv2v_reg ,\piso.data_r_3784_sv2v_reg ,\piso.data_r_3783_sv2v_reg ,
  \piso.data_r_3782_sv2v_reg ,\piso.data_r_3781_sv2v_reg ,\piso.data_r_3780_sv2v_reg ,
  \piso.data_r_3779_sv2v_reg ,\piso.data_r_3778_sv2v_reg ,\piso.data_r_3777_sv2v_reg ,
  \piso.data_r_3776_sv2v_reg ,\piso.data_r_3775_sv2v_reg ,\piso.data_r_3774_sv2v_reg ,
  \piso.data_r_3773_sv2v_reg ,\piso.data_r_3772_sv2v_reg ,\piso.data_r_3771_sv2v_reg ,
  \piso.data_r_3770_sv2v_reg ,\piso.data_r_3769_sv2v_reg ,
  \piso.data_r_3768_sv2v_reg ,\piso.data_r_3767_sv2v_reg ,\piso.data_r_3766_sv2v_reg ,
  \piso.data_r_3765_sv2v_reg ,\piso.data_r_3764_sv2v_reg ,\piso.data_r_3763_sv2v_reg ,
  \piso.data_r_3762_sv2v_reg ,\piso.data_r_3761_sv2v_reg ,\piso.data_r_3760_sv2v_reg ,
  \piso.data_r_3759_sv2v_reg ,\piso.data_r_3758_sv2v_reg ,\piso.data_r_3757_sv2v_reg ,
  \piso.data_r_3756_sv2v_reg ,\piso.data_r_3755_sv2v_reg ,\piso.data_r_3754_sv2v_reg ,
  \piso.data_r_3753_sv2v_reg ,\piso.data_r_3752_sv2v_reg ,\piso.data_r_3751_sv2v_reg ,
  \piso.data_r_3750_sv2v_reg ,\piso.data_r_3749_sv2v_reg ,
  \piso.data_r_3748_sv2v_reg ,\piso.data_r_3747_sv2v_reg ,\piso.data_r_3746_sv2v_reg ,
  \piso.data_r_3745_sv2v_reg ,\piso.data_r_3744_sv2v_reg ,\piso.data_r_3743_sv2v_reg ,
  \piso.data_r_3742_sv2v_reg ,\piso.data_r_3741_sv2v_reg ,\piso.data_r_3740_sv2v_reg ,
  \piso.data_r_3739_sv2v_reg ,\piso.data_r_3738_sv2v_reg ,\piso.data_r_3737_sv2v_reg ,
  \piso.data_r_3736_sv2v_reg ,\piso.data_r_3735_sv2v_reg ,\piso.data_r_3734_sv2v_reg ,
  \piso.data_r_3733_sv2v_reg ,\piso.data_r_3732_sv2v_reg ,\piso.data_r_3731_sv2v_reg ,
  \piso.data_r_3730_sv2v_reg ,\piso.data_r_3729_sv2v_reg ,
  \piso.data_r_3728_sv2v_reg ,\piso.data_r_3727_sv2v_reg ,\piso.data_r_3726_sv2v_reg ,
  \piso.data_r_3725_sv2v_reg ,\piso.data_r_3724_sv2v_reg ,\piso.data_r_3723_sv2v_reg ,
  \piso.data_r_3722_sv2v_reg ,\piso.data_r_3721_sv2v_reg ,\piso.data_r_3720_sv2v_reg ,
  \piso.data_r_3719_sv2v_reg ,\piso.data_r_3718_sv2v_reg ,\piso.data_r_3717_sv2v_reg ,
  \piso.data_r_3716_sv2v_reg ,\piso.data_r_3715_sv2v_reg ,\piso.data_r_3714_sv2v_reg ,
  \piso.data_r_3713_sv2v_reg ,\piso.data_r_3712_sv2v_reg ,\piso.data_r_3711_sv2v_reg ,
  \piso.data_r_3710_sv2v_reg ,\piso.data_r_3709_sv2v_reg ,
  \piso.data_r_3708_sv2v_reg ,\piso.data_r_3707_sv2v_reg ,\piso.data_r_3706_sv2v_reg ,
  \piso.data_r_3705_sv2v_reg ,\piso.data_r_3704_sv2v_reg ,\piso.data_r_3703_sv2v_reg ,
  \piso.data_r_3702_sv2v_reg ,\piso.data_r_3701_sv2v_reg ,\piso.data_r_3700_sv2v_reg ,
  \piso.data_r_3699_sv2v_reg ,\piso.data_r_3698_sv2v_reg ,\piso.data_r_3697_sv2v_reg ,
  \piso.data_r_3696_sv2v_reg ,\piso.data_r_3695_sv2v_reg ,\piso.data_r_3694_sv2v_reg ,
  \piso.data_r_3693_sv2v_reg ,\piso.data_r_3692_sv2v_reg ,\piso.data_r_3691_sv2v_reg ,
  \piso.data_r_3690_sv2v_reg ,\piso.data_r_3689_sv2v_reg ,
  \piso.data_r_3688_sv2v_reg ,\piso.data_r_3687_sv2v_reg ,\piso.data_r_3686_sv2v_reg ,
  \piso.data_r_3685_sv2v_reg ,\piso.data_r_3684_sv2v_reg ,\piso.data_r_3683_sv2v_reg ,
  \piso.data_r_3682_sv2v_reg ,\piso.data_r_3681_sv2v_reg ,\piso.data_r_3680_sv2v_reg ,
  \piso.data_r_3679_sv2v_reg ,\piso.data_r_3678_sv2v_reg ,\piso.data_r_3677_sv2v_reg ,
  \piso.data_r_3676_sv2v_reg ,\piso.data_r_3675_sv2v_reg ,\piso.data_r_3674_sv2v_reg ,
  \piso.data_r_3673_sv2v_reg ,\piso.data_r_3672_sv2v_reg ,\piso.data_r_3671_sv2v_reg ,
  \piso.data_r_3670_sv2v_reg ,\piso.data_r_3669_sv2v_reg ,
  \piso.data_r_3668_sv2v_reg ,\piso.data_r_3667_sv2v_reg ,\piso.data_r_3666_sv2v_reg ,
  \piso.data_r_3665_sv2v_reg ,\piso.data_r_3664_sv2v_reg ,\piso.data_r_3663_sv2v_reg ,
  \piso.data_r_3662_sv2v_reg ,\piso.data_r_3661_sv2v_reg ,\piso.data_r_3660_sv2v_reg ,
  \piso.data_r_3659_sv2v_reg ,\piso.data_r_3658_sv2v_reg ,\piso.data_r_3657_sv2v_reg ,
  \piso.data_r_3656_sv2v_reg ,\piso.data_r_3655_sv2v_reg ,\piso.data_r_3654_sv2v_reg ,
  \piso.data_r_3653_sv2v_reg ,\piso.data_r_3652_sv2v_reg ,\piso.data_r_3651_sv2v_reg ,
  \piso.data_r_3650_sv2v_reg ,\piso.data_r_3649_sv2v_reg ,
  \piso.data_r_3648_sv2v_reg ,\piso.data_r_3647_sv2v_reg ,\piso.data_r_3646_sv2v_reg ,
  \piso.data_r_3645_sv2v_reg ,\piso.data_r_3644_sv2v_reg ,\piso.data_r_3643_sv2v_reg ,
  \piso.data_r_3642_sv2v_reg ,\piso.data_r_3641_sv2v_reg ,\piso.data_r_3640_sv2v_reg ,
  \piso.data_r_3639_sv2v_reg ,\piso.data_r_3638_sv2v_reg ,\piso.data_r_3637_sv2v_reg ,
  \piso.data_r_3636_sv2v_reg ,\piso.data_r_3635_sv2v_reg ,\piso.data_r_3634_sv2v_reg ,
  \piso.data_r_3633_sv2v_reg ,\piso.data_r_3632_sv2v_reg ,\piso.data_r_3631_sv2v_reg ,
  \piso.data_r_3630_sv2v_reg ,\piso.data_r_3629_sv2v_reg ,
  \piso.data_r_3628_sv2v_reg ,\piso.data_r_3627_sv2v_reg ,\piso.data_r_3626_sv2v_reg ,
  \piso.data_r_3625_sv2v_reg ,\piso.data_r_3624_sv2v_reg ,\piso.data_r_3623_sv2v_reg ,
  \piso.data_r_3622_sv2v_reg ,\piso.data_r_3621_sv2v_reg ,\piso.data_r_3620_sv2v_reg ,
  \piso.data_r_3619_sv2v_reg ,\piso.data_r_3618_sv2v_reg ,\piso.data_r_3617_sv2v_reg ,
  \piso.data_r_3616_sv2v_reg ,\piso.data_r_3615_sv2v_reg ,\piso.data_r_3614_sv2v_reg ,
  \piso.data_r_3613_sv2v_reg ,\piso.data_r_3612_sv2v_reg ,\piso.data_r_3611_sv2v_reg ,
  \piso.data_r_3610_sv2v_reg ,\piso.data_r_3609_sv2v_reg ,
  \piso.data_r_3608_sv2v_reg ,\piso.data_r_3607_sv2v_reg ,\piso.data_r_3606_sv2v_reg ,
  \piso.data_r_3605_sv2v_reg ,\piso.data_r_3604_sv2v_reg ,\piso.data_r_3603_sv2v_reg ,
  \piso.data_r_3602_sv2v_reg ,\piso.data_r_3601_sv2v_reg ,\piso.data_r_3600_sv2v_reg ,
  \piso.data_r_3599_sv2v_reg ,\piso.data_r_3598_sv2v_reg ,\piso.data_r_3597_sv2v_reg ,
  \piso.data_r_3596_sv2v_reg ,\piso.data_r_3595_sv2v_reg ,\piso.data_r_3594_sv2v_reg ,
  \piso.data_r_3593_sv2v_reg ,\piso.data_r_3592_sv2v_reg ,\piso.data_r_3591_sv2v_reg ,
  \piso.data_r_3590_sv2v_reg ,\piso.data_r_3589_sv2v_reg ,
  \piso.data_r_3588_sv2v_reg ,\piso.data_r_3587_sv2v_reg ,\piso.data_r_3586_sv2v_reg ,
  \piso.data_r_3585_sv2v_reg ,\piso.data_r_3584_sv2v_reg ,\piso.data_r_3583_sv2v_reg ,
  \piso.data_r_3582_sv2v_reg ,\piso.data_r_3581_sv2v_reg ,\piso.data_r_3580_sv2v_reg ,
  \piso.data_r_3579_sv2v_reg ,\piso.data_r_3578_sv2v_reg ,\piso.data_r_3577_sv2v_reg ,
  \piso.data_r_3576_sv2v_reg ,\piso.data_r_3575_sv2v_reg ,\piso.data_r_3574_sv2v_reg ,
  \piso.data_r_3573_sv2v_reg ,\piso.data_r_3572_sv2v_reg ,\piso.data_r_3571_sv2v_reg ,
  \piso.data_r_3570_sv2v_reg ,\piso.data_r_3569_sv2v_reg ,
  \piso.data_r_3568_sv2v_reg ,\piso.data_r_3567_sv2v_reg ,\piso.data_r_3566_sv2v_reg ,
  \piso.data_r_3565_sv2v_reg ,\piso.data_r_3564_sv2v_reg ,\piso.data_r_3563_sv2v_reg ,
  \piso.data_r_3562_sv2v_reg ,\piso.data_r_3561_sv2v_reg ,\piso.data_r_3560_sv2v_reg ,
  \piso.data_r_3559_sv2v_reg ,\piso.data_r_3558_sv2v_reg ,\piso.data_r_3557_sv2v_reg ,
  \piso.data_r_3556_sv2v_reg ,\piso.data_r_3555_sv2v_reg ,\piso.data_r_3554_sv2v_reg ,
  \piso.data_r_3553_sv2v_reg ,\piso.data_r_3552_sv2v_reg ,\piso.data_r_3551_sv2v_reg ,
  \piso.data_r_3550_sv2v_reg ,\piso.data_r_3549_sv2v_reg ,
  \piso.data_r_3548_sv2v_reg ,\piso.data_r_3547_sv2v_reg ,\piso.data_r_3546_sv2v_reg ,
  \piso.data_r_3545_sv2v_reg ,\piso.data_r_3544_sv2v_reg ,\piso.data_r_3543_sv2v_reg ,
  \piso.data_r_3542_sv2v_reg ,\piso.data_r_3541_sv2v_reg ,\piso.data_r_3540_sv2v_reg ,
  \piso.data_r_3539_sv2v_reg ,\piso.data_r_3538_sv2v_reg ,\piso.data_r_3537_sv2v_reg ,
  \piso.data_r_3536_sv2v_reg ,\piso.data_r_3535_sv2v_reg ,\piso.data_r_3534_sv2v_reg ,
  \piso.data_r_3533_sv2v_reg ,\piso.data_r_3532_sv2v_reg ,\piso.data_r_3531_sv2v_reg ,
  \piso.data_r_3530_sv2v_reg ,\piso.data_r_3529_sv2v_reg ,
  \piso.data_r_3528_sv2v_reg ,\piso.data_r_3527_sv2v_reg ,\piso.data_r_3526_sv2v_reg ,
  \piso.data_r_3525_sv2v_reg ,\piso.data_r_3524_sv2v_reg ,\piso.data_r_3523_sv2v_reg ,
  \piso.data_r_3522_sv2v_reg ,\piso.data_r_3521_sv2v_reg ,\piso.data_r_3520_sv2v_reg ,
  \piso.data_r_3519_sv2v_reg ,\piso.data_r_3518_sv2v_reg ,\piso.data_r_3517_sv2v_reg ,
  \piso.data_r_3516_sv2v_reg ,\piso.data_r_3515_sv2v_reg ,\piso.data_r_3514_sv2v_reg ,
  \piso.data_r_3513_sv2v_reg ,\piso.data_r_3512_sv2v_reg ,\piso.data_r_3511_sv2v_reg ,
  \piso.data_r_3510_sv2v_reg ,\piso.data_r_3509_sv2v_reg ,
  \piso.data_r_3508_sv2v_reg ,\piso.data_r_3507_sv2v_reg ,\piso.data_r_3506_sv2v_reg ,
  \piso.data_r_3505_sv2v_reg ,\piso.data_r_3504_sv2v_reg ,\piso.data_r_3503_sv2v_reg ,
  \piso.data_r_3502_sv2v_reg ,\piso.data_r_3501_sv2v_reg ,\piso.data_r_3500_sv2v_reg ,
  \piso.data_r_3499_sv2v_reg ,\piso.data_r_3498_sv2v_reg ,\piso.data_r_3497_sv2v_reg ,
  \piso.data_r_3496_sv2v_reg ,\piso.data_r_3495_sv2v_reg ,\piso.data_r_3494_sv2v_reg ,
  \piso.data_r_3493_sv2v_reg ,\piso.data_r_3492_sv2v_reg ,\piso.data_r_3491_sv2v_reg ,
  \piso.data_r_3490_sv2v_reg ,\piso.data_r_3489_sv2v_reg ,
  \piso.data_r_3488_sv2v_reg ,\piso.data_r_3487_sv2v_reg ,\piso.data_r_3486_sv2v_reg ,
  \piso.data_r_3485_sv2v_reg ,\piso.data_r_3484_sv2v_reg ,\piso.data_r_3483_sv2v_reg ,
  \piso.data_r_3482_sv2v_reg ,\piso.data_r_3481_sv2v_reg ,\piso.data_r_3480_sv2v_reg ,
  \piso.data_r_3479_sv2v_reg ,\piso.data_r_3478_sv2v_reg ,\piso.data_r_3477_sv2v_reg ,
  \piso.data_r_3476_sv2v_reg ,\piso.data_r_3475_sv2v_reg ,\piso.data_r_3474_sv2v_reg ,
  \piso.data_r_3473_sv2v_reg ,\piso.data_r_3472_sv2v_reg ,\piso.data_r_3471_sv2v_reg ,
  \piso.data_r_3470_sv2v_reg ,\piso.data_r_3469_sv2v_reg ,
  \piso.data_r_3468_sv2v_reg ,\piso.data_r_3467_sv2v_reg ,\piso.data_r_3466_sv2v_reg ,
  \piso.data_r_3465_sv2v_reg ,\piso.data_r_3464_sv2v_reg ,\piso.data_r_3463_sv2v_reg ,
  \piso.data_r_3462_sv2v_reg ,\piso.data_r_3461_sv2v_reg ,\piso.data_r_3460_sv2v_reg ,
  \piso.data_r_3459_sv2v_reg ,\piso.data_r_3458_sv2v_reg ,\piso.data_r_3457_sv2v_reg ,
  \piso.data_r_3456_sv2v_reg ,\piso.data_r_3455_sv2v_reg ,\piso.data_r_3454_sv2v_reg ,
  \piso.data_r_3453_sv2v_reg ,\piso.data_r_3452_sv2v_reg ,\piso.data_r_3451_sv2v_reg ,
  \piso.data_r_3450_sv2v_reg ,\piso.data_r_3449_sv2v_reg ,
  \piso.data_r_3448_sv2v_reg ,\piso.data_r_3447_sv2v_reg ,\piso.data_r_3446_sv2v_reg ,
  \piso.data_r_3445_sv2v_reg ,\piso.data_r_3444_sv2v_reg ,\piso.data_r_3443_sv2v_reg ,
  \piso.data_r_3442_sv2v_reg ,\piso.data_r_3441_sv2v_reg ,\piso.data_r_3440_sv2v_reg ,
  \piso.data_r_3439_sv2v_reg ,\piso.data_r_3438_sv2v_reg ,\piso.data_r_3437_sv2v_reg ,
  \piso.data_r_3436_sv2v_reg ,\piso.data_r_3435_sv2v_reg ,\piso.data_r_3434_sv2v_reg ,
  \piso.data_r_3433_sv2v_reg ,\piso.data_r_3432_sv2v_reg ,\piso.data_r_3431_sv2v_reg ,
  \piso.data_r_3430_sv2v_reg ,\piso.data_r_3429_sv2v_reg ,
  \piso.data_r_3428_sv2v_reg ,\piso.data_r_3427_sv2v_reg ,\piso.data_r_3426_sv2v_reg ,
  \piso.data_r_3425_sv2v_reg ,\piso.data_r_3424_sv2v_reg ,\piso.data_r_3423_sv2v_reg ,
  \piso.data_r_3422_sv2v_reg ,\piso.data_r_3421_sv2v_reg ,\piso.data_r_3420_sv2v_reg ,
  \piso.data_r_3419_sv2v_reg ,\piso.data_r_3418_sv2v_reg ,\piso.data_r_3417_sv2v_reg ,
  \piso.data_r_3416_sv2v_reg ,\piso.data_r_3415_sv2v_reg ,\piso.data_r_3414_sv2v_reg ,
  \piso.data_r_3413_sv2v_reg ,\piso.data_r_3412_sv2v_reg ,\piso.data_r_3411_sv2v_reg ,
  \piso.data_r_3410_sv2v_reg ,\piso.data_r_3409_sv2v_reg ,
  \piso.data_r_3408_sv2v_reg ,\piso.data_r_3407_sv2v_reg ,\piso.data_r_3406_sv2v_reg ,
  \piso.data_r_3405_sv2v_reg ,\piso.data_r_3404_sv2v_reg ,\piso.data_r_3403_sv2v_reg ,
  \piso.data_r_3402_sv2v_reg ,\piso.data_r_3401_sv2v_reg ,\piso.data_r_3400_sv2v_reg ,
  \piso.data_r_3399_sv2v_reg ,\piso.data_r_3398_sv2v_reg ,\piso.data_r_3397_sv2v_reg ,
  \piso.data_r_3396_sv2v_reg ,\piso.data_r_3395_sv2v_reg ,\piso.data_r_3394_sv2v_reg ,
  \piso.data_r_3393_sv2v_reg ,\piso.data_r_3392_sv2v_reg ,\piso.data_r_3391_sv2v_reg ,
  \piso.data_r_3390_sv2v_reg ,\piso.data_r_3389_sv2v_reg ,
  \piso.data_r_3388_sv2v_reg ,\piso.data_r_3387_sv2v_reg ,\piso.data_r_3386_sv2v_reg ,
  \piso.data_r_3385_sv2v_reg ,\piso.data_r_3384_sv2v_reg ,\piso.data_r_3383_sv2v_reg ,
  \piso.data_r_3382_sv2v_reg ,\piso.data_r_3381_sv2v_reg ,\piso.data_r_3380_sv2v_reg ,
  \piso.data_r_3379_sv2v_reg ,\piso.data_r_3378_sv2v_reg ,\piso.data_r_3377_sv2v_reg ,
  \piso.data_r_3376_sv2v_reg ,\piso.data_r_3375_sv2v_reg ,\piso.data_r_3374_sv2v_reg ,
  \piso.data_r_3373_sv2v_reg ,\piso.data_r_3372_sv2v_reg ,\piso.data_r_3371_sv2v_reg ,
  \piso.data_r_3370_sv2v_reg ,\piso.data_r_3369_sv2v_reg ,
  \piso.data_r_3368_sv2v_reg ,\piso.data_r_3367_sv2v_reg ,\piso.data_r_3366_sv2v_reg ,
  \piso.data_r_3365_sv2v_reg ,\piso.data_r_3364_sv2v_reg ,\piso.data_r_3363_sv2v_reg ,
  \piso.data_r_3362_sv2v_reg ,\piso.data_r_3361_sv2v_reg ,\piso.data_r_3360_sv2v_reg ,
  \piso.data_r_3359_sv2v_reg ,\piso.data_r_3358_sv2v_reg ,\piso.data_r_3357_sv2v_reg ,
  \piso.data_r_3356_sv2v_reg ,\piso.data_r_3355_sv2v_reg ,\piso.data_r_3354_sv2v_reg ,
  \piso.data_r_3353_sv2v_reg ,\piso.data_r_3352_sv2v_reg ,\piso.data_r_3351_sv2v_reg ,
  \piso.data_r_3350_sv2v_reg ,\piso.data_r_3349_sv2v_reg ,
  \piso.data_r_3348_sv2v_reg ,\piso.data_r_3347_sv2v_reg ,\piso.data_r_3346_sv2v_reg ,
  \piso.data_r_3345_sv2v_reg ,\piso.data_r_3344_sv2v_reg ,\piso.data_r_3343_sv2v_reg ,
  \piso.data_r_3342_sv2v_reg ,\piso.data_r_3341_sv2v_reg ,\piso.data_r_3340_sv2v_reg ,
  \piso.data_r_3339_sv2v_reg ,\piso.data_r_3338_sv2v_reg ,\piso.data_r_3337_sv2v_reg ,
  \piso.data_r_3336_sv2v_reg ,\piso.data_r_3335_sv2v_reg ,\piso.data_r_3334_sv2v_reg ,
  \piso.data_r_3333_sv2v_reg ,\piso.data_r_3332_sv2v_reg ,\piso.data_r_3331_sv2v_reg ,
  \piso.data_r_3330_sv2v_reg ,\piso.data_r_3329_sv2v_reg ,
  \piso.data_r_3328_sv2v_reg ,\piso.data_r_3327_sv2v_reg ,\piso.data_r_3326_sv2v_reg ,
  \piso.data_r_3325_sv2v_reg ,\piso.data_r_3324_sv2v_reg ,\piso.data_r_3323_sv2v_reg ,
  \piso.data_r_3322_sv2v_reg ,\piso.data_r_3321_sv2v_reg ,\piso.data_r_3320_sv2v_reg ,
  \piso.data_r_3319_sv2v_reg ,\piso.data_r_3318_sv2v_reg ,\piso.data_r_3317_sv2v_reg ,
  \piso.data_r_3316_sv2v_reg ,\piso.data_r_3315_sv2v_reg ,\piso.data_r_3314_sv2v_reg ,
  \piso.data_r_3313_sv2v_reg ,\piso.data_r_3312_sv2v_reg ,\piso.data_r_3311_sv2v_reg ,
  \piso.data_r_3310_sv2v_reg ,\piso.data_r_3309_sv2v_reg ,
  \piso.data_r_3308_sv2v_reg ,\piso.data_r_3307_sv2v_reg ,\piso.data_r_3306_sv2v_reg ,
  \piso.data_r_3305_sv2v_reg ,\piso.data_r_3304_sv2v_reg ,\piso.data_r_3303_sv2v_reg ,
  \piso.data_r_3302_sv2v_reg ,\piso.data_r_3301_sv2v_reg ,\piso.data_r_3300_sv2v_reg ,
  \piso.data_r_3299_sv2v_reg ,\piso.data_r_3298_sv2v_reg ,\piso.data_r_3297_sv2v_reg ,
  \piso.data_r_3296_sv2v_reg ,\piso.data_r_3295_sv2v_reg ,\piso.data_r_3294_sv2v_reg ,
  \piso.data_r_3293_sv2v_reg ,\piso.data_r_3292_sv2v_reg ,\piso.data_r_3291_sv2v_reg ,
  \piso.data_r_3290_sv2v_reg ,\piso.data_r_3289_sv2v_reg ,
  \piso.data_r_3288_sv2v_reg ,\piso.data_r_3287_sv2v_reg ,\piso.data_r_3286_sv2v_reg ,
  \piso.data_r_3285_sv2v_reg ,\piso.data_r_3284_sv2v_reg ,\piso.data_r_3283_sv2v_reg ,
  \piso.data_r_3282_sv2v_reg ,\piso.data_r_3281_sv2v_reg ,\piso.data_r_3280_sv2v_reg ,
  \piso.data_r_3279_sv2v_reg ,\piso.data_r_3278_sv2v_reg ,\piso.data_r_3277_sv2v_reg ,
  \piso.data_r_3276_sv2v_reg ,\piso.data_r_3275_sv2v_reg ,\piso.data_r_3274_sv2v_reg ,
  \piso.data_r_3273_sv2v_reg ,\piso.data_r_3272_sv2v_reg ,\piso.data_r_3271_sv2v_reg ,
  \piso.data_r_3270_sv2v_reg ,\piso.data_r_3269_sv2v_reg ,
  \piso.data_r_3268_sv2v_reg ,\piso.data_r_3267_sv2v_reg ,\piso.data_r_3266_sv2v_reg ,
  \piso.data_r_3265_sv2v_reg ,\piso.data_r_3264_sv2v_reg ,\piso.data_r_3263_sv2v_reg ,
  \piso.data_r_3262_sv2v_reg ,\piso.data_r_3261_sv2v_reg ,\piso.data_r_3260_sv2v_reg ,
  \piso.data_r_3259_sv2v_reg ,\piso.data_r_3258_sv2v_reg ,\piso.data_r_3257_sv2v_reg ,
  \piso.data_r_3256_sv2v_reg ,\piso.data_r_3255_sv2v_reg ,\piso.data_r_3254_sv2v_reg ,
  \piso.data_r_3253_sv2v_reg ,\piso.data_r_3252_sv2v_reg ,\piso.data_r_3251_sv2v_reg ,
  \piso.data_r_3250_sv2v_reg ,\piso.data_r_3249_sv2v_reg ,
  \piso.data_r_3248_sv2v_reg ,\piso.data_r_3247_sv2v_reg ,\piso.data_r_3246_sv2v_reg ,
  \piso.data_r_3245_sv2v_reg ,\piso.data_r_3244_sv2v_reg ,\piso.data_r_3243_sv2v_reg ,
  \piso.data_r_3242_sv2v_reg ,\piso.data_r_3241_sv2v_reg ,\piso.data_r_3240_sv2v_reg ,
  \piso.data_r_3239_sv2v_reg ,\piso.data_r_3238_sv2v_reg ,\piso.data_r_3237_sv2v_reg ,
  \piso.data_r_3236_sv2v_reg ,\piso.data_r_3235_sv2v_reg ,\piso.data_r_3234_sv2v_reg ,
  \piso.data_r_3233_sv2v_reg ,\piso.data_r_3232_sv2v_reg ,\piso.data_r_3231_sv2v_reg ,
  \piso.data_r_3230_sv2v_reg ,\piso.data_r_3229_sv2v_reg ,
  \piso.data_r_3228_sv2v_reg ,\piso.data_r_3227_sv2v_reg ,\piso.data_r_3226_sv2v_reg ,
  \piso.data_r_3225_sv2v_reg ,\piso.data_r_3224_sv2v_reg ,\piso.data_r_3223_sv2v_reg ,
  \piso.data_r_3222_sv2v_reg ,\piso.data_r_3221_sv2v_reg ,\piso.data_r_3220_sv2v_reg ,
  \piso.data_r_3219_sv2v_reg ,\piso.data_r_3218_sv2v_reg ,\piso.data_r_3217_sv2v_reg ,
  \piso.data_r_3216_sv2v_reg ,\piso.data_r_3215_sv2v_reg ,\piso.data_r_3214_sv2v_reg ,
  \piso.data_r_3213_sv2v_reg ,\piso.data_r_3212_sv2v_reg ,\piso.data_r_3211_sv2v_reg ,
  \piso.data_r_3210_sv2v_reg ,\piso.data_r_3209_sv2v_reg ,
  \piso.data_r_3208_sv2v_reg ,\piso.data_r_3207_sv2v_reg ,\piso.data_r_3206_sv2v_reg ,
  \piso.data_r_3205_sv2v_reg ,\piso.data_r_3204_sv2v_reg ,\piso.data_r_3203_sv2v_reg ,
  \piso.data_r_3202_sv2v_reg ,\piso.data_r_3201_sv2v_reg ,\piso.data_r_3200_sv2v_reg ,
  \piso.data_r_3199_sv2v_reg ,\piso.data_r_3198_sv2v_reg ,\piso.data_r_3197_sv2v_reg ,
  \piso.data_r_3196_sv2v_reg ,\piso.data_r_3195_sv2v_reg ,\piso.data_r_3194_sv2v_reg ,
  \piso.data_r_3193_sv2v_reg ,\piso.data_r_3192_sv2v_reg ,\piso.data_r_3191_sv2v_reg ,
  \piso.data_r_3190_sv2v_reg ,\piso.data_r_3189_sv2v_reg ,
  \piso.data_r_3188_sv2v_reg ,\piso.data_r_3187_sv2v_reg ,\piso.data_r_3186_sv2v_reg ,
  \piso.data_r_3185_sv2v_reg ,\piso.data_r_3184_sv2v_reg ,\piso.data_r_3183_sv2v_reg ,
  \piso.data_r_3182_sv2v_reg ,\piso.data_r_3181_sv2v_reg ,\piso.data_r_3180_sv2v_reg ,
  \piso.data_r_3179_sv2v_reg ,\piso.data_r_3178_sv2v_reg ,\piso.data_r_3177_sv2v_reg ,
  \piso.data_r_3176_sv2v_reg ,\piso.data_r_3175_sv2v_reg ,\piso.data_r_3174_sv2v_reg ,
  \piso.data_r_3173_sv2v_reg ,\piso.data_r_3172_sv2v_reg ,\piso.data_r_3171_sv2v_reg ,
  \piso.data_r_3170_sv2v_reg ,\piso.data_r_3169_sv2v_reg ,
  \piso.data_r_3168_sv2v_reg ,\piso.data_r_3167_sv2v_reg ,\piso.data_r_3166_sv2v_reg ,
  \piso.data_r_3165_sv2v_reg ,\piso.data_r_3164_sv2v_reg ,\piso.data_r_3163_sv2v_reg ,
  \piso.data_r_3162_sv2v_reg ,\piso.data_r_3161_sv2v_reg ,\piso.data_r_3160_sv2v_reg ,
  \piso.data_r_3159_sv2v_reg ,\piso.data_r_3158_sv2v_reg ,\piso.data_r_3157_sv2v_reg ,
  \piso.data_r_3156_sv2v_reg ,\piso.data_r_3155_sv2v_reg ,\piso.data_r_3154_sv2v_reg ,
  \piso.data_r_3153_sv2v_reg ,\piso.data_r_3152_sv2v_reg ,\piso.data_r_3151_sv2v_reg ,
  \piso.data_r_3150_sv2v_reg ,\piso.data_r_3149_sv2v_reg ,
  \piso.data_r_3148_sv2v_reg ,\piso.data_r_3147_sv2v_reg ,\piso.data_r_3146_sv2v_reg ,
  \piso.data_r_3145_sv2v_reg ,\piso.data_r_3144_sv2v_reg ,\piso.data_r_3143_sv2v_reg ,
  \piso.data_r_3142_sv2v_reg ,\piso.data_r_3141_sv2v_reg ,\piso.data_r_3140_sv2v_reg ,
  \piso.data_r_3139_sv2v_reg ,\piso.data_r_3138_sv2v_reg ,\piso.data_r_3137_sv2v_reg ,
  \piso.data_r_3136_sv2v_reg ,\piso.data_r_3135_sv2v_reg ,\piso.data_r_3134_sv2v_reg ,
  \piso.data_r_3133_sv2v_reg ,\piso.data_r_3132_sv2v_reg ,\piso.data_r_3131_sv2v_reg ,
  \piso.data_r_3130_sv2v_reg ,\piso.data_r_3129_sv2v_reg ,
  \piso.data_r_3128_sv2v_reg ,\piso.data_r_3127_sv2v_reg ,\piso.data_r_3126_sv2v_reg ,
  \piso.data_r_3125_sv2v_reg ,\piso.data_r_3124_sv2v_reg ,\piso.data_r_3123_sv2v_reg ,
  \piso.data_r_3122_sv2v_reg ,\piso.data_r_3121_sv2v_reg ,\piso.data_r_3120_sv2v_reg ,
  \piso.data_r_3119_sv2v_reg ,\piso.data_r_3118_sv2v_reg ,\piso.data_r_3117_sv2v_reg ,
  \piso.data_r_3116_sv2v_reg ,\piso.data_r_3115_sv2v_reg ,\piso.data_r_3114_sv2v_reg ,
  \piso.data_r_3113_sv2v_reg ,\piso.data_r_3112_sv2v_reg ,\piso.data_r_3111_sv2v_reg ,
  \piso.data_r_3110_sv2v_reg ,\piso.data_r_3109_sv2v_reg ,
  \piso.data_r_3108_sv2v_reg ,\piso.data_r_3107_sv2v_reg ,\piso.data_r_3106_sv2v_reg ,
  \piso.data_r_3105_sv2v_reg ,\piso.data_r_3104_sv2v_reg ,\piso.data_r_3103_sv2v_reg ,
  \piso.data_r_3102_sv2v_reg ,\piso.data_r_3101_sv2v_reg ,\piso.data_r_3100_sv2v_reg ,
  \piso.data_r_3099_sv2v_reg ,\piso.data_r_3098_sv2v_reg ,\piso.data_r_3097_sv2v_reg ,
  \piso.data_r_3096_sv2v_reg ,\piso.data_r_3095_sv2v_reg ,\piso.data_r_3094_sv2v_reg ,
  \piso.data_r_3093_sv2v_reg ,\piso.data_r_3092_sv2v_reg ,\piso.data_r_3091_sv2v_reg ,
  \piso.data_r_3090_sv2v_reg ,\piso.data_r_3089_sv2v_reg ,
  \piso.data_r_3088_sv2v_reg ,\piso.data_r_3087_sv2v_reg ,\piso.data_r_3086_sv2v_reg ,
  \piso.data_r_3085_sv2v_reg ,\piso.data_r_3084_sv2v_reg ,\piso.data_r_3083_sv2v_reg ,
  \piso.data_r_3082_sv2v_reg ,\piso.data_r_3081_sv2v_reg ,\piso.data_r_3080_sv2v_reg ,
  \piso.data_r_3079_sv2v_reg ,\piso.data_r_3078_sv2v_reg ,\piso.data_r_3077_sv2v_reg ,
  \piso.data_r_3076_sv2v_reg ,\piso.data_r_3075_sv2v_reg ,\piso.data_r_3074_sv2v_reg ,
  \piso.data_r_3073_sv2v_reg ,\piso.data_r_3072_sv2v_reg ,\piso.data_r_3071_sv2v_reg ,
  \piso.data_r_3070_sv2v_reg ,\piso.data_r_3069_sv2v_reg ,
  \piso.data_r_3068_sv2v_reg ,\piso.data_r_3067_sv2v_reg ,\piso.data_r_3066_sv2v_reg ,
  \piso.data_r_3065_sv2v_reg ,\piso.data_r_3064_sv2v_reg ,\piso.data_r_3063_sv2v_reg ,
  \piso.data_r_3062_sv2v_reg ,\piso.data_r_3061_sv2v_reg ,\piso.data_r_3060_sv2v_reg ,
  \piso.data_r_3059_sv2v_reg ,\piso.data_r_3058_sv2v_reg ,\piso.data_r_3057_sv2v_reg ,
  \piso.data_r_3056_sv2v_reg ,\piso.data_r_3055_sv2v_reg ,\piso.data_r_3054_sv2v_reg ,
  \piso.data_r_3053_sv2v_reg ,\piso.data_r_3052_sv2v_reg ,\piso.data_r_3051_sv2v_reg ,
  \piso.data_r_3050_sv2v_reg ,\piso.data_r_3049_sv2v_reg ,
  \piso.data_r_3048_sv2v_reg ,\piso.data_r_3047_sv2v_reg ,\piso.data_r_3046_sv2v_reg ,
  \piso.data_r_3045_sv2v_reg ,\piso.data_r_3044_sv2v_reg ,\piso.data_r_3043_sv2v_reg ,
  \piso.data_r_3042_sv2v_reg ,\piso.data_r_3041_sv2v_reg ,\piso.data_r_3040_sv2v_reg ,
  \piso.data_r_3039_sv2v_reg ,\piso.data_r_3038_sv2v_reg ,\piso.data_r_3037_sv2v_reg ,
  \piso.data_r_3036_sv2v_reg ,\piso.data_r_3035_sv2v_reg ,\piso.data_r_3034_sv2v_reg ,
  \piso.data_r_3033_sv2v_reg ,\piso.data_r_3032_sv2v_reg ,\piso.data_r_3031_sv2v_reg ,
  \piso.data_r_3030_sv2v_reg ,\piso.data_r_3029_sv2v_reg ,
  \piso.data_r_3028_sv2v_reg ,\piso.data_r_3027_sv2v_reg ,\piso.data_r_3026_sv2v_reg ,
  \piso.data_r_3025_sv2v_reg ,\piso.data_r_3024_sv2v_reg ,\piso.data_r_3023_sv2v_reg ,
  \piso.data_r_3022_sv2v_reg ,\piso.data_r_3021_sv2v_reg ,\piso.data_r_3020_sv2v_reg ,
  \piso.data_r_3019_sv2v_reg ,\piso.data_r_3018_sv2v_reg ,\piso.data_r_3017_sv2v_reg ,
  \piso.data_r_3016_sv2v_reg ,\piso.data_r_3015_sv2v_reg ,\piso.data_r_3014_sv2v_reg ,
  \piso.data_r_3013_sv2v_reg ,\piso.data_r_3012_sv2v_reg ,\piso.data_r_3011_sv2v_reg ,
  \piso.data_r_3010_sv2v_reg ,\piso.data_r_3009_sv2v_reg ,
  \piso.data_r_3008_sv2v_reg ,\piso.data_r_3007_sv2v_reg ,\piso.data_r_3006_sv2v_reg ,
  \piso.data_r_3005_sv2v_reg ,\piso.data_r_3004_sv2v_reg ,\piso.data_r_3003_sv2v_reg ,
  \piso.data_r_3002_sv2v_reg ,\piso.data_r_3001_sv2v_reg ,\piso.data_r_3000_sv2v_reg ,
  \piso.data_r_2999_sv2v_reg ,\piso.data_r_2998_sv2v_reg ,\piso.data_r_2997_sv2v_reg ,
  \piso.data_r_2996_sv2v_reg ,\piso.data_r_2995_sv2v_reg ,\piso.data_r_2994_sv2v_reg ,
  \piso.data_r_2993_sv2v_reg ,\piso.data_r_2992_sv2v_reg ,\piso.data_r_2991_sv2v_reg ,
  \piso.data_r_2990_sv2v_reg ,\piso.data_r_2989_sv2v_reg ,
  \piso.data_r_2988_sv2v_reg ,\piso.data_r_2987_sv2v_reg ,\piso.data_r_2986_sv2v_reg ,
  \piso.data_r_2985_sv2v_reg ,\piso.data_r_2984_sv2v_reg ,\piso.data_r_2983_sv2v_reg ,
  \piso.data_r_2982_sv2v_reg ,\piso.data_r_2981_sv2v_reg ,\piso.data_r_2980_sv2v_reg ,
  \piso.data_r_2979_sv2v_reg ,\piso.data_r_2978_sv2v_reg ,\piso.data_r_2977_sv2v_reg ,
  \piso.data_r_2976_sv2v_reg ,\piso.data_r_2975_sv2v_reg ,\piso.data_r_2974_sv2v_reg ,
  \piso.data_r_2973_sv2v_reg ,\piso.data_r_2972_sv2v_reg ,\piso.data_r_2971_sv2v_reg ,
  \piso.data_r_2970_sv2v_reg ,\piso.data_r_2969_sv2v_reg ,
  \piso.data_r_2968_sv2v_reg ,\piso.data_r_2967_sv2v_reg ,\piso.data_r_2966_sv2v_reg ,
  \piso.data_r_2965_sv2v_reg ,\piso.data_r_2964_sv2v_reg ,\piso.data_r_2963_sv2v_reg ,
  \piso.data_r_2962_sv2v_reg ,\piso.data_r_2961_sv2v_reg ,\piso.data_r_2960_sv2v_reg ,
  \piso.data_r_2959_sv2v_reg ,\piso.data_r_2958_sv2v_reg ,\piso.data_r_2957_sv2v_reg ,
  \piso.data_r_2956_sv2v_reg ,\piso.data_r_2955_sv2v_reg ,\piso.data_r_2954_sv2v_reg ,
  \piso.data_r_2953_sv2v_reg ,\piso.data_r_2952_sv2v_reg ,\piso.data_r_2951_sv2v_reg ,
  \piso.data_r_2950_sv2v_reg ,\piso.data_r_2949_sv2v_reg ,
  \piso.data_r_2948_sv2v_reg ,\piso.data_r_2947_sv2v_reg ,\piso.data_r_2946_sv2v_reg ,
  \piso.data_r_2945_sv2v_reg ,\piso.data_r_2944_sv2v_reg ,\piso.data_r_2943_sv2v_reg ,
  \piso.data_r_2942_sv2v_reg ,\piso.data_r_2941_sv2v_reg ,\piso.data_r_2940_sv2v_reg ,
  \piso.data_r_2939_sv2v_reg ,\piso.data_r_2938_sv2v_reg ,\piso.data_r_2937_sv2v_reg ,
  \piso.data_r_2936_sv2v_reg ,\piso.data_r_2935_sv2v_reg ,\piso.data_r_2934_sv2v_reg ,
  \piso.data_r_2933_sv2v_reg ,\piso.data_r_2932_sv2v_reg ,\piso.data_r_2931_sv2v_reg ,
  \piso.data_r_2930_sv2v_reg ,\piso.data_r_2929_sv2v_reg ,
  \piso.data_r_2928_sv2v_reg ,\piso.data_r_2927_sv2v_reg ,\piso.data_r_2926_sv2v_reg ,
  \piso.data_r_2925_sv2v_reg ,\piso.data_r_2924_sv2v_reg ,\piso.data_r_2923_sv2v_reg ,
  \piso.data_r_2922_sv2v_reg ,\piso.data_r_2921_sv2v_reg ,\piso.data_r_2920_sv2v_reg ,
  \piso.data_r_2919_sv2v_reg ,\piso.data_r_2918_sv2v_reg ,\piso.data_r_2917_sv2v_reg ,
  \piso.data_r_2916_sv2v_reg ,\piso.data_r_2915_sv2v_reg ,\piso.data_r_2914_sv2v_reg ,
  \piso.data_r_2913_sv2v_reg ,\piso.data_r_2912_sv2v_reg ,\piso.data_r_2911_sv2v_reg ,
  \piso.data_r_2910_sv2v_reg ,\piso.data_r_2909_sv2v_reg ,
  \piso.data_r_2908_sv2v_reg ,\piso.data_r_2907_sv2v_reg ,\piso.data_r_2906_sv2v_reg ,
  \piso.data_r_2905_sv2v_reg ,\piso.data_r_2904_sv2v_reg ,\piso.data_r_2903_sv2v_reg ,
  \piso.data_r_2902_sv2v_reg ,\piso.data_r_2901_sv2v_reg ,\piso.data_r_2900_sv2v_reg ,
  \piso.data_r_2899_sv2v_reg ,\piso.data_r_2898_sv2v_reg ,\piso.data_r_2897_sv2v_reg ,
  \piso.data_r_2896_sv2v_reg ,\piso.data_r_2895_sv2v_reg ,\piso.data_r_2894_sv2v_reg ,
  \piso.data_r_2893_sv2v_reg ,\piso.data_r_2892_sv2v_reg ,\piso.data_r_2891_sv2v_reg ,
  \piso.data_r_2890_sv2v_reg ,\piso.data_r_2889_sv2v_reg ,
  \piso.data_r_2888_sv2v_reg ,\piso.data_r_2887_sv2v_reg ,\piso.data_r_2886_sv2v_reg ,
  \piso.data_r_2885_sv2v_reg ,\piso.data_r_2884_sv2v_reg ,\piso.data_r_2883_sv2v_reg ,
  \piso.data_r_2882_sv2v_reg ,\piso.data_r_2881_sv2v_reg ,\piso.data_r_2880_sv2v_reg ,
  \piso.data_r_2879_sv2v_reg ,\piso.data_r_2878_sv2v_reg ,\piso.data_r_2877_sv2v_reg ,
  \piso.data_r_2876_sv2v_reg ,\piso.data_r_2875_sv2v_reg ,\piso.data_r_2874_sv2v_reg ,
  \piso.data_r_2873_sv2v_reg ,\piso.data_r_2872_sv2v_reg ,\piso.data_r_2871_sv2v_reg ,
  \piso.data_r_2870_sv2v_reg ,\piso.data_r_2869_sv2v_reg ,
  \piso.data_r_2868_sv2v_reg ,\piso.data_r_2867_sv2v_reg ,\piso.data_r_2866_sv2v_reg ,
  \piso.data_r_2865_sv2v_reg ,\piso.data_r_2864_sv2v_reg ,\piso.data_r_2863_sv2v_reg ,
  \piso.data_r_2862_sv2v_reg ,\piso.data_r_2861_sv2v_reg ,\piso.data_r_2860_sv2v_reg ,
  \piso.data_r_2859_sv2v_reg ,\piso.data_r_2858_sv2v_reg ,\piso.data_r_2857_sv2v_reg ,
  \piso.data_r_2856_sv2v_reg ,\piso.data_r_2855_sv2v_reg ,\piso.data_r_2854_sv2v_reg ,
  \piso.data_r_2853_sv2v_reg ,\piso.data_r_2852_sv2v_reg ,\piso.data_r_2851_sv2v_reg ,
  \piso.data_r_2850_sv2v_reg ,\piso.data_r_2849_sv2v_reg ,
  \piso.data_r_2848_sv2v_reg ,\piso.data_r_2847_sv2v_reg ,\piso.data_r_2846_sv2v_reg ,
  \piso.data_r_2845_sv2v_reg ,\piso.data_r_2844_sv2v_reg ,\piso.data_r_2843_sv2v_reg ,
  \piso.data_r_2842_sv2v_reg ,\piso.data_r_2841_sv2v_reg ,\piso.data_r_2840_sv2v_reg ,
  \piso.data_r_2839_sv2v_reg ,\piso.data_r_2838_sv2v_reg ,\piso.data_r_2837_sv2v_reg ,
  \piso.data_r_2836_sv2v_reg ,\piso.data_r_2835_sv2v_reg ,\piso.data_r_2834_sv2v_reg ,
  \piso.data_r_2833_sv2v_reg ,\piso.data_r_2832_sv2v_reg ,\piso.data_r_2831_sv2v_reg ,
  \piso.data_r_2830_sv2v_reg ,\piso.data_r_2829_sv2v_reg ,
  \piso.data_r_2828_sv2v_reg ,\piso.data_r_2827_sv2v_reg ,\piso.data_r_2826_sv2v_reg ,
  \piso.data_r_2825_sv2v_reg ,\piso.data_r_2824_sv2v_reg ,\piso.data_r_2823_sv2v_reg ,
  \piso.data_r_2822_sv2v_reg ,\piso.data_r_2821_sv2v_reg ,\piso.data_r_2820_sv2v_reg ,
  \piso.data_r_2819_sv2v_reg ,\piso.data_r_2818_sv2v_reg ,\piso.data_r_2817_sv2v_reg ,
  \piso.data_r_2816_sv2v_reg ,\piso.data_r_2815_sv2v_reg ,\piso.data_r_2814_sv2v_reg ,
  \piso.data_r_2813_sv2v_reg ,\piso.data_r_2812_sv2v_reg ,\piso.data_r_2811_sv2v_reg ,
  \piso.data_r_2810_sv2v_reg ,\piso.data_r_2809_sv2v_reg ,
  \piso.data_r_2808_sv2v_reg ,\piso.data_r_2807_sv2v_reg ,\piso.data_r_2806_sv2v_reg ,
  \piso.data_r_2805_sv2v_reg ,\piso.data_r_2804_sv2v_reg ,\piso.data_r_2803_sv2v_reg ,
  \piso.data_r_2802_sv2v_reg ,\piso.data_r_2801_sv2v_reg ,\piso.data_r_2800_sv2v_reg ,
  \piso.data_r_2799_sv2v_reg ,\piso.data_r_2798_sv2v_reg ,\piso.data_r_2797_sv2v_reg ,
  \piso.data_r_2796_sv2v_reg ,\piso.data_r_2795_sv2v_reg ,\piso.data_r_2794_sv2v_reg ,
  \piso.data_r_2793_sv2v_reg ,\piso.data_r_2792_sv2v_reg ,\piso.data_r_2791_sv2v_reg ,
  \piso.data_r_2790_sv2v_reg ,\piso.data_r_2789_sv2v_reg ,
  \piso.data_r_2788_sv2v_reg ,\piso.data_r_2787_sv2v_reg ,\piso.data_r_2786_sv2v_reg ,
  \piso.data_r_2785_sv2v_reg ,\piso.data_r_2784_sv2v_reg ,\piso.data_r_2783_sv2v_reg ,
  \piso.data_r_2782_sv2v_reg ,\piso.data_r_2781_sv2v_reg ,\piso.data_r_2780_sv2v_reg ,
  \piso.data_r_2779_sv2v_reg ,\piso.data_r_2778_sv2v_reg ,\piso.data_r_2777_sv2v_reg ,
  \piso.data_r_2776_sv2v_reg ,\piso.data_r_2775_sv2v_reg ,\piso.data_r_2774_sv2v_reg ,
  \piso.data_r_2773_sv2v_reg ,\piso.data_r_2772_sv2v_reg ,\piso.data_r_2771_sv2v_reg ,
  \piso.data_r_2770_sv2v_reg ,\piso.data_r_2769_sv2v_reg ,
  \piso.data_r_2768_sv2v_reg ,\piso.data_r_2767_sv2v_reg ,\piso.data_r_2766_sv2v_reg ,
  \piso.data_r_2765_sv2v_reg ,\piso.data_r_2764_sv2v_reg ,\piso.data_r_2763_sv2v_reg ,
  \piso.data_r_2762_sv2v_reg ,\piso.data_r_2761_sv2v_reg ,\piso.data_r_2760_sv2v_reg ,
  \piso.data_r_2759_sv2v_reg ,\piso.data_r_2758_sv2v_reg ,\piso.data_r_2757_sv2v_reg ,
  \piso.data_r_2756_sv2v_reg ,\piso.data_r_2755_sv2v_reg ,\piso.data_r_2754_sv2v_reg ,
  \piso.data_r_2753_sv2v_reg ,\piso.data_r_2752_sv2v_reg ,\piso.data_r_2751_sv2v_reg ,
  \piso.data_r_2750_sv2v_reg ,\piso.data_r_2749_sv2v_reg ,
  \piso.data_r_2748_sv2v_reg ,\piso.data_r_2747_sv2v_reg ,\piso.data_r_2746_sv2v_reg ,
  \piso.data_r_2745_sv2v_reg ,\piso.data_r_2744_sv2v_reg ,\piso.data_r_2743_sv2v_reg ,
  \piso.data_r_2742_sv2v_reg ,\piso.data_r_2741_sv2v_reg ,\piso.data_r_2740_sv2v_reg ,
  \piso.data_r_2739_sv2v_reg ,\piso.data_r_2738_sv2v_reg ,\piso.data_r_2737_sv2v_reg ,
  \piso.data_r_2736_sv2v_reg ,\piso.data_r_2735_sv2v_reg ,\piso.data_r_2734_sv2v_reg ,
  \piso.data_r_2733_sv2v_reg ,\piso.data_r_2732_sv2v_reg ,\piso.data_r_2731_sv2v_reg ,
  \piso.data_r_2730_sv2v_reg ,\piso.data_r_2729_sv2v_reg ,
  \piso.data_r_2728_sv2v_reg ,\piso.data_r_2727_sv2v_reg ,\piso.data_r_2726_sv2v_reg ,
  \piso.data_r_2725_sv2v_reg ,\piso.data_r_2724_sv2v_reg ,\piso.data_r_2723_sv2v_reg ,
  \piso.data_r_2722_sv2v_reg ,\piso.data_r_2721_sv2v_reg ,\piso.data_r_2720_sv2v_reg ,
  \piso.data_r_2719_sv2v_reg ,\piso.data_r_2718_sv2v_reg ,\piso.data_r_2717_sv2v_reg ,
  \piso.data_r_2716_sv2v_reg ,\piso.data_r_2715_sv2v_reg ,\piso.data_r_2714_sv2v_reg ,
  \piso.data_r_2713_sv2v_reg ,\piso.data_r_2712_sv2v_reg ,\piso.data_r_2711_sv2v_reg ,
  \piso.data_r_2710_sv2v_reg ,\piso.data_r_2709_sv2v_reg ,
  \piso.data_r_2708_sv2v_reg ,\piso.data_r_2707_sv2v_reg ,\piso.data_r_2706_sv2v_reg ,
  \piso.data_r_2705_sv2v_reg ,\piso.data_r_2704_sv2v_reg ,\piso.data_r_2703_sv2v_reg ,
  \piso.data_r_2702_sv2v_reg ,\piso.data_r_2701_sv2v_reg ,\piso.data_r_2700_sv2v_reg ,
  \piso.data_r_2699_sv2v_reg ,\piso.data_r_2698_sv2v_reg ,\piso.data_r_2697_sv2v_reg ,
  \piso.data_r_2696_sv2v_reg ,\piso.data_r_2695_sv2v_reg ,\piso.data_r_2694_sv2v_reg ,
  \piso.data_r_2693_sv2v_reg ,\piso.data_r_2692_sv2v_reg ,\piso.data_r_2691_sv2v_reg ,
  \piso.data_r_2690_sv2v_reg ,\piso.data_r_2689_sv2v_reg ,
  \piso.data_r_2688_sv2v_reg ,\piso.data_r_2687_sv2v_reg ,\piso.data_r_2686_sv2v_reg ,
  \piso.data_r_2685_sv2v_reg ,\piso.data_r_2684_sv2v_reg ,\piso.data_r_2683_sv2v_reg ,
  \piso.data_r_2682_sv2v_reg ,\piso.data_r_2681_sv2v_reg ,\piso.data_r_2680_sv2v_reg ,
  \piso.data_r_2679_sv2v_reg ,\piso.data_r_2678_sv2v_reg ,\piso.data_r_2677_sv2v_reg ,
  \piso.data_r_2676_sv2v_reg ,\piso.data_r_2675_sv2v_reg ,\piso.data_r_2674_sv2v_reg ,
  \piso.data_r_2673_sv2v_reg ,\piso.data_r_2672_sv2v_reg ,\piso.data_r_2671_sv2v_reg ,
  \piso.data_r_2670_sv2v_reg ,\piso.data_r_2669_sv2v_reg ,
  \piso.data_r_2668_sv2v_reg ,\piso.data_r_2667_sv2v_reg ,\piso.data_r_2666_sv2v_reg ,
  \piso.data_r_2665_sv2v_reg ,\piso.data_r_2664_sv2v_reg ,\piso.data_r_2663_sv2v_reg ,
  \piso.data_r_2662_sv2v_reg ,\piso.data_r_2661_sv2v_reg ,\piso.data_r_2660_sv2v_reg ,
  \piso.data_r_2659_sv2v_reg ,\piso.data_r_2658_sv2v_reg ,\piso.data_r_2657_sv2v_reg ,
  \piso.data_r_2656_sv2v_reg ,\piso.data_r_2655_sv2v_reg ,\piso.data_r_2654_sv2v_reg ,
  \piso.data_r_2653_sv2v_reg ,\piso.data_r_2652_sv2v_reg ,\piso.data_r_2651_sv2v_reg ,
  \piso.data_r_2650_sv2v_reg ,\piso.data_r_2649_sv2v_reg ,
  \piso.data_r_2648_sv2v_reg ,\piso.data_r_2647_sv2v_reg ,\piso.data_r_2646_sv2v_reg ,
  \piso.data_r_2645_sv2v_reg ,\piso.data_r_2644_sv2v_reg ,\piso.data_r_2643_sv2v_reg ,
  \piso.data_r_2642_sv2v_reg ,\piso.data_r_2641_sv2v_reg ,\piso.data_r_2640_sv2v_reg ,
  \piso.data_r_2639_sv2v_reg ,\piso.data_r_2638_sv2v_reg ,\piso.data_r_2637_sv2v_reg ,
  \piso.data_r_2636_sv2v_reg ,\piso.data_r_2635_sv2v_reg ,\piso.data_r_2634_sv2v_reg ,
  \piso.data_r_2633_sv2v_reg ,\piso.data_r_2632_sv2v_reg ,\piso.data_r_2631_sv2v_reg ,
  \piso.data_r_2630_sv2v_reg ,\piso.data_r_2629_sv2v_reg ,
  \piso.data_r_2628_sv2v_reg ,\piso.data_r_2627_sv2v_reg ,\piso.data_r_2626_sv2v_reg ,
  \piso.data_r_2625_sv2v_reg ,\piso.data_r_2624_sv2v_reg ,\piso.data_r_2623_sv2v_reg ,
  \piso.data_r_2622_sv2v_reg ,\piso.data_r_2621_sv2v_reg ,\piso.data_r_2620_sv2v_reg ,
  \piso.data_r_2619_sv2v_reg ,\piso.data_r_2618_sv2v_reg ,\piso.data_r_2617_sv2v_reg ,
  \piso.data_r_2616_sv2v_reg ,\piso.data_r_2615_sv2v_reg ,\piso.data_r_2614_sv2v_reg ,
  \piso.data_r_2613_sv2v_reg ,\piso.data_r_2612_sv2v_reg ,\piso.data_r_2611_sv2v_reg ,
  \piso.data_r_2610_sv2v_reg ,\piso.data_r_2609_sv2v_reg ,
  \piso.data_r_2608_sv2v_reg ,\piso.data_r_2607_sv2v_reg ,\piso.data_r_2606_sv2v_reg ,
  \piso.data_r_2605_sv2v_reg ,\piso.data_r_2604_sv2v_reg ,\piso.data_r_2603_sv2v_reg ,
  \piso.data_r_2602_sv2v_reg ,\piso.data_r_2601_sv2v_reg ,\piso.data_r_2600_sv2v_reg ,
  \piso.data_r_2599_sv2v_reg ,\piso.data_r_2598_sv2v_reg ,\piso.data_r_2597_sv2v_reg ,
  \piso.data_r_2596_sv2v_reg ,\piso.data_r_2595_sv2v_reg ,\piso.data_r_2594_sv2v_reg ,
  \piso.data_r_2593_sv2v_reg ,\piso.data_r_2592_sv2v_reg ,\piso.data_r_2591_sv2v_reg ,
  \piso.data_r_2590_sv2v_reg ,\piso.data_r_2589_sv2v_reg ,
  \piso.data_r_2588_sv2v_reg ,\piso.data_r_2587_sv2v_reg ,\piso.data_r_2586_sv2v_reg ,
  \piso.data_r_2585_sv2v_reg ,\piso.data_r_2584_sv2v_reg ,\piso.data_r_2583_sv2v_reg ,
  \piso.data_r_2582_sv2v_reg ,\piso.data_r_2581_sv2v_reg ,\piso.data_r_2580_sv2v_reg ,
  \piso.data_r_2579_sv2v_reg ,\piso.data_r_2578_sv2v_reg ,\piso.data_r_2577_sv2v_reg ,
  \piso.data_r_2576_sv2v_reg ,\piso.data_r_2575_sv2v_reg ,\piso.data_r_2574_sv2v_reg ,
  \piso.data_r_2573_sv2v_reg ,\piso.data_r_2572_sv2v_reg ,\piso.data_r_2571_sv2v_reg ,
  \piso.data_r_2570_sv2v_reg ,\piso.data_r_2569_sv2v_reg ,
  \piso.data_r_2568_sv2v_reg ,\piso.data_r_2567_sv2v_reg ,\piso.data_r_2566_sv2v_reg ,
  \piso.data_r_2565_sv2v_reg ,\piso.data_r_2564_sv2v_reg ,\piso.data_r_2563_sv2v_reg ,
  \piso.data_r_2562_sv2v_reg ,\piso.data_r_2561_sv2v_reg ,\piso.data_r_2560_sv2v_reg ,
  \piso.data_r_2559_sv2v_reg ,\piso.data_r_2558_sv2v_reg ,\piso.data_r_2557_sv2v_reg ,
  \piso.data_r_2556_sv2v_reg ,\piso.data_r_2555_sv2v_reg ,\piso.data_r_2554_sv2v_reg ,
  \piso.data_r_2553_sv2v_reg ,\piso.data_r_2552_sv2v_reg ,\piso.data_r_2551_sv2v_reg ,
  \piso.data_r_2550_sv2v_reg ,\piso.data_r_2549_sv2v_reg ,
  \piso.data_r_2548_sv2v_reg ,\piso.data_r_2547_sv2v_reg ,\piso.data_r_2546_sv2v_reg ,
  \piso.data_r_2545_sv2v_reg ,\piso.data_r_2544_sv2v_reg ,\piso.data_r_2543_sv2v_reg ,
  \piso.data_r_2542_sv2v_reg ,\piso.data_r_2541_sv2v_reg ,\piso.data_r_2540_sv2v_reg ,
  \piso.data_r_2539_sv2v_reg ,\piso.data_r_2538_sv2v_reg ,\piso.data_r_2537_sv2v_reg ,
  \piso.data_r_2536_sv2v_reg ,\piso.data_r_2535_sv2v_reg ,\piso.data_r_2534_sv2v_reg ,
  \piso.data_r_2533_sv2v_reg ,\piso.data_r_2532_sv2v_reg ,\piso.data_r_2531_sv2v_reg ,
  \piso.data_r_2530_sv2v_reg ,\piso.data_r_2529_sv2v_reg ,
  \piso.data_r_2528_sv2v_reg ,\piso.data_r_2527_sv2v_reg ,\piso.data_r_2526_sv2v_reg ,
  \piso.data_r_2525_sv2v_reg ,\piso.data_r_2524_sv2v_reg ,\piso.data_r_2523_sv2v_reg ,
  \piso.data_r_2522_sv2v_reg ,\piso.data_r_2521_sv2v_reg ,\piso.data_r_2520_sv2v_reg ,
  \piso.data_r_2519_sv2v_reg ,\piso.data_r_2518_sv2v_reg ,\piso.data_r_2517_sv2v_reg ,
  \piso.data_r_2516_sv2v_reg ,\piso.data_r_2515_sv2v_reg ,\piso.data_r_2514_sv2v_reg ,
  \piso.data_r_2513_sv2v_reg ,\piso.data_r_2512_sv2v_reg ,\piso.data_r_2511_sv2v_reg ,
  \piso.data_r_2510_sv2v_reg ,\piso.data_r_2509_sv2v_reg ,
  \piso.data_r_2508_sv2v_reg ,\piso.data_r_2507_sv2v_reg ,\piso.data_r_2506_sv2v_reg ,
  \piso.data_r_2505_sv2v_reg ,\piso.data_r_2504_sv2v_reg ,\piso.data_r_2503_sv2v_reg ,
  \piso.data_r_2502_sv2v_reg ,\piso.data_r_2501_sv2v_reg ,\piso.data_r_2500_sv2v_reg ,
  \piso.data_r_2499_sv2v_reg ,\piso.data_r_2498_sv2v_reg ,\piso.data_r_2497_sv2v_reg ,
  \piso.data_r_2496_sv2v_reg ,\piso.data_r_2495_sv2v_reg ,\piso.data_r_2494_sv2v_reg ,
  \piso.data_r_2493_sv2v_reg ,\piso.data_r_2492_sv2v_reg ,\piso.data_r_2491_sv2v_reg ,
  \piso.data_r_2490_sv2v_reg ,\piso.data_r_2489_sv2v_reg ,
  \piso.data_r_2488_sv2v_reg ,\piso.data_r_2487_sv2v_reg ,\piso.data_r_2486_sv2v_reg ,
  \piso.data_r_2485_sv2v_reg ,\piso.data_r_2484_sv2v_reg ,\piso.data_r_2483_sv2v_reg ,
  \piso.data_r_2482_sv2v_reg ,\piso.data_r_2481_sv2v_reg ,\piso.data_r_2480_sv2v_reg ,
  \piso.data_r_2479_sv2v_reg ,\piso.data_r_2478_sv2v_reg ,\piso.data_r_2477_sv2v_reg ,
  \piso.data_r_2476_sv2v_reg ,\piso.data_r_2475_sv2v_reg ,\piso.data_r_2474_sv2v_reg ,
  \piso.data_r_2473_sv2v_reg ,\piso.data_r_2472_sv2v_reg ,\piso.data_r_2471_sv2v_reg ,
  \piso.data_r_2470_sv2v_reg ,\piso.data_r_2469_sv2v_reg ,
  \piso.data_r_2468_sv2v_reg ,\piso.data_r_2467_sv2v_reg ,\piso.data_r_2466_sv2v_reg ,
  \piso.data_r_2465_sv2v_reg ,\piso.data_r_2464_sv2v_reg ,\piso.data_r_2463_sv2v_reg ,
  \piso.data_r_2462_sv2v_reg ,\piso.data_r_2461_sv2v_reg ,\piso.data_r_2460_sv2v_reg ,
  \piso.data_r_2459_sv2v_reg ,\piso.data_r_2458_sv2v_reg ,\piso.data_r_2457_sv2v_reg ,
  \piso.data_r_2456_sv2v_reg ,\piso.data_r_2455_sv2v_reg ,\piso.data_r_2454_sv2v_reg ,
  \piso.data_r_2453_sv2v_reg ,\piso.data_r_2452_sv2v_reg ,\piso.data_r_2451_sv2v_reg ,
  \piso.data_r_2450_sv2v_reg ,\piso.data_r_2449_sv2v_reg ,
  \piso.data_r_2448_sv2v_reg ,\piso.data_r_2447_sv2v_reg ,\piso.data_r_2446_sv2v_reg ,
  \piso.data_r_2445_sv2v_reg ,\piso.data_r_2444_sv2v_reg ,\piso.data_r_2443_sv2v_reg ,
  \piso.data_r_2442_sv2v_reg ,\piso.data_r_2441_sv2v_reg ,\piso.data_r_2440_sv2v_reg ,
  \piso.data_r_2439_sv2v_reg ,\piso.data_r_2438_sv2v_reg ,\piso.data_r_2437_sv2v_reg ,
  \piso.data_r_2436_sv2v_reg ,\piso.data_r_2435_sv2v_reg ,\piso.data_r_2434_sv2v_reg ,
  \piso.data_r_2433_sv2v_reg ,\piso.data_r_2432_sv2v_reg ,\piso.data_r_2431_sv2v_reg ,
  \piso.data_r_2430_sv2v_reg ,\piso.data_r_2429_sv2v_reg ,
  \piso.data_r_2428_sv2v_reg ,\piso.data_r_2427_sv2v_reg ,\piso.data_r_2426_sv2v_reg ,
  \piso.data_r_2425_sv2v_reg ,\piso.data_r_2424_sv2v_reg ,\piso.data_r_2423_sv2v_reg ,
  \piso.data_r_2422_sv2v_reg ,\piso.data_r_2421_sv2v_reg ,\piso.data_r_2420_sv2v_reg ,
  \piso.data_r_2419_sv2v_reg ,\piso.data_r_2418_sv2v_reg ,\piso.data_r_2417_sv2v_reg ,
  \piso.data_r_2416_sv2v_reg ,\piso.data_r_2415_sv2v_reg ,\piso.data_r_2414_sv2v_reg ,
  \piso.data_r_2413_sv2v_reg ,\piso.data_r_2412_sv2v_reg ,\piso.data_r_2411_sv2v_reg ,
  \piso.data_r_2410_sv2v_reg ,\piso.data_r_2409_sv2v_reg ,
  \piso.data_r_2408_sv2v_reg ,\piso.data_r_2407_sv2v_reg ,\piso.data_r_2406_sv2v_reg ,
  \piso.data_r_2405_sv2v_reg ,\piso.data_r_2404_sv2v_reg ,\piso.data_r_2403_sv2v_reg ,
  \piso.data_r_2402_sv2v_reg ,\piso.data_r_2401_sv2v_reg ,\piso.data_r_2400_sv2v_reg ,
  \piso.data_r_2399_sv2v_reg ,\piso.data_r_2398_sv2v_reg ,\piso.data_r_2397_sv2v_reg ,
  \piso.data_r_2396_sv2v_reg ,\piso.data_r_2395_sv2v_reg ,\piso.data_r_2394_sv2v_reg ,
  \piso.data_r_2393_sv2v_reg ,\piso.data_r_2392_sv2v_reg ,\piso.data_r_2391_sv2v_reg ,
  \piso.data_r_2390_sv2v_reg ,\piso.data_r_2389_sv2v_reg ,
  \piso.data_r_2388_sv2v_reg ,\piso.data_r_2387_sv2v_reg ,\piso.data_r_2386_sv2v_reg ,
  \piso.data_r_2385_sv2v_reg ,\piso.data_r_2384_sv2v_reg ,\piso.data_r_2383_sv2v_reg ,
  \piso.data_r_2382_sv2v_reg ,\piso.data_r_2381_sv2v_reg ,\piso.data_r_2380_sv2v_reg ,
  \piso.data_r_2379_sv2v_reg ,\piso.data_r_2378_sv2v_reg ,\piso.data_r_2377_sv2v_reg ,
  \piso.data_r_2376_sv2v_reg ,\piso.data_r_2375_sv2v_reg ,\piso.data_r_2374_sv2v_reg ,
  \piso.data_r_2373_sv2v_reg ,\piso.data_r_2372_sv2v_reg ,\piso.data_r_2371_sv2v_reg ,
  \piso.data_r_2370_sv2v_reg ,\piso.data_r_2369_sv2v_reg ,
  \piso.data_r_2368_sv2v_reg ,\piso.data_r_2367_sv2v_reg ,\piso.data_r_2366_sv2v_reg ,
  \piso.data_r_2365_sv2v_reg ,\piso.data_r_2364_sv2v_reg ,\piso.data_r_2363_sv2v_reg ,
  \piso.data_r_2362_sv2v_reg ,\piso.data_r_2361_sv2v_reg ,\piso.data_r_2360_sv2v_reg ,
  \piso.data_r_2359_sv2v_reg ,\piso.data_r_2358_sv2v_reg ,\piso.data_r_2357_sv2v_reg ,
  \piso.data_r_2356_sv2v_reg ,\piso.data_r_2355_sv2v_reg ,\piso.data_r_2354_sv2v_reg ,
  \piso.data_r_2353_sv2v_reg ,\piso.data_r_2352_sv2v_reg ,\piso.data_r_2351_sv2v_reg ,
  \piso.data_r_2350_sv2v_reg ,\piso.data_r_2349_sv2v_reg ,
  \piso.data_r_2348_sv2v_reg ,\piso.data_r_2347_sv2v_reg ,\piso.data_r_2346_sv2v_reg ,
  \piso.data_r_2345_sv2v_reg ,\piso.data_r_2344_sv2v_reg ,\piso.data_r_2343_sv2v_reg ,
  \piso.data_r_2342_sv2v_reg ,\piso.data_r_2341_sv2v_reg ,\piso.data_r_2340_sv2v_reg ,
  \piso.data_r_2339_sv2v_reg ,\piso.data_r_2338_sv2v_reg ,\piso.data_r_2337_sv2v_reg ,
  \piso.data_r_2336_sv2v_reg ,\piso.data_r_2335_sv2v_reg ,\piso.data_r_2334_sv2v_reg ,
  \piso.data_r_2333_sv2v_reg ,\piso.data_r_2332_sv2v_reg ,\piso.data_r_2331_sv2v_reg ,
  \piso.data_r_2330_sv2v_reg ,\piso.data_r_2329_sv2v_reg ,
  \piso.data_r_2328_sv2v_reg ,\piso.data_r_2327_sv2v_reg ,\piso.data_r_2326_sv2v_reg ,
  \piso.data_r_2325_sv2v_reg ,\piso.data_r_2324_sv2v_reg ,\piso.data_r_2323_sv2v_reg ,
  \piso.data_r_2322_sv2v_reg ,\piso.data_r_2321_sv2v_reg ,\piso.data_r_2320_sv2v_reg ,
  \piso.data_r_2319_sv2v_reg ,\piso.data_r_2318_sv2v_reg ,\piso.data_r_2317_sv2v_reg ,
  \piso.data_r_2316_sv2v_reg ,\piso.data_r_2315_sv2v_reg ,\piso.data_r_2314_sv2v_reg ,
  \piso.data_r_2313_sv2v_reg ,\piso.data_r_2312_sv2v_reg ,\piso.data_r_2311_sv2v_reg ,
  \piso.data_r_2310_sv2v_reg ,\piso.data_r_2309_sv2v_reg ,
  \piso.data_r_2308_sv2v_reg ,\piso.data_r_2307_sv2v_reg ,\piso.data_r_2306_sv2v_reg ,
  \piso.data_r_2305_sv2v_reg ,\piso.data_r_2304_sv2v_reg ,\piso.data_r_2303_sv2v_reg ,
  \piso.data_r_2302_sv2v_reg ,\piso.data_r_2301_sv2v_reg ,\piso.data_r_2300_sv2v_reg ,
  \piso.data_r_2299_sv2v_reg ,\piso.data_r_2298_sv2v_reg ,\piso.data_r_2297_sv2v_reg ,
  \piso.data_r_2296_sv2v_reg ,\piso.data_r_2295_sv2v_reg ,\piso.data_r_2294_sv2v_reg ,
  \piso.data_r_2293_sv2v_reg ,\piso.data_r_2292_sv2v_reg ,\piso.data_r_2291_sv2v_reg ,
  \piso.data_r_2290_sv2v_reg ,\piso.data_r_2289_sv2v_reg ,
  \piso.data_r_2288_sv2v_reg ,\piso.data_r_2287_sv2v_reg ,\piso.data_r_2286_sv2v_reg ,
  \piso.data_r_2285_sv2v_reg ,\piso.data_r_2284_sv2v_reg ,\piso.data_r_2283_sv2v_reg ,
  \piso.data_r_2282_sv2v_reg ,\piso.data_r_2281_sv2v_reg ,\piso.data_r_2280_sv2v_reg ,
  \piso.data_r_2279_sv2v_reg ,\piso.data_r_2278_sv2v_reg ,\piso.data_r_2277_sv2v_reg ,
  \piso.data_r_2276_sv2v_reg ,\piso.data_r_2275_sv2v_reg ,\piso.data_r_2274_sv2v_reg ,
  \piso.data_r_2273_sv2v_reg ,\piso.data_r_2272_sv2v_reg ,\piso.data_r_2271_sv2v_reg ,
  \piso.data_r_2270_sv2v_reg ,\piso.data_r_2269_sv2v_reg ,
  \piso.data_r_2268_sv2v_reg ,\piso.data_r_2267_sv2v_reg ,\piso.data_r_2266_sv2v_reg ,
  \piso.data_r_2265_sv2v_reg ,\piso.data_r_2264_sv2v_reg ,\piso.data_r_2263_sv2v_reg ,
  \piso.data_r_2262_sv2v_reg ,\piso.data_r_2261_sv2v_reg ,\piso.data_r_2260_sv2v_reg ,
  \piso.data_r_2259_sv2v_reg ,\piso.data_r_2258_sv2v_reg ,\piso.data_r_2257_sv2v_reg ,
  \piso.data_r_2256_sv2v_reg ,\piso.data_r_2255_sv2v_reg ,\piso.data_r_2254_sv2v_reg ,
  \piso.data_r_2253_sv2v_reg ,\piso.data_r_2252_sv2v_reg ,\piso.data_r_2251_sv2v_reg ,
  \piso.data_r_2250_sv2v_reg ,\piso.data_r_2249_sv2v_reg ,
  \piso.data_r_2248_sv2v_reg ,\piso.data_r_2247_sv2v_reg ,\piso.data_r_2246_sv2v_reg ,
  \piso.data_r_2245_sv2v_reg ,\piso.data_r_2244_sv2v_reg ,\piso.data_r_2243_sv2v_reg ,
  \piso.data_r_2242_sv2v_reg ,\piso.data_r_2241_sv2v_reg ,\piso.data_r_2240_sv2v_reg ,
  \piso.data_r_2239_sv2v_reg ,\piso.data_r_2238_sv2v_reg ,\piso.data_r_2237_sv2v_reg ,
  \piso.data_r_2236_sv2v_reg ,\piso.data_r_2235_sv2v_reg ,\piso.data_r_2234_sv2v_reg ,
  \piso.data_r_2233_sv2v_reg ,\piso.data_r_2232_sv2v_reg ,\piso.data_r_2231_sv2v_reg ,
  \piso.data_r_2230_sv2v_reg ,\piso.data_r_2229_sv2v_reg ,
  \piso.data_r_2228_sv2v_reg ,\piso.data_r_2227_sv2v_reg ,\piso.data_r_2226_sv2v_reg ,
  \piso.data_r_2225_sv2v_reg ,\piso.data_r_2224_sv2v_reg ,\piso.data_r_2223_sv2v_reg ,
  \piso.data_r_2222_sv2v_reg ,\piso.data_r_2221_sv2v_reg ,\piso.data_r_2220_sv2v_reg ,
  \piso.data_r_2219_sv2v_reg ,\piso.data_r_2218_sv2v_reg ,\piso.data_r_2217_sv2v_reg ,
  \piso.data_r_2216_sv2v_reg ,\piso.data_r_2215_sv2v_reg ,\piso.data_r_2214_sv2v_reg ,
  \piso.data_r_2213_sv2v_reg ,\piso.data_r_2212_sv2v_reg ,\piso.data_r_2211_sv2v_reg ,
  \piso.data_r_2210_sv2v_reg ,\piso.data_r_2209_sv2v_reg ,
  \piso.data_r_2208_sv2v_reg ,\piso.data_r_2207_sv2v_reg ,\piso.data_r_2206_sv2v_reg ,
  \piso.data_r_2205_sv2v_reg ,\piso.data_r_2204_sv2v_reg ,\piso.data_r_2203_sv2v_reg ,
  \piso.data_r_2202_sv2v_reg ,\piso.data_r_2201_sv2v_reg ,\piso.data_r_2200_sv2v_reg ,
  \piso.data_r_2199_sv2v_reg ,\piso.data_r_2198_sv2v_reg ,\piso.data_r_2197_sv2v_reg ,
  \piso.data_r_2196_sv2v_reg ,\piso.data_r_2195_sv2v_reg ,\piso.data_r_2194_sv2v_reg ,
  \piso.data_r_2193_sv2v_reg ,\piso.data_r_2192_sv2v_reg ,\piso.data_r_2191_sv2v_reg ,
  \piso.data_r_2190_sv2v_reg ,\piso.data_r_2189_sv2v_reg ,
  \piso.data_r_2188_sv2v_reg ,\piso.data_r_2187_sv2v_reg ,\piso.data_r_2186_sv2v_reg ,
  \piso.data_r_2185_sv2v_reg ,\piso.data_r_2184_sv2v_reg ,\piso.data_r_2183_sv2v_reg ,
  \piso.data_r_2182_sv2v_reg ,\piso.data_r_2181_sv2v_reg ,\piso.data_r_2180_sv2v_reg ,
  \piso.data_r_2179_sv2v_reg ,\piso.data_r_2178_sv2v_reg ,\piso.data_r_2177_sv2v_reg ,
  \piso.data_r_2176_sv2v_reg ,\piso.data_r_2175_sv2v_reg ,\piso.data_r_2174_sv2v_reg ,
  \piso.data_r_2173_sv2v_reg ,\piso.data_r_2172_sv2v_reg ,\piso.data_r_2171_sv2v_reg ,
  \piso.data_r_2170_sv2v_reg ,\piso.data_r_2169_sv2v_reg ,
  \piso.data_r_2168_sv2v_reg ,\piso.data_r_2167_sv2v_reg ,\piso.data_r_2166_sv2v_reg ,
  \piso.data_r_2165_sv2v_reg ,\piso.data_r_2164_sv2v_reg ,\piso.data_r_2163_sv2v_reg ,
  \piso.data_r_2162_sv2v_reg ,\piso.data_r_2161_sv2v_reg ,\piso.data_r_2160_sv2v_reg ,
  \piso.data_r_2159_sv2v_reg ,\piso.data_r_2158_sv2v_reg ,\piso.data_r_2157_sv2v_reg ,
  \piso.data_r_2156_sv2v_reg ,\piso.data_r_2155_sv2v_reg ,\piso.data_r_2154_sv2v_reg ,
  \piso.data_r_2153_sv2v_reg ,\piso.data_r_2152_sv2v_reg ,\piso.data_r_2151_sv2v_reg ,
  \piso.data_r_2150_sv2v_reg ,\piso.data_r_2149_sv2v_reg ,
  \piso.data_r_2148_sv2v_reg ,\piso.data_r_2147_sv2v_reg ,\piso.data_r_2146_sv2v_reg ,
  \piso.data_r_2145_sv2v_reg ,\piso.data_r_2144_sv2v_reg ,\piso.data_r_2143_sv2v_reg ,
  \piso.data_r_2142_sv2v_reg ,\piso.data_r_2141_sv2v_reg ,\piso.data_r_2140_sv2v_reg ,
  \piso.data_r_2139_sv2v_reg ,\piso.data_r_2138_sv2v_reg ,\piso.data_r_2137_sv2v_reg ,
  \piso.data_r_2136_sv2v_reg ,\piso.data_r_2135_sv2v_reg ,\piso.data_r_2134_sv2v_reg ,
  \piso.data_r_2133_sv2v_reg ,\piso.data_r_2132_sv2v_reg ,\piso.data_r_2131_sv2v_reg ,
  \piso.data_r_2130_sv2v_reg ,\piso.data_r_2129_sv2v_reg ,
  \piso.data_r_2128_sv2v_reg ,\piso.data_r_2127_sv2v_reg ,\piso.data_r_2126_sv2v_reg ,
  \piso.data_r_2125_sv2v_reg ,\piso.data_r_2124_sv2v_reg ,\piso.data_r_2123_sv2v_reg ,
  \piso.data_r_2122_sv2v_reg ,\piso.data_r_2121_sv2v_reg ,\piso.data_r_2120_sv2v_reg ,
  \piso.data_r_2119_sv2v_reg ,\piso.data_r_2118_sv2v_reg ,\piso.data_r_2117_sv2v_reg ,
  \piso.data_r_2116_sv2v_reg ,\piso.data_r_2115_sv2v_reg ,\piso.data_r_2114_sv2v_reg ,
  \piso.data_r_2113_sv2v_reg ,\piso.data_r_2112_sv2v_reg ,\piso.data_r_2111_sv2v_reg ,
  \piso.data_r_2110_sv2v_reg ,\piso.data_r_2109_sv2v_reg ,
  \piso.data_r_2108_sv2v_reg ,\piso.data_r_2107_sv2v_reg ,\piso.data_r_2106_sv2v_reg ,
  \piso.data_r_2105_sv2v_reg ,\piso.data_r_2104_sv2v_reg ,\piso.data_r_2103_sv2v_reg ,
  \piso.data_r_2102_sv2v_reg ,\piso.data_r_2101_sv2v_reg ,\piso.data_r_2100_sv2v_reg ,
  \piso.data_r_2099_sv2v_reg ,\piso.data_r_2098_sv2v_reg ,\piso.data_r_2097_sv2v_reg ,
  \piso.data_r_2096_sv2v_reg ,\piso.data_r_2095_sv2v_reg ,\piso.data_r_2094_sv2v_reg ,
  \piso.data_r_2093_sv2v_reg ,\piso.data_r_2092_sv2v_reg ,\piso.data_r_2091_sv2v_reg ,
  \piso.data_r_2090_sv2v_reg ,\piso.data_r_2089_sv2v_reg ,
  \piso.data_r_2088_sv2v_reg ,\piso.data_r_2087_sv2v_reg ,\piso.data_r_2086_sv2v_reg ,
  \piso.data_r_2085_sv2v_reg ,\piso.data_r_2084_sv2v_reg ,\piso.data_r_2083_sv2v_reg ,
  \piso.data_r_2082_sv2v_reg ,\piso.data_r_2081_sv2v_reg ,\piso.data_r_2080_sv2v_reg ,
  \piso.data_r_2079_sv2v_reg ,\piso.data_r_2078_sv2v_reg ,\piso.data_r_2077_sv2v_reg ,
  \piso.data_r_2076_sv2v_reg ,\piso.data_r_2075_sv2v_reg ,\piso.data_r_2074_sv2v_reg ,
  \piso.data_r_2073_sv2v_reg ,\piso.data_r_2072_sv2v_reg ,\piso.data_r_2071_sv2v_reg ,
  \piso.data_r_2070_sv2v_reg ,\piso.data_r_2069_sv2v_reg ,
  \piso.data_r_2068_sv2v_reg ,\piso.data_r_2067_sv2v_reg ,\piso.data_r_2066_sv2v_reg ,
  \piso.data_r_2065_sv2v_reg ,\piso.data_r_2064_sv2v_reg ,\piso.data_r_2063_sv2v_reg ,
  \piso.data_r_2062_sv2v_reg ,\piso.data_r_2061_sv2v_reg ,\piso.data_r_2060_sv2v_reg ,
  \piso.data_r_2059_sv2v_reg ,\piso.data_r_2058_sv2v_reg ,\piso.data_r_2057_sv2v_reg ,
  \piso.data_r_2056_sv2v_reg ,\piso.data_r_2055_sv2v_reg ,\piso.data_r_2054_sv2v_reg ,
  \piso.data_r_2053_sv2v_reg ,\piso.data_r_2052_sv2v_reg ,\piso.data_r_2051_sv2v_reg ,
  \piso.data_r_2050_sv2v_reg ,\piso.data_r_2049_sv2v_reg ,
  \piso.data_r_2048_sv2v_reg ,\piso.data_r_2047_sv2v_reg ,\piso.data_r_2046_sv2v_reg ,
  \piso.data_r_2045_sv2v_reg ,\piso.data_r_2044_sv2v_reg ,\piso.data_r_2043_sv2v_reg ,
  \piso.data_r_2042_sv2v_reg ,\piso.data_r_2041_sv2v_reg ,\piso.data_r_2040_sv2v_reg ,
  \piso.data_r_2039_sv2v_reg ,\piso.data_r_2038_sv2v_reg ,\piso.data_r_2037_sv2v_reg ,
  \piso.data_r_2036_sv2v_reg ,\piso.data_r_2035_sv2v_reg ,\piso.data_r_2034_sv2v_reg ,
  \piso.data_r_2033_sv2v_reg ,\piso.data_r_2032_sv2v_reg ,\piso.data_r_2031_sv2v_reg ,
  \piso.data_r_2030_sv2v_reg ,\piso.data_r_2029_sv2v_reg ,
  \piso.data_r_2028_sv2v_reg ,\piso.data_r_2027_sv2v_reg ,\piso.data_r_2026_sv2v_reg ,
  \piso.data_r_2025_sv2v_reg ,\piso.data_r_2024_sv2v_reg ,\piso.data_r_2023_sv2v_reg ,
  \piso.data_r_2022_sv2v_reg ,\piso.data_r_2021_sv2v_reg ,\piso.data_r_2020_sv2v_reg ,
  \piso.data_r_2019_sv2v_reg ,\piso.data_r_2018_sv2v_reg ,\piso.data_r_2017_sv2v_reg ,
  \piso.data_r_2016_sv2v_reg ,\piso.data_r_2015_sv2v_reg ,\piso.data_r_2014_sv2v_reg ,
  \piso.data_r_2013_sv2v_reg ,\piso.data_r_2012_sv2v_reg ,\piso.data_r_2011_sv2v_reg ,
  \piso.data_r_2010_sv2v_reg ,\piso.data_r_2009_sv2v_reg ,
  \piso.data_r_2008_sv2v_reg ,\piso.data_r_2007_sv2v_reg ,\piso.data_r_2006_sv2v_reg ,
  \piso.data_r_2005_sv2v_reg ,\piso.data_r_2004_sv2v_reg ,\piso.data_r_2003_sv2v_reg ,
  \piso.data_r_2002_sv2v_reg ,\piso.data_r_2001_sv2v_reg ,\piso.data_r_2000_sv2v_reg ,
  \piso.data_r_1999_sv2v_reg ,\piso.data_r_1998_sv2v_reg ,\piso.data_r_1997_sv2v_reg ,
  \piso.data_r_1996_sv2v_reg ,\piso.data_r_1995_sv2v_reg ,\piso.data_r_1994_sv2v_reg ,
  \piso.data_r_1993_sv2v_reg ,\piso.data_r_1992_sv2v_reg ,\piso.data_r_1991_sv2v_reg ,
  \piso.data_r_1990_sv2v_reg ,\piso.data_r_1989_sv2v_reg ,
  \piso.data_r_1988_sv2v_reg ,\piso.data_r_1987_sv2v_reg ,\piso.data_r_1986_sv2v_reg ,
  \piso.data_r_1985_sv2v_reg ,\piso.data_r_1984_sv2v_reg ,\piso.data_r_1983_sv2v_reg ,
  \piso.data_r_1982_sv2v_reg ,\piso.data_r_1981_sv2v_reg ,\piso.data_r_1980_sv2v_reg ,
  \piso.data_r_1979_sv2v_reg ,\piso.data_r_1978_sv2v_reg ,\piso.data_r_1977_sv2v_reg ,
  \piso.data_r_1976_sv2v_reg ,\piso.data_r_1975_sv2v_reg ,\piso.data_r_1974_sv2v_reg ,
  \piso.data_r_1973_sv2v_reg ,\piso.data_r_1972_sv2v_reg ,\piso.data_r_1971_sv2v_reg ,
  \piso.data_r_1970_sv2v_reg ,\piso.data_r_1969_sv2v_reg ,
  \piso.data_r_1968_sv2v_reg ,\piso.data_r_1967_sv2v_reg ,\piso.data_r_1966_sv2v_reg ,
  \piso.data_r_1965_sv2v_reg ,\piso.data_r_1964_sv2v_reg ,\piso.data_r_1963_sv2v_reg ,
  \piso.data_r_1962_sv2v_reg ,\piso.data_r_1961_sv2v_reg ,\piso.data_r_1960_sv2v_reg ,
  \piso.data_r_1959_sv2v_reg ,\piso.data_r_1958_sv2v_reg ,\piso.data_r_1957_sv2v_reg ,
  \piso.data_r_1956_sv2v_reg ,\piso.data_r_1955_sv2v_reg ,\piso.data_r_1954_sv2v_reg ,
  \piso.data_r_1953_sv2v_reg ,\piso.data_r_1952_sv2v_reg ,\piso.data_r_1951_sv2v_reg ,
  \piso.data_r_1950_sv2v_reg ,\piso.data_r_1949_sv2v_reg ,
  \piso.data_r_1948_sv2v_reg ,\piso.data_r_1947_sv2v_reg ,\piso.data_r_1946_sv2v_reg ,
  \piso.data_r_1945_sv2v_reg ,\piso.data_r_1944_sv2v_reg ,\piso.data_r_1943_sv2v_reg ,
  \piso.data_r_1942_sv2v_reg ,\piso.data_r_1941_sv2v_reg ,\piso.data_r_1940_sv2v_reg ,
  \piso.data_r_1939_sv2v_reg ,\piso.data_r_1938_sv2v_reg ,\piso.data_r_1937_sv2v_reg ,
  \piso.data_r_1936_sv2v_reg ,\piso.data_r_1935_sv2v_reg ,\piso.data_r_1934_sv2v_reg ,
  \piso.data_r_1933_sv2v_reg ,\piso.data_r_1932_sv2v_reg ,\piso.data_r_1931_sv2v_reg ,
  \piso.data_r_1930_sv2v_reg ,\piso.data_r_1929_sv2v_reg ,
  \piso.data_r_1928_sv2v_reg ,\piso.data_r_1927_sv2v_reg ,\piso.data_r_1926_sv2v_reg ,
  \piso.data_r_1925_sv2v_reg ,\piso.data_r_1924_sv2v_reg ,\piso.data_r_1923_sv2v_reg ,
  \piso.data_r_1922_sv2v_reg ,\piso.data_r_1921_sv2v_reg ,\piso.data_r_1920_sv2v_reg ,
  \piso.data_r_1919_sv2v_reg ,\piso.data_r_1918_sv2v_reg ,\piso.data_r_1917_sv2v_reg ,
  \piso.data_r_1916_sv2v_reg ,\piso.data_r_1915_sv2v_reg ,\piso.data_r_1914_sv2v_reg ,
  \piso.data_r_1913_sv2v_reg ,\piso.data_r_1912_sv2v_reg ,\piso.data_r_1911_sv2v_reg ,
  \piso.data_r_1910_sv2v_reg ,\piso.data_r_1909_sv2v_reg ,
  \piso.data_r_1908_sv2v_reg ,\piso.data_r_1907_sv2v_reg ,\piso.data_r_1906_sv2v_reg ,
  \piso.data_r_1905_sv2v_reg ,\piso.data_r_1904_sv2v_reg ,\piso.data_r_1903_sv2v_reg ,
  \piso.data_r_1902_sv2v_reg ,\piso.data_r_1901_sv2v_reg ,\piso.data_r_1900_sv2v_reg ,
  \piso.data_r_1899_sv2v_reg ,\piso.data_r_1898_sv2v_reg ,\piso.data_r_1897_sv2v_reg ,
  \piso.data_r_1896_sv2v_reg ,\piso.data_r_1895_sv2v_reg ,\piso.data_r_1894_sv2v_reg ,
  \piso.data_r_1893_sv2v_reg ,\piso.data_r_1892_sv2v_reg ,\piso.data_r_1891_sv2v_reg ,
  \piso.data_r_1890_sv2v_reg ,\piso.data_r_1889_sv2v_reg ,
  \piso.data_r_1888_sv2v_reg ,\piso.data_r_1887_sv2v_reg ,\piso.data_r_1886_sv2v_reg ,
  \piso.data_r_1885_sv2v_reg ,\piso.data_r_1884_sv2v_reg ,\piso.data_r_1883_sv2v_reg ,
  \piso.data_r_1882_sv2v_reg ,\piso.data_r_1881_sv2v_reg ,\piso.data_r_1880_sv2v_reg ,
  \piso.data_r_1879_sv2v_reg ,\piso.data_r_1878_sv2v_reg ,\piso.data_r_1877_sv2v_reg ,
  \piso.data_r_1876_sv2v_reg ,\piso.data_r_1875_sv2v_reg ,\piso.data_r_1874_sv2v_reg ,
  \piso.data_r_1873_sv2v_reg ,\piso.data_r_1872_sv2v_reg ,\piso.data_r_1871_sv2v_reg ,
  \piso.data_r_1870_sv2v_reg ,\piso.data_r_1869_sv2v_reg ,
  \piso.data_r_1868_sv2v_reg ,\piso.data_r_1867_sv2v_reg ,\piso.data_r_1866_sv2v_reg ,
  \piso.data_r_1865_sv2v_reg ,\piso.data_r_1864_sv2v_reg ,\piso.data_r_1863_sv2v_reg ,
  \piso.data_r_1862_sv2v_reg ,\piso.data_r_1861_sv2v_reg ,\piso.data_r_1860_sv2v_reg ,
  \piso.data_r_1859_sv2v_reg ,\piso.data_r_1858_sv2v_reg ,\piso.data_r_1857_sv2v_reg ,
  \piso.data_r_1856_sv2v_reg ,\piso.data_r_1855_sv2v_reg ,\piso.data_r_1854_sv2v_reg ,
  \piso.data_r_1853_sv2v_reg ,\piso.data_r_1852_sv2v_reg ,\piso.data_r_1851_sv2v_reg ,
  \piso.data_r_1850_sv2v_reg ,\piso.data_r_1849_sv2v_reg ,
  \piso.data_r_1848_sv2v_reg ,\piso.data_r_1847_sv2v_reg ,\piso.data_r_1846_sv2v_reg ,
  \piso.data_r_1845_sv2v_reg ,\piso.data_r_1844_sv2v_reg ,\piso.data_r_1843_sv2v_reg ,
  \piso.data_r_1842_sv2v_reg ,\piso.data_r_1841_sv2v_reg ,\piso.data_r_1840_sv2v_reg ,
  \piso.data_r_1839_sv2v_reg ,\piso.data_r_1838_sv2v_reg ,\piso.data_r_1837_sv2v_reg ,
  \piso.data_r_1836_sv2v_reg ,\piso.data_r_1835_sv2v_reg ,\piso.data_r_1834_sv2v_reg ,
  \piso.data_r_1833_sv2v_reg ,\piso.data_r_1832_sv2v_reg ,\piso.data_r_1831_sv2v_reg ,
  \piso.data_r_1830_sv2v_reg ,\piso.data_r_1829_sv2v_reg ,
  \piso.data_r_1828_sv2v_reg ,\piso.data_r_1827_sv2v_reg ,\piso.data_r_1826_sv2v_reg ,
  \piso.data_r_1825_sv2v_reg ,\piso.data_r_1824_sv2v_reg ,\piso.data_r_1823_sv2v_reg ,
  \piso.data_r_1822_sv2v_reg ,\piso.data_r_1821_sv2v_reg ,\piso.data_r_1820_sv2v_reg ,
  \piso.data_r_1819_sv2v_reg ,\piso.data_r_1818_sv2v_reg ,\piso.data_r_1817_sv2v_reg ,
  \piso.data_r_1816_sv2v_reg ,\piso.data_r_1815_sv2v_reg ,\piso.data_r_1814_sv2v_reg ,
  \piso.data_r_1813_sv2v_reg ,\piso.data_r_1812_sv2v_reg ,\piso.data_r_1811_sv2v_reg ,
  \piso.data_r_1810_sv2v_reg ,\piso.data_r_1809_sv2v_reg ,
  \piso.data_r_1808_sv2v_reg ,\piso.data_r_1807_sv2v_reg ,\piso.data_r_1806_sv2v_reg ,
  \piso.data_r_1805_sv2v_reg ,\piso.data_r_1804_sv2v_reg ,\piso.data_r_1803_sv2v_reg ,
  \piso.data_r_1802_sv2v_reg ,\piso.data_r_1801_sv2v_reg ,\piso.data_r_1800_sv2v_reg ,
  \piso.data_r_1799_sv2v_reg ,\piso.data_r_1798_sv2v_reg ,\piso.data_r_1797_sv2v_reg ,
  \piso.data_r_1796_sv2v_reg ,\piso.data_r_1795_sv2v_reg ,\piso.data_r_1794_sv2v_reg ,
  \piso.data_r_1793_sv2v_reg ,\piso.data_r_1792_sv2v_reg ,\piso.data_r_1791_sv2v_reg ,
  \piso.data_r_1790_sv2v_reg ,\piso.data_r_1789_sv2v_reg ,
  \piso.data_r_1788_sv2v_reg ,\piso.data_r_1787_sv2v_reg ,\piso.data_r_1786_sv2v_reg ,
  \piso.data_r_1785_sv2v_reg ,\piso.data_r_1784_sv2v_reg ,\piso.data_r_1783_sv2v_reg ,
  \piso.data_r_1782_sv2v_reg ,\piso.data_r_1781_sv2v_reg ,\piso.data_r_1780_sv2v_reg ,
  \piso.data_r_1779_sv2v_reg ,\piso.data_r_1778_sv2v_reg ,\piso.data_r_1777_sv2v_reg ,
  \piso.data_r_1776_sv2v_reg ,\piso.data_r_1775_sv2v_reg ,\piso.data_r_1774_sv2v_reg ,
  \piso.data_r_1773_sv2v_reg ,\piso.data_r_1772_sv2v_reg ,\piso.data_r_1771_sv2v_reg ,
  \piso.data_r_1770_sv2v_reg ,\piso.data_r_1769_sv2v_reg ,
  \piso.data_r_1768_sv2v_reg ,\piso.data_r_1767_sv2v_reg ,\piso.data_r_1766_sv2v_reg ,
  \piso.data_r_1765_sv2v_reg ,\piso.data_r_1764_sv2v_reg ,\piso.data_r_1763_sv2v_reg ,
  \piso.data_r_1762_sv2v_reg ,\piso.data_r_1761_sv2v_reg ,\piso.data_r_1760_sv2v_reg ,
  \piso.data_r_1759_sv2v_reg ,\piso.data_r_1758_sv2v_reg ,\piso.data_r_1757_sv2v_reg ,
  \piso.data_r_1756_sv2v_reg ,\piso.data_r_1755_sv2v_reg ,\piso.data_r_1754_sv2v_reg ,
  \piso.data_r_1753_sv2v_reg ,\piso.data_r_1752_sv2v_reg ,\piso.data_r_1751_sv2v_reg ,
  \piso.data_r_1750_sv2v_reg ,\piso.data_r_1749_sv2v_reg ,
  \piso.data_r_1748_sv2v_reg ,\piso.data_r_1747_sv2v_reg ,\piso.data_r_1746_sv2v_reg ,
  \piso.data_r_1745_sv2v_reg ,\piso.data_r_1744_sv2v_reg ,\piso.data_r_1743_sv2v_reg ,
  \piso.data_r_1742_sv2v_reg ,\piso.data_r_1741_sv2v_reg ,\piso.data_r_1740_sv2v_reg ,
  \piso.data_r_1739_sv2v_reg ,\piso.data_r_1738_sv2v_reg ,\piso.data_r_1737_sv2v_reg ,
  \piso.data_r_1736_sv2v_reg ,\piso.data_r_1735_sv2v_reg ,\piso.data_r_1734_sv2v_reg ,
  \piso.data_r_1733_sv2v_reg ,\piso.data_r_1732_sv2v_reg ,\piso.data_r_1731_sv2v_reg ,
  \piso.data_r_1730_sv2v_reg ,\piso.data_r_1729_sv2v_reg ,
  \piso.data_r_1728_sv2v_reg ,\piso.data_r_1727_sv2v_reg ,\piso.data_r_1726_sv2v_reg ,
  \piso.data_r_1725_sv2v_reg ,\piso.data_r_1724_sv2v_reg ,\piso.data_r_1723_sv2v_reg ,
  \piso.data_r_1722_sv2v_reg ,\piso.data_r_1721_sv2v_reg ,\piso.data_r_1720_sv2v_reg ,
  \piso.data_r_1719_sv2v_reg ,\piso.data_r_1718_sv2v_reg ,\piso.data_r_1717_sv2v_reg ,
  \piso.data_r_1716_sv2v_reg ,\piso.data_r_1715_sv2v_reg ,\piso.data_r_1714_sv2v_reg ,
  \piso.data_r_1713_sv2v_reg ,\piso.data_r_1712_sv2v_reg ,\piso.data_r_1711_sv2v_reg ,
  \piso.data_r_1710_sv2v_reg ,\piso.data_r_1709_sv2v_reg ,
  \piso.data_r_1708_sv2v_reg ,\piso.data_r_1707_sv2v_reg ,\piso.data_r_1706_sv2v_reg ,
  \piso.data_r_1705_sv2v_reg ,\piso.data_r_1704_sv2v_reg ,\piso.data_r_1703_sv2v_reg ,
  \piso.data_r_1702_sv2v_reg ,\piso.data_r_1701_sv2v_reg ,\piso.data_r_1700_sv2v_reg ,
  \piso.data_r_1699_sv2v_reg ,\piso.data_r_1698_sv2v_reg ,\piso.data_r_1697_sv2v_reg ,
  \piso.data_r_1696_sv2v_reg ,\piso.data_r_1695_sv2v_reg ,\piso.data_r_1694_sv2v_reg ,
  \piso.data_r_1693_sv2v_reg ,\piso.data_r_1692_sv2v_reg ,\piso.data_r_1691_sv2v_reg ,
  \piso.data_r_1690_sv2v_reg ,\piso.data_r_1689_sv2v_reg ,
  \piso.data_r_1688_sv2v_reg ,\piso.data_r_1687_sv2v_reg ,\piso.data_r_1686_sv2v_reg ,
  \piso.data_r_1685_sv2v_reg ,\piso.data_r_1684_sv2v_reg ,\piso.data_r_1683_sv2v_reg ,
  \piso.data_r_1682_sv2v_reg ,\piso.data_r_1681_sv2v_reg ,\piso.data_r_1680_sv2v_reg ,
  \piso.data_r_1679_sv2v_reg ,\piso.data_r_1678_sv2v_reg ,\piso.data_r_1677_sv2v_reg ,
  \piso.data_r_1676_sv2v_reg ,\piso.data_r_1675_sv2v_reg ,\piso.data_r_1674_sv2v_reg ,
  \piso.data_r_1673_sv2v_reg ,\piso.data_r_1672_sv2v_reg ,\piso.data_r_1671_sv2v_reg ,
  \piso.data_r_1670_sv2v_reg ,\piso.data_r_1669_sv2v_reg ,
  \piso.data_r_1668_sv2v_reg ,\piso.data_r_1667_sv2v_reg ,\piso.data_r_1666_sv2v_reg ,
  \piso.data_r_1665_sv2v_reg ,\piso.data_r_1664_sv2v_reg ,\piso.data_r_1663_sv2v_reg ,
  \piso.data_r_1662_sv2v_reg ,\piso.data_r_1661_sv2v_reg ,\piso.data_r_1660_sv2v_reg ,
  \piso.data_r_1659_sv2v_reg ,\piso.data_r_1658_sv2v_reg ,\piso.data_r_1657_sv2v_reg ,
  \piso.data_r_1656_sv2v_reg ,\piso.data_r_1655_sv2v_reg ,\piso.data_r_1654_sv2v_reg ,
  \piso.data_r_1653_sv2v_reg ,\piso.data_r_1652_sv2v_reg ,\piso.data_r_1651_sv2v_reg ,
  \piso.data_r_1650_sv2v_reg ,\piso.data_r_1649_sv2v_reg ,
  \piso.data_r_1648_sv2v_reg ,\piso.data_r_1647_sv2v_reg ,\piso.data_r_1646_sv2v_reg ,
  \piso.data_r_1645_sv2v_reg ,\piso.data_r_1644_sv2v_reg ,\piso.data_r_1643_sv2v_reg ,
  \piso.data_r_1642_sv2v_reg ,\piso.data_r_1641_sv2v_reg ,\piso.data_r_1640_sv2v_reg ,
  \piso.data_r_1639_sv2v_reg ,\piso.data_r_1638_sv2v_reg ,\piso.data_r_1637_sv2v_reg ,
  \piso.data_r_1636_sv2v_reg ,\piso.data_r_1635_sv2v_reg ,\piso.data_r_1634_sv2v_reg ,
  \piso.data_r_1633_sv2v_reg ,\piso.data_r_1632_sv2v_reg ,\piso.data_r_1631_sv2v_reg ,
  \piso.data_r_1630_sv2v_reg ,\piso.data_r_1629_sv2v_reg ,
  \piso.data_r_1628_sv2v_reg ,\piso.data_r_1627_sv2v_reg ,\piso.data_r_1626_sv2v_reg ,
  \piso.data_r_1625_sv2v_reg ,\piso.data_r_1624_sv2v_reg ,\piso.data_r_1623_sv2v_reg ,
  \piso.data_r_1622_sv2v_reg ,\piso.data_r_1621_sv2v_reg ,\piso.data_r_1620_sv2v_reg ,
  \piso.data_r_1619_sv2v_reg ,\piso.data_r_1618_sv2v_reg ,\piso.data_r_1617_sv2v_reg ,
  \piso.data_r_1616_sv2v_reg ,\piso.data_r_1615_sv2v_reg ,\piso.data_r_1614_sv2v_reg ,
  \piso.data_r_1613_sv2v_reg ,\piso.data_r_1612_sv2v_reg ,\piso.data_r_1611_sv2v_reg ,
  \piso.data_r_1610_sv2v_reg ,\piso.data_r_1609_sv2v_reg ,
  \piso.data_r_1608_sv2v_reg ,\piso.data_r_1607_sv2v_reg ,\piso.data_r_1606_sv2v_reg ,
  \piso.data_r_1605_sv2v_reg ,\piso.data_r_1604_sv2v_reg ,\piso.data_r_1603_sv2v_reg ,
  \piso.data_r_1602_sv2v_reg ,\piso.data_r_1601_sv2v_reg ,\piso.data_r_1600_sv2v_reg ,
  \piso.data_r_1599_sv2v_reg ,\piso.data_r_1598_sv2v_reg ,\piso.data_r_1597_sv2v_reg ,
  \piso.data_r_1596_sv2v_reg ,\piso.data_r_1595_sv2v_reg ,\piso.data_r_1594_sv2v_reg ,
  \piso.data_r_1593_sv2v_reg ,\piso.data_r_1592_sv2v_reg ,\piso.data_r_1591_sv2v_reg ,
  \piso.data_r_1590_sv2v_reg ,\piso.data_r_1589_sv2v_reg ,
  \piso.data_r_1588_sv2v_reg ,\piso.data_r_1587_sv2v_reg ,\piso.data_r_1586_sv2v_reg ,
  \piso.data_r_1585_sv2v_reg ,\piso.data_r_1584_sv2v_reg ,\piso.data_r_1583_sv2v_reg ,
  \piso.data_r_1582_sv2v_reg ,\piso.data_r_1581_sv2v_reg ,\piso.data_r_1580_sv2v_reg ,
  \piso.data_r_1579_sv2v_reg ,\piso.data_r_1578_sv2v_reg ,\piso.data_r_1577_sv2v_reg ,
  \piso.data_r_1576_sv2v_reg ,\piso.data_r_1575_sv2v_reg ,\piso.data_r_1574_sv2v_reg ,
  \piso.data_r_1573_sv2v_reg ,\piso.data_r_1572_sv2v_reg ,\piso.data_r_1571_sv2v_reg ,
  \piso.data_r_1570_sv2v_reg ,\piso.data_r_1569_sv2v_reg ,
  \piso.data_r_1568_sv2v_reg ,\piso.data_r_1567_sv2v_reg ,\piso.data_r_1566_sv2v_reg ,
  \piso.data_r_1565_sv2v_reg ,\piso.data_r_1564_sv2v_reg ,\piso.data_r_1563_sv2v_reg ,
  \piso.data_r_1562_sv2v_reg ,\piso.data_r_1561_sv2v_reg ,\piso.data_r_1560_sv2v_reg ,
  \piso.data_r_1559_sv2v_reg ,\piso.data_r_1558_sv2v_reg ,\piso.data_r_1557_sv2v_reg ,
  \piso.data_r_1556_sv2v_reg ,\piso.data_r_1555_sv2v_reg ,\piso.data_r_1554_sv2v_reg ,
  \piso.data_r_1553_sv2v_reg ,\piso.data_r_1552_sv2v_reg ,\piso.data_r_1551_sv2v_reg ,
  \piso.data_r_1550_sv2v_reg ,\piso.data_r_1549_sv2v_reg ,
  \piso.data_r_1548_sv2v_reg ,\piso.data_r_1547_sv2v_reg ,\piso.data_r_1546_sv2v_reg ,
  \piso.data_r_1545_sv2v_reg ,\piso.data_r_1544_sv2v_reg ,\piso.data_r_1543_sv2v_reg ,
  \piso.data_r_1542_sv2v_reg ,\piso.data_r_1541_sv2v_reg ,\piso.data_r_1540_sv2v_reg ,
  \piso.data_r_1539_sv2v_reg ,\piso.data_r_1538_sv2v_reg ,\piso.data_r_1537_sv2v_reg ,
  \piso.data_r_1536_sv2v_reg ,\piso.data_r_1535_sv2v_reg ,\piso.data_r_1534_sv2v_reg ,
  \piso.data_r_1533_sv2v_reg ,\piso.data_r_1532_sv2v_reg ,\piso.data_r_1531_sv2v_reg ,
  \piso.data_r_1530_sv2v_reg ,\piso.data_r_1529_sv2v_reg ,
  \piso.data_r_1528_sv2v_reg ,\piso.data_r_1527_sv2v_reg ,\piso.data_r_1526_sv2v_reg ,
  \piso.data_r_1525_sv2v_reg ,\piso.data_r_1524_sv2v_reg ,\piso.data_r_1523_sv2v_reg ,
  \piso.data_r_1522_sv2v_reg ,\piso.data_r_1521_sv2v_reg ,\piso.data_r_1520_sv2v_reg ,
  \piso.data_r_1519_sv2v_reg ,\piso.data_r_1518_sv2v_reg ,\piso.data_r_1517_sv2v_reg ,
  \piso.data_r_1516_sv2v_reg ,\piso.data_r_1515_sv2v_reg ,\piso.data_r_1514_sv2v_reg ,
  \piso.data_r_1513_sv2v_reg ,\piso.data_r_1512_sv2v_reg ,\piso.data_r_1511_sv2v_reg ,
  \piso.data_r_1510_sv2v_reg ,\piso.data_r_1509_sv2v_reg ,
  \piso.data_r_1508_sv2v_reg ,\piso.data_r_1507_sv2v_reg ,\piso.data_r_1506_sv2v_reg ,
  \piso.data_r_1505_sv2v_reg ,\piso.data_r_1504_sv2v_reg ,\piso.data_r_1503_sv2v_reg ,
  \piso.data_r_1502_sv2v_reg ,\piso.data_r_1501_sv2v_reg ,\piso.data_r_1500_sv2v_reg ,
  \piso.data_r_1499_sv2v_reg ,\piso.data_r_1498_sv2v_reg ,\piso.data_r_1497_sv2v_reg ,
  \piso.data_r_1496_sv2v_reg ,\piso.data_r_1495_sv2v_reg ,\piso.data_r_1494_sv2v_reg ,
  \piso.data_r_1493_sv2v_reg ,\piso.data_r_1492_sv2v_reg ,\piso.data_r_1491_sv2v_reg ,
  \piso.data_r_1490_sv2v_reg ,\piso.data_r_1489_sv2v_reg ,
  \piso.data_r_1488_sv2v_reg ,\piso.data_r_1487_sv2v_reg ,\piso.data_r_1486_sv2v_reg ,
  \piso.data_r_1485_sv2v_reg ,\piso.data_r_1484_sv2v_reg ,\piso.data_r_1483_sv2v_reg ,
  \piso.data_r_1482_sv2v_reg ,\piso.data_r_1481_sv2v_reg ,\piso.data_r_1480_sv2v_reg ,
  \piso.data_r_1479_sv2v_reg ,\piso.data_r_1478_sv2v_reg ,\piso.data_r_1477_sv2v_reg ,
  \piso.data_r_1476_sv2v_reg ,\piso.data_r_1475_sv2v_reg ,\piso.data_r_1474_sv2v_reg ,
  \piso.data_r_1473_sv2v_reg ,\piso.data_r_1472_sv2v_reg ,\piso.data_r_1471_sv2v_reg ,
  \piso.data_r_1470_sv2v_reg ,\piso.data_r_1469_sv2v_reg ,
  \piso.data_r_1468_sv2v_reg ,\piso.data_r_1467_sv2v_reg ,\piso.data_r_1466_sv2v_reg ,
  \piso.data_r_1465_sv2v_reg ,\piso.data_r_1464_sv2v_reg ,\piso.data_r_1463_sv2v_reg ,
  \piso.data_r_1462_sv2v_reg ,\piso.data_r_1461_sv2v_reg ,\piso.data_r_1460_sv2v_reg ,
  \piso.data_r_1459_sv2v_reg ,\piso.data_r_1458_sv2v_reg ,\piso.data_r_1457_sv2v_reg ,
  \piso.data_r_1456_sv2v_reg ,\piso.data_r_1455_sv2v_reg ,\piso.data_r_1454_sv2v_reg ,
  \piso.data_r_1453_sv2v_reg ,\piso.data_r_1452_sv2v_reg ,\piso.data_r_1451_sv2v_reg ,
  \piso.data_r_1450_sv2v_reg ,\piso.data_r_1449_sv2v_reg ,
  \piso.data_r_1448_sv2v_reg ,\piso.data_r_1447_sv2v_reg ,\piso.data_r_1446_sv2v_reg ,
  \piso.data_r_1445_sv2v_reg ,\piso.data_r_1444_sv2v_reg ,\piso.data_r_1443_sv2v_reg ,
  \piso.data_r_1442_sv2v_reg ,\piso.data_r_1441_sv2v_reg ,\piso.data_r_1440_sv2v_reg ,
  \piso.data_r_1439_sv2v_reg ,\piso.data_r_1438_sv2v_reg ,\piso.data_r_1437_sv2v_reg ,
  \piso.data_r_1436_sv2v_reg ,\piso.data_r_1435_sv2v_reg ,\piso.data_r_1434_sv2v_reg ,
  \piso.data_r_1433_sv2v_reg ,\piso.data_r_1432_sv2v_reg ,\piso.data_r_1431_sv2v_reg ,
  \piso.data_r_1430_sv2v_reg ,\piso.data_r_1429_sv2v_reg ,
  \piso.data_r_1428_sv2v_reg ,\piso.data_r_1427_sv2v_reg ,\piso.data_r_1426_sv2v_reg ,
  \piso.data_r_1425_sv2v_reg ,\piso.data_r_1424_sv2v_reg ,\piso.data_r_1423_sv2v_reg ,
  \piso.data_r_1422_sv2v_reg ,\piso.data_r_1421_sv2v_reg ,\piso.data_r_1420_sv2v_reg ,
  \piso.data_r_1419_sv2v_reg ,\piso.data_r_1418_sv2v_reg ,\piso.data_r_1417_sv2v_reg ,
  \piso.data_r_1416_sv2v_reg ,\piso.data_r_1415_sv2v_reg ,\piso.data_r_1414_sv2v_reg ,
  \piso.data_r_1413_sv2v_reg ,\piso.data_r_1412_sv2v_reg ,\piso.data_r_1411_sv2v_reg ,
  \piso.data_r_1410_sv2v_reg ,\piso.data_r_1409_sv2v_reg ,
  \piso.data_r_1408_sv2v_reg ,\piso.data_r_1407_sv2v_reg ,\piso.data_r_1406_sv2v_reg ,
  \piso.data_r_1405_sv2v_reg ,\piso.data_r_1404_sv2v_reg ,\piso.data_r_1403_sv2v_reg ,
  \piso.data_r_1402_sv2v_reg ,\piso.data_r_1401_sv2v_reg ,\piso.data_r_1400_sv2v_reg ,
  \piso.data_r_1399_sv2v_reg ,\piso.data_r_1398_sv2v_reg ,\piso.data_r_1397_sv2v_reg ,
  \piso.data_r_1396_sv2v_reg ,\piso.data_r_1395_sv2v_reg ,\piso.data_r_1394_sv2v_reg ,
  \piso.data_r_1393_sv2v_reg ,\piso.data_r_1392_sv2v_reg ,\piso.data_r_1391_sv2v_reg ,
  \piso.data_r_1390_sv2v_reg ,\piso.data_r_1389_sv2v_reg ,
  \piso.data_r_1388_sv2v_reg ,\piso.data_r_1387_sv2v_reg ,\piso.data_r_1386_sv2v_reg ,
  \piso.data_r_1385_sv2v_reg ,\piso.data_r_1384_sv2v_reg ,\piso.data_r_1383_sv2v_reg ,
  \piso.data_r_1382_sv2v_reg ,\piso.data_r_1381_sv2v_reg ,\piso.data_r_1380_sv2v_reg ,
  \piso.data_r_1379_sv2v_reg ,\piso.data_r_1378_sv2v_reg ,\piso.data_r_1377_sv2v_reg ,
  \piso.data_r_1376_sv2v_reg ,\piso.data_r_1375_sv2v_reg ,\piso.data_r_1374_sv2v_reg ,
  \piso.data_r_1373_sv2v_reg ,\piso.data_r_1372_sv2v_reg ,\piso.data_r_1371_sv2v_reg ,
  \piso.data_r_1370_sv2v_reg ,\piso.data_r_1369_sv2v_reg ,
  \piso.data_r_1368_sv2v_reg ,\piso.data_r_1367_sv2v_reg ,\piso.data_r_1366_sv2v_reg ,
  \piso.data_r_1365_sv2v_reg ,\piso.data_r_1364_sv2v_reg ,\piso.data_r_1363_sv2v_reg ,
  \piso.data_r_1362_sv2v_reg ,\piso.data_r_1361_sv2v_reg ,\piso.data_r_1360_sv2v_reg ,
  \piso.data_r_1359_sv2v_reg ,\piso.data_r_1358_sv2v_reg ,\piso.data_r_1357_sv2v_reg ,
  \piso.data_r_1356_sv2v_reg ,\piso.data_r_1355_sv2v_reg ,\piso.data_r_1354_sv2v_reg ,
  \piso.data_r_1353_sv2v_reg ,\piso.data_r_1352_sv2v_reg ,\piso.data_r_1351_sv2v_reg ,
  \piso.data_r_1350_sv2v_reg ,\piso.data_r_1349_sv2v_reg ,
  \piso.data_r_1348_sv2v_reg ,\piso.data_r_1347_sv2v_reg ,\piso.data_r_1346_sv2v_reg ,
  \piso.data_r_1345_sv2v_reg ,\piso.data_r_1344_sv2v_reg ,\piso.data_r_1343_sv2v_reg ,
  \piso.data_r_1342_sv2v_reg ,\piso.data_r_1341_sv2v_reg ,\piso.data_r_1340_sv2v_reg ,
  \piso.data_r_1339_sv2v_reg ,\piso.data_r_1338_sv2v_reg ,\piso.data_r_1337_sv2v_reg ,
  \piso.data_r_1336_sv2v_reg ,\piso.data_r_1335_sv2v_reg ,\piso.data_r_1334_sv2v_reg ,
  \piso.data_r_1333_sv2v_reg ,\piso.data_r_1332_sv2v_reg ,\piso.data_r_1331_sv2v_reg ,
  \piso.data_r_1330_sv2v_reg ,\piso.data_r_1329_sv2v_reg ,
  \piso.data_r_1328_sv2v_reg ,\piso.data_r_1327_sv2v_reg ,\piso.data_r_1326_sv2v_reg ,
  \piso.data_r_1325_sv2v_reg ,\piso.data_r_1324_sv2v_reg ,\piso.data_r_1323_sv2v_reg ,
  \piso.data_r_1322_sv2v_reg ,\piso.data_r_1321_sv2v_reg ,\piso.data_r_1320_sv2v_reg ,
  \piso.data_r_1319_sv2v_reg ,\piso.data_r_1318_sv2v_reg ,\piso.data_r_1317_sv2v_reg ,
  \piso.data_r_1316_sv2v_reg ,\piso.data_r_1315_sv2v_reg ,\piso.data_r_1314_sv2v_reg ,
  \piso.data_r_1313_sv2v_reg ,\piso.data_r_1312_sv2v_reg ,\piso.data_r_1311_sv2v_reg ,
  \piso.data_r_1310_sv2v_reg ,\piso.data_r_1309_sv2v_reg ,
  \piso.data_r_1308_sv2v_reg ,\piso.data_r_1307_sv2v_reg ,\piso.data_r_1306_sv2v_reg ,
  \piso.data_r_1305_sv2v_reg ,\piso.data_r_1304_sv2v_reg ,\piso.data_r_1303_sv2v_reg ,
  \piso.data_r_1302_sv2v_reg ,\piso.data_r_1301_sv2v_reg ,\piso.data_r_1300_sv2v_reg ,
  \piso.data_r_1299_sv2v_reg ,\piso.data_r_1298_sv2v_reg ,\piso.data_r_1297_sv2v_reg ,
  \piso.data_r_1296_sv2v_reg ,\piso.data_r_1295_sv2v_reg ,\piso.data_r_1294_sv2v_reg ,
  \piso.data_r_1293_sv2v_reg ,\piso.data_r_1292_sv2v_reg ,\piso.data_r_1291_sv2v_reg ,
  \piso.data_r_1290_sv2v_reg ,\piso.data_r_1289_sv2v_reg ,
  \piso.data_r_1288_sv2v_reg ,\piso.data_r_1287_sv2v_reg ,\piso.data_r_1286_sv2v_reg ,
  \piso.data_r_1285_sv2v_reg ,\piso.data_r_1284_sv2v_reg ,\piso.data_r_1283_sv2v_reg ,
  \piso.data_r_1282_sv2v_reg ,\piso.data_r_1281_sv2v_reg ,\piso.data_r_1280_sv2v_reg ,
  \piso.data_r_1279_sv2v_reg ,\piso.data_r_1278_sv2v_reg ,\piso.data_r_1277_sv2v_reg ,
  \piso.data_r_1276_sv2v_reg ,\piso.data_r_1275_sv2v_reg ,\piso.data_r_1274_sv2v_reg ,
  \piso.data_r_1273_sv2v_reg ,\piso.data_r_1272_sv2v_reg ,\piso.data_r_1271_sv2v_reg ,
  \piso.data_r_1270_sv2v_reg ,\piso.data_r_1269_sv2v_reg ,
  \piso.data_r_1268_sv2v_reg ,\piso.data_r_1267_sv2v_reg ,\piso.data_r_1266_sv2v_reg ,
  \piso.data_r_1265_sv2v_reg ,\piso.data_r_1264_sv2v_reg ,\piso.data_r_1263_sv2v_reg ,
  \piso.data_r_1262_sv2v_reg ,\piso.data_r_1261_sv2v_reg ,\piso.data_r_1260_sv2v_reg ,
  \piso.data_r_1259_sv2v_reg ,\piso.data_r_1258_sv2v_reg ,\piso.data_r_1257_sv2v_reg ,
  \piso.data_r_1256_sv2v_reg ,\piso.data_r_1255_sv2v_reg ,\piso.data_r_1254_sv2v_reg ,
  \piso.data_r_1253_sv2v_reg ,\piso.data_r_1252_sv2v_reg ,\piso.data_r_1251_sv2v_reg ,
  \piso.data_r_1250_sv2v_reg ,\piso.data_r_1249_sv2v_reg ,
  \piso.data_r_1248_sv2v_reg ,\piso.data_r_1247_sv2v_reg ,\piso.data_r_1246_sv2v_reg ,
  \piso.data_r_1245_sv2v_reg ,\piso.data_r_1244_sv2v_reg ,\piso.data_r_1243_sv2v_reg ,
  \piso.data_r_1242_sv2v_reg ,\piso.data_r_1241_sv2v_reg ,\piso.data_r_1240_sv2v_reg ,
  \piso.data_r_1239_sv2v_reg ,\piso.data_r_1238_sv2v_reg ,\piso.data_r_1237_sv2v_reg ,
  \piso.data_r_1236_sv2v_reg ,\piso.data_r_1235_sv2v_reg ,\piso.data_r_1234_sv2v_reg ,
  \piso.data_r_1233_sv2v_reg ,\piso.data_r_1232_sv2v_reg ,\piso.data_r_1231_sv2v_reg ,
  \piso.data_r_1230_sv2v_reg ,\piso.data_r_1229_sv2v_reg ,
  \piso.data_r_1228_sv2v_reg ,\piso.data_r_1227_sv2v_reg ,\piso.data_r_1226_sv2v_reg ,
  \piso.data_r_1225_sv2v_reg ,\piso.data_r_1224_sv2v_reg ,\piso.data_r_1223_sv2v_reg ,
  \piso.data_r_1222_sv2v_reg ,\piso.data_r_1221_sv2v_reg ,\piso.data_r_1220_sv2v_reg ,
  \piso.data_r_1219_sv2v_reg ,\piso.data_r_1218_sv2v_reg ,\piso.data_r_1217_sv2v_reg ,
  \piso.data_r_1216_sv2v_reg ,\piso.data_r_1215_sv2v_reg ,\piso.data_r_1214_sv2v_reg ,
  \piso.data_r_1213_sv2v_reg ,\piso.data_r_1212_sv2v_reg ,\piso.data_r_1211_sv2v_reg ,
  \piso.data_r_1210_sv2v_reg ,\piso.data_r_1209_sv2v_reg ,
  \piso.data_r_1208_sv2v_reg ,\piso.data_r_1207_sv2v_reg ,\piso.data_r_1206_sv2v_reg ,
  \piso.data_r_1205_sv2v_reg ,\piso.data_r_1204_sv2v_reg ,\piso.data_r_1203_sv2v_reg ,
  \piso.data_r_1202_sv2v_reg ,\piso.data_r_1201_sv2v_reg ,\piso.data_r_1200_sv2v_reg ,
  \piso.data_r_1199_sv2v_reg ,\piso.data_r_1198_sv2v_reg ,\piso.data_r_1197_sv2v_reg ,
  \piso.data_r_1196_sv2v_reg ,\piso.data_r_1195_sv2v_reg ,\piso.data_r_1194_sv2v_reg ,
  \piso.data_r_1193_sv2v_reg ,\piso.data_r_1192_sv2v_reg ,\piso.data_r_1191_sv2v_reg ,
  \piso.data_r_1190_sv2v_reg ,\piso.data_r_1189_sv2v_reg ,
  \piso.data_r_1188_sv2v_reg ,\piso.data_r_1187_sv2v_reg ,\piso.data_r_1186_sv2v_reg ,
  \piso.data_r_1185_sv2v_reg ,\piso.data_r_1184_sv2v_reg ,\piso.data_r_1183_sv2v_reg ,
  \piso.data_r_1182_sv2v_reg ,\piso.data_r_1181_sv2v_reg ,\piso.data_r_1180_sv2v_reg ,
  \piso.data_r_1179_sv2v_reg ,\piso.data_r_1178_sv2v_reg ,\piso.data_r_1177_sv2v_reg ,
  \piso.data_r_1176_sv2v_reg ,\piso.data_r_1175_sv2v_reg ,\piso.data_r_1174_sv2v_reg ,
  \piso.data_r_1173_sv2v_reg ,\piso.data_r_1172_sv2v_reg ,\piso.data_r_1171_sv2v_reg ,
  \piso.data_r_1170_sv2v_reg ,\piso.data_r_1169_sv2v_reg ,
  \piso.data_r_1168_sv2v_reg ,\piso.data_r_1167_sv2v_reg ,\piso.data_r_1166_sv2v_reg ,
  \piso.data_r_1165_sv2v_reg ,\piso.data_r_1164_sv2v_reg ,\piso.data_r_1163_sv2v_reg ,
  \piso.data_r_1162_sv2v_reg ,\piso.data_r_1161_sv2v_reg ,\piso.data_r_1160_sv2v_reg ,
  \piso.data_r_1159_sv2v_reg ,\piso.data_r_1158_sv2v_reg ,\piso.data_r_1157_sv2v_reg ,
  \piso.data_r_1156_sv2v_reg ,\piso.data_r_1155_sv2v_reg ,\piso.data_r_1154_sv2v_reg ,
  \piso.data_r_1153_sv2v_reg ,\piso.data_r_1152_sv2v_reg ,\piso.data_r_1151_sv2v_reg ,
  \piso.data_r_1150_sv2v_reg ,\piso.data_r_1149_sv2v_reg ,
  \piso.data_r_1148_sv2v_reg ,\piso.data_r_1147_sv2v_reg ,\piso.data_r_1146_sv2v_reg ,
  \piso.data_r_1145_sv2v_reg ,\piso.data_r_1144_sv2v_reg ,\piso.data_r_1143_sv2v_reg ,
  \piso.data_r_1142_sv2v_reg ,\piso.data_r_1141_sv2v_reg ,\piso.data_r_1140_sv2v_reg ,
  \piso.data_r_1139_sv2v_reg ,\piso.data_r_1138_sv2v_reg ,\piso.data_r_1137_sv2v_reg ,
  \piso.data_r_1136_sv2v_reg ,\piso.data_r_1135_sv2v_reg ,\piso.data_r_1134_sv2v_reg ,
  \piso.data_r_1133_sv2v_reg ,\piso.data_r_1132_sv2v_reg ,\piso.data_r_1131_sv2v_reg ,
  \piso.data_r_1130_sv2v_reg ,\piso.data_r_1129_sv2v_reg ,
  \piso.data_r_1128_sv2v_reg ,\piso.data_r_1127_sv2v_reg ,\piso.data_r_1126_sv2v_reg ,
  \piso.data_r_1125_sv2v_reg ,\piso.data_r_1124_sv2v_reg ,\piso.data_r_1123_sv2v_reg ,
  \piso.data_r_1122_sv2v_reg ,\piso.data_r_1121_sv2v_reg ,\piso.data_r_1120_sv2v_reg ,
  \piso.data_r_1119_sv2v_reg ,\piso.data_r_1118_sv2v_reg ,\piso.data_r_1117_sv2v_reg ,
  \piso.data_r_1116_sv2v_reg ,\piso.data_r_1115_sv2v_reg ,\piso.data_r_1114_sv2v_reg ,
  \piso.data_r_1113_sv2v_reg ,\piso.data_r_1112_sv2v_reg ,\piso.data_r_1111_sv2v_reg ,
  \piso.data_r_1110_sv2v_reg ,\piso.data_r_1109_sv2v_reg ,
  \piso.data_r_1108_sv2v_reg ,\piso.data_r_1107_sv2v_reg ,\piso.data_r_1106_sv2v_reg ,
  \piso.data_r_1105_sv2v_reg ,\piso.data_r_1104_sv2v_reg ,\piso.data_r_1103_sv2v_reg ,
  \piso.data_r_1102_sv2v_reg ,\piso.data_r_1101_sv2v_reg ,\piso.data_r_1100_sv2v_reg ,
  \piso.data_r_1099_sv2v_reg ,\piso.data_r_1098_sv2v_reg ,\piso.data_r_1097_sv2v_reg ,
  \piso.data_r_1096_sv2v_reg ,\piso.data_r_1095_sv2v_reg ,\piso.data_r_1094_sv2v_reg ,
  \piso.data_r_1093_sv2v_reg ,\piso.data_r_1092_sv2v_reg ,\piso.data_r_1091_sv2v_reg ,
  \piso.data_r_1090_sv2v_reg ,\piso.data_r_1089_sv2v_reg ,
  \piso.data_r_1088_sv2v_reg ,\piso.data_r_1087_sv2v_reg ,\piso.data_r_1086_sv2v_reg ,
  \piso.data_r_1085_sv2v_reg ,\piso.data_r_1084_sv2v_reg ,\piso.data_r_1083_sv2v_reg ,
  \piso.data_r_1082_sv2v_reg ,\piso.data_r_1081_sv2v_reg ,\piso.data_r_1080_sv2v_reg ,
  \piso.data_r_1079_sv2v_reg ,\piso.data_r_1078_sv2v_reg ,\piso.data_r_1077_sv2v_reg ,
  \piso.data_r_1076_sv2v_reg ,\piso.data_r_1075_sv2v_reg ,\piso.data_r_1074_sv2v_reg ,
  \piso.data_r_1073_sv2v_reg ,\piso.data_r_1072_sv2v_reg ,\piso.data_r_1071_sv2v_reg ,
  \piso.data_r_1070_sv2v_reg ,\piso.data_r_1069_sv2v_reg ,
  \piso.data_r_1068_sv2v_reg ,\piso.data_r_1067_sv2v_reg ,\piso.data_r_1066_sv2v_reg ,
  \piso.data_r_1065_sv2v_reg ,\piso.data_r_1064_sv2v_reg ,\piso.data_r_1063_sv2v_reg ,
  \piso.data_r_1062_sv2v_reg ,\piso.data_r_1061_sv2v_reg ,\piso.data_r_1060_sv2v_reg ,
  \piso.data_r_1059_sv2v_reg ,\piso.data_r_1058_sv2v_reg ,\piso.data_r_1057_sv2v_reg ,
  \piso.data_r_1056_sv2v_reg ,\piso.data_r_1055_sv2v_reg ,\piso.data_r_1054_sv2v_reg ,
  \piso.data_r_1053_sv2v_reg ,\piso.data_r_1052_sv2v_reg ,\piso.data_r_1051_sv2v_reg ,
  \piso.data_r_1050_sv2v_reg ,\piso.data_r_1049_sv2v_reg ,
  \piso.data_r_1048_sv2v_reg ,\piso.data_r_1047_sv2v_reg ,\piso.data_r_1046_sv2v_reg ,
  \piso.data_r_1045_sv2v_reg ,\piso.data_r_1044_sv2v_reg ,\piso.data_r_1043_sv2v_reg ,
  \piso.data_r_1042_sv2v_reg ,\piso.data_r_1041_sv2v_reg ,\piso.data_r_1040_sv2v_reg ,
  \piso.data_r_1039_sv2v_reg ,\piso.data_r_1038_sv2v_reg ,\piso.data_r_1037_sv2v_reg ,
  \piso.data_r_1036_sv2v_reg ,\piso.data_r_1035_sv2v_reg ,\piso.data_r_1034_sv2v_reg ,
  \piso.data_r_1033_sv2v_reg ,\piso.data_r_1032_sv2v_reg ,\piso.data_r_1031_sv2v_reg ,
  \piso.data_r_1030_sv2v_reg ,\piso.data_r_1029_sv2v_reg ,
  \piso.data_r_1028_sv2v_reg ,\piso.data_r_1027_sv2v_reg ,\piso.data_r_1026_sv2v_reg ,
  \piso.data_r_1025_sv2v_reg ,\piso.data_r_1024_sv2v_reg ,\piso.data_r_1023_sv2v_reg ,
  \piso.data_r_1022_sv2v_reg ,\piso.data_r_1021_sv2v_reg ,\piso.data_r_1020_sv2v_reg ,
  \piso.data_r_1019_sv2v_reg ,\piso.data_r_1018_sv2v_reg ,\piso.data_r_1017_sv2v_reg ,
  \piso.data_r_1016_sv2v_reg ,\piso.data_r_1015_sv2v_reg ,\piso.data_r_1014_sv2v_reg ,
  \piso.data_r_1013_sv2v_reg ,\piso.data_r_1012_sv2v_reg ,\piso.data_r_1011_sv2v_reg ,
  \piso.data_r_1010_sv2v_reg ,\piso.data_r_1009_sv2v_reg ,
  \piso.data_r_1008_sv2v_reg ,\piso.data_r_1007_sv2v_reg ,\piso.data_r_1006_sv2v_reg ,
  \piso.data_r_1005_sv2v_reg ,\piso.data_r_1004_sv2v_reg ,\piso.data_r_1003_sv2v_reg ,
  \piso.data_r_1002_sv2v_reg ,\piso.data_r_1001_sv2v_reg ,\piso.data_r_1000_sv2v_reg ,
  \piso.data_r_999_sv2v_reg ,\piso.data_r_998_sv2v_reg ,\piso.data_r_997_sv2v_reg ,
  \piso.data_r_996_sv2v_reg ,\piso.data_r_995_sv2v_reg ,\piso.data_r_994_sv2v_reg ,
  \piso.data_r_993_sv2v_reg ,\piso.data_r_992_sv2v_reg ,\piso.data_r_991_sv2v_reg ,
  \piso.data_r_990_sv2v_reg ,\piso.data_r_989_sv2v_reg ,\piso.data_r_988_sv2v_reg ,
  \piso.data_r_987_sv2v_reg ,\piso.data_r_986_sv2v_reg ,\piso.data_r_985_sv2v_reg ,
  \piso.data_r_984_sv2v_reg ,\piso.data_r_983_sv2v_reg ,\piso.data_r_982_sv2v_reg ,
  \piso.data_r_981_sv2v_reg ,\piso.data_r_980_sv2v_reg ,\piso.data_r_979_sv2v_reg ,
  \piso.data_r_978_sv2v_reg ,\piso.data_r_977_sv2v_reg ,\piso.data_r_976_sv2v_reg ,
  \piso.data_r_975_sv2v_reg ,\piso.data_r_974_sv2v_reg ,\piso.data_r_973_sv2v_reg ,
  \piso.data_r_972_sv2v_reg ,\piso.data_r_971_sv2v_reg ,\piso.data_r_970_sv2v_reg ,
  \piso.data_r_969_sv2v_reg ,\piso.data_r_968_sv2v_reg ,\piso.data_r_967_sv2v_reg ,
  \piso.data_r_966_sv2v_reg ,\piso.data_r_965_sv2v_reg ,\piso.data_r_964_sv2v_reg ,
  \piso.data_r_963_sv2v_reg ,\piso.data_r_962_sv2v_reg ,\piso.data_r_961_sv2v_reg ,
  \piso.data_r_960_sv2v_reg ,\piso.data_r_959_sv2v_reg ,\piso.data_r_958_sv2v_reg ,
  \piso.data_r_957_sv2v_reg ,\piso.data_r_956_sv2v_reg ,\piso.data_r_955_sv2v_reg ,
  \piso.data_r_954_sv2v_reg ,\piso.data_r_953_sv2v_reg ,
  \piso.data_r_952_sv2v_reg ,\piso.data_r_951_sv2v_reg ,\piso.data_r_950_sv2v_reg ,
  \piso.data_r_949_sv2v_reg ,\piso.data_r_948_sv2v_reg ,\piso.data_r_947_sv2v_reg ,
  \piso.data_r_946_sv2v_reg ,\piso.data_r_945_sv2v_reg ,\piso.data_r_944_sv2v_reg ,
  \piso.data_r_943_sv2v_reg ,\piso.data_r_942_sv2v_reg ,\piso.data_r_941_sv2v_reg ,
  \piso.data_r_940_sv2v_reg ,\piso.data_r_939_sv2v_reg ,\piso.data_r_938_sv2v_reg ,
  \piso.data_r_937_sv2v_reg ,\piso.data_r_936_sv2v_reg ,\piso.data_r_935_sv2v_reg ,
  \piso.data_r_934_sv2v_reg ,\piso.data_r_933_sv2v_reg ,\piso.data_r_932_sv2v_reg ,
  \piso.data_r_931_sv2v_reg ,\piso.data_r_930_sv2v_reg ,\piso.data_r_929_sv2v_reg ,
  \piso.data_r_928_sv2v_reg ,\piso.data_r_927_sv2v_reg ,\piso.data_r_926_sv2v_reg ,
  \piso.data_r_925_sv2v_reg ,\piso.data_r_924_sv2v_reg ,\piso.data_r_923_sv2v_reg ,
  \piso.data_r_922_sv2v_reg ,\piso.data_r_921_sv2v_reg ,\piso.data_r_920_sv2v_reg ,
  \piso.data_r_919_sv2v_reg ,\piso.data_r_918_sv2v_reg ,\piso.data_r_917_sv2v_reg ,
  \piso.data_r_916_sv2v_reg ,\piso.data_r_915_sv2v_reg ,\piso.data_r_914_sv2v_reg ,
  \piso.data_r_913_sv2v_reg ,\piso.data_r_912_sv2v_reg ,\piso.data_r_911_sv2v_reg ,
  \piso.data_r_910_sv2v_reg ,\piso.data_r_909_sv2v_reg ,\piso.data_r_908_sv2v_reg ,
  \piso.data_r_907_sv2v_reg ,\piso.data_r_906_sv2v_reg ,\piso.data_r_905_sv2v_reg ,
  \piso.data_r_904_sv2v_reg ,\piso.data_r_903_sv2v_reg ,\piso.data_r_902_sv2v_reg ,
  \piso.data_r_901_sv2v_reg ,\piso.data_r_900_sv2v_reg ,\piso.data_r_899_sv2v_reg ,
  \piso.data_r_898_sv2v_reg ,\piso.data_r_897_sv2v_reg ,\piso.data_r_896_sv2v_reg ,
  \piso.data_r_895_sv2v_reg ,\piso.data_r_894_sv2v_reg ,\piso.data_r_893_sv2v_reg ,
  \piso.data_r_892_sv2v_reg ,\piso.data_r_891_sv2v_reg ,\piso.data_r_890_sv2v_reg ,
  \piso.data_r_889_sv2v_reg ,\piso.data_r_888_sv2v_reg ,\piso.data_r_887_sv2v_reg ,
  \piso.data_r_886_sv2v_reg ,\piso.data_r_885_sv2v_reg ,\piso.data_r_884_sv2v_reg ,
  \piso.data_r_883_sv2v_reg ,\piso.data_r_882_sv2v_reg ,\piso.data_r_881_sv2v_reg ,
  \piso.data_r_880_sv2v_reg ,\piso.data_r_879_sv2v_reg ,\piso.data_r_878_sv2v_reg ,
  \piso.data_r_877_sv2v_reg ,\piso.data_r_876_sv2v_reg ,\piso.data_r_875_sv2v_reg ,
  \piso.data_r_874_sv2v_reg ,\piso.data_r_873_sv2v_reg ,
  \piso.data_r_872_sv2v_reg ,\piso.data_r_871_sv2v_reg ,\piso.data_r_870_sv2v_reg ,
  \piso.data_r_869_sv2v_reg ,\piso.data_r_868_sv2v_reg ,\piso.data_r_867_sv2v_reg ,
  \piso.data_r_866_sv2v_reg ,\piso.data_r_865_sv2v_reg ,\piso.data_r_864_sv2v_reg ,
  \piso.data_r_863_sv2v_reg ,\piso.data_r_862_sv2v_reg ,\piso.data_r_861_sv2v_reg ,
  \piso.data_r_860_sv2v_reg ,\piso.data_r_859_sv2v_reg ,\piso.data_r_858_sv2v_reg ,
  \piso.data_r_857_sv2v_reg ,\piso.data_r_856_sv2v_reg ,\piso.data_r_855_sv2v_reg ,
  \piso.data_r_854_sv2v_reg ,\piso.data_r_853_sv2v_reg ,\piso.data_r_852_sv2v_reg ,
  \piso.data_r_851_sv2v_reg ,\piso.data_r_850_sv2v_reg ,\piso.data_r_849_sv2v_reg ,
  \piso.data_r_848_sv2v_reg ,\piso.data_r_847_sv2v_reg ,\piso.data_r_846_sv2v_reg ,
  \piso.data_r_845_sv2v_reg ,\piso.data_r_844_sv2v_reg ,\piso.data_r_843_sv2v_reg ,
  \piso.data_r_842_sv2v_reg ,\piso.data_r_841_sv2v_reg ,\piso.data_r_840_sv2v_reg ,
  \piso.data_r_839_sv2v_reg ,\piso.data_r_838_sv2v_reg ,\piso.data_r_837_sv2v_reg ,
  \piso.data_r_836_sv2v_reg ,\piso.data_r_835_sv2v_reg ,\piso.data_r_834_sv2v_reg ,
  \piso.data_r_833_sv2v_reg ,\piso.data_r_832_sv2v_reg ,\piso.data_r_831_sv2v_reg ,
  \piso.data_r_830_sv2v_reg ,\piso.data_r_829_sv2v_reg ,\piso.data_r_828_sv2v_reg ,
  \piso.data_r_827_sv2v_reg ,\piso.data_r_826_sv2v_reg ,\piso.data_r_825_sv2v_reg ,
  \piso.data_r_824_sv2v_reg ,\piso.data_r_823_sv2v_reg ,\piso.data_r_822_sv2v_reg ,
  \piso.data_r_821_sv2v_reg ,\piso.data_r_820_sv2v_reg ,\piso.data_r_819_sv2v_reg ,
  \piso.data_r_818_sv2v_reg ,\piso.data_r_817_sv2v_reg ,\piso.data_r_816_sv2v_reg ,
  \piso.data_r_815_sv2v_reg ,\piso.data_r_814_sv2v_reg ,\piso.data_r_813_sv2v_reg ,
  \piso.data_r_812_sv2v_reg ,\piso.data_r_811_sv2v_reg ,\piso.data_r_810_sv2v_reg ,
  \piso.data_r_809_sv2v_reg ,\piso.data_r_808_sv2v_reg ,\piso.data_r_807_sv2v_reg ,
  \piso.data_r_806_sv2v_reg ,\piso.data_r_805_sv2v_reg ,\piso.data_r_804_sv2v_reg ,
  \piso.data_r_803_sv2v_reg ,\piso.data_r_802_sv2v_reg ,\piso.data_r_801_sv2v_reg ,
  \piso.data_r_800_sv2v_reg ,\piso.data_r_799_sv2v_reg ,\piso.data_r_798_sv2v_reg ,
  \piso.data_r_797_sv2v_reg ,\piso.data_r_796_sv2v_reg ,\piso.data_r_795_sv2v_reg ,
  \piso.data_r_794_sv2v_reg ,\piso.data_r_793_sv2v_reg ,
  \piso.data_r_792_sv2v_reg ,\piso.data_r_791_sv2v_reg ,\piso.data_r_790_sv2v_reg ,
  \piso.data_r_789_sv2v_reg ,\piso.data_r_788_sv2v_reg ,\piso.data_r_787_sv2v_reg ,
  \piso.data_r_786_sv2v_reg ,\piso.data_r_785_sv2v_reg ,\piso.data_r_784_sv2v_reg ,
  \piso.data_r_783_sv2v_reg ,\piso.data_r_782_sv2v_reg ,\piso.data_r_781_sv2v_reg ,
  \piso.data_r_780_sv2v_reg ,\piso.data_r_779_sv2v_reg ,\piso.data_r_778_sv2v_reg ,
  \piso.data_r_777_sv2v_reg ,\piso.data_r_776_sv2v_reg ,\piso.data_r_775_sv2v_reg ,
  \piso.data_r_774_sv2v_reg ,\piso.data_r_773_sv2v_reg ,\piso.data_r_772_sv2v_reg ,
  \piso.data_r_771_sv2v_reg ,\piso.data_r_770_sv2v_reg ,\piso.data_r_769_sv2v_reg ,
  \piso.data_r_768_sv2v_reg ,\piso.data_r_767_sv2v_reg ,\piso.data_r_766_sv2v_reg ,
  \piso.data_r_765_sv2v_reg ,\piso.data_r_764_sv2v_reg ,\piso.data_r_763_sv2v_reg ,
  \piso.data_r_762_sv2v_reg ,\piso.data_r_761_sv2v_reg ,\piso.data_r_760_sv2v_reg ,
  \piso.data_r_759_sv2v_reg ,\piso.data_r_758_sv2v_reg ,\piso.data_r_757_sv2v_reg ,
  \piso.data_r_756_sv2v_reg ,\piso.data_r_755_sv2v_reg ,\piso.data_r_754_sv2v_reg ,
  \piso.data_r_753_sv2v_reg ,\piso.data_r_752_sv2v_reg ,\piso.data_r_751_sv2v_reg ,
  \piso.data_r_750_sv2v_reg ,\piso.data_r_749_sv2v_reg ,\piso.data_r_748_sv2v_reg ,
  \piso.data_r_747_sv2v_reg ,\piso.data_r_746_sv2v_reg ,\piso.data_r_745_sv2v_reg ,
  \piso.data_r_744_sv2v_reg ,\piso.data_r_743_sv2v_reg ,\piso.data_r_742_sv2v_reg ,
  \piso.data_r_741_sv2v_reg ,\piso.data_r_740_sv2v_reg ,\piso.data_r_739_sv2v_reg ,
  \piso.data_r_738_sv2v_reg ,\piso.data_r_737_sv2v_reg ,\piso.data_r_736_sv2v_reg ,
  \piso.data_r_735_sv2v_reg ,\piso.data_r_734_sv2v_reg ,\piso.data_r_733_sv2v_reg ,
  \piso.data_r_732_sv2v_reg ,\piso.data_r_731_sv2v_reg ,\piso.data_r_730_sv2v_reg ,
  \piso.data_r_729_sv2v_reg ,\piso.data_r_728_sv2v_reg ,\piso.data_r_727_sv2v_reg ,
  \piso.data_r_726_sv2v_reg ,\piso.data_r_725_sv2v_reg ,\piso.data_r_724_sv2v_reg ,
  \piso.data_r_723_sv2v_reg ,\piso.data_r_722_sv2v_reg ,\piso.data_r_721_sv2v_reg ,
  \piso.data_r_720_sv2v_reg ,\piso.data_r_719_sv2v_reg ,\piso.data_r_718_sv2v_reg ,
  \piso.data_r_717_sv2v_reg ,\piso.data_r_716_sv2v_reg ,\piso.data_r_715_sv2v_reg ,
  \piso.data_r_714_sv2v_reg ,\piso.data_r_713_sv2v_reg ,
  \piso.data_r_712_sv2v_reg ,\piso.data_r_711_sv2v_reg ,\piso.data_r_710_sv2v_reg ,
  \piso.data_r_709_sv2v_reg ,\piso.data_r_708_sv2v_reg ,\piso.data_r_707_sv2v_reg ,
  \piso.data_r_706_sv2v_reg ,\piso.data_r_705_sv2v_reg ,\piso.data_r_704_sv2v_reg ,
  \piso.data_r_703_sv2v_reg ,\piso.data_r_702_sv2v_reg ,\piso.data_r_701_sv2v_reg ,
  \piso.data_r_700_sv2v_reg ,\piso.data_r_699_sv2v_reg ,\piso.data_r_698_sv2v_reg ,
  \piso.data_r_697_sv2v_reg ,\piso.data_r_696_sv2v_reg ,\piso.data_r_695_sv2v_reg ,
  \piso.data_r_694_sv2v_reg ,\piso.data_r_693_sv2v_reg ,\piso.data_r_692_sv2v_reg ,
  \piso.data_r_691_sv2v_reg ,\piso.data_r_690_sv2v_reg ,\piso.data_r_689_sv2v_reg ,
  \piso.data_r_688_sv2v_reg ,\piso.data_r_687_sv2v_reg ,\piso.data_r_686_sv2v_reg ,
  \piso.data_r_685_sv2v_reg ,\piso.data_r_684_sv2v_reg ,\piso.data_r_683_sv2v_reg ,
  \piso.data_r_682_sv2v_reg ,\piso.data_r_681_sv2v_reg ,\piso.data_r_680_sv2v_reg ,
  \piso.data_r_679_sv2v_reg ,\piso.data_r_678_sv2v_reg ,\piso.data_r_677_sv2v_reg ,
  \piso.data_r_676_sv2v_reg ,\piso.data_r_675_sv2v_reg ,\piso.data_r_674_sv2v_reg ,
  \piso.data_r_673_sv2v_reg ,\piso.data_r_672_sv2v_reg ,\piso.data_r_671_sv2v_reg ,
  \piso.data_r_670_sv2v_reg ,\piso.data_r_669_sv2v_reg ,\piso.data_r_668_sv2v_reg ,
  \piso.data_r_667_sv2v_reg ,\piso.data_r_666_sv2v_reg ,\piso.data_r_665_sv2v_reg ,
  \piso.data_r_664_sv2v_reg ,\piso.data_r_663_sv2v_reg ,\piso.data_r_662_sv2v_reg ,
  \piso.data_r_661_sv2v_reg ,\piso.data_r_660_sv2v_reg ,\piso.data_r_659_sv2v_reg ,
  \piso.data_r_658_sv2v_reg ,\piso.data_r_657_sv2v_reg ,\piso.data_r_656_sv2v_reg ,
  \piso.data_r_655_sv2v_reg ,\piso.data_r_654_sv2v_reg ,\piso.data_r_653_sv2v_reg ,
  \piso.data_r_652_sv2v_reg ,\piso.data_r_651_sv2v_reg ,\piso.data_r_650_sv2v_reg ,
  \piso.data_r_649_sv2v_reg ,\piso.data_r_648_sv2v_reg ,\piso.data_r_647_sv2v_reg ,
  \piso.data_r_646_sv2v_reg ,\piso.data_r_645_sv2v_reg ,\piso.data_r_644_sv2v_reg ,
  \piso.data_r_643_sv2v_reg ,\piso.data_r_642_sv2v_reg ,\piso.data_r_641_sv2v_reg ,
  \piso.data_r_640_sv2v_reg ,\piso.data_r_639_sv2v_reg ,\piso.data_r_638_sv2v_reg ,
  \piso.data_r_637_sv2v_reg ,\piso.data_r_636_sv2v_reg ,\piso.data_r_635_sv2v_reg ,
  \piso.data_r_634_sv2v_reg ,\piso.data_r_633_sv2v_reg ,
  \piso.data_r_632_sv2v_reg ,\piso.data_r_631_sv2v_reg ,\piso.data_r_630_sv2v_reg ,
  \piso.data_r_629_sv2v_reg ,\piso.data_r_628_sv2v_reg ,\piso.data_r_627_sv2v_reg ,
  \piso.data_r_626_sv2v_reg ,\piso.data_r_625_sv2v_reg ,\piso.data_r_624_sv2v_reg ,
  \piso.data_r_623_sv2v_reg ,\piso.data_r_622_sv2v_reg ,\piso.data_r_621_sv2v_reg ,
  \piso.data_r_620_sv2v_reg ,\piso.data_r_619_sv2v_reg ,\piso.data_r_618_sv2v_reg ,
  \piso.data_r_617_sv2v_reg ,\piso.data_r_616_sv2v_reg ,\piso.data_r_615_sv2v_reg ,
  \piso.data_r_614_sv2v_reg ,\piso.data_r_613_sv2v_reg ,\piso.data_r_612_sv2v_reg ,
  \piso.data_r_611_sv2v_reg ,\piso.data_r_610_sv2v_reg ,\piso.data_r_609_sv2v_reg ,
  \piso.data_r_608_sv2v_reg ,\piso.data_r_607_sv2v_reg ,\piso.data_r_606_sv2v_reg ,
  \piso.data_r_605_sv2v_reg ,\piso.data_r_604_sv2v_reg ,\piso.data_r_603_sv2v_reg ,
  \piso.data_r_602_sv2v_reg ,\piso.data_r_601_sv2v_reg ,\piso.data_r_600_sv2v_reg ,
  \piso.data_r_599_sv2v_reg ,\piso.data_r_598_sv2v_reg ,\piso.data_r_597_sv2v_reg ,
  \piso.data_r_596_sv2v_reg ,\piso.data_r_595_sv2v_reg ,\piso.data_r_594_sv2v_reg ,
  \piso.data_r_593_sv2v_reg ,\piso.data_r_592_sv2v_reg ,\piso.data_r_591_sv2v_reg ,
  \piso.data_r_590_sv2v_reg ,\piso.data_r_589_sv2v_reg ,\piso.data_r_588_sv2v_reg ,
  \piso.data_r_587_sv2v_reg ,\piso.data_r_586_sv2v_reg ,\piso.data_r_585_sv2v_reg ,
  \piso.data_r_584_sv2v_reg ,\piso.data_r_583_sv2v_reg ,\piso.data_r_582_sv2v_reg ,
  \piso.data_r_581_sv2v_reg ,\piso.data_r_580_sv2v_reg ,\piso.data_r_579_sv2v_reg ,
  \piso.data_r_578_sv2v_reg ,\piso.data_r_577_sv2v_reg ,\piso.data_r_576_sv2v_reg ,
  \piso.data_r_575_sv2v_reg ,\piso.data_r_574_sv2v_reg ,\piso.data_r_573_sv2v_reg ,
  \piso.data_r_572_sv2v_reg ,\piso.data_r_571_sv2v_reg ,\piso.data_r_570_sv2v_reg ,
  \piso.data_r_569_sv2v_reg ,\piso.data_r_568_sv2v_reg ,\piso.data_r_567_sv2v_reg ,
  \piso.data_r_566_sv2v_reg ,\piso.data_r_565_sv2v_reg ,\piso.data_r_564_sv2v_reg ,
  \piso.data_r_563_sv2v_reg ,\piso.data_r_562_sv2v_reg ,\piso.data_r_561_sv2v_reg ,
  \piso.data_r_560_sv2v_reg ,\piso.data_r_559_sv2v_reg ,\piso.data_r_558_sv2v_reg ,
  \piso.data_r_557_sv2v_reg ,\piso.data_r_556_sv2v_reg ,\piso.data_r_555_sv2v_reg ,
  \piso.data_r_554_sv2v_reg ,\piso.data_r_553_sv2v_reg ,
  \piso.data_r_552_sv2v_reg ,\piso.data_r_551_sv2v_reg ,\piso.data_r_550_sv2v_reg ,
  \piso.data_r_549_sv2v_reg ,\piso.data_r_548_sv2v_reg ,\piso.data_r_547_sv2v_reg ,
  \piso.data_r_546_sv2v_reg ,\piso.data_r_545_sv2v_reg ,\piso.data_r_544_sv2v_reg ,
  \piso.data_r_543_sv2v_reg ,\piso.data_r_542_sv2v_reg ,\piso.data_r_541_sv2v_reg ,
  \piso.data_r_540_sv2v_reg ,\piso.data_r_539_sv2v_reg ,\piso.data_r_538_sv2v_reg ,
  \piso.data_r_537_sv2v_reg ,\piso.data_r_536_sv2v_reg ,\piso.data_r_535_sv2v_reg ,
  \piso.data_r_534_sv2v_reg ,\piso.data_r_533_sv2v_reg ,\piso.data_r_532_sv2v_reg ,
  \piso.data_r_531_sv2v_reg ,\piso.data_r_530_sv2v_reg ,\piso.data_r_529_sv2v_reg ,
  \piso.data_r_528_sv2v_reg ,\piso.data_r_527_sv2v_reg ,\piso.data_r_526_sv2v_reg ,
  \piso.data_r_525_sv2v_reg ,\piso.data_r_524_sv2v_reg ,\piso.data_r_523_sv2v_reg ,
  \piso.data_r_522_sv2v_reg ,\piso.data_r_521_sv2v_reg ,\piso.data_r_520_sv2v_reg ,
  \piso.data_r_519_sv2v_reg ,\piso.data_r_518_sv2v_reg ,\piso.data_r_517_sv2v_reg ,
  \piso.data_r_516_sv2v_reg ,\piso.data_r_515_sv2v_reg ,\piso.data_r_514_sv2v_reg ,
  \piso.data_r_513_sv2v_reg ,\piso.data_r_512_sv2v_reg ,\piso.data_r_511_sv2v_reg ,
  \piso.data_r_510_sv2v_reg ,\piso.data_r_509_sv2v_reg ,\piso.data_r_508_sv2v_reg ,
  \piso.data_r_507_sv2v_reg ,\piso.data_r_506_sv2v_reg ,\piso.data_r_505_sv2v_reg ,
  \piso.data_r_504_sv2v_reg ,\piso.data_r_503_sv2v_reg ,\piso.data_r_502_sv2v_reg ,
  \piso.data_r_501_sv2v_reg ,\piso.data_r_500_sv2v_reg ,\piso.data_r_499_sv2v_reg ,
  \piso.data_r_498_sv2v_reg ,\piso.data_r_497_sv2v_reg ,\piso.data_r_496_sv2v_reg ,
  \piso.data_r_495_sv2v_reg ,\piso.data_r_494_sv2v_reg ,\piso.data_r_493_sv2v_reg ,
  \piso.data_r_492_sv2v_reg ,\piso.data_r_491_sv2v_reg ,\piso.data_r_490_sv2v_reg ,
  \piso.data_r_489_sv2v_reg ,\piso.data_r_488_sv2v_reg ,\piso.data_r_487_sv2v_reg ,
  \piso.data_r_486_sv2v_reg ,\piso.data_r_485_sv2v_reg ,\piso.data_r_484_sv2v_reg ,
  \piso.data_r_483_sv2v_reg ,\piso.data_r_482_sv2v_reg ,\piso.data_r_481_sv2v_reg ,
  \piso.data_r_480_sv2v_reg ,\piso.data_r_479_sv2v_reg ,\piso.data_r_478_sv2v_reg ,
  \piso.data_r_477_sv2v_reg ,\piso.data_r_476_sv2v_reg ,\piso.data_r_475_sv2v_reg ,
  \piso.data_r_474_sv2v_reg ,\piso.data_r_473_sv2v_reg ,
  \piso.data_r_472_sv2v_reg ,\piso.data_r_471_sv2v_reg ,\piso.data_r_470_sv2v_reg ,
  \piso.data_r_469_sv2v_reg ,\piso.data_r_468_sv2v_reg ,\piso.data_r_467_sv2v_reg ,
  \piso.data_r_466_sv2v_reg ,\piso.data_r_465_sv2v_reg ,\piso.data_r_464_sv2v_reg ,
  \piso.data_r_463_sv2v_reg ,\piso.data_r_462_sv2v_reg ,\piso.data_r_461_sv2v_reg ,
  \piso.data_r_460_sv2v_reg ,\piso.data_r_459_sv2v_reg ,\piso.data_r_458_sv2v_reg ,
  \piso.data_r_457_sv2v_reg ,\piso.data_r_456_sv2v_reg ,\piso.data_r_455_sv2v_reg ,
  \piso.data_r_454_sv2v_reg ,\piso.data_r_453_sv2v_reg ,\piso.data_r_452_sv2v_reg ,
  \piso.data_r_451_sv2v_reg ,\piso.data_r_450_sv2v_reg ,\piso.data_r_449_sv2v_reg ,
  \piso.data_r_448_sv2v_reg ,\piso.data_r_447_sv2v_reg ,\piso.data_r_446_sv2v_reg ,
  \piso.data_r_445_sv2v_reg ,\piso.data_r_444_sv2v_reg ,\piso.data_r_443_sv2v_reg ,
  \piso.data_r_442_sv2v_reg ,\piso.data_r_441_sv2v_reg ,\piso.data_r_440_sv2v_reg ,
  \piso.data_r_439_sv2v_reg ,\piso.data_r_438_sv2v_reg ,\piso.data_r_437_sv2v_reg ,
  \piso.data_r_436_sv2v_reg ,\piso.data_r_435_sv2v_reg ,\piso.data_r_434_sv2v_reg ,
  \piso.data_r_433_sv2v_reg ,\piso.data_r_432_sv2v_reg ,\piso.data_r_431_sv2v_reg ,
  \piso.data_r_430_sv2v_reg ,\piso.data_r_429_sv2v_reg ,\piso.data_r_428_sv2v_reg ,
  \piso.data_r_427_sv2v_reg ,\piso.data_r_426_sv2v_reg ,\piso.data_r_425_sv2v_reg ,
  \piso.data_r_424_sv2v_reg ,\piso.data_r_423_sv2v_reg ,\piso.data_r_422_sv2v_reg ,
  \piso.data_r_421_sv2v_reg ,\piso.data_r_420_sv2v_reg ,\piso.data_r_419_sv2v_reg ,
  \piso.data_r_418_sv2v_reg ,\piso.data_r_417_sv2v_reg ,\piso.data_r_416_sv2v_reg ,
  \piso.data_r_415_sv2v_reg ,\piso.data_r_414_sv2v_reg ,\piso.data_r_413_sv2v_reg ,
  \piso.data_r_412_sv2v_reg ,\piso.data_r_411_sv2v_reg ,\piso.data_r_410_sv2v_reg ,
  \piso.data_r_409_sv2v_reg ,\piso.data_r_408_sv2v_reg ,\piso.data_r_407_sv2v_reg ,
  \piso.data_r_406_sv2v_reg ,\piso.data_r_405_sv2v_reg ,\piso.data_r_404_sv2v_reg ,
  \piso.data_r_403_sv2v_reg ,\piso.data_r_402_sv2v_reg ,\piso.data_r_401_sv2v_reg ,
  \piso.data_r_400_sv2v_reg ,\piso.data_r_399_sv2v_reg ,\piso.data_r_398_sv2v_reg ,
  \piso.data_r_397_sv2v_reg ,\piso.data_r_396_sv2v_reg ,\piso.data_r_395_sv2v_reg ,
  \piso.data_r_394_sv2v_reg ,\piso.data_r_393_sv2v_reg ,
  \piso.data_r_392_sv2v_reg ,\piso.data_r_391_sv2v_reg ,\piso.data_r_390_sv2v_reg ,
  \piso.data_r_389_sv2v_reg ,\piso.data_r_388_sv2v_reg ,\piso.data_r_387_sv2v_reg ,
  \piso.data_r_386_sv2v_reg ,\piso.data_r_385_sv2v_reg ,\piso.data_r_384_sv2v_reg ,
  \piso.data_r_383_sv2v_reg ,\piso.data_r_382_sv2v_reg ,\piso.data_r_381_sv2v_reg ,
  \piso.data_r_380_sv2v_reg ,\piso.data_r_379_sv2v_reg ,\piso.data_r_378_sv2v_reg ,
  \piso.data_r_377_sv2v_reg ,\piso.data_r_376_sv2v_reg ,\piso.data_r_375_sv2v_reg ,
  \piso.data_r_374_sv2v_reg ,\piso.data_r_373_sv2v_reg ,\piso.data_r_372_sv2v_reg ,
  \piso.data_r_371_sv2v_reg ,\piso.data_r_370_sv2v_reg ,\piso.data_r_369_sv2v_reg ,
  \piso.data_r_368_sv2v_reg ,\piso.data_r_367_sv2v_reg ,\piso.data_r_366_sv2v_reg ,
  \piso.data_r_365_sv2v_reg ,\piso.data_r_364_sv2v_reg ,\piso.data_r_363_sv2v_reg ,
  \piso.data_r_362_sv2v_reg ,\piso.data_r_361_sv2v_reg ,\piso.data_r_360_sv2v_reg ,
  \piso.data_r_359_sv2v_reg ,\piso.data_r_358_sv2v_reg ,\piso.data_r_357_sv2v_reg ,
  \piso.data_r_356_sv2v_reg ,\piso.data_r_355_sv2v_reg ,\piso.data_r_354_sv2v_reg ,
  \piso.data_r_353_sv2v_reg ,\piso.data_r_352_sv2v_reg ,\piso.data_r_351_sv2v_reg ,
  \piso.data_r_350_sv2v_reg ,\piso.data_r_349_sv2v_reg ,\piso.data_r_348_sv2v_reg ,
  \piso.data_r_347_sv2v_reg ,\piso.data_r_346_sv2v_reg ,\piso.data_r_345_sv2v_reg ,
  \piso.data_r_344_sv2v_reg ,\piso.data_r_343_sv2v_reg ,\piso.data_r_342_sv2v_reg ,
  \piso.data_r_341_sv2v_reg ,\piso.data_r_340_sv2v_reg ,\piso.data_r_339_sv2v_reg ,
  \piso.data_r_338_sv2v_reg ,\piso.data_r_337_sv2v_reg ,\piso.data_r_336_sv2v_reg ,
  \piso.data_r_335_sv2v_reg ,\piso.data_r_334_sv2v_reg ,\piso.data_r_333_sv2v_reg ,
  \piso.data_r_332_sv2v_reg ,\piso.data_r_331_sv2v_reg ,\piso.data_r_330_sv2v_reg ,
  \piso.data_r_329_sv2v_reg ,\piso.data_r_328_sv2v_reg ,\piso.data_r_327_sv2v_reg ,
  \piso.data_r_326_sv2v_reg ,\piso.data_r_325_sv2v_reg ,\piso.data_r_324_sv2v_reg ,
  \piso.data_r_323_sv2v_reg ,\piso.data_r_322_sv2v_reg ,\piso.data_r_321_sv2v_reg ,
  \piso.data_r_320_sv2v_reg ,\piso.data_r_319_sv2v_reg ,\piso.data_r_318_sv2v_reg ,
  \piso.data_r_317_sv2v_reg ,\piso.data_r_316_sv2v_reg ,\piso.data_r_315_sv2v_reg ,
  \piso.data_r_314_sv2v_reg ,\piso.data_r_313_sv2v_reg ,
  \piso.data_r_312_sv2v_reg ,\piso.data_r_311_sv2v_reg ,\piso.data_r_310_sv2v_reg ,
  \piso.data_r_309_sv2v_reg ,\piso.data_r_308_sv2v_reg ,\piso.data_r_307_sv2v_reg ,
  \piso.data_r_306_sv2v_reg ,\piso.data_r_305_sv2v_reg ,\piso.data_r_304_sv2v_reg ,
  \piso.data_r_303_sv2v_reg ,\piso.data_r_302_sv2v_reg ,\piso.data_r_301_sv2v_reg ,
  \piso.data_r_300_sv2v_reg ,\piso.data_r_299_sv2v_reg ,\piso.data_r_298_sv2v_reg ,
  \piso.data_r_297_sv2v_reg ,\piso.data_r_296_sv2v_reg ,\piso.data_r_295_sv2v_reg ,
  \piso.data_r_294_sv2v_reg ,\piso.data_r_293_sv2v_reg ,\piso.data_r_292_sv2v_reg ,
  \piso.data_r_291_sv2v_reg ,\piso.data_r_290_sv2v_reg ,\piso.data_r_289_sv2v_reg ,
  \piso.data_r_288_sv2v_reg ,\piso.data_r_287_sv2v_reg ,\piso.data_r_286_sv2v_reg ,
  \piso.data_r_285_sv2v_reg ,\piso.data_r_284_sv2v_reg ,\piso.data_r_283_sv2v_reg ,
  \piso.data_r_282_sv2v_reg ,\piso.data_r_281_sv2v_reg ,\piso.data_r_280_sv2v_reg ,
  \piso.data_r_279_sv2v_reg ,\piso.data_r_278_sv2v_reg ,\piso.data_r_277_sv2v_reg ,
  \piso.data_r_276_sv2v_reg ,\piso.data_r_275_sv2v_reg ,\piso.data_r_274_sv2v_reg ,
  \piso.data_r_273_sv2v_reg ,\piso.data_r_272_sv2v_reg ,\piso.data_r_271_sv2v_reg ,
  \piso.data_r_270_sv2v_reg ,\piso.data_r_269_sv2v_reg ,\piso.data_r_268_sv2v_reg ,
  \piso.data_r_267_sv2v_reg ,\piso.data_r_266_sv2v_reg ,\piso.data_r_265_sv2v_reg ,
  \piso.data_r_264_sv2v_reg ,\piso.data_r_263_sv2v_reg ,\piso.data_r_262_sv2v_reg ,
  \piso.data_r_261_sv2v_reg ,\piso.data_r_260_sv2v_reg ,\piso.data_r_259_sv2v_reg ,
  \piso.data_r_258_sv2v_reg ,\piso.data_r_257_sv2v_reg ,\piso.data_r_256_sv2v_reg ,
  \piso.data_r_255_sv2v_reg ,\piso.data_r_254_sv2v_reg ,\piso.data_r_253_sv2v_reg ,
  \piso.data_r_252_sv2v_reg ,\piso.data_r_251_sv2v_reg ,\piso.data_r_250_sv2v_reg ,
  \piso.data_r_249_sv2v_reg ,\piso.data_r_248_sv2v_reg ,\piso.data_r_247_sv2v_reg ,
  \piso.data_r_246_sv2v_reg ,\piso.data_r_245_sv2v_reg ,\piso.data_r_244_sv2v_reg ,
  \piso.data_r_243_sv2v_reg ,\piso.data_r_242_sv2v_reg ,\piso.data_r_241_sv2v_reg ,
  \piso.data_r_240_sv2v_reg ,\piso.data_r_239_sv2v_reg ,\piso.data_r_238_sv2v_reg ,
  \piso.data_r_237_sv2v_reg ,\piso.data_r_236_sv2v_reg ,\piso.data_r_235_sv2v_reg ,
  \piso.data_r_234_sv2v_reg ,\piso.data_r_233_sv2v_reg ,
  \piso.data_r_232_sv2v_reg ,\piso.data_r_231_sv2v_reg ,\piso.data_r_230_sv2v_reg ,
  \piso.data_r_229_sv2v_reg ,\piso.data_r_228_sv2v_reg ,\piso.data_r_227_sv2v_reg ,
  \piso.data_r_226_sv2v_reg ,\piso.data_r_225_sv2v_reg ,\piso.data_r_224_sv2v_reg ,
  \piso.data_r_223_sv2v_reg ,\piso.data_r_222_sv2v_reg ,\piso.data_r_221_sv2v_reg ,
  \piso.data_r_220_sv2v_reg ,\piso.data_r_219_sv2v_reg ,\piso.data_r_218_sv2v_reg ,
  \piso.data_r_217_sv2v_reg ,\piso.data_r_216_sv2v_reg ,\piso.data_r_215_sv2v_reg ,
  \piso.data_r_214_sv2v_reg ,\piso.data_r_213_sv2v_reg ,\piso.data_r_212_sv2v_reg ,
  \piso.data_r_211_sv2v_reg ,\piso.data_r_210_sv2v_reg ,\piso.data_r_209_sv2v_reg ,
  \piso.data_r_208_sv2v_reg ,\piso.data_r_207_sv2v_reg ,\piso.data_r_206_sv2v_reg ,
  \piso.data_r_205_sv2v_reg ,\piso.data_r_204_sv2v_reg ,\piso.data_r_203_sv2v_reg ,
  \piso.data_r_202_sv2v_reg ,\piso.data_r_201_sv2v_reg ,\piso.data_r_200_sv2v_reg ,
  \piso.data_r_199_sv2v_reg ,\piso.data_r_198_sv2v_reg ,\piso.data_r_197_sv2v_reg ,
  \piso.data_r_196_sv2v_reg ,\piso.data_r_195_sv2v_reg ,\piso.data_r_194_sv2v_reg ,
  \piso.data_r_193_sv2v_reg ,\piso.data_r_192_sv2v_reg ,\piso.data_r_191_sv2v_reg ,
  \piso.data_r_190_sv2v_reg ,\piso.data_r_189_sv2v_reg ,\piso.data_r_188_sv2v_reg ,
  \piso.data_r_187_sv2v_reg ,\piso.data_r_186_sv2v_reg ,\piso.data_r_185_sv2v_reg ,
  \piso.data_r_184_sv2v_reg ,\piso.data_r_183_sv2v_reg ,\piso.data_r_182_sv2v_reg ,
  \piso.data_r_181_sv2v_reg ,\piso.data_r_180_sv2v_reg ,\piso.data_r_179_sv2v_reg ,
  \piso.data_r_178_sv2v_reg ,\piso.data_r_177_sv2v_reg ,\piso.data_r_176_sv2v_reg ,
  \piso.data_r_175_sv2v_reg ,\piso.data_r_174_sv2v_reg ,\piso.data_r_173_sv2v_reg ,
  \piso.data_r_172_sv2v_reg ,\piso.data_r_171_sv2v_reg ,\piso.data_r_170_sv2v_reg ,
  \piso.data_r_169_sv2v_reg ,\piso.data_r_168_sv2v_reg ,\piso.data_r_167_sv2v_reg ,
  \piso.data_r_166_sv2v_reg ,\piso.data_r_165_sv2v_reg ,\piso.data_r_164_sv2v_reg ,
  \piso.data_r_163_sv2v_reg ,\piso.data_r_162_sv2v_reg ,\piso.data_r_161_sv2v_reg ,
  \piso.data_r_160_sv2v_reg ,\piso.data_r_159_sv2v_reg ,\piso.data_r_158_sv2v_reg ,
  \piso.data_r_157_sv2v_reg ,\piso.data_r_156_sv2v_reg ,\piso.data_r_155_sv2v_reg ,
  \piso.data_r_154_sv2v_reg ,\piso.data_r_153_sv2v_reg ,
  \piso.data_r_152_sv2v_reg ,\piso.data_r_151_sv2v_reg ,\piso.data_r_150_sv2v_reg ,
  \piso.data_r_149_sv2v_reg ,\piso.data_r_148_sv2v_reg ,\piso.data_r_147_sv2v_reg ,
  \piso.data_r_146_sv2v_reg ,\piso.data_r_145_sv2v_reg ,\piso.data_r_144_sv2v_reg ,
  \piso.data_r_143_sv2v_reg ,\piso.data_r_142_sv2v_reg ,\piso.data_r_141_sv2v_reg ,
  \piso.data_r_140_sv2v_reg ,\piso.data_r_139_sv2v_reg ,\piso.data_r_138_sv2v_reg ,
  \piso.data_r_137_sv2v_reg ,\piso.data_r_136_sv2v_reg ,\piso.data_r_135_sv2v_reg ,
  \piso.data_r_134_sv2v_reg ,\piso.data_r_133_sv2v_reg ,\piso.data_r_132_sv2v_reg ,
  \piso.data_r_131_sv2v_reg ,\piso.data_r_130_sv2v_reg ,\piso.data_r_129_sv2v_reg ,
  \piso.data_r_128_sv2v_reg ,\piso.data_r_127_sv2v_reg ,\piso.data_r_126_sv2v_reg ,
  \piso.data_r_125_sv2v_reg ,\piso.data_r_124_sv2v_reg ,\piso.data_r_123_sv2v_reg ,
  \piso.data_r_122_sv2v_reg ,\piso.data_r_121_sv2v_reg ,\piso.data_r_120_sv2v_reg ,
  \piso.data_r_119_sv2v_reg ,\piso.data_r_118_sv2v_reg ,\piso.data_r_117_sv2v_reg ,
  \piso.data_r_116_sv2v_reg ,\piso.data_r_115_sv2v_reg ,\piso.data_r_114_sv2v_reg ,
  \piso.data_r_113_sv2v_reg ,\piso.data_r_112_sv2v_reg ,\piso.data_r_111_sv2v_reg ,
  \piso.data_r_110_sv2v_reg ,\piso.data_r_109_sv2v_reg ,\piso.data_r_108_sv2v_reg ,
  \piso.data_r_107_sv2v_reg ,\piso.data_r_106_sv2v_reg ,\piso.data_r_105_sv2v_reg ,
  \piso.data_r_104_sv2v_reg ,\piso.data_r_103_sv2v_reg ,\piso.data_r_102_sv2v_reg ,
  \piso.data_r_101_sv2v_reg ,\piso.data_r_100_sv2v_reg ,\piso.data_r_99_sv2v_reg ,
  \piso.data_r_98_sv2v_reg ,\piso.data_r_97_sv2v_reg ,\piso.data_r_96_sv2v_reg ,
  \piso.data_r_95_sv2v_reg ,\piso.data_r_94_sv2v_reg ,\piso.data_r_93_sv2v_reg ,
  \piso.data_r_92_sv2v_reg ,\piso.data_r_91_sv2v_reg ,\piso.data_r_90_sv2v_reg ,
  \piso.data_r_89_sv2v_reg ,\piso.data_r_88_sv2v_reg ,\piso.data_r_87_sv2v_reg ,
  \piso.data_r_86_sv2v_reg ,\piso.data_r_85_sv2v_reg ,\piso.data_r_84_sv2v_reg ,
  \piso.data_r_83_sv2v_reg ,\piso.data_r_82_sv2v_reg ,\piso.data_r_81_sv2v_reg ,
  \piso.data_r_80_sv2v_reg ,\piso.data_r_79_sv2v_reg ,\piso.data_r_78_sv2v_reg ,
  \piso.data_r_77_sv2v_reg ,\piso.data_r_76_sv2v_reg ,\piso.data_r_75_sv2v_reg ,
  \piso.data_r_74_sv2v_reg ,\piso.data_r_73_sv2v_reg ,\piso.data_r_72_sv2v_reg ,\piso.data_r_71_sv2v_reg ,
  \piso.data_r_70_sv2v_reg ,\piso.data_r_69_sv2v_reg ,\piso.data_r_68_sv2v_reg ,
  \piso.data_r_67_sv2v_reg ,\piso.data_r_66_sv2v_reg ,\piso.data_r_65_sv2v_reg ,
  \piso.data_r_64_sv2v_reg ,\piso.data_r_63_sv2v_reg ,\piso.data_r_62_sv2v_reg ,
  \piso.data_r_61_sv2v_reg ,\piso.data_r_60_sv2v_reg ,\piso.data_r_59_sv2v_reg ,
  \piso.data_r_58_sv2v_reg ,\piso.data_r_57_sv2v_reg ,\piso.data_r_56_sv2v_reg ,
  \piso.data_r_55_sv2v_reg ,\piso.data_r_54_sv2v_reg ,\piso.data_r_53_sv2v_reg ,
  \piso.data_r_52_sv2v_reg ,\piso.data_r_51_sv2v_reg ,\piso.data_r_50_sv2v_reg ,
  \piso.data_r_49_sv2v_reg ,\piso.data_r_48_sv2v_reg ,\piso.data_r_47_sv2v_reg ,
  \piso.data_r_46_sv2v_reg ,\piso.data_r_45_sv2v_reg ,\piso.data_r_44_sv2v_reg ,
  \piso.data_r_43_sv2v_reg ,\piso.data_r_42_sv2v_reg ,\piso.data_r_41_sv2v_reg ,
  \piso.data_r_40_sv2v_reg ,\piso.data_r_39_sv2v_reg ,\piso.data_r_38_sv2v_reg ,
  \piso.data_r_37_sv2v_reg ,\piso.data_r_36_sv2v_reg ,\piso.data_r_35_sv2v_reg ,
  \piso.data_r_34_sv2v_reg ,\piso.data_r_33_sv2v_reg ,\piso.data_r_32_sv2v_reg ,\piso.data_r_31_sv2v_reg ,
  \piso.data_r_30_sv2v_reg ,\piso.data_r_29_sv2v_reg ,\piso.data_r_28_sv2v_reg ,
  \piso.data_r_27_sv2v_reg ,\piso.data_r_26_sv2v_reg ,\piso.data_r_25_sv2v_reg ,
  \piso.data_r_24_sv2v_reg ,\piso.data_r_23_sv2v_reg ,\piso.data_r_22_sv2v_reg ,
  \piso.data_r_21_sv2v_reg ,\piso.data_r_20_sv2v_reg ,\piso.data_r_19_sv2v_reg ,
  \piso.data_r_18_sv2v_reg ,\piso.data_r_17_sv2v_reg ,\piso.data_r_16_sv2v_reg ,
  \piso.data_r_15_sv2v_reg ,\piso.data_r_14_sv2v_reg ,\piso.data_r_13_sv2v_reg ,
  \piso.data_r_12_sv2v_reg ,\piso.data_r_11_sv2v_reg ,\piso.data_r_10_sv2v_reg ,
  \piso.data_r_9_sv2v_reg ,\piso.data_r_8_sv2v_reg ,\piso.data_r_7_sv2v_reg ,
  \piso.data_r_6_sv2v_reg ,\piso.data_r_5_sv2v_reg ,\piso.data_r_4_sv2v_reg ,\piso.data_r_3_sv2v_reg ,
  \piso.data_r_2_sv2v_reg ,\piso.data_r_1_sv2v_reg ,\piso.data_r_0_sv2v_reg ,
  \piso.shift_ctr_r_6_sv2v_reg ,\piso.shift_ctr_r_5_sv2v_reg ,
  \piso.shift_ctr_r_4_sv2v_reg ,\piso.shift_ctr_r_3_sv2v_reg ,\piso.shift_ctr_r_2_sv2v_reg ,
  \piso.shift_ctr_r_1_sv2v_reg ,\piso.shift_ctr_r_0_sv2v_reg ;
  assign valid_o = valid_o_sv2v_reg;
  assign \piso.data_r [4095] = \piso.data_r_4095_sv2v_reg ;
  assign \piso.data_r [4094] = \piso.data_r_4094_sv2v_reg ;
  assign \piso.data_r [4093] = \piso.data_r_4093_sv2v_reg ;
  assign \piso.data_r [4092] = \piso.data_r_4092_sv2v_reg ;
  assign \piso.data_r [4091] = \piso.data_r_4091_sv2v_reg ;
  assign \piso.data_r [4090] = \piso.data_r_4090_sv2v_reg ;
  assign \piso.data_r [4089] = \piso.data_r_4089_sv2v_reg ;
  assign \piso.data_r [4088] = \piso.data_r_4088_sv2v_reg ;
  assign \piso.data_r [4087] = \piso.data_r_4087_sv2v_reg ;
  assign \piso.data_r [4086] = \piso.data_r_4086_sv2v_reg ;
  assign \piso.data_r [4085] = \piso.data_r_4085_sv2v_reg ;
  assign \piso.data_r [4084] = \piso.data_r_4084_sv2v_reg ;
  assign \piso.data_r [4083] = \piso.data_r_4083_sv2v_reg ;
  assign \piso.data_r [4082] = \piso.data_r_4082_sv2v_reg ;
  assign \piso.data_r [4081] = \piso.data_r_4081_sv2v_reg ;
  assign \piso.data_r [4080] = \piso.data_r_4080_sv2v_reg ;
  assign \piso.data_r [4079] = \piso.data_r_4079_sv2v_reg ;
  assign \piso.data_r [4078] = \piso.data_r_4078_sv2v_reg ;
  assign \piso.data_r [4077] = \piso.data_r_4077_sv2v_reg ;
  assign \piso.data_r [4076] = \piso.data_r_4076_sv2v_reg ;
  assign \piso.data_r [4075] = \piso.data_r_4075_sv2v_reg ;
  assign \piso.data_r [4074] = \piso.data_r_4074_sv2v_reg ;
  assign \piso.data_r [4073] = \piso.data_r_4073_sv2v_reg ;
  assign \piso.data_r [4072] = \piso.data_r_4072_sv2v_reg ;
  assign \piso.data_r [4071] = \piso.data_r_4071_sv2v_reg ;
  assign \piso.data_r [4070] = \piso.data_r_4070_sv2v_reg ;
  assign \piso.data_r [4069] = \piso.data_r_4069_sv2v_reg ;
  assign \piso.data_r [4068] = \piso.data_r_4068_sv2v_reg ;
  assign \piso.data_r [4067] = \piso.data_r_4067_sv2v_reg ;
  assign \piso.data_r [4066] = \piso.data_r_4066_sv2v_reg ;
  assign \piso.data_r [4065] = \piso.data_r_4065_sv2v_reg ;
  assign \piso.data_r [4064] = \piso.data_r_4064_sv2v_reg ;
  assign \piso.data_r [4063] = \piso.data_r_4063_sv2v_reg ;
  assign \piso.data_r [4062] = \piso.data_r_4062_sv2v_reg ;
  assign \piso.data_r [4061] = \piso.data_r_4061_sv2v_reg ;
  assign \piso.data_r [4060] = \piso.data_r_4060_sv2v_reg ;
  assign \piso.data_r [4059] = \piso.data_r_4059_sv2v_reg ;
  assign \piso.data_r [4058] = \piso.data_r_4058_sv2v_reg ;
  assign \piso.data_r [4057] = \piso.data_r_4057_sv2v_reg ;
  assign \piso.data_r [4056] = \piso.data_r_4056_sv2v_reg ;
  assign \piso.data_r [4055] = \piso.data_r_4055_sv2v_reg ;
  assign \piso.data_r [4054] = \piso.data_r_4054_sv2v_reg ;
  assign \piso.data_r [4053] = \piso.data_r_4053_sv2v_reg ;
  assign \piso.data_r [4052] = \piso.data_r_4052_sv2v_reg ;
  assign \piso.data_r [4051] = \piso.data_r_4051_sv2v_reg ;
  assign \piso.data_r [4050] = \piso.data_r_4050_sv2v_reg ;
  assign \piso.data_r [4049] = \piso.data_r_4049_sv2v_reg ;
  assign \piso.data_r [4048] = \piso.data_r_4048_sv2v_reg ;
  assign \piso.data_r [4047] = \piso.data_r_4047_sv2v_reg ;
  assign \piso.data_r [4046] = \piso.data_r_4046_sv2v_reg ;
  assign \piso.data_r [4045] = \piso.data_r_4045_sv2v_reg ;
  assign \piso.data_r [4044] = \piso.data_r_4044_sv2v_reg ;
  assign \piso.data_r [4043] = \piso.data_r_4043_sv2v_reg ;
  assign \piso.data_r [4042] = \piso.data_r_4042_sv2v_reg ;
  assign \piso.data_r [4041] = \piso.data_r_4041_sv2v_reg ;
  assign \piso.data_r [4040] = \piso.data_r_4040_sv2v_reg ;
  assign \piso.data_r [4039] = \piso.data_r_4039_sv2v_reg ;
  assign \piso.data_r [4038] = \piso.data_r_4038_sv2v_reg ;
  assign \piso.data_r [4037] = \piso.data_r_4037_sv2v_reg ;
  assign \piso.data_r [4036] = \piso.data_r_4036_sv2v_reg ;
  assign \piso.data_r [4035] = \piso.data_r_4035_sv2v_reg ;
  assign \piso.data_r [4034] = \piso.data_r_4034_sv2v_reg ;
  assign \piso.data_r [4033] = \piso.data_r_4033_sv2v_reg ;
  assign \piso.data_r [4032] = \piso.data_r_4032_sv2v_reg ;
  assign \piso.data_r [4031] = \piso.data_r_4031_sv2v_reg ;
  assign \piso.data_r [4030] = \piso.data_r_4030_sv2v_reg ;
  assign \piso.data_r [4029] = \piso.data_r_4029_sv2v_reg ;
  assign \piso.data_r [4028] = \piso.data_r_4028_sv2v_reg ;
  assign \piso.data_r [4027] = \piso.data_r_4027_sv2v_reg ;
  assign \piso.data_r [4026] = \piso.data_r_4026_sv2v_reg ;
  assign \piso.data_r [4025] = \piso.data_r_4025_sv2v_reg ;
  assign \piso.data_r [4024] = \piso.data_r_4024_sv2v_reg ;
  assign \piso.data_r [4023] = \piso.data_r_4023_sv2v_reg ;
  assign \piso.data_r [4022] = \piso.data_r_4022_sv2v_reg ;
  assign \piso.data_r [4021] = \piso.data_r_4021_sv2v_reg ;
  assign \piso.data_r [4020] = \piso.data_r_4020_sv2v_reg ;
  assign \piso.data_r [4019] = \piso.data_r_4019_sv2v_reg ;
  assign \piso.data_r [4018] = \piso.data_r_4018_sv2v_reg ;
  assign \piso.data_r [4017] = \piso.data_r_4017_sv2v_reg ;
  assign \piso.data_r [4016] = \piso.data_r_4016_sv2v_reg ;
  assign \piso.data_r [4015] = \piso.data_r_4015_sv2v_reg ;
  assign \piso.data_r [4014] = \piso.data_r_4014_sv2v_reg ;
  assign \piso.data_r [4013] = \piso.data_r_4013_sv2v_reg ;
  assign \piso.data_r [4012] = \piso.data_r_4012_sv2v_reg ;
  assign \piso.data_r [4011] = \piso.data_r_4011_sv2v_reg ;
  assign \piso.data_r [4010] = \piso.data_r_4010_sv2v_reg ;
  assign \piso.data_r [4009] = \piso.data_r_4009_sv2v_reg ;
  assign \piso.data_r [4008] = \piso.data_r_4008_sv2v_reg ;
  assign \piso.data_r [4007] = \piso.data_r_4007_sv2v_reg ;
  assign \piso.data_r [4006] = \piso.data_r_4006_sv2v_reg ;
  assign \piso.data_r [4005] = \piso.data_r_4005_sv2v_reg ;
  assign \piso.data_r [4004] = \piso.data_r_4004_sv2v_reg ;
  assign \piso.data_r [4003] = \piso.data_r_4003_sv2v_reg ;
  assign \piso.data_r [4002] = \piso.data_r_4002_sv2v_reg ;
  assign \piso.data_r [4001] = \piso.data_r_4001_sv2v_reg ;
  assign \piso.data_r [4000] = \piso.data_r_4000_sv2v_reg ;
  assign \piso.data_r [3999] = \piso.data_r_3999_sv2v_reg ;
  assign \piso.data_r [3998] = \piso.data_r_3998_sv2v_reg ;
  assign \piso.data_r [3997] = \piso.data_r_3997_sv2v_reg ;
  assign \piso.data_r [3996] = \piso.data_r_3996_sv2v_reg ;
  assign \piso.data_r [3995] = \piso.data_r_3995_sv2v_reg ;
  assign \piso.data_r [3994] = \piso.data_r_3994_sv2v_reg ;
  assign \piso.data_r [3993] = \piso.data_r_3993_sv2v_reg ;
  assign \piso.data_r [3992] = \piso.data_r_3992_sv2v_reg ;
  assign \piso.data_r [3991] = \piso.data_r_3991_sv2v_reg ;
  assign \piso.data_r [3990] = \piso.data_r_3990_sv2v_reg ;
  assign \piso.data_r [3989] = \piso.data_r_3989_sv2v_reg ;
  assign \piso.data_r [3988] = \piso.data_r_3988_sv2v_reg ;
  assign \piso.data_r [3987] = \piso.data_r_3987_sv2v_reg ;
  assign \piso.data_r [3986] = \piso.data_r_3986_sv2v_reg ;
  assign \piso.data_r [3985] = \piso.data_r_3985_sv2v_reg ;
  assign \piso.data_r [3984] = \piso.data_r_3984_sv2v_reg ;
  assign \piso.data_r [3983] = \piso.data_r_3983_sv2v_reg ;
  assign \piso.data_r [3982] = \piso.data_r_3982_sv2v_reg ;
  assign \piso.data_r [3981] = \piso.data_r_3981_sv2v_reg ;
  assign \piso.data_r [3980] = \piso.data_r_3980_sv2v_reg ;
  assign \piso.data_r [3979] = \piso.data_r_3979_sv2v_reg ;
  assign \piso.data_r [3978] = \piso.data_r_3978_sv2v_reg ;
  assign \piso.data_r [3977] = \piso.data_r_3977_sv2v_reg ;
  assign \piso.data_r [3976] = \piso.data_r_3976_sv2v_reg ;
  assign \piso.data_r [3975] = \piso.data_r_3975_sv2v_reg ;
  assign \piso.data_r [3974] = \piso.data_r_3974_sv2v_reg ;
  assign \piso.data_r [3973] = \piso.data_r_3973_sv2v_reg ;
  assign \piso.data_r [3972] = \piso.data_r_3972_sv2v_reg ;
  assign \piso.data_r [3971] = \piso.data_r_3971_sv2v_reg ;
  assign \piso.data_r [3970] = \piso.data_r_3970_sv2v_reg ;
  assign \piso.data_r [3969] = \piso.data_r_3969_sv2v_reg ;
  assign \piso.data_r [3968] = \piso.data_r_3968_sv2v_reg ;
  assign \piso.data_r [3967] = \piso.data_r_3967_sv2v_reg ;
  assign \piso.data_r [3966] = \piso.data_r_3966_sv2v_reg ;
  assign \piso.data_r [3965] = \piso.data_r_3965_sv2v_reg ;
  assign \piso.data_r [3964] = \piso.data_r_3964_sv2v_reg ;
  assign \piso.data_r [3963] = \piso.data_r_3963_sv2v_reg ;
  assign \piso.data_r [3962] = \piso.data_r_3962_sv2v_reg ;
  assign \piso.data_r [3961] = \piso.data_r_3961_sv2v_reg ;
  assign \piso.data_r [3960] = \piso.data_r_3960_sv2v_reg ;
  assign \piso.data_r [3959] = \piso.data_r_3959_sv2v_reg ;
  assign \piso.data_r [3958] = \piso.data_r_3958_sv2v_reg ;
  assign \piso.data_r [3957] = \piso.data_r_3957_sv2v_reg ;
  assign \piso.data_r [3956] = \piso.data_r_3956_sv2v_reg ;
  assign \piso.data_r [3955] = \piso.data_r_3955_sv2v_reg ;
  assign \piso.data_r [3954] = \piso.data_r_3954_sv2v_reg ;
  assign \piso.data_r [3953] = \piso.data_r_3953_sv2v_reg ;
  assign \piso.data_r [3952] = \piso.data_r_3952_sv2v_reg ;
  assign \piso.data_r [3951] = \piso.data_r_3951_sv2v_reg ;
  assign \piso.data_r [3950] = \piso.data_r_3950_sv2v_reg ;
  assign \piso.data_r [3949] = \piso.data_r_3949_sv2v_reg ;
  assign \piso.data_r [3948] = \piso.data_r_3948_sv2v_reg ;
  assign \piso.data_r [3947] = \piso.data_r_3947_sv2v_reg ;
  assign \piso.data_r [3946] = \piso.data_r_3946_sv2v_reg ;
  assign \piso.data_r [3945] = \piso.data_r_3945_sv2v_reg ;
  assign \piso.data_r [3944] = \piso.data_r_3944_sv2v_reg ;
  assign \piso.data_r [3943] = \piso.data_r_3943_sv2v_reg ;
  assign \piso.data_r [3942] = \piso.data_r_3942_sv2v_reg ;
  assign \piso.data_r [3941] = \piso.data_r_3941_sv2v_reg ;
  assign \piso.data_r [3940] = \piso.data_r_3940_sv2v_reg ;
  assign \piso.data_r [3939] = \piso.data_r_3939_sv2v_reg ;
  assign \piso.data_r [3938] = \piso.data_r_3938_sv2v_reg ;
  assign \piso.data_r [3937] = \piso.data_r_3937_sv2v_reg ;
  assign \piso.data_r [3936] = \piso.data_r_3936_sv2v_reg ;
  assign \piso.data_r [3935] = \piso.data_r_3935_sv2v_reg ;
  assign \piso.data_r [3934] = \piso.data_r_3934_sv2v_reg ;
  assign \piso.data_r [3933] = \piso.data_r_3933_sv2v_reg ;
  assign \piso.data_r [3932] = \piso.data_r_3932_sv2v_reg ;
  assign \piso.data_r [3931] = \piso.data_r_3931_sv2v_reg ;
  assign \piso.data_r [3930] = \piso.data_r_3930_sv2v_reg ;
  assign \piso.data_r [3929] = \piso.data_r_3929_sv2v_reg ;
  assign \piso.data_r [3928] = \piso.data_r_3928_sv2v_reg ;
  assign \piso.data_r [3927] = \piso.data_r_3927_sv2v_reg ;
  assign \piso.data_r [3926] = \piso.data_r_3926_sv2v_reg ;
  assign \piso.data_r [3925] = \piso.data_r_3925_sv2v_reg ;
  assign \piso.data_r [3924] = \piso.data_r_3924_sv2v_reg ;
  assign \piso.data_r [3923] = \piso.data_r_3923_sv2v_reg ;
  assign \piso.data_r [3922] = \piso.data_r_3922_sv2v_reg ;
  assign \piso.data_r [3921] = \piso.data_r_3921_sv2v_reg ;
  assign \piso.data_r [3920] = \piso.data_r_3920_sv2v_reg ;
  assign \piso.data_r [3919] = \piso.data_r_3919_sv2v_reg ;
  assign \piso.data_r [3918] = \piso.data_r_3918_sv2v_reg ;
  assign \piso.data_r [3917] = \piso.data_r_3917_sv2v_reg ;
  assign \piso.data_r [3916] = \piso.data_r_3916_sv2v_reg ;
  assign \piso.data_r [3915] = \piso.data_r_3915_sv2v_reg ;
  assign \piso.data_r [3914] = \piso.data_r_3914_sv2v_reg ;
  assign \piso.data_r [3913] = \piso.data_r_3913_sv2v_reg ;
  assign \piso.data_r [3912] = \piso.data_r_3912_sv2v_reg ;
  assign \piso.data_r [3911] = \piso.data_r_3911_sv2v_reg ;
  assign \piso.data_r [3910] = \piso.data_r_3910_sv2v_reg ;
  assign \piso.data_r [3909] = \piso.data_r_3909_sv2v_reg ;
  assign \piso.data_r [3908] = \piso.data_r_3908_sv2v_reg ;
  assign \piso.data_r [3907] = \piso.data_r_3907_sv2v_reg ;
  assign \piso.data_r [3906] = \piso.data_r_3906_sv2v_reg ;
  assign \piso.data_r [3905] = \piso.data_r_3905_sv2v_reg ;
  assign \piso.data_r [3904] = \piso.data_r_3904_sv2v_reg ;
  assign \piso.data_r [3903] = \piso.data_r_3903_sv2v_reg ;
  assign \piso.data_r [3902] = \piso.data_r_3902_sv2v_reg ;
  assign \piso.data_r [3901] = \piso.data_r_3901_sv2v_reg ;
  assign \piso.data_r [3900] = \piso.data_r_3900_sv2v_reg ;
  assign \piso.data_r [3899] = \piso.data_r_3899_sv2v_reg ;
  assign \piso.data_r [3898] = \piso.data_r_3898_sv2v_reg ;
  assign \piso.data_r [3897] = \piso.data_r_3897_sv2v_reg ;
  assign \piso.data_r [3896] = \piso.data_r_3896_sv2v_reg ;
  assign \piso.data_r [3895] = \piso.data_r_3895_sv2v_reg ;
  assign \piso.data_r [3894] = \piso.data_r_3894_sv2v_reg ;
  assign \piso.data_r [3893] = \piso.data_r_3893_sv2v_reg ;
  assign \piso.data_r [3892] = \piso.data_r_3892_sv2v_reg ;
  assign \piso.data_r [3891] = \piso.data_r_3891_sv2v_reg ;
  assign \piso.data_r [3890] = \piso.data_r_3890_sv2v_reg ;
  assign \piso.data_r [3889] = \piso.data_r_3889_sv2v_reg ;
  assign \piso.data_r [3888] = \piso.data_r_3888_sv2v_reg ;
  assign \piso.data_r [3887] = \piso.data_r_3887_sv2v_reg ;
  assign \piso.data_r [3886] = \piso.data_r_3886_sv2v_reg ;
  assign \piso.data_r [3885] = \piso.data_r_3885_sv2v_reg ;
  assign \piso.data_r [3884] = \piso.data_r_3884_sv2v_reg ;
  assign \piso.data_r [3883] = \piso.data_r_3883_sv2v_reg ;
  assign \piso.data_r [3882] = \piso.data_r_3882_sv2v_reg ;
  assign \piso.data_r [3881] = \piso.data_r_3881_sv2v_reg ;
  assign \piso.data_r [3880] = \piso.data_r_3880_sv2v_reg ;
  assign \piso.data_r [3879] = \piso.data_r_3879_sv2v_reg ;
  assign \piso.data_r [3878] = \piso.data_r_3878_sv2v_reg ;
  assign \piso.data_r [3877] = \piso.data_r_3877_sv2v_reg ;
  assign \piso.data_r [3876] = \piso.data_r_3876_sv2v_reg ;
  assign \piso.data_r [3875] = \piso.data_r_3875_sv2v_reg ;
  assign \piso.data_r [3874] = \piso.data_r_3874_sv2v_reg ;
  assign \piso.data_r [3873] = \piso.data_r_3873_sv2v_reg ;
  assign \piso.data_r [3872] = \piso.data_r_3872_sv2v_reg ;
  assign \piso.data_r [3871] = \piso.data_r_3871_sv2v_reg ;
  assign \piso.data_r [3870] = \piso.data_r_3870_sv2v_reg ;
  assign \piso.data_r [3869] = \piso.data_r_3869_sv2v_reg ;
  assign \piso.data_r [3868] = \piso.data_r_3868_sv2v_reg ;
  assign \piso.data_r [3867] = \piso.data_r_3867_sv2v_reg ;
  assign \piso.data_r [3866] = \piso.data_r_3866_sv2v_reg ;
  assign \piso.data_r [3865] = \piso.data_r_3865_sv2v_reg ;
  assign \piso.data_r [3864] = \piso.data_r_3864_sv2v_reg ;
  assign \piso.data_r [3863] = \piso.data_r_3863_sv2v_reg ;
  assign \piso.data_r [3862] = \piso.data_r_3862_sv2v_reg ;
  assign \piso.data_r [3861] = \piso.data_r_3861_sv2v_reg ;
  assign \piso.data_r [3860] = \piso.data_r_3860_sv2v_reg ;
  assign \piso.data_r [3859] = \piso.data_r_3859_sv2v_reg ;
  assign \piso.data_r [3858] = \piso.data_r_3858_sv2v_reg ;
  assign \piso.data_r [3857] = \piso.data_r_3857_sv2v_reg ;
  assign \piso.data_r [3856] = \piso.data_r_3856_sv2v_reg ;
  assign \piso.data_r [3855] = \piso.data_r_3855_sv2v_reg ;
  assign \piso.data_r [3854] = \piso.data_r_3854_sv2v_reg ;
  assign \piso.data_r [3853] = \piso.data_r_3853_sv2v_reg ;
  assign \piso.data_r [3852] = \piso.data_r_3852_sv2v_reg ;
  assign \piso.data_r [3851] = \piso.data_r_3851_sv2v_reg ;
  assign \piso.data_r [3850] = \piso.data_r_3850_sv2v_reg ;
  assign \piso.data_r [3849] = \piso.data_r_3849_sv2v_reg ;
  assign \piso.data_r [3848] = \piso.data_r_3848_sv2v_reg ;
  assign \piso.data_r [3847] = \piso.data_r_3847_sv2v_reg ;
  assign \piso.data_r [3846] = \piso.data_r_3846_sv2v_reg ;
  assign \piso.data_r [3845] = \piso.data_r_3845_sv2v_reg ;
  assign \piso.data_r [3844] = \piso.data_r_3844_sv2v_reg ;
  assign \piso.data_r [3843] = \piso.data_r_3843_sv2v_reg ;
  assign \piso.data_r [3842] = \piso.data_r_3842_sv2v_reg ;
  assign \piso.data_r [3841] = \piso.data_r_3841_sv2v_reg ;
  assign \piso.data_r [3840] = \piso.data_r_3840_sv2v_reg ;
  assign \piso.data_r [3839] = \piso.data_r_3839_sv2v_reg ;
  assign \piso.data_r [3838] = \piso.data_r_3838_sv2v_reg ;
  assign \piso.data_r [3837] = \piso.data_r_3837_sv2v_reg ;
  assign \piso.data_r [3836] = \piso.data_r_3836_sv2v_reg ;
  assign \piso.data_r [3835] = \piso.data_r_3835_sv2v_reg ;
  assign \piso.data_r [3834] = \piso.data_r_3834_sv2v_reg ;
  assign \piso.data_r [3833] = \piso.data_r_3833_sv2v_reg ;
  assign \piso.data_r [3832] = \piso.data_r_3832_sv2v_reg ;
  assign \piso.data_r [3831] = \piso.data_r_3831_sv2v_reg ;
  assign \piso.data_r [3830] = \piso.data_r_3830_sv2v_reg ;
  assign \piso.data_r [3829] = \piso.data_r_3829_sv2v_reg ;
  assign \piso.data_r [3828] = \piso.data_r_3828_sv2v_reg ;
  assign \piso.data_r [3827] = \piso.data_r_3827_sv2v_reg ;
  assign \piso.data_r [3826] = \piso.data_r_3826_sv2v_reg ;
  assign \piso.data_r [3825] = \piso.data_r_3825_sv2v_reg ;
  assign \piso.data_r [3824] = \piso.data_r_3824_sv2v_reg ;
  assign \piso.data_r [3823] = \piso.data_r_3823_sv2v_reg ;
  assign \piso.data_r [3822] = \piso.data_r_3822_sv2v_reg ;
  assign \piso.data_r [3821] = \piso.data_r_3821_sv2v_reg ;
  assign \piso.data_r [3820] = \piso.data_r_3820_sv2v_reg ;
  assign \piso.data_r [3819] = \piso.data_r_3819_sv2v_reg ;
  assign \piso.data_r [3818] = \piso.data_r_3818_sv2v_reg ;
  assign \piso.data_r [3817] = \piso.data_r_3817_sv2v_reg ;
  assign \piso.data_r [3816] = \piso.data_r_3816_sv2v_reg ;
  assign \piso.data_r [3815] = \piso.data_r_3815_sv2v_reg ;
  assign \piso.data_r [3814] = \piso.data_r_3814_sv2v_reg ;
  assign \piso.data_r [3813] = \piso.data_r_3813_sv2v_reg ;
  assign \piso.data_r [3812] = \piso.data_r_3812_sv2v_reg ;
  assign \piso.data_r [3811] = \piso.data_r_3811_sv2v_reg ;
  assign \piso.data_r [3810] = \piso.data_r_3810_sv2v_reg ;
  assign \piso.data_r [3809] = \piso.data_r_3809_sv2v_reg ;
  assign \piso.data_r [3808] = \piso.data_r_3808_sv2v_reg ;
  assign \piso.data_r [3807] = \piso.data_r_3807_sv2v_reg ;
  assign \piso.data_r [3806] = \piso.data_r_3806_sv2v_reg ;
  assign \piso.data_r [3805] = \piso.data_r_3805_sv2v_reg ;
  assign \piso.data_r [3804] = \piso.data_r_3804_sv2v_reg ;
  assign \piso.data_r [3803] = \piso.data_r_3803_sv2v_reg ;
  assign \piso.data_r [3802] = \piso.data_r_3802_sv2v_reg ;
  assign \piso.data_r [3801] = \piso.data_r_3801_sv2v_reg ;
  assign \piso.data_r [3800] = \piso.data_r_3800_sv2v_reg ;
  assign \piso.data_r [3799] = \piso.data_r_3799_sv2v_reg ;
  assign \piso.data_r [3798] = \piso.data_r_3798_sv2v_reg ;
  assign \piso.data_r [3797] = \piso.data_r_3797_sv2v_reg ;
  assign \piso.data_r [3796] = \piso.data_r_3796_sv2v_reg ;
  assign \piso.data_r [3795] = \piso.data_r_3795_sv2v_reg ;
  assign \piso.data_r [3794] = \piso.data_r_3794_sv2v_reg ;
  assign \piso.data_r [3793] = \piso.data_r_3793_sv2v_reg ;
  assign \piso.data_r [3792] = \piso.data_r_3792_sv2v_reg ;
  assign \piso.data_r [3791] = \piso.data_r_3791_sv2v_reg ;
  assign \piso.data_r [3790] = \piso.data_r_3790_sv2v_reg ;
  assign \piso.data_r [3789] = \piso.data_r_3789_sv2v_reg ;
  assign \piso.data_r [3788] = \piso.data_r_3788_sv2v_reg ;
  assign \piso.data_r [3787] = \piso.data_r_3787_sv2v_reg ;
  assign \piso.data_r [3786] = \piso.data_r_3786_sv2v_reg ;
  assign \piso.data_r [3785] = \piso.data_r_3785_sv2v_reg ;
  assign \piso.data_r [3784] = \piso.data_r_3784_sv2v_reg ;
  assign \piso.data_r [3783] = \piso.data_r_3783_sv2v_reg ;
  assign \piso.data_r [3782] = \piso.data_r_3782_sv2v_reg ;
  assign \piso.data_r [3781] = \piso.data_r_3781_sv2v_reg ;
  assign \piso.data_r [3780] = \piso.data_r_3780_sv2v_reg ;
  assign \piso.data_r [3779] = \piso.data_r_3779_sv2v_reg ;
  assign \piso.data_r [3778] = \piso.data_r_3778_sv2v_reg ;
  assign \piso.data_r [3777] = \piso.data_r_3777_sv2v_reg ;
  assign \piso.data_r [3776] = \piso.data_r_3776_sv2v_reg ;
  assign \piso.data_r [3775] = \piso.data_r_3775_sv2v_reg ;
  assign \piso.data_r [3774] = \piso.data_r_3774_sv2v_reg ;
  assign \piso.data_r [3773] = \piso.data_r_3773_sv2v_reg ;
  assign \piso.data_r [3772] = \piso.data_r_3772_sv2v_reg ;
  assign \piso.data_r [3771] = \piso.data_r_3771_sv2v_reg ;
  assign \piso.data_r [3770] = \piso.data_r_3770_sv2v_reg ;
  assign \piso.data_r [3769] = \piso.data_r_3769_sv2v_reg ;
  assign \piso.data_r [3768] = \piso.data_r_3768_sv2v_reg ;
  assign \piso.data_r [3767] = \piso.data_r_3767_sv2v_reg ;
  assign \piso.data_r [3766] = \piso.data_r_3766_sv2v_reg ;
  assign \piso.data_r [3765] = \piso.data_r_3765_sv2v_reg ;
  assign \piso.data_r [3764] = \piso.data_r_3764_sv2v_reg ;
  assign \piso.data_r [3763] = \piso.data_r_3763_sv2v_reg ;
  assign \piso.data_r [3762] = \piso.data_r_3762_sv2v_reg ;
  assign \piso.data_r [3761] = \piso.data_r_3761_sv2v_reg ;
  assign \piso.data_r [3760] = \piso.data_r_3760_sv2v_reg ;
  assign \piso.data_r [3759] = \piso.data_r_3759_sv2v_reg ;
  assign \piso.data_r [3758] = \piso.data_r_3758_sv2v_reg ;
  assign \piso.data_r [3757] = \piso.data_r_3757_sv2v_reg ;
  assign \piso.data_r [3756] = \piso.data_r_3756_sv2v_reg ;
  assign \piso.data_r [3755] = \piso.data_r_3755_sv2v_reg ;
  assign \piso.data_r [3754] = \piso.data_r_3754_sv2v_reg ;
  assign \piso.data_r [3753] = \piso.data_r_3753_sv2v_reg ;
  assign \piso.data_r [3752] = \piso.data_r_3752_sv2v_reg ;
  assign \piso.data_r [3751] = \piso.data_r_3751_sv2v_reg ;
  assign \piso.data_r [3750] = \piso.data_r_3750_sv2v_reg ;
  assign \piso.data_r [3749] = \piso.data_r_3749_sv2v_reg ;
  assign \piso.data_r [3748] = \piso.data_r_3748_sv2v_reg ;
  assign \piso.data_r [3747] = \piso.data_r_3747_sv2v_reg ;
  assign \piso.data_r [3746] = \piso.data_r_3746_sv2v_reg ;
  assign \piso.data_r [3745] = \piso.data_r_3745_sv2v_reg ;
  assign \piso.data_r [3744] = \piso.data_r_3744_sv2v_reg ;
  assign \piso.data_r [3743] = \piso.data_r_3743_sv2v_reg ;
  assign \piso.data_r [3742] = \piso.data_r_3742_sv2v_reg ;
  assign \piso.data_r [3741] = \piso.data_r_3741_sv2v_reg ;
  assign \piso.data_r [3740] = \piso.data_r_3740_sv2v_reg ;
  assign \piso.data_r [3739] = \piso.data_r_3739_sv2v_reg ;
  assign \piso.data_r [3738] = \piso.data_r_3738_sv2v_reg ;
  assign \piso.data_r [3737] = \piso.data_r_3737_sv2v_reg ;
  assign \piso.data_r [3736] = \piso.data_r_3736_sv2v_reg ;
  assign \piso.data_r [3735] = \piso.data_r_3735_sv2v_reg ;
  assign \piso.data_r [3734] = \piso.data_r_3734_sv2v_reg ;
  assign \piso.data_r [3733] = \piso.data_r_3733_sv2v_reg ;
  assign \piso.data_r [3732] = \piso.data_r_3732_sv2v_reg ;
  assign \piso.data_r [3731] = \piso.data_r_3731_sv2v_reg ;
  assign \piso.data_r [3730] = \piso.data_r_3730_sv2v_reg ;
  assign \piso.data_r [3729] = \piso.data_r_3729_sv2v_reg ;
  assign \piso.data_r [3728] = \piso.data_r_3728_sv2v_reg ;
  assign \piso.data_r [3727] = \piso.data_r_3727_sv2v_reg ;
  assign \piso.data_r [3726] = \piso.data_r_3726_sv2v_reg ;
  assign \piso.data_r [3725] = \piso.data_r_3725_sv2v_reg ;
  assign \piso.data_r [3724] = \piso.data_r_3724_sv2v_reg ;
  assign \piso.data_r [3723] = \piso.data_r_3723_sv2v_reg ;
  assign \piso.data_r [3722] = \piso.data_r_3722_sv2v_reg ;
  assign \piso.data_r [3721] = \piso.data_r_3721_sv2v_reg ;
  assign \piso.data_r [3720] = \piso.data_r_3720_sv2v_reg ;
  assign \piso.data_r [3719] = \piso.data_r_3719_sv2v_reg ;
  assign \piso.data_r [3718] = \piso.data_r_3718_sv2v_reg ;
  assign \piso.data_r [3717] = \piso.data_r_3717_sv2v_reg ;
  assign \piso.data_r [3716] = \piso.data_r_3716_sv2v_reg ;
  assign \piso.data_r [3715] = \piso.data_r_3715_sv2v_reg ;
  assign \piso.data_r [3714] = \piso.data_r_3714_sv2v_reg ;
  assign \piso.data_r [3713] = \piso.data_r_3713_sv2v_reg ;
  assign \piso.data_r [3712] = \piso.data_r_3712_sv2v_reg ;
  assign \piso.data_r [3711] = \piso.data_r_3711_sv2v_reg ;
  assign \piso.data_r [3710] = \piso.data_r_3710_sv2v_reg ;
  assign \piso.data_r [3709] = \piso.data_r_3709_sv2v_reg ;
  assign \piso.data_r [3708] = \piso.data_r_3708_sv2v_reg ;
  assign \piso.data_r [3707] = \piso.data_r_3707_sv2v_reg ;
  assign \piso.data_r [3706] = \piso.data_r_3706_sv2v_reg ;
  assign \piso.data_r [3705] = \piso.data_r_3705_sv2v_reg ;
  assign \piso.data_r [3704] = \piso.data_r_3704_sv2v_reg ;
  assign \piso.data_r [3703] = \piso.data_r_3703_sv2v_reg ;
  assign \piso.data_r [3702] = \piso.data_r_3702_sv2v_reg ;
  assign \piso.data_r [3701] = \piso.data_r_3701_sv2v_reg ;
  assign \piso.data_r [3700] = \piso.data_r_3700_sv2v_reg ;
  assign \piso.data_r [3699] = \piso.data_r_3699_sv2v_reg ;
  assign \piso.data_r [3698] = \piso.data_r_3698_sv2v_reg ;
  assign \piso.data_r [3697] = \piso.data_r_3697_sv2v_reg ;
  assign \piso.data_r [3696] = \piso.data_r_3696_sv2v_reg ;
  assign \piso.data_r [3695] = \piso.data_r_3695_sv2v_reg ;
  assign \piso.data_r [3694] = \piso.data_r_3694_sv2v_reg ;
  assign \piso.data_r [3693] = \piso.data_r_3693_sv2v_reg ;
  assign \piso.data_r [3692] = \piso.data_r_3692_sv2v_reg ;
  assign \piso.data_r [3691] = \piso.data_r_3691_sv2v_reg ;
  assign \piso.data_r [3690] = \piso.data_r_3690_sv2v_reg ;
  assign \piso.data_r [3689] = \piso.data_r_3689_sv2v_reg ;
  assign \piso.data_r [3688] = \piso.data_r_3688_sv2v_reg ;
  assign \piso.data_r [3687] = \piso.data_r_3687_sv2v_reg ;
  assign \piso.data_r [3686] = \piso.data_r_3686_sv2v_reg ;
  assign \piso.data_r [3685] = \piso.data_r_3685_sv2v_reg ;
  assign \piso.data_r [3684] = \piso.data_r_3684_sv2v_reg ;
  assign \piso.data_r [3683] = \piso.data_r_3683_sv2v_reg ;
  assign \piso.data_r [3682] = \piso.data_r_3682_sv2v_reg ;
  assign \piso.data_r [3681] = \piso.data_r_3681_sv2v_reg ;
  assign \piso.data_r [3680] = \piso.data_r_3680_sv2v_reg ;
  assign \piso.data_r [3679] = \piso.data_r_3679_sv2v_reg ;
  assign \piso.data_r [3678] = \piso.data_r_3678_sv2v_reg ;
  assign \piso.data_r [3677] = \piso.data_r_3677_sv2v_reg ;
  assign \piso.data_r [3676] = \piso.data_r_3676_sv2v_reg ;
  assign \piso.data_r [3675] = \piso.data_r_3675_sv2v_reg ;
  assign \piso.data_r [3674] = \piso.data_r_3674_sv2v_reg ;
  assign \piso.data_r [3673] = \piso.data_r_3673_sv2v_reg ;
  assign \piso.data_r [3672] = \piso.data_r_3672_sv2v_reg ;
  assign \piso.data_r [3671] = \piso.data_r_3671_sv2v_reg ;
  assign \piso.data_r [3670] = \piso.data_r_3670_sv2v_reg ;
  assign \piso.data_r [3669] = \piso.data_r_3669_sv2v_reg ;
  assign \piso.data_r [3668] = \piso.data_r_3668_sv2v_reg ;
  assign \piso.data_r [3667] = \piso.data_r_3667_sv2v_reg ;
  assign \piso.data_r [3666] = \piso.data_r_3666_sv2v_reg ;
  assign \piso.data_r [3665] = \piso.data_r_3665_sv2v_reg ;
  assign \piso.data_r [3664] = \piso.data_r_3664_sv2v_reg ;
  assign \piso.data_r [3663] = \piso.data_r_3663_sv2v_reg ;
  assign \piso.data_r [3662] = \piso.data_r_3662_sv2v_reg ;
  assign \piso.data_r [3661] = \piso.data_r_3661_sv2v_reg ;
  assign \piso.data_r [3660] = \piso.data_r_3660_sv2v_reg ;
  assign \piso.data_r [3659] = \piso.data_r_3659_sv2v_reg ;
  assign \piso.data_r [3658] = \piso.data_r_3658_sv2v_reg ;
  assign \piso.data_r [3657] = \piso.data_r_3657_sv2v_reg ;
  assign \piso.data_r [3656] = \piso.data_r_3656_sv2v_reg ;
  assign \piso.data_r [3655] = \piso.data_r_3655_sv2v_reg ;
  assign \piso.data_r [3654] = \piso.data_r_3654_sv2v_reg ;
  assign \piso.data_r [3653] = \piso.data_r_3653_sv2v_reg ;
  assign \piso.data_r [3652] = \piso.data_r_3652_sv2v_reg ;
  assign \piso.data_r [3651] = \piso.data_r_3651_sv2v_reg ;
  assign \piso.data_r [3650] = \piso.data_r_3650_sv2v_reg ;
  assign \piso.data_r [3649] = \piso.data_r_3649_sv2v_reg ;
  assign \piso.data_r [3648] = \piso.data_r_3648_sv2v_reg ;
  assign \piso.data_r [3647] = \piso.data_r_3647_sv2v_reg ;
  assign \piso.data_r [3646] = \piso.data_r_3646_sv2v_reg ;
  assign \piso.data_r [3645] = \piso.data_r_3645_sv2v_reg ;
  assign \piso.data_r [3644] = \piso.data_r_3644_sv2v_reg ;
  assign \piso.data_r [3643] = \piso.data_r_3643_sv2v_reg ;
  assign \piso.data_r [3642] = \piso.data_r_3642_sv2v_reg ;
  assign \piso.data_r [3641] = \piso.data_r_3641_sv2v_reg ;
  assign \piso.data_r [3640] = \piso.data_r_3640_sv2v_reg ;
  assign \piso.data_r [3639] = \piso.data_r_3639_sv2v_reg ;
  assign \piso.data_r [3638] = \piso.data_r_3638_sv2v_reg ;
  assign \piso.data_r [3637] = \piso.data_r_3637_sv2v_reg ;
  assign \piso.data_r [3636] = \piso.data_r_3636_sv2v_reg ;
  assign \piso.data_r [3635] = \piso.data_r_3635_sv2v_reg ;
  assign \piso.data_r [3634] = \piso.data_r_3634_sv2v_reg ;
  assign \piso.data_r [3633] = \piso.data_r_3633_sv2v_reg ;
  assign \piso.data_r [3632] = \piso.data_r_3632_sv2v_reg ;
  assign \piso.data_r [3631] = \piso.data_r_3631_sv2v_reg ;
  assign \piso.data_r [3630] = \piso.data_r_3630_sv2v_reg ;
  assign \piso.data_r [3629] = \piso.data_r_3629_sv2v_reg ;
  assign \piso.data_r [3628] = \piso.data_r_3628_sv2v_reg ;
  assign \piso.data_r [3627] = \piso.data_r_3627_sv2v_reg ;
  assign \piso.data_r [3626] = \piso.data_r_3626_sv2v_reg ;
  assign \piso.data_r [3625] = \piso.data_r_3625_sv2v_reg ;
  assign \piso.data_r [3624] = \piso.data_r_3624_sv2v_reg ;
  assign \piso.data_r [3623] = \piso.data_r_3623_sv2v_reg ;
  assign \piso.data_r [3622] = \piso.data_r_3622_sv2v_reg ;
  assign \piso.data_r [3621] = \piso.data_r_3621_sv2v_reg ;
  assign \piso.data_r [3620] = \piso.data_r_3620_sv2v_reg ;
  assign \piso.data_r [3619] = \piso.data_r_3619_sv2v_reg ;
  assign \piso.data_r [3618] = \piso.data_r_3618_sv2v_reg ;
  assign \piso.data_r [3617] = \piso.data_r_3617_sv2v_reg ;
  assign \piso.data_r [3616] = \piso.data_r_3616_sv2v_reg ;
  assign \piso.data_r [3615] = \piso.data_r_3615_sv2v_reg ;
  assign \piso.data_r [3614] = \piso.data_r_3614_sv2v_reg ;
  assign \piso.data_r [3613] = \piso.data_r_3613_sv2v_reg ;
  assign \piso.data_r [3612] = \piso.data_r_3612_sv2v_reg ;
  assign \piso.data_r [3611] = \piso.data_r_3611_sv2v_reg ;
  assign \piso.data_r [3610] = \piso.data_r_3610_sv2v_reg ;
  assign \piso.data_r [3609] = \piso.data_r_3609_sv2v_reg ;
  assign \piso.data_r [3608] = \piso.data_r_3608_sv2v_reg ;
  assign \piso.data_r [3607] = \piso.data_r_3607_sv2v_reg ;
  assign \piso.data_r [3606] = \piso.data_r_3606_sv2v_reg ;
  assign \piso.data_r [3605] = \piso.data_r_3605_sv2v_reg ;
  assign \piso.data_r [3604] = \piso.data_r_3604_sv2v_reg ;
  assign \piso.data_r [3603] = \piso.data_r_3603_sv2v_reg ;
  assign \piso.data_r [3602] = \piso.data_r_3602_sv2v_reg ;
  assign \piso.data_r [3601] = \piso.data_r_3601_sv2v_reg ;
  assign \piso.data_r [3600] = \piso.data_r_3600_sv2v_reg ;
  assign \piso.data_r [3599] = \piso.data_r_3599_sv2v_reg ;
  assign \piso.data_r [3598] = \piso.data_r_3598_sv2v_reg ;
  assign \piso.data_r [3597] = \piso.data_r_3597_sv2v_reg ;
  assign \piso.data_r [3596] = \piso.data_r_3596_sv2v_reg ;
  assign \piso.data_r [3595] = \piso.data_r_3595_sv2v_reg ;
  assign \piso.data_r [3594] = \piso.data_r_3594_sv2v_reg ;
  assign \piso.data_r [3593] = \piso.data_r_3593_sv2v_reg ;
  assign \piso.data_r [3592] = \piso.data_r_3592_sv2v_reg ;
  assign \piso.data_r [3591] = \piso.data_r_3591_sv2v_reg ;
  assign \piso.data_r [3590] = \piso.data_r_3590_sv2v_reg ;
  assign \piso.data_r [3589] = \piso.data_r_3589_sv2v_reg ;
  assign \piso.data_r [3588] = \piso.data_r_3588_sv2v_reg ;
  assign \piso.data_r [3587] = \piso.data_r_3587_sv2v_reg ;
  assign \piso.data_r [3586] = \piso.data_r_3586_sv2v_reg ;
  assign \piso.data_r [3585] = \piso.data_r_3585_sv2v_reg ;
  assign \piso.data_r [3584] = \piso.data_r_3584_sv2v_reg ;
  assign \piso.data_r [3583] = \piso.data_r_3583_sv2v_reg ;
  assign \piso.data_r [3582] = \piso.data_r_3582_sv2v_reg ;
  assign \piso.data_r [3581] = \piso.data_r_3581_sv2v_reg ;
  assign \piso.data_r [3580] = \piso.data_r_3580_sv2v_reg ;
  assign \piso.data_r [3579] = \piso.data_r_3579_sv2v_reg ;
  assign \piso.data_r [3578] = \piso.data_r_3578_sv2v_reg ;
  assign \piso.data_r [3577] = \piso.data_r_3577_sv2v_reg ;
  assign \piso.data_r [3576] = \piso.data_r_3576_sv2v_reg ;
  assign \piso.data_r [3575] = \piso.data_r_3575_sv2v_reg ;
  assign \piso.data_r [3574] = \piso.data_r_3574_sv2v_reg ;
  assign \piso.data_r [3573] = \piso.data_r_3573_sv2v_reg ;
  assign \piso.data_r [3572] = \piso.data_r_3572_sv2v_reg ;
  assign \piso.data_r [3571] = \piso.data_r_3571_sv2v_reg ;
  assign \piso.data_r [3570] = \piso.data_r_3570_sv2v_reg ;
  assign \piso.data_r [3569] = \piso.data_r_3569_sv2v_reg ;
  assign \piso.data_r [3568] = \piso.data_r_3568_sv2v_reg ;
  assign \piso.data_r [3567] = \piso.data_r_3567_sv2v_reg ;
  assign \piso.data_r [3566] = \piso.data_r_3566_sv2v_reg ;
  assign \piso.data_r [3565] = \piso.data_r_3565_sv2v_reg ;
  assign \piso.data_r [3564] = \piso.data_r_3564_sv2v_reg ;
  assign \piso.data_r [3563] = \piso.data_r_3563_sv2v_reg ;
  assign \piso.data_r [3562] = \piso.data_r_3562_sv2v_reg ;
  assign \piso.data_r [3561] = \piso.data_r_3561_sv2v_reg ;
  assign \piso.data_r [3560] = \piso.data_r_3560_sv2v_reg ;
  assign \piso.data_r [3559] = \piso.data_r_3559_sv2v_reg ;
  assign \piso.data_r [3558] = \piso.data_r_3558_sv2v_reg ;
  assign \piso.data_r [3557] = \piso.data_r_3557_sv2v_reg ;
  assign \piso.data_r [3556] = \piso.data_r_3556_sv2v_reg ;
  assign \piso.data_r [3555] = \piso.data_r_3555_sv2v_reg ;
  assign \piso.data_r [3554] = \piso.data_r_3554_sv2v_reg ;
  assign \piso.data_r [3553] = \piso.data_r_3553_sv2v_reg ;
  assign \piso.data_r [3552] = \piso.data_r_3552_sv2v_reg ;
  assign \piso.data_r [3551] = \piso.data_r_3551_sv2v_reg ;
  assign \piso.data_r [3550] = \piso.data_r_3550_sv2v_reg ;
  assign \piso.data_r [3549] = \piso.data_r_3549_sv2v_reg ;
  assign \piso.data_r [3548] = \piso.data_r_3548_sv2v_reg ;
  assign \piso.data_r [3547] = \piso.data_r_3547_sv2v_reg ;
  assign \piso.data_r [3546] = \piso.data_r_3546_sv2v_reg ;
  assign \piso.data_r [3545] = \piso.data_r_3545_sv2v_reg ;
  assign \piso.data_r [3544] = \piso.data_r_3544_sv2v_reg ;
  assign \piso.data_r [3543] = \piso.data_r_3543_sv2v_reg ;
  assign \piso.data_r [3542] = \piso.data_r_3542_sv2v_reg ;
  assign \piso.data_r [3541] = \piso.data_r_3541_sv2v_reg ;
  assign \piso.data_r [3540] = \piso.data_r_3540_sv2v_reg ;
  assign \piso.data_r [3539] = \piso.data_r_3539_sv2v_reg ;
  assign \piso.data_r [3538] = \piso.data_r_3538_sv2v_reg ;
  assign \piso.data_r [3537] = \piso.data_r_3537_sv2v_reg ;
  assign \piso.data_r [3536] = \piso.data_r_3536_sv2v_reg ;
  assign \piso.data_r [3535] = \piso.data_r_3535_sv2v_reg ;
  assign \piso.data_r [3534] = \piso.data_r_3534_sv2v_reg ;
  assign \piso.data_r [3533] = \piso.data_r_3533_sv2v_reg ;
  assign \piso.data_r [3532] = \piso.data_r_3532_sv2v_reg ;
  assign \piso.data_r [3531] = \piso.data_r_3531_sv2v_reg ;
  assign \piso.data_r [3530] = \piso.data_r_3530_sv2v_reg ;
  assign \piso.data_r [3529] = \piso.data_r_3529_sv2v_reg ;
  assign \piso.data_r [3528] = \piso.data_r_3528_sv2v_reg ;
  assign \piso.data_r [3527] = \piso.data_r_3527_sv2v_reg ;
  assign \piso.data_r [3526] = \piso.data_r_3526_sv2v_reg ;
  assign \piso.data_r [3525] = \piso.data_r_3525_sv2v_reg ;
  assign \piso.data_r [3524] = \piso.data_r_3524_sv2v_reg ;
  assign \piso.data_r [3523] = \piso.data_r_3523_sv2v_reg ;
  assign \piso.data_r [3522] = \piso.data_r_3522_sv2v_reg ;
  assign \piso.data_r [3521] = \piso.data_r_3521_sv2v_reg ;
  assign \piso.data_r [3520] = \piso.data_r_3520_sv2v_reg ;
  assign \piso.data_r [3519] = \piso.data_r_3519_sv2v_reg ;
  assign \piso.data_r [3518] = \piso.data_r_3518_sv2v_reg ;
  assign \piso.data_r [3517] = \piso.data_r_3517_sv2v_reg ;
  assign \piso.data_r [3516] = \piso.data_r_3516_sv2v_reg ;
  assign \piso.data_r [3515] = \piso.data_r_3515_sv2v_reg ;
  assign \piso.data_r [3514] = \piso.data_r_3514_sv2v_reg ;
  assign \piso.data_r [3513] = \piso.data_r_3513_sv2v_reg ;
  assign \piso.data_r [3512] = \piso.data_r_3512_sv2v_reg ;
  assign \piso.data_r [3511] = \piso.data_r_3511_sv2v_reg ;
  assign \piso.data_r [3510] = \piso.data_r_3510_sv2v_reg ;
  assign \piso.data_r [3509] = \piso.data_r_3509_sv2v_reg ;
  assign \piso.data_r [3508] = \piso.data_r_3508_sv2v_reg ;
  assign \piso.data_r [3507] = \piso.data_r_3507_sv2v_reg ;
  assign \piso.data_r [3506] = \piso.data_r_3506_sv2v_reg ;
  assign \piso.data_r [3505] = \piso.data_r_3505_sv2v_reg ;
  assign \piso.data_r [3504] = \piso.data_r_3504_sv2v_reg ;
  assign \piso.data_r [3503] = \piso.data_r_3503_sv2v_reg ;
  assign \piso.data_r [3502] = \piso.data_r_3502_sv2v_reg ;
  assign \piso.data_r [3501] = \piso.data_r_3501_sv2v_reg ;
  assign \piso.data_r [3500] = \piso.data_r_3500_sv2v_reg ;
  assign \piso.data_r [3499] = \piso.data_r_3499_sv2v_reg ;
  assign \piso.data_r [3498] = \piso.data_r_3498_sv2v_reg ;
  assign \piso.data_r [3497] = \piso.data_r_3497_sv2v_reg ;
  assign \piso.data_r [3496] = \piso.data_r_3496_sv2v_reg ;
  assign \piso.data_r [3495] = \piso.data_r_3495_sv2v_reg ;
  assign \piso.data_r [3494] = \piso.data_r_3494_sv2v_reg ;
  assign \piso.data_r [3493] = \piso.data_r_3493_sv2v_reg ;
  assign \piso.data_r [3492] = \piso.data_r_3492_sv2v_reg ;
  assign \piso.data_r [3491] = \piso.data_r_3491_sv2v_reg ;
  assign \piso.data_r [3490] = \piso.data_r_3490_sv2v_reg ;
  assign \piso.data_r [3489] = \piso.data_r_3489_sv2v_reg ;
  assign \piso.data_r [3488] = \piso.data_r_3488_sv2v_reg ;
  assign \piso.data_r [3487] = \piso.data_r_3487_sv2v_reg ;
  assign \piso.data_r [3486] = \piso.data_r_3486_sv2v_reg ;
  assign \piso.data_r [3485] = \piso.data_r_3485_sv2v_reg ;
  assign \piso.data_r [3484] = \piso.data_r_3484_sv2v_reg ;
  assign \piso.data_r [3483] = \piso.data_r_3483_sv2v_reg ;
  assign \piso.data_r [3482] = \piso.data_r_3482_sv2v_reg ;
  assign \piso.data_r [3481] = \piso.data_r_3481_sv2v_reg ;
  assign \piso.data_r [3480] = \piso.data_r_3480_sv2v_reg ;
  assign \piso.data_r [3479] = \piso.data_r_3479_sv2v_reg ;
  assign \piso.data_r [3478] = \piso.data_r_3478_sv2v_reg ;
  assign \piso.data_r [3477] = \piso.data_r_3477_sv2v_reg ;
  assign \piso.data_r [3476] = \piso.data_r_3476_sv2v_reg ;
  assign \piso.data_r [3475] = \piso.data_r_3475_sv2v_reg ;
  assign \piso.data_r [3474] = \piso.data_r_3474_sv2v_reg ;
  assign \piso.data_r [3473] = \piso.data_r_3473_sv2v_reg ;
  assign \piso.data_r [3472] = \piso.data_r_3472_sv2v_reg ;
  assign \piso.data_r [3471] = \piso.data_r_3471_sv2v_reg ;
  assign \piso.data_r [3470] = \piso.data_r_3470_sv2v_reg ;
  assign \piso.data_r [3469] = \piso.data_r_3469_sv2v_reg ;
  assign \piso.data_r [3468] = \piso.data_r_3468_sv2v_reg ;
  assign \piso.data_r [3467] = \piso.data_r_3467_sv2v_reg ;
  assign \piso.data_r [3466] = \piso.data_r_3466_sv2v_reg ;
  assign \piso.data_r [3465] = \piso.data_r_3465_sv2v_reg ;
  assign \piso.data_r [3464] = \piso.data_r_3464_sv2v_reg ;
  assign \piso.data_r [3463] = \piso.data_r_3463_sv2v_reg ;
  assign \piso.data_r [3462] = \piso.data_r_3462_sv2v_reg ;
  assign \piso.data_r [3461] = \piso.data_r_3461_sv2v_reg ;
  assign \piso.data_r [3460] = \piso.data_r_3460_sv2v_reg ;
  assign \piso.data_r [3459] = \piso.data_r_3459_sv2v_reg ;
  assign \piso.data_r [3458] = \piso.data_r_3458_sv2v_reg ;
  assign \piso.data_r [3457] = \piso.data_r_3457_sv2v_reg ;
  assign \piso.data_r [3456] = \piso.data_r_3456_sv2v_reg ;
  assign \piso.data_r [3455] = \piso.data_r_3455_sv2v_reg ;
  assign \piso.data_r [3454] = \piso.data_r_3454_sv2v_reg ;
  assign \piso.data_r [3453] = \piso.data_r_3453_sv2v_reg ;
  assign \piso.data_r [3452] = \piso.data_r_3452_sv2v_reg ;
  assign \piso.data_r [3451] = \piso.data_r_3451_sv2v_reg ;
  assign \piso.data_r [3450] = \piso.data_r_3450_sv2v_reg ;
  assign \piso.data_r [3449] = \piso.data_r_3449_sv2v_reg ;
  assign \piso.data_r [3448] = \piso.data_r_3448_sv2v_reg ;
  assign \piso.data_r [3447] = \piso.data_r_3447_sv2v_reg ;
  assign \piso.data_r [3446] = \piso.data_r_3446_sv2v_reg ;
  assign \piso.data_r [3445] = \piso.data_r_3445_sv2v_reg ;
  assign \piso.data_r [3444] = \piso.data_r_3444_sv2v_reg ;
  assign \piso.data_r [3443] = \piso.data_r_3443_sv2v_reg ;
  assign \piso.data_r [3442] = \piso.data_r_3442_sv2v_reg ;
  assign \piso.data_r [3441] = \piso.data_r_3441_sv2v_reg ;
  assign \piso.data_r [3440] = \piso.data_r_3440_sv2v_reg ;
  assign \piso.data_r [3439] = \piso.data_r_3439_sv2v_reg ;
  assign \piso.data_r [3438] = \piso.data_r_3438_sv2v_reg ;
  assign \piso.data_r [3437] = \piso.data_r_3437_sv2v_reg ;
  assign \piso.data_r [3436] = \piso.data_r_3436_sv2v_reg ;
  assign \piso.data_r [3435] = \piso.data_r_3435_sv2v_reg ;
  assign \piso.data_r [3434] = \piso.data_r_3434_sv2v_reg ;
  assign \piso.data_r [3433] = \piso.data_r_3433_sv2v_reg ;
  assign \piso.data_r [3432] = \piso.data_r_3432_sv2v_reg ;
  assign \piso.data_r [3431] = \piso.data_r_3431_sv2v_reg ;
  assign \piso.data_r [3430] = \piso.data_r_3430_sv2v_reg ;
  assign \piso.data_r [3429] = \piso.data_r_3429_sv2v_reg ;
  assign \piso.data_r [3428] = \piso.data_r_3428_sv2v_reg ;
  assign \piso.data_r [3427] = \piso.data_r_3427_sv2v_reg ;
  assign \piso.data_r [3426] = \piso.data_r_3426_sv2v_reg ;
  assign \piso.data_r [3425] = \piso.data_r_3425_sv2v_reg ;
  assign \piso.data_r [3424] = \piso.data_r_3424_sv2v_reg ;
  assign \piso.data_r [3423] = \piso.data_r_3423_sv2v_reg ;
  assign \piso.data_r [3422] = \piso.data_r_3422_sv2v_reg ;
  assign \piso.data_r [3421] = \piso.data_r_3421_sv2v_reg ;
  assign \piso.data_r [3420] = \piso.data_r_3420_sv2v_reg ;
  assign \piso.data_r [3419] = \piso.data_r_3419_sv2v_reg ;
  assign \piso.data_r [3418] = \piso.data_r_3418_sv2v_reg ;
  assign \piso.data_r [3417] = \piso.data_r_3417_sv2v_reg ;
  assign \piso.data_r [3416] = \piso.data_r_3416_sv2v_reg ;
  assign \piso.data_r [3415] = \piso.data_r_3415_sv2v_reg ;
  assign \piso.data_r [3414] = \piso.data_r_3414_sv2v_reg ;
  assign \piso.data_r [3413] = \piso.data_r_3413_sv2v_reg ;
  assign \piso.data_r [3412] = \piso.data_r_3412_sv2v_reg ;
  assign \piso.data_r [3411] = \piso.data_r_3411_sv2v_reg ;
  assign \piso.data_r [3410] = \piso.data_r_3410_sv2v_reg ;
  assign \piso.data_r [3409] = \piso.data_r_3409_sv2v_reg ;
  assign \piso.data_r [3408] = \piso.data_r_3408_sv2v_reg ;
  assign \piso.data_r [3407] = \piso.data_r_3407_sv2v_reg ;
  assign \piso.data_r [3406] = \piso.data_r_3406_sv2v_reg ;
  assign \piso.data_r [3405] = \piso.data_r_3405_sv2v_reg ;
  assign \piso.data_r [3404] = \piso.data_r_3404_sv2v_reg ;
  assign \piso.data_r [3403] = \piso.data_r_3403_sv2v_reg ;
  assign \piso.data_r [3402] = \piso.data_r_3402_sv2v_reg ;
  assign \piso.data_r [3401] = \piso.data_r_3401_sv2v_reg ;
  assign \piso.data_r [3400] = \piso.data_r_3400_sv2v_reg ;
  assign \piso.data_r [3399] = \piso.data_r_3399_sv2v_reg ;
  assign \piso.data_r [3398] = \piso.data_r_3398_sv2v_reg ;
  assign \piso.data_r [3397] = \piso.data_r_3397_sv2v_reg ;
  assign \piso.data_r [3396] = \piso.data_r_3396_sv2v_reg ;
  assign \piso.data_r [3395] = \piso.data_r_3395_sv2v_reg ;
  assign \piso.data_r [3394] = \piso.data_r_3394_sv2v_reg ;
  assign \piso.data_r [3393] = \piso.data_r_3393_sv2v_reg ;
  assign \piso.data_r [3392] = \piso.data_r_3392_sv2v_reg ;
  assign \piso.data_r [3391] = \piso.data_r_3391_sv2v_reg ;
  assign \piso.data_r [3390] = \piso.data_r_3390_sv2v_reg ;
  assign \piso.data_r [3389] = \piso.data_r_3389_sv2v_reg ;
  assign \piso.data_r [3388] = \piso.data_r_3388_sv2v_reg ;
  assign \piso.data_r [3387] = \piso.data_r_3387_sv2v_reg ;
  assign \piso.data_r [3386] = \piso.data_r_3386_sv2v_reg ;
  assign \piso.data_r [3385] = \piso.data_r_3385_sv2v_reg ;
  assign \piso.data_r [3384] = \piso.data_r_3384_sv2v_reg ;
  assign \piso.data_r [3383] = \piso.data_r_3383_sv2v_reg ;
  assign \piso.data_r [3382] = \piso.data_r_3382_sv2v_reg ;
  assign \piso.data_r [3381] = \piso.data_r_3381_sv2v_reg ;
  assign \piso.data_r [3380] = \piso.data_r_3380_sv2v_reg ;
  assign \piso.data_r [3379] = \piso.data_r_3379_sv2v_reg ;
  assign \piso.data_r [3378] = \piso.data_r_3378_sv2v_reg ;
  assign \piso.data_r [3377] = \piso.data_r_3377_sv2v_reg ;
  assign \piso.data_r [3376] = \piso.data_r_3376_sv2v_reg ;
  assign \piso.data_r [3375] = \piso.data_r_3375_sv2v_reg ;
  assign \piso.data_r [3374] = \piso.data_r_3374_sv2v_reg ;
  assign \piso.data_r [3373] = \piso.data_r_3373_sv2v_reg ;
  assign \piso.data_r [3372] = \piso.data_r_3372_sv2v_reg ;
  assign \piso.data_r [3371] = \piso.data_r_3371_sv2v_reg ;
  assign \piso.data_r [3370] = \piso.data_r_3370_sv2v_reg ;
  assign \piso.data_r [3369] = \piso.data_r_3369_sv2v_reg ;
  assign \piso.data_r [3368] = \piso.data_r_3368_sv2v_reg ;
  assign \piso.data_r [3367] = \piso.data_r_3367_sv2v_reg ;
  assign \piso.data_r [3366] = \piso.data_r_3366_sv2v_reg ;
  assign \piso.data_r [3365] = \piso.data_r_3365_sv2v_reg ;
  assign \piso.data_r [3364] = \piso.data_r_3364_sv2v_reg ;
  assign \piso.data_r [3363] = \piso.data_r_3363_sv2v_reg ;
  assign \piso.data_r [3362] = \piso.data_r_3362_sv2v_reg ;
  assign \piso.data_r [3361] = \piso.data_r_3361_sv2v_reg ;
  assign \piso.data_r [3360] = \piso.data_r_3360_sv2v_reg ;
  assign \piso.data_r [3359] = \piso.data_r_3359_sv2v_reg ;
  assign \piso.data_r [3358] = \piso.data_r_3358_sv2v_reg ;
  assign \piso.data_r [3357] = \piso.data_r_3357_sv2v_reg ;
  assign \piso.data_r [3356] = \piso.data_r_3356_sv2v_reg ;
  assign \piso.data_r [3355] = \piso.data_r_3355_sv2v_reg ;
  assign \piso.data_r [3354] = \piso.data_r_3354_sv2v_reg ;
  assign \piso.data_r [3353] = \piso.data_r_3353_sv2v_reg ;
  assign \piso.data_r [3352] = \piso.data_r_3352_sv2v_reg ;
  assign \piso.data_r [3351] = \piso.data_r_3351_sv2v_reg ;
  assign \piso.data_r [3350] = \piso.data_r_3350_sv2v_reg ;
  assign \piso.data_r [3349] = \piso.data_r_3349_sv2v_reg ;
  assign \piso.data_r [3348] = \piso.data_r_3348_sv2v_reg ;
  assign \piso.data_r [3347] = \piso.data_r_3347_sv2v_reg ;
  assign \piso.data_r [3346] = \piso.data_r_3346_sv2v_reg ;
  assign \piso.data_r [3345] = \piso.data_r_3345_sv2v_reg ;
  assign \piso.data_r [3344] = \piso.data_r_3344_sv2v_reg ;
  assign \piso.data_r [3343] = \piso.data_r_3343_sv2v_reg ;
  assign \piso.data_r [3342] = \piso.data_r_3342_sv2v_reg ;
  assign \piso.data_r [3341] = \piso.data_r_3341_sv2v_reg ;
  assign \piso.data_r [3340] = \piso.data_r_3340_sv2v_reg ;
  assign \piso.data_r [3339] = \piso.data_r_3339_sv2v_reg ;
  assign \piso.data_r [3338] = \piso.data_r_3338_sv2v_reg ;
  assign \piso.data_r [3337] = \piso.data_r_3337_sv2v_reg ;
  assign \piso.data_r [3336] = \piso.data_r_3336_sv2v_reg ;
  assign \piso.data_r [3335] = \piso.data_r_3335_sv2v_reg ;
  assign \piso.data_r [3334] = \piso.data_r_3334_sv2v_reg ;
  assign \piso.data_r [3333] = \piso.data_r_3333_sv2v_reg ;
  assign \piso.data_r [3332] = \piso.data_r_3332_sv2v_reg ;
  assign \piso.data_r [3331] = \piso.data_r_3331_sv2v_reg ;
  assign \piso.data_r [3330] = \piso.data_r_3330_sv2v_reg ;
  assign \piso.data_r [3329] = \piso.data_r_3329_sv2v_reg ;
  assign \piso.data_r [3328] = \piso.data_r_3328_sv2v_reg ;
  assign \piso.data_r [3327] = \piso.data_r_3327_sv2v_reg ;
  assign \piso.data_r [3326] = \piso.data_r_3326_sv2v_reg ;
  assign \piso.data_r [3325] = \piso.data_r_3325_sv2v_reg ;
  assign \piso.data_r [3324] = \piso.data_r_3324_sv2v_reg ;
  assign \piso.data_r [3323] = \piso.data_r_3323_sv2v_reg ;
  assign \piso.data_r [3322] = \piso.data_r_3322_sv2v_reg ;
  assign \piso.data_r [3321] = \piso.data_r_3321_sv2v_reg ;
  assign \piso.data_r [3320] = \piso.data_r_3320_sv2v_reg ;
  assign \piso.data_r [3319] = \piso.data_r_3319_sv2v_reg ;
  assign \piso.data_r [3318] = \piso.data_r_3318_sv2v_reg ;
  assign \piso.data_r [3317] = \piso.data_r_3317_sv2v_reg ;
  assign \piso.data_r [3316] = \piso.data_r_3316_sv2v_reg ;
  assign \piso.data_r [3315] = \piso.data_r_3315_sv2v_reg ;
  assign \piso.data_r [3314] = \piso.data_r_3314_sv2v_reg ;
  assign \piso.data_r [3313] = \piso.data_r_3313_sv2v_reg ;
  assign \piso.data_r [3312] = \piso.data_r_3312_sv2v_reg ;
  assign \piso.data_r [3311] = \piso.data_r_3311_sv2v_reg ;
  assign \piso.data_r [3310] = \piso.data_r_3310_sv2v_reg ;
  assign \piso.data_r [3309] = \piso.data_r_3309_sv2v_reg ;
  assign \piso.data_r [3308] = \piso.data_r_3308_sv2v_reg ;
  assign \piso.data_r [3307] = \piso.data_r_3307_sv2v_reg ;
  assign \piso.data_r [3306] = \piso.data_r_3306_sv2v_reg ;
  assign \piso.data_r [3305] = \piso.data_r_3305_sv2v_reg ;
  assign \piso.data_r [3304] = \piso.data_r_3304_sv2v_reg ;
  assign \piso.data_r [3303] = \piso.data_r_3303_sv2v_reg ;
  assign \piso.data_r [3302] = \piso.data_r_3302_sv2v_reg ;
  assign \piso.data_r [3301] = \piso.data_r_3301_sv2v_reg ;
  assign \piso.data_r [3300] = \piso.data_r_3300_sv2v_reg ;
  assign \piso.data_r [3299] = \piso.data_r_3299_sv2v_reg ;
  assign \piso.data_r [3298] = \piso.data_r_3298_sv2v_reg ;
  assign \piso.data_r [3297] = \piso.data_r_3297_sv2v_reg ;
  assign \piso.data_r [3296] = \piso.data_r_3296_sv2v_reg ;
  assign \piso.data_r [3295] = \piso.data_r_3295_sv2v_reg ;
  assign \piso.data_r [3294] = \piso.data_r_3294_sv2v_reg ;
  assign \piso.data_r [3293] = \piso.data_r_3293_sv2v_reg ;
  assign \piso.data_r [3292] = \piso.data_r_3292_sv2v_reg ;
  assign \piso.data_r [3291] = \piso.data_r_3291_sv2v_reg ;
  assign \piso.data_r [3290] = \piso.data_r_3290_sv2v_reg ;
  assign \piso.data_r [3289] = \piso.data_r_3289_sv2v_reg ;
  assign \piso.data_r [3288] = \piso.data_r_3288_sv2v_reg ;
  assign \piso.data_r [3287] = \piso.data_r_3287_sv2v_reg ;
  assign \piso.data_r [3286] = \piso.data_r_3286_sv2v_reg ;
  assign \piso.data_r [3285] = \piso.data_r_3285_sv2v_reg ;
  assign \piso.data_r [3284] = \piso.data_r_3284_sv2v_reg ;
  assign \piso.data_r [3283] = \piso.data_r_3283_sv2v_reg ;
  assign \piso.data_r [3282] = \piso.data_r_3282_sv2v_reg ;
  assign \piso.data_r [3281] = \piso.data_r_3281_sv2v_reg ;
  assign \piso.data_r [3280] = \piso.data_r_3280_sv2v_reg ;
  assign \piso.data_r [3279] = \piso.data_r_3279_sv2v_reg ;
  assign \piso.data_r [3278] = \piso.data_r_3278_sv2v_reg ;
  assign \piso.data_r [3277] = \piso.data_r_3277_sv2v_reg ;
  assign \piso.data_r [3276] = \piso.data_r_3276_sv2v_reg ;
  assign \piso.data_r [3275] = \piso.data_r_3275_sv2v_reg ;
  assign \piso.data_r [3274] = \piso.data_r_3274_sv2v_reg ;
  assign \piso.data_r [3273] = \piso.data_r_3273_sv2v_reg ;
  assign \piso.data_r [3272] = \piso.data_r_3272_sv2v_reg ;
  assign \piso.data_r [3271] = \piso.data_r_3271_sv2v_reg ;
  assign \piso.data_r [3270] = \piso.data_r_3270_sv2v_reg ;
  assign \piso.data_r [3269] = \piso.data_r_3269_sv2v_reg ;
  assign \piso.data_r [3268] = \piso.data_r_3268_sv2v_reg ;
  assign \piso.data_r [3267] = \piso.data_r_3267_sv2v_reg ;
  assign \piso.data_r [3266] = \piso.data_r_3266_sv2v_reg ;
  assign \piso.data_r [3265] = \piso.data_r_3265_sv2v_reg ;
  assign \piso.data_r [3264] = \piso.data_r_3264_sv2v_reg ;
  assign \piso.data_r [3263] = \piso.data_r_3263_sv2v_reg ;
  assign \piso.data_r [3262] = \piso.data_r_3262_sv2v_reg ;
  assign \piso.data_r [3261] = \piso.data_r_3261_sv2v_reg ;
  assign \piso.data_r [3260] = \piso.data_r_3260_sv2v_reg ;
  assign \piso.data_r [3259] = \piso.data_r_3259_sv2v_reg ;
  assign \piso.data_r [3258] = \piso.data_r_3258_sv2v_reg ;
  assign \piso.data_r [3257] = \piso.data_r_3257_sv2v_reg ;
  assign \piso.data_r [3256] = \piso.data_r_3256_sv2v_reg ;
  assign \piso.data_r [3255] = \piso.data_r_3255_sv2v_reg ;
  assign \piso.data_r [3254] = \piso.data_r_3254_sv2v_reg ;
  assign \piso.data_r [3253] = \piso.data_r_3253_sv2v_reg ;
  assign \piso.data_r [3252] = \piso.data_r_3252_sv2v_reg ;
  assign \piso.data_r [3251] = \piso.data_r_3251_sv2v_reg ;
  assign \piso.data_r [3250] = \piso.data_r_3250_sv2v_reg ;
  assign \piso.data_r [3249] = \piso.data_r_3249_sv2v_reg ;
  assign \piso.data_r [3248] = \piso.data_r_3248_sv2v_reg ;
  assign \piso.data_r [3247] = \piso.data_r_3247_sv2v_reg ;
  assign \piso.data_r [3246] = \piso.data_r_3246_sv2v_reg ;
  assign \piso.data_r [3245] = \piso.data_r_3245_sv2v_reg ;
  assign \piso.data_r [3244] = \piso.data_r_3244_sv2v_reg ;
  assign \piso.data_r [3243] = \piso.data_r_3243_sv2v_reg ;
  assign \piso.data_r [3242] = \piso.data_r_3242_sv2v_reg ;
  assign \piso.data_r [3241] = \piso.data_r_3241_sv2v_reg ;
  assign \piso.data_r [3240] = \piso.data_r_3240_sv2v_reg ;
  assign \piso.data_r [3239] = \piso.data_r_3239_sv2v_reg ;
  assign \piso.data_r [3238] = \piso.data_r_3238_sv2v_reg ;
  assign \piso.data_r [3237] = \piso.data_r_3237_sv2v_reg ;
  assign \piso.data_r [3236] = \piso.data_r_3236_sv2v_reg ;
  assign \piso.data_r [3235] = \piso.data_r_3235_sv2v_reg ;
  assign \piso.data_r [3234] = \piso.data_r_3234_sv2v_reg ;
  assign \piso.data_r [3233] = \piso.data_r_3233_sv2v_reg ;
  assign \piso.data_r [3232] = \piso.data_r_3232_sv2v_reg ;
  assign \piso.data_r [3231] = \piso.data_r_3231_sv2v_reg ;
  assign \piso.data_r [3230] = \piso.data_r_3230_sv2v_reg ;
  assign \piso.data_r [3229] = \piso.data_r_3229_sv2v_reg ;
  assign \piso.data_r [3228] = \piso.data_r_3228_sv2v_reg ;
  assign \piso.data_r [3227] = \piso.data_r_3227_sv2v_reg ;
  assign \piso.data_r [3226] = \piso.data_r_3226_sv2v_reg ;
  assign \piso.data_r [3225] = \piso.data_r_3225_sv2v_reg ;
  assign \piso.data_r [3224] = \piso.data_r_3224_sv2v_reg ;
  assign \piso.data_r [3223] = \piso.data_r_3223_sv2v_reg ;
  assign \piso.data_r [3222] = \piso.data_r_3222_sv2v_reg ;
  assign \piso.data_r [3221] = \piso.data_r_3221_sv2v_reg ;
  assign \piso.data_r [3220] = \piso.data_r_3220_sv2v_reg ;
  assign \piso.data_r [3219] = \piso.data_r_3219_sv2v_reg ;
  assign \piso.data_r [3218] = \piso.data_r_3218_sv2v_reg ;
  assign \piso.data_r [3217] = \piso.data_r_3217_sv2v_reg ;
  assign \piso.data_r [3216] = \piso.data_r_3216_sv2v_reg ;
  assign \piso.data_r [3215] = \piso.data_r_3215_sv2v_reg ;
  assign \piso.data_r [3214] = \piso.data_r_3214_sv2v_reg ;
  assign \piso.data_r [3213] = \piso.data_r_3213_sv2v_reg ;
  assign \piso.data_r [3212] = \piso.data_r_3212_sv2v_reg ;
  assign \piso.data_r [3211] = \piso.data_r_3211_sv2v_reg ;
  assign \piso.data_r [3210] = \piso.data_r_3210_sv2v_reg ;
  assign \piso.data_r [3209] = \piso.data_r_3209_sv2v_reg ;
  assign \piso.data_r [3208] = \piso.data_r_3208_sv2v_reg ;
  assign \piso.data_r [3207] = \piso.data_r_3207_sv2v_reg ;
  assign \piso.data_r [3206] = \piso.data_r_3206_sv2v_reg ;
  assign \piso.data_r [3205] = \piso.data_r_3205_sv2v_reg ;
  assign \piso.data_r [3204] = \piso.data_r_3204_sv2v_reg ;
  assign \piso.data_r [3203] = \piso.data_r_3203_sv2v_reg ;
  assign \piso.data_r [3202] = \piso.data_r_3202_sv2v_reg ;
  assign \piso.data_r [3201] = \piso.data_r_3201_sv2v_reg ;
  assign \piso.data_r [3200] = \piso.data_r_3200_sv2v_reg ;
  assign \piso.data_r [3199] = \piso.data_r_3199_sv2v_reg ;
  assign \piso.data_r [3198] = \piso.data_r_3198_sv2v_reg ;
  assign \piso.data_r [3197] = \piso.data_r_3197_sv2v_reg ;
  assign \piso.data_r [3196] = \piso.data_r_3196_sv2v_reg ;
  assign \piso.data_r [3195] = \piso.data_r_3195_sv2v_reg ;
  assign \piso.data_r [3194] = \piso.data_r_3194_sv2v_reg ;
  assign \piso.data_r [3193] = \piso.data_r_3193_sv2v_reg ;
  assign \piso.data_r [3192] = \piso.data_r_3192_sv2v_reg ;
  assign \piso.data_r [3191] = \piso.data_r_3191_sv2v_reg ;
  assign \piso.data_r [3190] = \piso.data_r_3190_sv2v_reg ;
  assign \piso.data_r [3189] = \piso.data_r_3189_sv2v_reg ;
  assign \piso.data_r [3188] = \piso.data_r_3188_sv2v_reg ;
  assign \piso.data_r [3187] = \piso.data_r_3187_sv2v_reg ;
  assign \piso.data_r [3186] = \piso.data_r_3186_sv2v_reg ;
  assign \piso.data_r [3185] = \piso.data_r_3185_sv2v_reg ;
  assign \piso.data_r [3184] = \piso.data_r_3184_sv2v_reg ;
  assign \piso.data_r [3183] = \piso.data_r_3183_sv2v_reg ;
  assign \piso.data_r [3182] = \piso.data_r_3182_sv2v_reg ;
  assign \piso.data_r [3181] = \piso.data_r_3181_sv2v_reg ;
  assign \piso.data_r [3180] = \piso.data_r_3180_sv2v_reg ;
  assign \piso.data_r [3179] = \piso.data_r_3179_sv2v_reg ;
  assign \piso.data_r [3178] = \piso.data_r_3178_sv2v_reg ;
  assign \piso.data_r [3177] = \piso.data_r_3177_sv2v_reg ;
  assign \piso.data_r [3176] = \piso.data_r_3176_sv2v_reg ;
  assign \piso.data_r [3175] = \piso.data_r_3175_sv2v_reg ;
  assign \piso.data_r [3174] = \piso.data_r_3174_sv2v_reg ;
  assign \piso.data_r [3173] = \piso.data_r_3173_sv2v_reg ;
  assign \piso.data_r [3172] = \piso.data_r_3172_sv2v_reg ;
  assign \piso.data_r [3171] = \piso.data_r_3171_sv2v_reg ;
  assign \piso.data_r [3170] = \piso.data_r_3170_sv2v_reg ;
  assign \piso.data_r [3169] = \piso.data_r_3169_sv2v_reg ;
  assign \piso.data_r [3168] = \piso.data_r_3168_sv2v_reg ;
  assign \piso.data_r [3167] = \piso.data_r_3167_sv2v_reg ;
  assign \piso.data_r [3166] = \piso.data_r_3166_sv2v_reg ;
  assign \piso.data_r [3165] = \piso.data_r_3165_sv2v_reg ;
  assign \piso.data_r [3164] = \piso.data_r_3164_sv2v_reg ;
  assign \piso.data_r [3163] = \piso.data_r_3163_sv2v_reg ;
  assign \piso.data_r [3162] = \piso.data_r_3162_sv2v_reg ;
  assign \piso.data_r [3161] = \piso.data_r_3161_sv2v_reg ;
  assign \piso.data_r [3160] = \piso.data_r_3160_sv2v_reg ;
  assign \piso.data_r [3159] = \piso.data_r_3159_sv2v_reg ;
  assign \piso.data_r [3158] = \piso.data_r_3158_sv2v_reg ;
  assign \piso.data_r [3157] = \piso.data_r_3157_sv2v_reg ;
  assign \piso.data_r [3156] = \piso.data_r_3156_sv2v_reg ;
  assign \piso.data_r [3155] = \piso.data_r_3155_sv2v_reg ;
  assign \piso.data_r [3154] = \piso.data_r_3154_sv2v_reg ;
  assign \piso.data_r [3153] = \piso.data_r_3153_sv2v_reg ;
  assign \piso.data_r [3152] = \piso.data_r_3152_sv2v_reg ;
  assign \piso.data_r [3151] = \piso.data_r_3151_sv2v_reg ;
  assign \piso.data_r [3150] = \piso.data_r_3150_sv2v_reg ;
  assign \piso.data_r [3149] = \piso.data_r_3149_sv2v_reg ;
  assign \piso.data_r [3148] = \piso.data_r_3148_sv2v_reg ;
  assign \piso.data_r [3147] = \piso.data_r_3147_sv2v_reg ;
  assign \piso.data_r [3146] = \piso.data_r_3146_sv2v_reg ;
  assign \piso.data_r [3145] = \piso.data_r_3145_sv2v_reg ;
  assign \piso.data_r [3144] = \piso.data_r_3144_sv2v_reg ;
  assign \piso.data_r [3143] = \piso.data_r_3143_sv2v_reg ;
  assign \piso.data_r [3142] = \piso.data_r_3142_sv2v_reg ;
  assign \piso.data_r [3141] = \piso.data_r_3141_sv2v_reg ;
  assign \piso.data_r [3140] = \piso.data_r_3140_sv2v_reg ;
  assign \piso.data_r [3139] = \piso.data_r_3139_sv2v_reg ;
  assign \piso.data_r [3138] = \piso.data_r_3138_sv2v_reg ;
  assign \piso.data_r [3137] = \piso.data_r_3137_sv2v_reg ;
  assign \piso.data_r [3136] = \piso.data_r_3136_sv2v_reg ;
  assign \piso.data_r [3135] = \piso.data_r_3135_sv2v_reg ;
  assign \piso.data_r [3134] = \piso.data_r_3134_sv2v_reg ;
  assign \piso.data_r [3133] = \piso.data_r_3133_sv2v_reg ;
  assign \piso.data_r [3132] = \piso.data_r_3132_sv2v_reg ;
  assign \piso.data_r [3131] = \piso.data_r_3131_sv2v_reg ;
  assign \piso.data_r [3130] = \piso.data_r_3130_sv2v_reg ;
  assign \piso.data_r [3129] = \piso.data_r_3129_sv2v_reg ;
  assign \piso.data_r [3128] = \piso.data_r_3128_sv2v_reg ;
  assign \piso.data_r [3127] = \piso.data_r_3127_sv2v_reg ;
  assign \piso.data_r [3126] = \piso.data_r_3126_sv2v_reg ;
  assign \piso.data_r [3125] = \piso.data_r_3125_sv2v_reg ;
  assign \piso.data_r [3124] = \piso.data_r_3124_sv2v_reg ;
  assign \piso.data_r [3123] = \piso.data_r_3123_sv2v_reg ;
  assign \piso.data_r [3122] = \piso.data_r_3122_sv2v_reg ;
  assign \piso.data_r [3121] = \piso.data_r_3121_sv2v_reg ;
  assign \piso.data_r [3120] = \piso.data_r_3120_sv2v_reg ;
  assign \piso.data_r [3119] = \piso.data_r_3119_sv2v_reg ;
  assign \piso.data_r [3118] = \piso.data_r_3118_sv2v_reg ;
  assign \piso.data_r [3117] = \piso.data_r_3117_sv2v_reg ;
  assign \piso.data_r [3116] = \piso.data_r_3116_sv2v_reg ;
  assign \piso.data_r [3115] = \piso.data_r_3115_sv2v_reg ;
  assign \piso.data_r [3114] = \piso.data_r_3114_sv2v_reg ;
  assign \piso.data_r [3113] = \piso.data_r_3113_sv2v_reg ;
  assign \piso.data_r [3112] = \piso.data_r_3112_sv2v_reg ;
  assign \piso.data_r [3111] = \piso.data_r_3111_sv2v_reg ;
  assign \piso.data_r [3110] = \piso.data_r_3110_sv2v_reg ;
  assign \piso.data_r [3109] = \piso.data_r_3109_sv2v_reg ;
  assign \piso.data_r [3108] = \piso.data_r_3108_sv2v_reg ;
  assign \piso.data_r [3107] = \piso.data_r_3107_sv2v_reg ;
  assign \piso.data_r [3106] = \piso.data_r_3106_sv2v_reg ;
  assign \piso.data_r [3105] = \piso.data_r_3105_sv2v_reg ;
  assign \piso.data_r [3104] = \piso.data_r_3104_sv2v_reg ;
  assign \piso.data_r [3103] = \piso.data_r_3103_sv2v_reg ;
  assign \piso.data_r [3102] = \piso.data_r_3102_sv2v_reg ;
  assign \piso.data_r [3101] = \piso.data_r_3101_sv2v_reg ;
  assign \piso.data_r [3100] = \piso.data_r_3100_sv2v_reg ;
  assign \piso.data_r [3099] = \piso.data_r_3099_sv2v_reg ;
  assign \piso.data_r [3098] = \piso.data_r_3098_sv2v_reg ;
  assign \piso.data_r [3097] = \piso.data_r_3097_sv2v_reg ;
  assign \piso.data_r [3096] = \piso.data_r_3096_sv2v_reg ;
  assign \piso.data_r [3095] = \piso.data_r_3095_sv2v_reg ;
  assign \piso.data_r [3094] = \piso.data_r_3094_sv2v_reg ;
  assign \piso.data_r [3093] = \piso.data_r_3093_sv2v_reg ;
  assign \piso.data_r [3092] = \piso.data_r_3092_sv2v_reg ;
  assign \piso.data_r [3091] = \piso.data_r_3091_sv2v_reg ;
  assign \piso.data_r [3090] = \piso.data_r_3090_sv2v_reg ;
  assign \piso.data_r [3089] = \piso.data_r_3089_sv2v_reg ;
  assign \piso.data_r [3088] = \piso.data_r_3088_sv2v_reg ;
  assign \piso.data_r [3087] = \piso.data_r_3087_sv2v_reg ;
  assign \piso.data_r [3086] = \piso.data_r_3086_sv2v_reg ;
  assign \piso.data_r [3085] = \piso.data_r_3085_sv2v_reg ;
  assign \piso.data_r [3084] = \piso.data_r_3084_sv2v_reg ;
  assign \piso.data_r [3083] = \piso.data_r_3083_sv2v_reg ;
  assign \piso.data_r [3082] = \piso.data_r_3082_sv2v_reg ;
  assign \piso.data_r [3081] = \piso.data_r_3081_sv2v_reg ;
  assign \piso.data_r [3080] = \piso.data_r_3080_sv2v_reg ;
  assign \piso.data_r [3079] = \piso.data_r_3079_sv2v_reg ;
  assign \piso.data_r [3078] = \piso.data_r_3078_sv2v_reg ;
  assign \piso.data_r [3077] = \piso.data_r_3077_sv2v_reg ;
  assign \piso.data_r [3076] = \piso.data_r_3076_sv2v_reg ;
  assign \piso.data_r [3075] = \piso.data_r_3075_sv2v_reg ;
  assign \piso.data_r [3074] = \piso.data_r_3074_sv2v_reg ;
  assign \piso.data_r [3073] = \piso.data_r_3073_sv2v_reg ;
  assign \piso.data_r [3072] = \piso.data_r_3072_sv2v_reg ;
  assign \piso.data_r [3071] = \piso.data_r_3071_sv2v_reg ;
  assign \piso.data_r [3070] = \piso.data_r_3070_sv2v_reg ;
  assign \piso.data_r [3069] = \piso.data_r_3069_sv2v_reg ;
  assign \piso.data_r [3068] = \piso.data_r_3068_sv2v_reg ;
  assign \piso.data_r [3067] = \piso.data_r_3067_sv2v_reg ;
  assign \piso.data_r [3066] = \piso.data_r_3066_sv2v_reg ;
  assign \piso.data_r [3065] = \piso.data_r_3065_sv2v_reg ;
  assign \piso.data_r [3064] = \piso.data_r_3064_sv2v_reg ;
  assign \piso.data_r [3063] = \piso.data_r_3063_sv2v_reg ;
  assign \piso.data_r [3062] = \piso.data_r_3062_sv2v_reg ;
  assign \piso.data_r [3061] = \piso.data_r_3061_sv2v_reg ;
  assign \piso.data_r [3060] = \piso.data_r_3060_sv2v_reg ;
  assign \piso.data_r [3059] = \piso.data_r_3059_sv2v_reg ;
  assign \piso.data_r [3058] = \piso.data_r_3058_sv2v_reg ;
  assign \piso.data_r [3057] = \piso.data_r_3057_sv2v_reg ;
  assign \piso.data_r [3056] = \piso.data_r_3056_sv2v_reg ;
  assign \piso.data_r [3055] = \piso.data_r_3055_sv2v_reg ;
  assign \piso.data_r [3054] = \piso.data_r_3054_sv2v_reg ;
  assign \piso.data_r [3053] = \piso.data_r_3053_sv2v_reg ;
  assign \piso.data_r [3052] = \piso.data_r_3052_sv2v_reg ;
  assign \piso.data_r [3051] = \piso.data_r_3051_sv2v_reg ;
  assign \piso.data_r [3050] = \piso.data_r_3050_sv2v_reg ;
  assign \piso.data_r [3049] = \piso.data_r_3049_sv2v_reg ;
  assign \piso.data_r [3048] = \piso.data_r_3048_sv2v_reg ;
  assign \piso.data_r [3047] = \piso.data_r_3047_sv2v_reg ;
  assign \piso.data_r [3046] = \piso.data_r_3046_sv2v_reg ;
  assign \piso.data_r [3045] = \piso.data_r_3045_sv2v_reg ;
  assign \piso.data_r [3044] = \piso.data_r_3044_sv2v_reg ;
  assign \piso.data_r [3043] = \piso.data_r_3043_sv2v_reg ;
  assign \piso.data_r [3042] = \piso.data_r_3042_sv2v_reg ;
  assign \piso.data_r [3041] = \piso.data_r_3041_sv2v_reg ;
  assign \piso.data_r [3040] = \piso.data_r_3040_sv2v_reg ;
  assign \piso.data_r [3039] = \piso.data_r_3039_sv2v_reg ;
  assign \piso.data_r [3038] = \piso.data_r_3038_sv2v_reg ;
  assign \piso.data_r [3037] = \piso.data_r_3037_sv2v_reg ;
  assign \piso.data_r [3036] = \piso.data_r_3036_sv2v_reg ;
  assign \piso.data_r [3035] = \piso.data_r_3035_sv2v_reg ;
  assign \piso.data_r [3034] = \piso.data_r_3034_sv2v_reg ;
  assign \piso.data_r [3033] = \piso.data_r_3033_sv2v_reg ;
  assign \piso.data_r [3032] = \piso.data_r_3032_sv2v_reg ;
  assign \piso.data_r [3031] = \piso.data_r_3031_sv2v_reg ;
  assign \piso.data_r [3030] = \piso.data_r_3030_sv2v_reg ;
  assign \piso.data_r [3029] = \piso.data_r_3029_sv2v_reg ;
  assign \piso.data_r [3028] = \piso.data_r_3028_sv2v_reg ;
  assign \piso.data_r [3027] = \piso.data_r_3027_sv2v_reg ;
  assign \piso.data_r [3026] = \piso.data_r_3026_sv2v_reg ;
  assign \piso.data_r [3025] = \piso.data_r_3025_sv2v_reg ;
  assign \piso.data_r [3024] = \piso.data_r_3024_sv2v_reg ;
  assign \piso.data_r [3023] = \piso.data_r_3023_sv2v_reg ;
  assign \piso.data_r [3022] = \piso.data_r_3022_sv2v_reg ;
  assign \piso.data_r [3021] = \piso.data_r_3021_sv2v_reg ;
  assign \piso.data_r [3020] = \piso.data_r_3020_sv2v_reg ;
  assign \piso.data_r [3019] = \piso.data_r_3019_sv2v_reg ;
  assign \piso.data_r [3018] = \piso.data_r_3018_sv2v_reg ;
  assign \piso.data_r [3017] = \piso.data_r_3017_sv2v_reg ;
  assign \piso.data_r [3016] = \piso.data_r_3016_sv2v_reg ;
  assign \piso.data_r [3015] = \piso.data_r_3015_sv2v_reg ;
  assign \piso.data_r [3014] = \piso.data_r_3014_sv2v_reg ;
  assign \piso.data_r [3013] = \piso.data_r_3013_sv2v_reg ;
  assign \piso.data_r [3012] = \piso.data_r_3012_sv2v_reg ;
  assign \piso.data_r [3011] = \piso.data_r_3011_sv2v_reg ;
  assign \piso.data_r [3010] = \piso.data_r_3010_sv2v_reg ;
  assign \piso.data_r [3009] = \piso.data_r_3009_sv2v_reg ;
  assign \piso.data_r [3008] = \piso.data_r_3008_sv2v_reg ;
  assign \piso.data_r [3007] = \piso.data_r_3007_sv2v_reg ;
  assign \piso.data_r [3006] = \piso.data_r_3006_sv2v_reg ;
  assign \piso.data_r [3005] = \piso.data_r_3005_sv2v_reg ;
  assign \piso.data_r [3004] = \piso.data_r_3004_sv2v_reg ;
  assign \piso.data_r [3003] = \piso.data_r_3003_sv2v_reg ;
  assign \piso.data_r [3002] = \piso.data_r_3002_sv2v_reg ;
  assign \piso.data_r [3001] = \piso.data_r_3001_sv2v_reg ;
  assign \piso.data_r [3000] = \piso.data_r_3000_sv2v_reg ;
  assign \piso.data_r [2999] = \piso.data_r_2999_sv2v_reg ;
  assign \piso.data_r [2998] = \piso.data_r_2998_sv2v_reg ;
  assign \piso.data_r [2997] = \piso.data_r_2997_sv2v_reg ;
  assign \piso.data_r [2996] = \piso.data_r_2996_sv2v_reg ;
  assign \piso.data_r [2995] = \piso.data_r_2995_sv2v_reg ;
  assign \piso.data_r [2994] = \piso.data_r_2994_sv2v_reg ;
  assign \piso.data_r [2993] = \piso.data_r_2993_sv2v_reg ;
  assign \piso.data_r [2992] = \piso.data_r_2992_sv2v_reg ;
  assign \piso.data_r [2991] = \piso.data_r_2991_sv2v_reg ;
  assign \piso.data_r [2990] = \piso.data_r_2990_sv2v_reg ;
  assign \piso.data_r [2989] = \piso.data_r_2989_sv2v_reg ;
  assign \piso.data_r [2988] = \piso.data_r_2988_sv2v_reg ;
  assign \piso.data_r [2987] = \piso.data_r_2987_sv2v_reg ;
  assign \piso.data_r [2986] = \piso.data_r_2986_sv2v_reg ;
  assign \piso.data_r [2985] = \piso.data_r_2985_sv2v_reg ;
  assign \piso.data_r [2984] = \piso.data_r_2984_sv2v_reg ;
  assign \piso.data_r [2983] = \piso.data_r_2983_sv2v_reg ;
  assign \piso.data_r [2982] = \piso.data_r_2982_sv2v_reg ;
  assign \piso.data_r [2981] = \piso.data_r_2981_sv2v_reg ;
  assign \piso.data_r [2980] = \piso.data_r_2980_sv2v_reg ;
  assign \piso.data_r [2979] = \piso.data_r_2979_sv2v_reg ;
  assign \piso.data_r [2978] = \piso.data_r_2978_sv2v_reg ;
  assign \piso.data_r [2977] = \piso.data_r_2977_sv2v_reg ;
  assign \piso.data_r [2976] = \piso.data_r_2976_sv2v_reg ;
  assign \piso.data_r [2975] = \piso.data_r_2975_sv2v_reg ;
  assign \piso.data_r [2974] = \piso.data_r_2974_sv2v_reg ;
  assign \piso.data_r [2973] = \piso.data_r_2973_sv2v_reg ;
  assign \piso.data_r [2972] = \piso.data_r_2972_sv2v_reg ;
  assign \piso.data_r [2971] = \piso.data_r_2971_sv2v_reg ;
  assign \piso.data_r [2970] = \piso.data_r_2970_sv2v_reg ;
  assign \piso.data_r [2969] = \piso.data_r_2969_sv2v_reg ;
  assign \piso.data_r [2968] = \piso.data_r_2968_sv2v_reg ;
  assign \piso.data_r [2967] = \piso.data_r_2967_sv2v_reg ;
  assign \piso.data_r [2966] = \piso.data_r_2966_sv2v_reg ;
  assign \piso.data_r [2965] = \piso.data_r_2965_sv2v_reg ;
  assign \piso.data_r [2964] = \piso.data_r_2964_sv2v_reg ;
  assign \piso.data_r [2963] = \piso.data_r_2963_sv2v_reg ;
  assign \piso.data_r [2962] = \piso.data_r_2962_sv2v_reg ;
  assign \piso.data_r [2961] = \piso.data_r_2961_sv2v_reg ;
  assign \piso.data_r [2960] = \piso.data_r_2960_sv2v_reg ;
  assign \piso.data_r [2959] = \piso.data_r_2959_sv2v_reg ;
  assign \piso.data_r [2958] = \piso.data_r_2958_sv2v_reg ;
  assign \piso.data_r [2957] = \piso.data_r_2957_sv2v_reg ;
  assign \piso.data_r [2956] = \piso.data_r_2956_sv2v_reg ;
  assign \piso.data_r [2955] = \piso.data_r_2955_sv2v_reg ;
  assign \piso.data_r [2954] = \piso.data_r_2954_sv2v_reg ;
  assign \piso.data_r [2953] = \piso.data_r_2953_sv2v_reg ;
  assign \piso.data_r [2952] = \piso.data_r_2952_sv2v_reg ;
  assign \piso.data_r [2951] = \piso.data_r_2951_sv2v_reg ;
  assign \piso.data_r [2950] = \piso.data_r_2950_sv2v_reg ;
  assign \piso.data_r [2949] = \piso.data_r_2949_sv2v_reg ;
  assign \piso.data_r [2948] = \piso.data_r_2948_sv2v_reg ;
  assign \piso.data_r [2947] = \piso.data_r_2947_sv2v_reg ;
  assign \piso.data_r [2946] = \piso.data_r_2946_sv2v_reg ;
  assign \piso.data_r [2945] = \piso.data_r_2945_sv2v_reg ;
  assign \piso.data_r [2944] = \piso.data_r_2944_sv2v_reg ;
  assign \piso.data_r [2943] = \piso.data_r_2943_sv2v_reg ;
  assign \piso.data_r [2942] = \piso.data_r_2942_sv2v_reg ;
  assign \piso.data_r [2941] = \piso.data_r_2941_sv2v_reg ;
  assign \piso.data_r [2940] = \piso.data_r_2940_sv2v_reg ;
  assign \piso.data_r [2939] = \piso.data_r_2939_sv2v_reg ;
  assign \piso.data_r [2938] = \piso.data_r_2938_sv2v_reg ;
  assign \piso.data_r [2937] = \piso.data_r_2937_sv2v_reg ;
  assign \piso.data_r [2936] = \piso.data_r_2936_sv2v_reg ;
  assign \piso.data_r [2935] = \piso.data_r_2935_sv2v_reg ;
  assign \piso.data_r [2934] = \piso.data_r_2934_sv2v_reg ;
  assign \piso.data_r [2933] = \piso.data_r_2933_sv2v_reg ;
  assign \piso.data_r [2932] = \piso.data_r_2932_sv2v_reg ;
  assign \piso.data_r [2931] = \piso.data_r_2931_sv2v_reg ;
  assign \piso.data_r [2930] = \piso.data_r_2930_sv2v_reg ;
  assign \piso.data_r [2929] = \piso.data_r_2929_sv2v_reg ;
  assign \piso.data_r [2928] = \piso.data_r_2928_sv2v_reg ;
  assign \piso.data_r [2927] = \piso.data_r_2927_sv2v_reg ;
  assign \piso.data_r [2926] = \piso.data_r_2926_sv2v_reg ;
  assign \piso.data_r [2925] = \piso.data_r_2925_sv2v_reg ;
  assign \piso.data_r [2924] = \piso.data_r_2924_sv2v_reg ;
  assign \piso.data_r [2923] = \piso.data_r_2923_sv2v_reg ;
  assign \piso.data_r [2922] = \piso.data_r_2922_sv2v_reg ;
  assign \piso.data_r [2921] = \piso.data_r_2921_sv2v_reg ;
  assign \piso.data_r [2920] = \piso.data_r_2920_sv2v_reg ;
  assign \piso.data_r [2919] = \piso.data_r_2919_sv2v_reg ;
  assign \piso.data_r [2918] = \piso.data_r_2918_sv2v_reg ;
  assign \piso.data_r [2917] = \piso.data_r_2917_sv2v_reg ;
  assign \piso.data_r [2916] = \piso.data_r_2916_sv2v_reg ;
  assign \piso.data_r [2915] = \piso.data_r_2915_sv2v_reg ;
  assign \piso.data_r [2914] = \piso.data_r_2914_sv2v_reg ;
  assign \piso.data_r [2913] = \piso.data_r_2913_sv2v_reg ;
  assign \piso.data_r [2912] = \piso.data_r_2912_sv2v_reg ;
  assign \piso.data_r [2911] = \piso.data_r_2911_sv2v_reg ;
  assign \piso.data_r [2910] = \piso.data_r_2910_sv2v_reg ;
  assign \piso.data_r [2909] = \piso.data_r_2909_sv2v_reg ;
  assign \piso.data_r [2908] = \piso.data_r_2908_sv2v_reg ;
  assign \piso.data_r [2907] = \piso.data_r_2907_sv2v_reg ;
  assign \piso.data_r [2906] = \piso.data_r_2906_sv2v_reg ;
  assign \piso.data_r [2905] = \piso.data_r_2905_sv2v_reg ;
  assign \piso.data_r [2904] = \piso.data_r_2904_sv2v_reg ;
  assign \piso.data_r [2903] = \piso.data_r_2903_sv2v_reg ;
  assign \piso.data_r [2902] = \piso.data_r_2902_sv2v_reg ;
  assign \piso.data_r [2901] = \piso.data_r_2901_sv2v_reg ;
  assign \piso.data_r [2900] = \piso.data_r_2900_sv2v_reg ;
  assign \piso.data_r [2899] = \piso.data_r_2899_sv2v_reg ;
  assign \piso.data_r [2898] = \piso.data_r_2898_sv2v_reg ;
  assign \piso.data_r [2897] = \piso.data_r_2897_sv2v_reg ;
  assign \piso.data_r [2896] = \piso.data_r_2896_sv2v_reg ;
  assign \piso.data_r [2895] = \piso.data_r_2895_sv2v_reg ;
  assign \piso.data_r [2894] = \piso.data_r_2894_sv2v_reg ;
  assign \piso.data_r [2893] = \piso.data_r_2893_sv2v_reg ;
  assign \piso.data_r [2892] = \piso.data_r_2892_sv2v_reg ;
  assign \piso.data_r [2891] = \piso.data_r_2891_sv2v_reg ;
  assign \piso.data_r [2890] = \piso.data_r_2890_sv2v_reg ;
  assign \piso.data_r [2889] = \piso.data_r_2889_sv2v_reg ;
  assign \piso.data_r [2888] = \piso.data_r_2888_sv2v_reg ;
  assign \piso.data_r [2887] = \piso.data_r_2887_sv2v_reg ;
  assign \piso.data_r [2886] = \piso.data_r_2886_sv2v_reg ;
  assign \piso.data_r [2885] = \piso.data_r_2885_sv2v_reg ;
  assign \piso.data_r [2884] = \piso.data_r_2884_sv2v_reg ;
  assign \piso.data_r [2883] = \piso.data_r_2883_sv2v_reg ;
  assign \piso.data_r [2882] = \piso.data_r_2882_sv2v_reg ;
  assign \piso.data_r [2881] = \piso.data_r_2881_sv2v_reg ;
  assign \piso.data_r [2880] = \piso.data_r_2880_sv2v_reg ;
  assign \piso.data_r [2879] = \piso.data_r_2879_sv2v_reg ;
  assign \piso.data_r [2878] = \piso.data_r_2878_sv2v_reg ;
  assign \piso.data_r [2877] = \piso.data_r_2877_sv2v_reg ;
  assign \piso.data_r [2876] = \piso.data_r_2876_sv2v_reg ;
  assign \piso.data_r [2875] = \piso.data_r_2875_sv2v_reg ;
  assign \piso.data_r [2874] = \piso.data_r_2874_sv2v_reg ;
  assign \piso.data_r [2873] = \piso.data_r_2873_sv2v_reg ;
  assign \piso.data_r [2872] = \piso.data_r_2872_sv2v_reg ;
  assign \piso.data_r [2871] = \piso.data_r_2871_sv2v_reg ;
  assign \piso.data_r [2870] = \piso.data_r_2870_sv2v_reg ;
  assign \piso.data_r [2869] = \piso.data_r_2869_sv2v_reg ;
  assign \piso.data_r [2868] = \piso.data_r_2868_sv2v_reg ;
  assign \piso.data_r [2867] = \piso.data_r_2867_sv2v_reg ;
  assign \piso.data_r [2866] = \piso.data_r_2866_sv2v_reg ;
  assign \piso.data_r [2865] = \piso.data_r_2865_sv2v_reg ;
  assign \piso.data_r [2864] = \piso.data_r_2864_sv2v_reg ;
  assign \piso.data_r [2863] = \piso.data_r_2863_sv2v_reg ;
  assign \piso.data_r [2862] = \piso.data_r_2862_sv2v_reg ;
  assign \piso.data_r [2861] = \piso.data_r_2861_sv2v_reg ;
  assign \piso.data_r [2860] = \piso.data_r_2860_sv2v_reg ;
  assign \piso.data_r [2859] = \piso.data_r_2859_sv2v_reg ;
  assign \piso.data_r [2858] = \piso.data_r_2858_sv2v_reg ;
  assign \piso.data_r [2857] = \piso.data_r_2857_sv2v_reg ;
  assign \piso.data_r [2856] = \piso.data_r_2856_sv2v_reg ;
  assign \piso.data_r [2855] = \piso.data_r_2855_sv2v_reg ;
  assign \piso.data_r [2854] = \piso.data_r_2854_sv2v_reg ;
  assign \piso.data_r [2853] = \piso.data_r_2853_sv2v_reg ;
  assign \piso.data_r [2852] = \piso.data_r_2852_sv2v_reg ;
  assign \piso.data_r [2851] = \piso.data_r_2851_sv2v_reg ;
  assign \piso.data_r [2850] = \piso.data_r_2850_sv2v_reg ;
  assign \piso.data_r [2849] = \piso.data_r_2849_sv2v_reg ;
  assign \piso.data_r [2848] = \piso.data_r_2848_sv2v_reg ;
  assign \piso.data_r [2847] = \piso.data_r_2847_sv2v_reg ;
  assign \piso.data_r [2846] = \piso.data_r_2846_sv2v_reg ;
  assign \piso.data_r [2845] = \piso.data_r_2845_sv2v_reg ;
  assign \piso.data_r [2844] = \piso.data_r_2844_sv2v_reg ;
  assign \piso.data_r [2843] = \piso.data_r_2843_sv2v_reg ;
  assign \piso.data_r [2842] = \piso.data_r_2842_sv2v_reg ;
  assign \piso.data_r [2841] = \piso.data_r_2841_sv2v_reg ;
  assign \piso.data_r [2840] = \piso.data_r_2840_sv2v_reg ;
  assign \piso.data_r [2839] = \piso.data_r_2839_sv2v_reg ;
  assign \piso.data_r [2838] = \piso.data_r_2838_sv2v_reg ;
  assign \piso.data_r [2837] = \piso.data_r_2837_sv2v_reg ;
  assign \piso.data_r [2836] = \piso.data_r_2836_sv2v_reg ;
  assign \piso.data_r [2835] = \piso.data_r_2835_sv2v_reg ;
  assign \piso.data_r [2834] = \piso.data_r_2834_sv2v_reg ;
  assign \piso.data_r [2833] = \piso.data_r_2833_sv2v_reg ;
  assign \piso.data_r [2832] = \piso.data_r_2832_sv2v_reg ;
  assign \piso.data_r [2831] = \piso.data_r_2831_sv2v_reg ;
  assign \piso.data_r [2830] = \piso.data_r_2830_sv2v_reg ;
  assign \piso.data_r [2829] = \piso.data_r_2829_sv2v_reg ;
  assign \piso.data_r [2828] = \piso.data_r_2828_sv2v_reg ;
  assign \piso.data_r [2827] = \piso.data_r_2827_sv2v_reg ;
  assign \piso.data_r [2826] = \piso.data_r_2826_sv2v_reg ;
  assign \piso.data_r [2825] = \piso.data_r_2825_sv2v_reg ;
  assign \piso.data_r [2824] = \piso.data_r_2824_sv2v_reg ;
  assign \piso.data_r [2823] = \piso.data_r_2823_sv2v_reg ;
  assign \piso.data_r [2822] = \piso.data_r_2822_sv2v_reg ;
  assign \piso.data_r [2821] = \piso.data_r_2821_sv2v_reg ;
  assign \piso.data_r [2820] = \piso.data_r_2820_sv2v_reg ;
  assign \piso.data_r [2819] = \piso.data_r_2819_sv2v_reg ;
  assign \piso.data_r [2818] = \piso.data_r_2818_sv2v_reg ;
  assign \piso.data_r [2817] = \piso.data_r_2817_sv2v_reg ;
  assign \piso.data_r [2816] = \piso.data_r_2816_sv2v_reg ;
  assign \piso.data_r [2815] = \piso.data_r_2815_sv2v_reg ;
  assign \piso.data_r [2814] = \piso.data_r_2814_sv2v_reg ;
  assign \piso.data_r [2813] = \piso.data_r_2813_sv2v_reg ;
  assign \piso.data_r [2812] = \piso.data_r_2812_sv2v_reg ;
  assign \piso.data_r [2811] = \piso.data_r_2811_sv2v_reg ;
  assign \piso.data_r [2810] = \piso.data_r_2810_sv2v_reg ;
  assign \piso.data_r [2809] = \piso.data_r_2809_sv2v_reg ;
  assign \piso.data_r [2808] = \piso.data_r_2808_sv2v_reg ;
  assign \piso.data_r [2807] = \piso.data_r_2807_sv2v_reg ;
  assign \piso.data_r [2806] = \piso.data_r_2806_sv2v_reg ;
  assign \piso.data_r [2805] = \piso.data_r_2805_sv2v_reg ;
  assign \piso.data_r [2804] = \piso.data_r_2804_sv2v_reg ;
  assign \piso.data_r [2803] = \piso.data_r_2803_sv2v_reg ;
  assign \piso.data_r [2802] = \piso.data_r_2802_sv2v_reg ;
  assign \piso.data_r [2801] = \piso.data_r_2801_sv2v_reg ;
  assign \piso.data_r [2800] = \piso.data_r_2800_sv2v_reg ;
  assign \piso.data_r [2799] = \piso.data_r_2799_sv2v_reg ;
  assign \piso.data_r [2798] = \piso.data_r_2798_sv2v_reg ;
  assign \piso.data_r [2797] = \piso.data_r_2797_sv2v_reg ;
  assign \piso.data_r [2796] = \piso.data_r_2796_sv2v_reg ;
  assign \piso.data_r [2795] = \piso.data_r_2795_sv2v_reg ;
  assign \piso.data_r [2794] = \piso.data_r_2794_sv2v_reg ;
  assign \piso.data_r [2793] = \piso.data_r_2793_sv2v_reg ;
  assign \piso.data_r [2792] = \piso.data_r_2792_sv2v_reg ;
  assign \piso.data_r [2791] = \piso.data_r_2791_sv2v_reg ;
  assign \piso.data_r [2790] = \piso.data_r_2790_sv2v_reg ;
  assign \piso.data_r [2789] = \piso.data_r_2789_sv2v_reg ;
  assign \piso.data_r [2788] = \piso.data_r_2788_sv2v_reg ;
  assign \piso.data_r [2787] = \piso.data_r_2787_sv2v_reg ;
  assign \piso.data_r [2786] = \piso.data_r_2786_sv2v_reg ;
  assign \piso.data_r [2785] = \piso.data_r_2785_sv2v_reg ;
  assign \piso.data_r [2784] = \piso.data_r_2784_sv2v_reg ;
  assign \piso.data_r [2783] = \piso.data_r_2783_sv2v_reg ;
  assign \piso.data_r [2782] = \piso.data_r_2782_sv2v_reg ;
  assign \piso.data_r [2781] = \piso.data_r_2781_sv2v_reg ;
  assign \piso.data_r [2780] = \piso.data_r_2780_sv2v_reg ;
  assign \piso.data_r [2779] = \piso.data_r_2779_sv2v_reg ;
  assign \piso.data_r [2778] = \piso.data_r_2778_sv2v_reg ;
  assign \piso.data_r [2777] = \piso.data_r_2777_sv2v_reg ;
  assign \piso.data_r [2776] = \piso.data_r_2776_sv2v_reg ;
  assign \piso.data_r [2775] = \piso.data_r_2775_sv2v_reg ;
  assign \piso.data_r [2774] = \piso.data_r_2774_sv2v_reg ;
  assign \piso.data_r [2773] = \piso.data_r_2773_sv2v_reg ;
  assign \piso.data_r [2772] = \piso.data_r_2772_sv2v_reg ;
  assign \piso.data_r [2771] = \piso.data_r_2771_sv2v_reg ;
  assign \piso.data_r [2770] = \piso.data_r_2770_sv2v_reg ;
  assign \piso.data_r [2769] = \piso.data_r_2769_sv2v_reg ;
  assign \piso.data_r [2768] = \piso.data_r_2768_sv2v_reg ;
  assign \piso.data_r [2767] = \piso.data_r_2767_sv2v_reg ;
  assign \piso.data_r [2766] = \piso.data_r_2766_sv2v_reg ;
  assign \piso.data_r [2765] = \piso.data_r_2765_sv2v_reg ;
  assign \piso.data_r [2764] = \piso.data_r_2764_sv2v_reg ;
  assign \piso.data_r [2763] = \piso.data_r_2763_sv2v_reg ;
  assign \piso.data_r [2762] = \piso.data_r_2762_sv2v_reg ;
  assign \piso.data_r [2761] = \piso.data_r_2761_sv2v_reg ;
  assign \piso.data_r [2760] = \piso.data_r_2760_sv2v_reg ;
  assign \piso.data_r [2759] = \piso.data_r_2759_sv2v_reg ;
  assign \piso.data_r [2758] = \piso.data_r_2758_sv2v_reg ;
  assign \piso.data_r [2757] = \piso.data_r_2757_sv2v_reg ;
  assign \piso.data_r [2756] = \piso.data_r_2756_sv2v_reg ;
  assign \piso.data_r [2755] = \piso.data_r_2755_sv2v_reg ;
  assign \piso.data_r [2754] = \piso.data_r_2754_sv2v_reg ;
  assign \piso.data_r [2753] = \piso.data_r_2753_sv2v_reg ;
  assign \piso.data_r [2752] = \piso.data_r_2752_sv2v_reg ;
  assign \piso.data_r [2751] = \piso.data_r_2751_sv2v_reg ;
  assign \piso.data_r [2750] = \piso.data_r_2750_sv2v_reg ;
  assign \piso.data_r [2749] = \piso.data_r_2749_sv2v_reg ;
  assign \piso.data_r [2748] = \piso.data_r_2748_sv2v_reg ;
  assign \piso.data_r [2747] = \piso.data_r_2747_sv2v_reg ;
  assign \piso.data_r [2746] = \piso.data_r_2746_sv2v_reg ;
  assign \piso.data_r [2745] = \piso.data_r_2745_sv2v_reg ;
  assign \piso.data_r [2744] = \piso.data_r_2744_sv2v_reg ;
  assign \piso.data_r [2743] = \piso.data_r_2743_sv2v_reg ;
  assign \piso.data_r [2742] = \piso.data_r_2742_sv2v_reg ;
  assign \piso.data_r [2741] = \piso.data_r_2741_sv2v_reg ;
  assign \piso.data_r [2740] = \piso.data_r_2740_sv2v_reg ;
  assign \piso.data_r [2739] = \piso.data_r_2739_sv2v_reg ;
  assign \piso.data_r [2738] = \piso.data_r_2738_sv2v_reg ;
  assign \piso.data_r [2737] = \piso.data_r_2737_sv2v_reg ;
  assign \piso.data_r [2736] = \piso.data_r_2736_sv2v_reg ;
  assign \piso.data_r [2735] = \piso.data_r_2735_sv2v_reg ;
  assign \piso.data_r [2734] = \piso.data_r_2734_sv2v_reg ;
  assign \piso.data_r [2733] = \piso.data_r_2733_sv2v_reg ;
  assign \piso.data_r [2732] = \piso.data_r_2732_sv2v_reg ;
  assign \piso.data_r [2731] = \piso.data_r_2731_sv2v_reg ;
  assign \piso.data_r [2730] = \piso.data_r_2730_sv2v_reg ;
  assign \piso.data_r [2729] = \piso.data_r_2729_sv2v_reg ;
  assign \piso.data_r [2728] = \piso.data_r_2728_sv2v_reg ;
  assign \piso.data_r [2727] = \piso.data_r_2727_sv2v_reg ;
  assign \piso.data_r [2726] = \piso.data_r_2726_sv2v_reg ;
  assign \piso.data_r [2725] = \piso.data_r_2725_sv2v_reg ;
  assign \piso.data_r [2724] = \piso.data_r_2724_sv2v_reg ;
  assign \piso.data_r [2723] = \piso.data_r_2723_sv2v_reg ;
  assign \piso.data_r [2722] = \piso.data_r_2722_sv2v_reg ;
  assign \piso.data_r [2721] = \piso.data_r_2721_sv2v_reg ;
  assign \piso.data_r [2720] = \piso.data_r_2720_sv2v_reg ;
  assign \piso.data_r [2719] = \piso.data_r_2719_sv2v_reg ;
  assign \piso.data_r [2718] = \piso.data_r_2718_sv2v_reg ;
  assign \piso.data_r [2717] = \piso.data_r_2717_sv2v_reg ;
  assign \piso.data_r [2716] = \piso.data_r_2716_sv2v_reg ;
  assign \piso.data_r [2715] = \piso.data_r_2715_sv2v_reg ;
  assign \piso.data_r [2714] = \piso.data_r_2714_sv2v_reg ;
  assign \piso.data_r [2713] = \piso.data_r_2713_sv2v_reg ;
  assign \piso.data_r [2712] = \piso.data_r_2712_sv2v_reg ;
  assign \piso.data_r [2711] = \piso.data_r_2711_sv2v_reg ;
  assign \piso.data_r [2710] = \piso.data_r_2710_sv2v_reg ;
  assign \piso.data_r [2709] = \piso.data_r_2709_sv2v_reg ;
  assign \piso.data_r [2708] = \piso.data_r_2708_sv2v_reg ;
  assign \piso.data_r [2707] = \piso.data_r_2707_sv2v_reg ;
  assign \piso.data_r [2706] = \piso.data_r_2706_sv2v_reg ;
  assign \piso.data_r [2705] = \piso.data_r_2705_sv2v_reg ;
  assign \piso.data_r [2704] = \piso.data_r_2704_sv2v_reg ;
  assign \piso.data_r [2703] = \piso.data_r_2703_sv2v_reg ;
  assign \piso.data_r [2702] = \piso.data_r_2702_sv2v_reg ;
  assign \piso.data_r [2701] = \piso.data_r_2701_sv2v_reg ;
  assign \piso.data_r [2700] = \piso.data_r_2700_sv2v_reg ;
  assign \piso.data_r [2699] = \piso.data_r_2699_sv2v_reg ;
  assign \piso.data_r [2698] = \piso.data_r_2698_sv2v_reg ;
  assign \piso.data_r [2697] = \piso.data_r_2697_sv2v_reg ;
  assign \piso.data_r [2696] = \piso.data_r_2696_sv2v_reg ;
  assign \piso.data_r [2695] = \piso.data_r_2695_sv2v_reg ;
  assign \piso.data_r [2694] = \piso.data_r_2694_sv2v_reg ;
  assign \piso.data_r [2693] = \piso.data_r_2693_sv2v_reg ;
  assign \piso.data_r [2692] = \piso.data_r_2692_sv2v_reg ;
  assign \piso.data_r [2691] = \piso.data_r_2691_sv2v_reg ;
  assign \piso.data_r [2690] = \piso.data_r_2690_sv2v_reg ;
  assign \piso.data_r [2689] = \piso.data_r_2689_sv2v_reg ;
  assign \piso.data_r [2688] = \piso.data_r_2688_sv2v_reg ;
  assign \piso.data_r [2687] = \piso.data_r_2687_sv2v_reg ;
  assign \piso.data_r [2686] = \piso.data_r_2686_sv2v_reg ;
  assign \piso.data_r [2685] = \piso.data_r_2685_sv2v_reg ;
  assign \piso.data_r [2684] = \piso.data_r_2684_sv2v_reg ;
  assign \piso.data_r [2683] = \piso.data_r_2683_sv2v_reg ;
  assign \piso.data_r [2682] = \piso.data_r_2682_sv2v_reg ;
  assign \piso.data_r [2681] = \piso.data_r_2681_sv2v_reg ;
  assign \piso.data_r [2680] = \piso.data_r_2680_sv2v_reg ;
  assign \piso.data_r [2679] = \piso.data_r_2679_sv2v_reg ;
  assign \piso.data_r [2678] = \piso.data_r_2678_sv2v_reg ;
  assign \piso.data_r [2677] = \piso.data_r_2677_sv2v_reg ;
  assign \piso.data_r [2676] = \piso.data_r_2676_sv2v_reg ;
  assign \piso.data_r [2675] = \piso.data_r_2675_sv2v_reg ;
  assign \piso.data_r [2674] = \piso.data_r_2674_sv2v_reg ;
  assign \piso.data_r [2673] = \piso.data_r_2673_sv2v_reg ;
  assign \piso.data_r [2672] = \piso.data_r_2672_sv2v_reg ;
  assign \piso.data_r [2671] = \piso.data_r_2671_sv2v_reg ;
  assign \piso.data_r [2670] = \piso.data_r_2670_sv2v_reg ;
  assign \piso.data_r [2669] = \piso.data_r_2669_sv2v_reg ;
  assign \piso.data_r [2668] = \piso.data_r_2668_sv2v_reg ;
  assign \piso.data_r [2667] = \piso.data_r_2667_sv2v_reg ;
  assign \piso.data_r [2666] = \piso.data_r_2666_sv2v_reg ;
  assign \piso.data_r [2665] = \piso.data_r_2665_sv2v_reg ;
  assign \piso.data_r [2664] = \piso.data_r_2664_sv2v_reg ;
  assign \piso.data_r [2663] = \piso.data_r_2663_sv2v_reg ;
  assign \piso.data_r [2662] = \piso.data_r_2662_sv2v_reg ;
  assign \piso.data_r [2661] = \piso.data_r_2661_sv2v_reg ;
  assign \piso.data_r [2660] = \piso.data_r_2660_sv2v_reg ;
  assign \piso.data_r [2659] = \piso.data_r_2659_sv2v_reg ;
  assign \piso.data_r [2658] = \piso.data_r_2658_sv2v_reg ;
  assign \piso.data_r [2657] = \piso.data_r_2657_sv2v_reg ;
  assign \piso.data_r [2656] = \piso.data_r_2656_sv2v_reg ;
  assign \piso.data_r [2655] = \piso.data_r_2655_sv2v_reg ;
  assign \piso.data_r [2654] = \piso.data_r_2654_sv2v_reg ;
  assign \piso.data_r [2653] = \piso.data_r_2653_sv2v_reg ;
  assign \piso.data_r [2652] = \piso.data_r_2652_sv2v_reg ;
  assign \piso.data_r [2651] = \piso.data_r_2651_sv2v_reg ;
  assign \piso.data_r [2650] = \piso.data_r_2650_sv2v_reg ;
  assign \piso.data_r [2649] = \piso.data_r_2649_sv2v_reg ;
  assign \piso.data_r [2648] = \piso.data_r_2648_sv2v_reg ;
  assign \piso.data_r [2647] = \piso.data_r_2647_sv2v_reg ;
  assign \piso.data_r [2646] = \piso.data_r_2646_sv2v_reg ;
  assign \piso.data_r [2645] = \piso.data_r_2645_sv2v_reg ;
  assign \piso.data_r [2644] = \piso.data_r_2644_sv2v_reg ;
  assign \piso.data_r [2643] = \piso.data_r_2643_sv2v_reg ;
  assign \piso.data_r [2642] = \piso.data_r_2642_sv2v_reg ;
  assign \piso.data_r [2641] = \piso.data_r_2641_sv2v_reg ;
  assign \piso.data_r [2640] = \piso.data_r_2640_sv2v_reg ;
  assign \piso.data_r [2639] = \piso.data_r_2639_sv2v_reg ;
  assign \piso.data_r [2638] = \piso.data_r_2638_sv2v_reg ;
  assign \piso.data_r [2637] = \piso.data_r_2637_sv2v_reg ;
  assign \piso.data_r [2636] = \piso.data_r_2636_sv2v_reg ;
  assign \piso.data_r [2635] = \piso.data_r_2635_sv2v_reg ;
  assign \piso.data_r [2634] = \piso.data_r_2634_sv2v_reg ;
  assign \piso.data_r [2633] = \piso.data_r_2633_sv2v_reg ;
  assign \piso.data_r [2632] = \piso.data_r_2632_sv2v_reg ;
  assign \piso.data_r [2631] = \piso.data_r_2631_sv2v_reg ;
  assign \piso.data_r [2630] = \piso.data_r_2630_sv2v_reg ;
  assign \piso.data_r [2629] = \piso.data_r_2629_sv2v_reg ;
  assign \piso.data_r [2628] = \piso.data_r_2628_sv2v_reg ;
  assign \piso.data_r [2627] = \piso.data_r_2627_sv2v_reg ;
  assign \piso.data_r [2626] = \piso.data_r_2626_sv2v_reg ;
  assign \piso.data_r [2625] = \piso.data_r_2625_sv2v_reg ;
  assign \piso.data_r [2624] = \piso.data_r_2624_sv2v_reg ;
  assign \piso.data_r [2623] = \piso.data_r_2623_sv2v_reg ;
  assign \piso.data_r [2622] = \piso.data_r_2622_sv2v_reg ;
  assign \piso.data_r [2621] = \piso.data_r_2621_sv2v_reg ;
  assign \piso.data_r [2620] = \piso.data_r_2620_sv2v_reg ;
  assign \piso.data_r [2619] = \piso.data_r_2619_sv2v_reg ;
  assign \piso.data_r [2618] = \piso.data_r_2618_sv2v_reg ;
  assign \piso.data_r [2617] = \piso.data_r_2617_sv2v_reg ;
  assign \piso.data_r [2616] = \piso.data_r_2616_sv2v_reg ;
  assign \piso.data_r [2615] = \piso.data_r_2615_sv2v_reg ;
  assign \piso.data_r [2614] = \piso.data_r_2614_sv2v_reg ;
  assign \piso.data_r [2613] = \piso.data_r_2613_sv2v_reg ;
  assign \piso.data_r [2612] = \piso.data_r_2612_sv2v_reg ;
  assign \piso.data_r [2611] = \piso.data_r_2611_sv2v_reg ;
  assign \piso.data_r [2610] = \piso.data_r_2610_sv2v_reg ;
  assign \piso.data_r [2609] = \piso.data_r_2609_sv2v_reg ;
  assign \piso.data_r [2608] = \piso.data_r_2608_sv2v_reg ;
  assign \piso.data_r [2607] = \piso.data_r_2607_sv2v_reg ;
  assign \piso.data_r [2606] = \piso.data_r_2606_sv2v_reg ;
  assign \piso.data_r [2605] = \piso.data_r_2605_sv2v_reg ;
  assign \piso.data_r [2604] = \piso.data_r_2604_sv2v_reg ;
  assign \piso.data_r [2603] = \piso.data_r_2603_sv2v_reg ;
  assign \piso.data_r [2602] = \piso.data_r_2602_sv2v_reg ;
  assign \piso.data_r [2601] = \piso.data_r_2601_sv2v_reg ;
  assign \piso.data_r [2600] = \piso.data_r_2600_sv2v_reg ;
  assign \piso.data_r [2599] = \piso.data_r_2599_sv2v_reg ;
  assign \piso.data_r [2598] = \piso.data_r_2598_sv2v_reg ;
  assign \piso.data_r [2597] = \piso.data_r_2597_sv2v_reg ;
  assign \piso.data_r [2596] = \piso.data_r_2596_sv2v_reg ;
  assign \piso.data_r [2595] = \piso.data_r_2595_sv2v_reg ;
  assign \piso.data_r [2594] = \piso.data_r_2594_sv2v_reg ;
  assign \piso.data_r [2593] = \piso.data_r_2593_sv2v_reg ;
  assign \piso.data_r [2592] = \piso.data_r_2592_sv2v_reg ;
  assign \piso.data_r [2591] = \piso.data_r_2591_sv2v_reg ;
  assign \piso.data_r [2590] = \piso.data_r_2590_sv2v_reg ;
  assign \piso.data_r [2589] = \piso.data_r_2589_sv2v_reg ;
  assign \piso.data_r [2588] = \piso.data_r_2588_sv2v_reg ;
  assign \piso.data_r [2587] = \piso.data_r_2587_sv2v_reg ;
  assign \piso.data_r [2586] = \piso.data_r_2586_sv2v_reg ;
  assign \piso.data_r [2585] = \piso.data_r_2585_sv2v_reg ;
  assign \piso.data_r [2584] = \piso.data_r_2584_sv2v_reg ;
  assign \piso.data_r [2583] = \piso.data_r_2583_sv2v_reg ;
  assign \piso.data_r [2582] = \piso.data_r_2582_sv2v_reg ;
  assign \piso.data_r [2581] = \piso.data_r_2581_sv2v_reg ;
  assign \piso.data_r [2580] = \piso.data_r_2580_sv2v_reg ;
  assign \piso.data_r [2579] = \piso.data_r_2579_sv2v_reg ;
  assign \piso.data_r [2578] = \piso.data_r_2578_sv2v_reg ;
  assign \piso.data_r [2577] = \piso.data_r_2577_sv2v_reg ;
  assign \piso.data_r [2576] = \piso.data_r_2576_sv2v_reg ;
  assign \piso.data_r [2575] = \piso.data_r_2575_sv2v_reg ;
  assign \piso.data_r [2574] = \piso.data_r_2574_sv2v_reg ;
  assign \piso.data_r [2573] = \piso.data_r_2573_sv2v_reg ;
  assign \piso.data_r [2572] = \piso.data_r_2572_sv2v_reg ;
  assign \piso.data_r [2571] = \piso.data_r_2571_sv2v_reg ;
  assign \piso.data_r [2570] = \piso.data_r_2570_sv2v_reg ;
  assign \piso.data_r [2569] = \piso.data_r_2569_sv2v_reg ;
  assign \piso.data_r [2568] = \piso.data_r_2568_sv2v_reg ;
  assign \piso.data_r [2567] = \piso.data_r_2567_sv2v_reg ;
  assign \piso.data_r [2566] = \piso.data_r_2566_sv2v_reg ;
  assign \piso.data_r [2565] = \piso.data_r_2565_sv2v_reg ;
  assign \piso.data_r [2564] = \piso.data_r_2564_sv2v_reg ;
  assign \piso.data_r [2563] = \piso.data_r_2563_sv2v_reg ;
  assign \piso.data_r [2562] = \piso.data_r_2562_sv2v_reg ;
  assign \piso.data_r [2561] = \piso.data_r_2561_sv2v_reg ;
  assign \piso.data_r [2560] = \piso.data_r_2560_sv2v_reg ;
  assign \piso.data_r [2559] = \piso.data_r_2559_sv2v_reg ;
  assign \piso.data_r [2558] = \piso.data_r_2558_sv2v_reg ;
  assign \piso.data_r [2557] = \piso.data_r_2557_sv2v_reg ;
  assign \piso.data_r [2556] = \piso.data_r_2556_sv2v_reg ;
  assign \piso.data_r [2555] = \piso.data_r_2555_sv2v_reg ;
  assign \piso.data_r [2554] = \piso.data_r_2554_sv2v_reg ;
  assign \piso.data_r [2553] = \piso.data_r_2553_sv2v_reg ;
  assign \piso.data_r [2552] = \piso.data_r_2552_sv2v_reg ;
  assign \piso.data_r [2551] = \piso.data_r_2551_sv2v_reg ;
  assign \piso.data_r [2550] = \piso.data_r_2550_sv2v_reg ;
  assign \piso.data_r [2549] = \piso.data_r_2549_sv2v_reg ;
  assign \piso.data_r [2548] = \piso.data_r_2548_sv2v_reg ;
  assign \piso.data_r [2547] = \piso.data_r_2547_sv2v_reg ;
  assign \piso.data_r [2546] = \piso.data_r_2546_sv2v_reg ;
  assign \piso.data_r [2545] = \piso.data_r_2545_sv2v_reg ;
  assign \piso.data_r [2544] = \piso.data_r_2544_sv2v_reg ;
  assign \piso.data_r [2543] = \piso.data_r_2543_sv2v_reg ;
  assign \piso.data_r [2542] = \piso.data_r_2542_sv2v_reg ;
  assign \piso.data_r [2541] = \piso.data_r_2541_sv2v_reg ;
  assign \piso.data_r [2540] = \piso.data_r_2540_sv2v_reg ;
  assign \piso.data_r [2539] = \piso.data_r_2539_sv2v_reg ;
  assign \piso.data_r [2538] = \piso.data_r_2538_sv2v_reg ;
  assign \piso.data_r [2537] = \piso.data_r_2537_sv2v_reg ;
  assign \piso.data_r [2536] = \piso.data_r_2536_sv2v_reg ;
  assign \piso.data_r [2535] = \piso.data_r_2535_sv2v_reg ;
  assign \piso.data_r [2534] = \piso.data_r_2534_sv2v_reg ;
  assign \piso.data_r [2533] = \piso.data_r_2533_sv2v_reg ;
  assign \piso.data_r [2532] = \piso.data_r_2532_sv2v_reg ;
  assign \piso.data_r [2531] = \piso.data_r_2531_sv2v_reg ;
  assign \piso.data_r [2530] = \piso.data_r_2530_sv2v_reg ;
  assign \piso.data_r [2529] = \piso.data_r_2529_sv2v_reg ;
  assign \piso.data_r [2528] = \piso.data_r_2528_sv2v_reg ;
  assign \piso.data_r [2527] = \piso.data_r_2527_sv2v_reg ;
  assign \piso.data_r [2526] = \piso.data_r_2526_sv2v_reg ;
  assign \piso.data_r [2525] = \piso.data_r_2525_sv2v_reg ;
  assign \piso.data_r [2524] = \piso.data_r_2524_sv2v_reg ;
  assign \piso.data_r [2523] = \piso.data_r_2523_sv2v_reg ;
  assign \piso.data_r [2522] = \piso.data_r_2522_sv2v_reg ;
  assign \piso.data_r [2521] = \piso.data_r_2521_sv2v_reg ;
  assign \piso.data_r [2520] = \piso.data_r_2520_sv2v_reg ;
  assign \piso.data_r [2519] = \piso.data_r_2519_sv2v_reg ;
  assign \piso.data_r [2518] = \piso.data_r_2518_sv2v_reg ;
  assign \piso.data_r [2517] = \piso.data_r_2517_sv2v_reg ;
  assign \piso.data_r [2516] = \piso.data_r_2516_sv2v_reg ;
  assign \piso.data_r [2515] = \piso.data_r_2515_sv2v_reg ;
  assign \piso.data_r [2514] = \piso.data_r_2514_sv2v_reg ;
  assign \piso.data_r [2513] = \piso.data_r_2513_sv2v_reg ;
  assign \piso.data_r [2512] = \piso.data_r_2512_sv2v_reg ;
  assign \piso.data_r [2511] = \piso.data_r_2511_sv2v_reg ;
  assign \piso.data_r [2510] = \piso.data_r_2510_sv2v_reg ;
  assign \piso.data_r [2509] = \piso.data_r_2509_sv2v_reg ;
  assign \piso.data_r [2508] = \piso.data_r_2508_sv2v_reg ;
  assign \piso.data_r [2507] = \piso.data_r_2507_sv2v_reg ;
  assign \piso.data_r [2506] = \piso.data_r_2506_sv2v_reg ;
  assign \piso.data_r [2505] = \piso.data_r_2505_sv2v_reg ;
  assign \piso.data_r [2504] = \piso.data_r_2504_sv2v_reg ;
  assign \piso.data_r [2503] = \piso.data_r_2503_sv2v_reg ;
  assign \piso.data_r [2502] = \piso.data_r_2502_sv2v_reg ;
  assign \piso.data_r [2501] = \piso.data_r_2501_sv2v_reg ;
  assign \piso.data_r [2500] = \piso.data_r_2500_sv2v_reg ;
  assign \piso.data_r [2499] = \piso.data_r_2499_sv2v_reg ;
  assign \piso.data_r [2498] = \piso.data_r_2498_sv2v_reg ;
  assign \piso.data_r [2497] = \piso.data_r_2497_sv2v_reg ;
  assign \piso.data_r [2496] = \piso.data_r_2496_sv2v_reg ;
  assign \piso.data_r [2495] = \piso.data_r_2495_sv2v_reg ;
  assign \piso.data_r [2494] = \piso.data_r_2494_sv2v_reg ;
  assign \piso.data_r [2493] = \piso.data_r_2493_sv2v_reg ;
  assign \piso.data_r [2492] = \piso.data_r_2492_sv2v_reg ;
  assign \piso.data_r [2491] = \piso.data_r_2491_sv2v_reg ;
  assign \piso.data_r [2490] = \piso.data_r_2490_sv2v_reg ;
  assign \piso.data_r [2489] = \piso.data_r_2489_sv2v_reg ;
  assign \piso.data_r [2488] = \piso.data_r_2488_sv2v_reg ;
  assign \piso.data_r [2487] = \piso.data_r_2487_sv2v_reg ;
  assign \piso.data_r [2486] = \piso.data_r_2486_sv2v_reg ;
  assign \piso.data_r [2485] = \piso.data_r_2485_sv2v_reg ;
  assign \piso.data_r [2484] = \piso.data_r_2484_sv2v_reg ;
  assign \piso.data_r [2483] = \piso.data_r_2483_sv2v_reg ;
  assign \piso.data_r [2482] = \piso.data_r_2482_sv2v_reg ;
  assign \piso.data_r [2481] = \piso.data_r_2481_sv2v_reg ;
  assign \piso.data_r [2480] = \piso.data_r_2480_sv2v_reg ;
  assign \piso.data_r [2479] = \piso.data_r_2479_sv2v_reg ;
  assign \piso.data_r [2478] = \piso.data_r_2478_sv2v_reg ;
  assign \piso.data_r [2477] = \piso.data_r_2477_sv2v_reg ;
  assign \piso.data_r [2476] = \piso.data_r_2476_sv2v_reg ;
  assign \piso.data_r [2475] = \piso.data_r_2475_sv2v_reg ;
  assign \piso.data_r [2474] = \piso.data_r_2474_sv2v_reg ;
  assign \piso.data_r [2473] = \piso.data_r_2473_sv2v_reg ;
  assign \piso.data_r [2472] = \piso.data_r_2472_sv2v_reg ;
  assign \piso.data_r [2471] = \piso.data_r_2471_sv2v_reg ;
  assign \piso.data_r [2470] = \piso.data_r_2470_sv2v_reg ;
  assign \piso.data_r [2469] = \piso.data_r_2469_sv2v_reg ;
  assign \piso.data_r [2468] = \piso.data_r_2468_sv2v_reg ;
  assign \piso.data_r [2467] = \piso.data_r_2467_sv2v_reg ;
  assign \piso.data_r [2466] = \piso.data_r_2466_sv2v_reg ;
  assign \piso.data_r [2465] = \piso.data_r_2465_sv2v_reg ;
  assign \piso.data_r [2464] = \piso.data_r_2464_sv2v_reg ;
  assign \piso.data_r [2463] = \piso.data_r_2463_sv2v_reg ;
  assign \piso.data_r [2462] = \piso.data_r_2462_sv2v_reg ;
  assign \piso.data_r [2461] = \piso.data_r_2461_sv2v_reg ;
  assign \piso.data_r [2460] = \piso.data_r_2460_sv2v_reg ;
  assign \piso.data_r [2459] = \piso.data_r_2459_sv2v_reg ;
  assign \piso.data_r [2458] = \piso.data_r_2458_sv2v_reg ;
  assign \piso.data_r [2457] = \piso.data_r_2457_sv2v_reg ;
  assign \piso.data_r [2456] = \piso.data_r_2456_sv2v_reg ;
  assign \piso.data_r [2455] = \piso.data_r_2455_sv2v_reg ;
  assign \piso.data_r [2454] = \piso.data_r_2454_sv2v_reg ;
  assign \piso.data_r [2453] = \piso.data_r_2453_sv2v_reg ;
  assign \piso.data_r [2452] = \piso.data_r_2452_sv2v_reg ;
  assign \piso.data_r [2451] = \piso.data_r_2451_sv2v_reg ;
  assign \piso.data_r [2450] = \piso.data_r_2450_sv2v_reg ;
  assign \piso.data_r [2449] = \piso.data_r_2449_sv2v_reg ;
  assign \piso.data_r [2448] = \piso.data_r_2448_sv2v_reg ;
  assign \piso.data_r [2447] = \piso.data_r_2447_sv2v_reg ;
  assign \piso.data_r [2446] = \piso.data_r_2446_sv2v_reg ;
  assign \piso.data_r [2445] = \piso.data_r_2445_sv2v_reg ;
  assign \piso.data_r [2444] = \piso.data_r_2444_sv2v_reg ;
  assign \piso.data_r [2443] = \piso.data_r_2443_sv2v_reg ;
  assign \piso.data_r [2442] = \piso.data_r_2442_sv2v_reg ;
  assign \piso.data_r [2441] = \piso.data_r_2441_sv2v_reg ;
  assign \piso.data_r [2440] = \piso.data_r_2440_sv2v_reg ;
  assign \piso.data_r [2439] = \piso.data_r_2439_sv2v_reg ;
  assign \piso.data_r [2438] = \piso.data_r_2438_sv2v_reg ;
  assign \piso.data_r [2437] = \piso.data_r_2437_sv2v_reg ;
  assign \piso.data_r [2436] = \piso.data_r_2436_sv2v_reg ;
  assign \piso.data_r [2435] = \piso.data_r_2435_sv2v_reg ;
  assign \piso.data_r [2434] = \piso.data_r_2434_sv2v_reg ;
  assign \piso.data_r [2433] = \piso.data_r_2433_sv2v_reg ;
  assign \piso.data_r [2432] = \piso.data_r_2432_sv2v_reg ;
  assign \piso.data_r [2431] = \piso.data_r_2431_sv2v_reg ;
  assign \piso.data_r [2430] = \piso.data_r_2430_sv2v_reg ;
  assign \piso.data_r [2429] = \piso.data_r_2429_sv2v_reg ;
  assign \piso.data_r [2428] = \piso.data_r_2428_sv2v_reg ;
  assign \piso.data_r [2427] = \piso.data_r_2427_sv2v_reg ;
  assign \piso.data_r [2426] = \piso.data_r_2426_sv2v_reg ;
  assign \piso.data_r [2425] = \piso.data_r_2425_sv2v_reg ;
  assign \piso.data_r [2424] = \piso.data_r_2424_sv2v_reg ;
  assign \piso.data_r [2423] = \piso.data_r_2423_sv2v_reg ;
  assign \piso.data_r [2422] = \piso.data_r_2422_sv2v_reg ;
  assign \piso.data_r [2421] = \piso.data_r_2421_sv2v_reg ;
  assign \piso.data_r [2420] = \piso.data_r_2420_sv2v_reg ;
  assign \piso.data_r [2419] = \piso.data_r_2419_sv2v_reg ;
  assign \piso.data_r [2418] = \piso.data_r_2418_sv2v_reg ;
  assign \piso.data_r [2417] = \piso.data_r_2417_sv2v_reg ;
  assign \piso.data_r [2416] = \piso.data_r_2416_sv2v_reg ;
  assign \piso.data_r [2415] = \piso.data_r_2415_sv2v_reg ;
  assign \piso.data_r [2414] = \piso.data_r_2414_sv2v_reg ;
  assign \piso.data_r [2413] = \piso.data_r_2413_sv2v_reg ;
  assign \piso.data_r [2412] = \piso.data_r_2412_sv2v_reg ;
  assign \piso.data_r [2411] = \piso.data_r_2411_sv2v_reg ;
  assign \piso.data_r [2410] = \piso.data_r_2410_sv2v_reg ;
  assign \piso.data_r [2409] = \piso.data_r_2409_sv2v_reg ;
  assign \piso.data_r [2408] = \piso.data_r_2408_sv2v_reg ;
  assign \piso.data_r [2407] = \piso.data_r_2407_sv2v_reg ;
  assign \piso.data_r [2406] = \piso.data_r_2406_sv2v_reg ;
  assign \piso.data_r [2405] = \piso.data_r_2405_sv2v_reg ;
  assign \piso.data_r [2404] = \piso.data_r_2404_sv2v_reg ;
  assign \piso.data_r [2403] = \piso.data_r_2403_sv2v_reg ;
  assign \piso.data_r [2402] = \piso.data_r_2402_sv2v_reg ;
  assign \piso.data_r [2401] = \piso.data_r_2401_sv2v_reg ;
  assign \piso.data_r [2400] = \piso.data_r_2400_sv2v_reg ;
  assign \piso.data_r [2399] = \piso.data_r_2399_sv2v_reg ;
  assign \piso.data_r [2398] = \piso.data_r_2398_sv2v_reg ;
  assign \piso.data_r [2397] = \piso.data_r_2397_sv2v_reg ;
  assign \piso.data_r [2396] = \piso.data_r_2396_sv2v_reg ;
  assign \piso.data_r [2395] = \piso.data_r_2395_sv2v_reg ;
  assign \piso.data_r [2394] = \piso.data_r_2394_sv2v_reg ;
  assign \piso.data_r [2393] = \piso.data_r_2393_sv2v_reg ;
  assign \piso.data_r [2392] = \piso.data_r_2392_sv2v_reg ;
  assign \piso.data_r [2391] = \piso.data_r_2391_sv2v_reg ;
  assign \piso.data_r [2390] = \piso.data_r_2390_sv2v_reg ;
  assign \piso.data_r [2389] = \piso.data_r_2389_sv2v_reg ;
  assign \piso.data_r [2388] = \piso.data_r_2388_sv2v_reg ;
  assign \piso.data_r [2387] = \piso.data_r_2387_sv2v_reg ;
  assign \piso.data_r [2386] = \piso.data_r_2386_sv2v_reg ;
  assign \piso.data_r [2385] = \piso.data_r_2385_sv2v_reg ;
  assign \piso.data_r [2384] = \piso.data_r_2384_sv2v_reg ;
  assign \piso.data_r [2383] = \piso.data_r_2383_sv2v_reg ;
  assign \piso.data_r [2382] = \piso.data_r_2382_sv2v_reg ;
  assign \piso.data_r [2381] = \piso.data_r_2381_sv2v_reg ;
  assign \piso.data_r [2380] = \piso.data_r_2380_sv2v_reg ;
  assign \piso.data_r [2379] = \piso.data_r_2379_sv2v_reg ;
  assign \piso.data_r [2378] = \piso.data_r_2378_sv2v_reg ;
  assign \piso.data_r [2377] = \piso.data_r_2377_sv2v_reg ;
  assign \piso.data_r [2376] = \piso.data_r_2376_sv2v_reg ;
  assign \piso.data_r [2375] = \piso.data_r_2375_sv2v_reg ;
  assign \piso.data_r [2374] = \piso.data_r_2374_sv2v_reg ;
  assign \piso.data_r [2373] = \piso.data_r_2373_sv2v_reg ;
  assign \piso.data_r [2372] = \piso.data_r_2372_sv2v_reg ;
  assign \piso.data_r [2371] = \piso.data_r_2371_sv2v_reg ;
  assign \piso.data_r [2370] = \piso.data_r_2370_sv2v_reg ;
  assign \piso.data_r [2369] = \piso.data_r_2369_sv2v_reg ;
  assign \piso.data_r [2368] = \piso.data_r_2368_sv2v_reg ;
  assign \piso.data_r [2367] = \piso.data_r_2367_sv2v_reg ;
  assign \piso.data_r [2366] = \piso.data_r_2366_sv2v_reg ;
  assign \piso.data_r [2365] = \piso.data_r_2365_sv2v_reg ;
  assign \piso.data_r [2364] = \piso.data_r_2364_sv2v_reg ;
  assign \piso.data_r [2363] = \piso.data_r_2363_sv2v_reg ;
  assign \piso.data_r [2362] = \piso.data_r_2362_sv2v_reg ;
  assign \piso.data_r [2361] = \piso.data_r_2361_sv2v_reg ;
  assign \piso.data_r [2360] = \piso.data_r_2360_sv2v_reg ;
  assign \piso.data_r [2359] = \piso.data_r_2359_sv2v_reg ;
  assign \piso.data_r [2358] = \piso.data_r_2358_sv2v_reg ;
  assign \piso.data_r [2357] = \piso.data_r_2357_sv2v_reg ;
  assign \piso.data_r [2356] = \piso.data_r_2356_sv2v_reg ;
  assign \piso.data_r [2355] = \piso.data_r_2355_sv2v_reg ;
  assign \piso.data_r [2354] = \piso.data_r_2354_sv2v_reg ;
  assign \piso.data_r [2353] = \piso.data_r_2353_sv2v_reg ;
  assign \piso.data_r [2352] = \piso.data_r_2352_sv2v_reg ;
  assign \piso.data_r [2351] = \piso.data_r_2351_sv2v_reg ;
  assign \piso.data_r [2350] = \piso.data_r_2350_sv2v_reg ;
  assign \piso.data_r [2349] = \piso.data_r_2349_sv2v_reg ;
  assign \piso.data_r [2348] = \piso.data_r_2348_sv2v_reg ;
  assign \piso.data_r [2347] = \piso.data_r_2347_sv2v_reg ;
  assign \piso.data_r [2346] = \piso.data_r_2346_sv2v_reg ;
  assign \piso.data_r [2345] = \piso.data_r_2345_sv2v_reg ;
  assign \piso.data_r [2344] = \piso.data_r_2344_sv2v_reg ;
  assign \piso.data_r [2343] = \piso.data_r_2343_sv2v_reg ;
  assign \piso.data_r [2342] = \piso.data_r_2342_sv2v_reg ;
  assign \piso.data_r [2341] = \piso.data_r_2341_sv2v_reg ;
  assign \piso.data_r [2340] = \piso.data_r_2340_sv2v_reg ;
  assign \piso.data_r [2339] = \piso.data_r_2339_sv2v_reg ;
  assign \piso.data_r [2338] = \piso.data_r_2338_sv2v_reg ;
  assign \piso.data_r [2337] = \piso.data_r_2337_sv2v_reg ;
  assign \piso.data_r [2336] = \piso.data_r_2336_sv2v_reg ;
  assign \piso.data_r [2335] = \piso.data_r_2335_sv2v_reg ;
  assign \piso.data_r [2334] = \piso.data_r_2334_sv2v_reg ;
  assign \piso.data_r [2333] = \piso.data_r_2333_sv2v_reg ;
  assign \piso.data_r [2332] = \piso.data_r_2332_sv2v_reg ;
  assign \piso.data_r [2331] = \piso.data_r_2331_sv2v_reg ;
  assign \piso.data_r [2330] = \piso.data_r_2330_sv2v_reg ;
  assign \piso.data_r [2329] = \piso.data_r_2329_sv2v_reg ;
  assign \piso.data_r [2328] = \piso.data_r_2328_sv2v_reg ;
  assign \piso.data_r [2327] = \piso.data_r_2327_sv2v_reg ;
  assign \piso.data_r [2326] = \piso.data_r_2326_sv2v_reg ;
  assign \piso.data_r [2325] = \piso.data_r_2325_sv2v_reg ;
  assign \piso.data_r [2324] = \piso.data_r_2324_sv2v_reg ;
  assign \piso.data_r [2323] = \piso.data_r_2323_sv2v_reg ;
  assign \piso.data_r [2322] = \piso.data_r_2322_sv2v_reg ;
  assign \piso.data_r [2321] = \piso.data_r_2321_sv2v_reg ;
  assign \piso.data_r [2320] = \piso.data_r_2320_sv2v_reg ;
  assign \piso.data_r [2319] = \piso.data_r_2319_sv2v_reg ;
  assign \piso.data_r [2318] = \piso.data_r_2318_sv2v_reg ;
  assign \piso.data_r [2317] = \piso.data_r_2317_sv2v_reg ;
  assign \piso.data_r [2316] = \piso.data_r_2316_sv2v_reg ;
  assign \piso.data_r [2315] = \piso.data_r_2315_sv2v_reg ;
  assign \piso.data_r [2314] = \piso.data_r_2314_sv2v_reg ;
  assign \piso.data_r [2313] = \piso.data_r_2313_sv2v_reg ;
  assign \piso.data_r [2312] = \piso.data_r_2312_sv2v_reg ;
  assign \piso.data_r [2311] = \piso.data_r_2311_sv2v_reg ;
  assign \piso.data_r [2310] = \piso.data_r_2310_sv2v_reg ;
  assign \piso.data_r [2309] = \piso.data_r_2309_sv2v_reg ;
  assign \piso.data_r [2308] = \piso.data_r_2308_sv2v_reg ;
  assign \piso.data_r [2307] = \piso.data_r_2307_sv2v_reg ;
  assign \piso.data_r [2306] = \piso.data_r_2306_sv2v_reg ;
  assign \piso.data_r [2305] = \piso.data_r_2305_sv2v_reg ;
  assign \piso.data_r [2304] = \piso.data_r_2304_sv2v_reg ;
  assign \piso.data_r [2303] = \piso.data_r_2303_sv2v_reg ;
  assign \piso.data_r [2302] = \piso.data_r_2302_sv2v_reg ;
  assign \piso.data_r [2301] = \piso.data_r_2301_sv2v_reg ;
  assign \piso.data_r [2300] = \piso.data_r_2300_sv2v_reg ;
  assign \piso.data_r [2299] = \piso.data_r_2299_sv2v_reg ;
  assign \piso.data_r [2298] = \piso.data_r_2298_sv2v_reg ;
  assign \piso.data_r [2297] = \piso.data_r_2297_sv2v_reg ;
  assign \piso.data_r [2296] = \piso.data_r_2296_sv2v_reg ;
  assign \piso.data_r [2295] = \piso.data_r_2295_sv2v_reg ;
  assign \piso.data_r [2294] = \piso.data_r_2294_sv2v_reg ;
  assign \piso.data_r [2293] = \piso.data_r_2293_sv2v_reg ;
  assign \piso.data_r [2292] = \piso.data_r_2292_sv2v_reg ;
  assign \piso.data_r [2291] = \piso.data_r_2291_sv2v_reg ;
  assign \piso.data_r [2290] = \piso.data_r_2290_sv2v_reg ;
  assign \piso.data_r [2289] = \piso.data_r_2289_sv2v_reg ;
  assign \piso.data_r [2288] = \piso.data_r_2288_sv2v_reg ;
  assign \piso.data_r [2287] = \piso.data_r_2287_sv2v_reg ;
  assign \piso.data_r [2286] = \piso.data_r_2286_sv2v_reg ;
  assign \piso.data_r [2285] = \piso.data_r_2285_sv2v_reg ;
  assign \piso.data_r [2284] = \piso.data_r_2284_sv2v_reg ;
  assign \piso.data_r [2283] = \piso.data_r_2283_sv2v_reg ;
  assign \piso.data_r [2282] = \piso.data_r_2282_sv2v_reg ;
  assign \piso.data_r [2281] = \piso.data_r_2281_sv2v_reg ;
  assign \piso.data_r [2280] = \piso.data_r_2280_sv2v_reg ;
  assign \piso.data_r [2279] = \piso.data_r_2279_sv2v_reg ;
  assign \piso.data_r [2278] = \piso.data_r_2278_sv2v_reg ;
  assign \piso.data_r [2277] = \piso.data_r_2277_sv2v_reg ;
  assign \piso.data_r [2276] = \piso.data_r_2276_sv2v_reg ;
  assign \piso.data_r [2275] = \piso.data_r_2275_sv2v_reg ;
  assign \piso.data_r [2274] = \piso.data_r_2274_sv2v_reg ;
  assign \piso.data_r [2273] = \piso.data_r_2273_sv2v_reg ;
  assign \piso.data_r [2272] = \piso.data_r_2272_sv2v_reg ;
  assign \piso.data_r [2271] = \piso.data_r_2271_sv2v_reg ;
  assign \piso.data_r [2270] = \piso.data_r_2270_sv2v_reg ;
  assign \piso.data_r [2269] = \piso.data_r_2269_sv2v_reg ;
  assign \piso.data_r [2268] = \piso.data_r_2268_sv2v_reg ;
  assign \piso.data_r [2267] = \piso.data_r_2267_sv2v_reg ;
  assign \piso.data_r [2266] = \piso.data_r_2266_sv2v_reg ;
  assign \piso.data_r [2265] = \piso.data_r_2265_sv2v_reg ;
  assign \piso.data_r [2264] = \piso.data_r_2264_sv2v_reg ;
  assign \piso.data_r [2263] = \piso.data_r_2263_sv2v_reg ;
  assign \piso.data_r [2262] = \piso.data_r_2262_sv2v_reg ;
  assign \piso.data_r [2261] = \piso.data_r_2261_sv2v_reg ;
  assign \piso.data_r [2260] = \piso.data_r_2260_sv2v_reg ;
  assign \piso.data_r [2259] = \piso.data_r_2259_sv2v_reg ;
  assign \piso.data_r [2258] = \piso.data_r_2258_sv2v_reg ;
  assign \piso.data_r [2257] = \piso.data_r_2257_sv2v_reg ;
  assign \piso.data_r [2256] = \piso.data_r_2256_sv2v_reg ;
  assign \piso.data_r [2255] = \piso.data_r_2255_sv2v_reg ;
  assign \piso.data_r [2254] = \piso.data_r_2254_sv2v_reg ;
  assign \piso.data_r [2253] = \piso.data_r_2253_sv2v_reg ;
  assign \piso.data_r [2252] = \piso.data_r_2252_sv2v_reg ;
  assign \piso.data_r [2251] = \piso.data_r_2251_sv2v_reg ;
  assign \piso.data_r [2250] = \piso.data_r_2250_sv2v_reg ;
  assign \piso.data_r [2249] = \piso.data_r_2249_sv2v_reg ;
  assign \piso.data_r [2248] = \piso.data_r_2248_sv2v_reg ;
  assign \piso.data_r [2247] = \piso.data_r_2247_sv2v_reg ;
  assign \piso.data_r [2246] = \piso.data_r_2246_sv2v_reg ;
  assign \piso.data_r [2245] = \piso.data_r_2245_sv2v_reg ;
  assign \piso.data_r [2244] = \piso.data_r_2244_sv2v_reg ;
  assign \piso.data_r [2243] = \piso.data_r_2243_sv2v_reg ;
  assign \piso.data_r [2242] = \piso.data_r_2242_sv2v_reg ;
  assign \piso.data_r [2241] = \piso.data_r_2241_sv2v_reg ;
  assign \piso.data_r [2240] = \piso.data_r_2240_sv2v_reg ;
  assign \piso.data_r [2239] = \piso.data_r_2239_sv2v_reg ;
  assign \piso.data_r [2238] = \piso.data_r_2238_sv2v_reg ;
  assign \piso.data_r [2237] = \piso.data_r_2237_sv2v_reg ;
  assign \piso.data_r [2236] = \piso.data_r_2236_sv2v_reg ;
  assign \piso.data_r [2235] = \piso.data_r_2235_sv2v_reg ;
  assign \piso.data_r [2234] = \piso.data_r_2234_sv2v_reg ;
  assign \piso.data_r [2233] = \piso.data_r_2233_sv2v_reg ;
  assign \piso.data_r [2232] = \piso.data_r_2232_sv2v_reg ;
  assign \piso.data_r [2231] = \piso.data_r_2231_sv2v_reg ;
  assign \piso.data_r [2230] = \piso.data_r_2230_sv2v_reg ;
  assign \piso.data_r [2229] = \piso.data_r_2229_sv2v_reg ;
  assign \piso.data_r [2228] = \piso.data_r_2228_sv2v_reg ;
  assign \piso.data_r [2227] = \piso.data_r_2227_sv2v_reg ;
  assign \piso.data_r [2226] = \piso.data_r_2226_sv2v_reg ;
  assign \piso.data_r [2225] = \piso.data_r_2225_sv2v_reg ;
  assign \piso.data_r [2224] = \piso.data_r_2224_sv2v_reg ;
  assign \piso.data_r [2223] = \piso.data_r_2223_sv2v_reg ;
  assign \piso.data_r [2222] = \piso.data_r_2222_sv2v_reg ;
  assign \piso.data_r [2221] = \piso.data_r_2221_sv2v_reg ;
  assign \piso.data_r [2220] = \piso.data_r_2220_sv2v_reg ;
  assign \piso.data_r [2219] = \piso.data_r_2219_sv2v_reg ;
  assign \piso.data_r [2218] = \piso.data_r_2218_sv2v_reg ;
  assign \piso.data_r [2217] = \piso.data_r_2217_sv2v_reg ;
  assign \piso.data_r [2216] = \piso.data_r_2216_sv2v_reg ;
  assign \piso.data_r [2215] = \piso.data_r_2215_sv2v_reg ;
  assign \piso.data_r [2214] = \piso.data_r_2214_sv2v_reg ;
  assign \piso.data_r [2213] = \piso.data_r_2213_sv2v_reg ;
  assign \piso.data_r [2212] = \piso.data_r_2212_sv2v_reg ;
  assign \piso.data_r [2211] = \piso.data_r_2211_sv2v_reg ;
  assign \piso.data_r [2210] = \piso.data_r_2210_sv2v_reg ;
  assign \piso.data_r [2209] = \piso.data_r_2209_sv2v_reg ;
  assign \piso.data_r [2208] = \piso.data_r_2208_sv2v_reg ;
  assign \piso.data_r [2207] = \piso.data_r_2207_sv2v_reg ;
  assign \piso.data_r [2206] = \piso.data_r_2206_sv2v_reg ;
  assign \piso.data_r [2205] = \piso.data_r_2205_sv2v_reg ;
  assign \piso.data_r [2204] = \piso.data_r_2204_sv2v_reg ;
  assign \piso.data_r [2203] = \piso.data_r_2203_sv2v_reg ;
  assign \piso.data_r [2202] = \piso.data_r_2202_sv2v_reg ;
  assign \piso.data_r [2201] = \piso.data_r_2201_sv2v_reg ;
  assign \piso.data_r [2200] = \piso.data_r_2200_sv2v_reg ;
  assign \piso.data_r [2199] = \piso.data_r_2199_sv2v_reg ;
  assign \piso.data_r [2198] = \piso.data_r_2198_sv2v_reg ;
  assign \piso.data_r [2197] = \piso.data_r_2197_sv2v_reg ;
  assign \piso.data_r [2196] = \piso.data_r_2196_sv2v_reg ;
  assign \piso.data_r [2195] = \piso.data_r_2195_sv2v_reg ;
  assign \piso.data_r [2194] = \piso.data_r_2194_sv2v_reg ;
  assign \piso.data_r [2193] = \piso.data_r_2193_sv2v_reg ;
  assign \piso.data_r [2192] = \piso.data_r_2192_sv2v_reg ;
  assign \piso.data_r [2191] = \piso.data_r_2191_sv2v_reg ;
  assign \piso.data_r [2190] = \piso.data_r_2190_sv2v_reg ;
  assign \piso.data_r [2189] = \piso.data_r_2189_sv2v_reg ;
  assign \piso.data_r [2188] = \piso.data_r_2188_sv2v_reg ;
  assign \piso.data_r [2187] = \piso.data_r_2187_sv2v_reg ;
  assign \piso.data_r [2186] = \piso.data_r_2186_sv2v_reg ;
  assign \piso.data_r [2185] = \piso.data_r_2185_sv2v_reg ;
  assign \piso.data_r [2184] = \piso.data_r_2184_sv2v_reg ;
  assign \piso.data_r [2183] = \piso.data_r_2183_sv2v_reg ;
  assign \piso.data_r [2182] = \piso.data_r_2182_sv2v_reg ;
  assign \piso.data_r [2181] = \piso.data_r_2181_sv2v_reg ;
  assign \piso.data_r [2180] = \piso.data_r_2180_sv2v_reg ;
  assign \piso.data_r [2179] = \piso.data_r_2179_sv2v_reg ;
  assign \piso.data_r [2178] = \piso.data_r_2178_sv2v_reg ;
  assign \piso.data_r [2177] = \piso.data_r_2177_sv2v_reg ;
  assign \piso.data_r [2176] = \piso.data_r_2176_sv2v_reg ;
  assign \piso.data_r [2175] = \piso.data_r_2175_sv2v_reg ;
  assign \piso.data_r [2174] = \piso.data_r_2174_sv2v_reg ;
  assign \piso.data_r [2173] = \piso.data_r_2173_sv2v_reg ;
  assign \piso.data_r [2172] = \piso.data_r_2172_sv2v_reg ;
  assign \piso.data_r [2171] = \piso.data_r_2171_sv2v_reg ;
  assign \piso.data_r [2170] = \piso.data_r_2170_sv2v_reg ;
  assign \piso.data_r [2169] = \piso.data_r_2169_sv2v_reg ;
  assign \piso.data_r [2168] = \piso.data_r_2168_sv2v_reg ;
  assign \piso.data_r [2167] = \piso.data_r_2167_sv2v_reg ;
  assign \piso.data_r [2166] = \piso.data_r_2166_sv2v_reg ;
  assign \piso.data_r [2165] = \piso.data_r_2165_sv2v_reg ;
  assign \piso.data_r [2164] = \piso.data_r_2164_sv2v_reg ;
  assign \piso.data_r [2163] = \piso.data_r_2163_sv2v_reg ;
  assign \piso.data_r [2162] = \piso.data_r_2162_sv2v_reg ;
  assign \piso.data_r [2161] = \piso.data_r_2161_sv2v_reg ;
  assign \piso.data_r [2160] = \piso.data_r_2160_sv2v_reg ;
  assign \piso.data_r [2159] = \piso.data_r_2159_sv2v_reg ;
  assign \piso.data_r [2158] = \piso.data_r_2158_sv2v_reg ;
  assign \piso.data_r [2157] = \piso.data_r_2157_sv2v_reg ;
  assign \piso.data_r [2156] = \piso.data_r_2156_sv2v_reg ;
  assign \piso.data_r [2155] = \piso.data_r_2155_sv2v_reg ;
  assign \piso.data_r [2154] = \piso.data_r_2154_sv2v_reg ;
  assign \piso.data_r [2153] = \piso.data_r_2153_sv2v_reg ;
  assign \piso.data_r [2152] = \piso.data_r_2152_sv2v_reg ;
  assign \piso.data_r [2151] = \piso.data_r_2151_sv2v_reg ;
  assign \piso.data_r [2150] = \piso.data_r_2150_sv2v_reg ;
  assign \piso.data_r [2149] = \piso.data_r_2149_sv2v_reg ;
  assign \piso.data_r [2148] = \piso.data_r_2148_sv2v_reg ;
  assign \piso.data_r [2147] = \piso.data_r_2147_sv2v_reg ;
  assign \piso.data_r [2146] = \piso.data_r_2146_sv2v_reg ;
  assign \piso.data_r [2145] = \piso.data_r_2145_sv2v_reg ;
  assign \piso.data_r [2144] = \piso.data_r_2144_sv2v_reg ;
  assign \piso.data_r [2143] = \piso.data_r_2143_sv2v_reg ;
  assign \piso.data_r [2142] = \piso.data_r_2142_sv2v_reg ;
  assign \piso.data_r [2141] = \piso.data_r_2141_sv2v_reg ;
  assign \piso.data_r [2140] = \piso.data_r_2140_sv2v_reg ;
  assign \piso.data_r [2139] = \piso.data_r_2139_sv2v_reg ;
  assign \piso.data_r [2138] = \piso.data_r_2138_sv2v_reg ;
  assign \piso.data_r [2137] = \piso.data_r_2137_sv2v_reg ;
  assign \piso.data_r [2136] = \piso.data_r_2136_sv2v_reg ;
  assign \piso.data_r [2135] = \piso.data_r_2135_sv2v_reg ;
  assign \piso.data_r [2134] = \piso.data_r_2134_sv2v_reg ;
  assign \piso.data_r [2133] = \piso.data_r_2133_sv2v_reg ;
  assign \piso.data_r [2132] = \piso.data_r_2132_sv2v_reg ;
  assign \piso.data_r [2131] = \piso.data_r_2131_sv2v_reg ;
  assign \piso.data_r [2130] = \piso.data_r_2130_sv2v_reg ;
  assign \piso.data_r [2129] = \piso.data_r_2129_sv2v_reg ;
  assign \piso.data_r [2128] = \piso.data_r_2128_sv2v_reg ;
  assign \piso.data_r [2127] = \piso.data_r_2127_sv2v_reg ;
  assign \piso.data_r [2126] = \piso.data_r_2126_sv2v_reg ;
  assign \piso.data_r [2125] = \piso.data_r_2125_sv2v_reg ;
  assign \piso.data_r [2124] = \piso.data_r_2124_sv2v_reg ;
  assign \piso.data_r [2123] = \piso.data_r_2123_sv2v_reg ;
  assign \piso.data_r [2122] = \piso.data_r_2122_sv2v_reg ;
  assign \piso.data_r [2121] = \piso.data_r_2121_sv2v_reg ;
  assign \piso.data_r [2120] = \piso.data_r_2120_sv2v_reg ;
  assign \piso.data_r [2119] = \piso.data_r_2119_sv2v_reg ;
  assign \piso.data_r [2118] = \piso.data_r_2118_sv2v_reg ;
  assign \piso.data_r [2117] = \piso.data_r_2117_sv2v_reg ;
  assign \piso.data_r [2116] = \piso.data_r_2116_sv2v_reg ;
  assign \piso.data_r [2115] = \piso.data_r_2115_sv2v_reg ;
  assign \piso.data_r [2114] = \piso.data_r_2114_sv2v_reg ;
  assign \piso.data_r [2113] = \piso.data_r_2113_sv2v_reg ;
  assign \piso.data_r [2112] = \piso.data_r_2112_sv2v_reg ;
  assign \piso.data_r [2111] = \piso.data_r_2111_sv2v_reg ;
  assign \piso.data_r [2110] = \piso.data_r_2110_sv2v_reg ;
  assign \piso.data_r [2109] = \piso.data_r_2109_sv2v_reg ;
  assign \piso.data_r [2108] = \piso.data_r_2108_sv2v_reg ;
  assign \piso.data_r [2107] = \piso.data_r_2107_sv2v_reg ;
  assign \piso.data_r [2106] = \piso.data_r_2106_sv2v_reg ;
  assign \piso.data_r [2105] = \piso.data_r_2105_sv2v_reg ;
  assign \piso.data_r [2104] = \piso.data_r_2104_sv2v_reg ;
  assign \piso.data_r [2103] = \piso.data_r_2103_sv2v_reg ;
  assign \piso.data_r [2102] = \piso.data_r_2102_sv2v_reg ;
  assign \piso.data_r [2101] = \piso.data_r_2101_sv2v_reg ;
  assign \piso.data_r [2100] = \piso.data_r_2100_sv2v_reg ;
  assign \piso.data_r [2099] = \piso.data_r_2099_sv2v_reg ;
  assign \piso.data_r [2098] = \piso.data_r_2098_sv2v_reg ;
  assign \piso.data_r [2097] = \piso.data_r_2097_sv2v_reg ;
  assign \piso.data_r [2096] = \piso.data_r_2096_sv2v_reg ;
  assign \piso.data_r [2095] = \piso.data_r_2095_sv2v_reg ;
  assign \piso.data_r [2094] = \piso.data_r_2094_sv2v_reg ;
  assign \piso.data_r [2093] = \piso.data_r_2093_sv2v_reg ;
  assign \piso.data_r [2092] = \piso.data_r_2092_sv2v_reg ;
  assign \piso.data_r [2091] = \piso.data_r_2091_sv2v_reg ;
  assign \piso.data_r [2090] = \piso.data_r_2090_sv2v_reg ;
  assign \piso.data_r [2089] = \piso.data_r_2089_sv2v_reg ;
  assign \piso.data_r [2088] = \piso.data_r_2088_sv2v_reg ;
  assign \piso.data_r [2087] = \piso.data_r_2087_sv2v_reg ;
  assign \piso.data_r [2086] = \piso.data_r_2086_sv2v_reg ;
  assign \piso.data_r [2085] = \piso.data_r_2085_sv2v_reg ;
  assign \piso.data_r [2084] = \piso.data_r_2084_sv2v_reg ;
  assign \piso.data_r [2083] = \piso.data_r_2083_sv2v_reg ;
  assign \piso.data_r [2082] = \piso.data_r_2082_sv2v_reg ;
  assign \piso.data_r [2081] = \piso.data_r_2081_sv2v_reg ;
  assign \piso.data_r [2080] = \piso.data_r_2080_sv2v_reg ;
  assign \piso.data_r [2079] = \piso.data_r_2079_sv2v_reg ;
  assign \piso.data_r [2078] = \piso.data_r_2078_sv2v_reg ;
  assign \piso.data_r [2077] = \piso.data_r_2077_sv2v_reg ;
  assign \piso.data_r [2076] = \piso.data_r_2076_sv2v_reg ;
  assign \piso.data_r [2075] = \piso.data_r_2075_sv2v_reg ;
  assign \piso.data_r [2074] = \piso.data_r_2074_sv2v_reg ;
  assign \piso.data_r [2073] = \piso.data_r_2073_sv2v_reg ;
  assign \piso.data_r [2072] = \piso.data_r_2072_sv2v_reg ;
  assign \piso.data_r [2071] = \piso.data_r_2071_sv2v_reg ;
  assign \piso.data_r [2070] = \piso.data_r_2070_sv2v_reg ;
  assign \piso.data_r [2069] = \piso.data_r_2069_sv2v_reg ;
  assign \piso.data_r [2068] = \piso.data_r_2068_sv2v_reg ;
  assign \piso.data_r [2067] = \piso.data_r_2067_sv2v_reg ;
  assign \piso.data_r [2066] = \piso.data_r_2066_sv2v_reg ;
  assign \piso.data_r [2065] = \piso.data_r_2065_sv2v_reg ;
  assign \piso.data_r [2064] = \piso.data_r_2064_sv2v_reg ;
  assign \piso.data_r [2063] = \piso.data_r_2063_sv2v_reg ;
  assign \piso.data_r [2062] = \piso.data_r_2062_sv2v_reg ;
  assign \piso.data_r [2061] = \piso.data_r_2061_sv2v_reg ;
  assign \piso.data_r [2060] = \piso.data_r_2060_sv2v_reg ;
  assign \piso.data_r [2059] = \piso.data_r_2059_sv2v_reg ;
  assign \piso.data_r [2058] = \piso.data_r_2058_sv2v_reg ;
  assign \piso.data_r [2057] = \piso.data_r_2057_sv2v_reg ;
  assign \piso.data_r [2056] = \piso.data_r_2056_sv2v_reg ;
  assign \piso.data_r [2055] = \piso.data_r_2055_sv2v_reg ;
  assign \piso.data_r [2054] = \piso.data_r_2054_sv2v_reg ;
  assign \piso.data_r [2053] = \piso.data_r_2053_sv2v_reg ;
  assign \piso.data_r [2052] = \piso.data_r_2052_sv2v_reg ;
  assign \piso.data_r [2051] = \piso.data_r_2051_sv2v_reg ;
  assign \piso.data_r [2050] = \piso.data_r_2050_sv2v_reg ;
  assign \piso.data_r [2049] = \piso.data_r_2049_sv2v_reg ;
  assign \piso.data_r [2048] = \piso.data_r_2048_sv2v_reg ;
  assign \piso.data_r [2047] = \piso.data_r_2047_sv2v_reg ;
  assign \piso.data_r [2046] = \piso.data_r_2046_sv2v_reg ;
  assign \piso.data_r [2045] = \piso.data_r_2045_sv2v_reg ;
  assign \piso.data_r [2044] = \piso.data_r_2044_sv2v_reg ;
  assign \piso.data_r [2043] = \piso.data_r_2043_sv2v_reg ;
  assign \piso.data_r [2042] = \piso.data_r_2042_sv2v_reg ;
  assign \piso.data_r [2041] = \piso.data_r_2041_sv2v_reg ;
  assign \piso.data_r [2040] = \piso.data_r_2040_sv2v_reg ;
  assign \piso.data_r [2039] = \piso.data_r_2039_sv2v_reg ;
  assign \piso.data_r [2038] = \piso.data_r_2038_sv2v_reg ;
  assign \piso.data_r [2037] = \piso.data_r_2037_sv2v_reg ;
  assign \piso.data_r [2036] = \piso.data_r_2036_sv2v_reg ;
  assign \piso.data_r [2035] = \piso.data_r_2035_sv2v_reg ;
  assign \piso.data_r [2034] = \piso.data_r_2034_sv2v_reg ;
  assign \piso.data_r [2033] = \piso.data_r_2033_sv2v_reg ;
  assign \piso.data_r [2032] = \piso.data_r_2032_sv2v_reg ;
  assign \piso.data_r [2031] = \piso.data_r_2031_sv2v_reg ;
  assign \piso.data_r [2030] = \piso.data_r_2030_sv2v_reg ;
  assign \piso.data_r [2029] = \piso.data_r_2029_sv2v_reg ;
  assign \piso.data_r [2028] = \piso.data_r_2028_sv2v_reg ;
  assign \piso.data_r [2027] = \piso.data_r_2027_sv2v_reg ;
  assign \piso.data_r [2026] = \piso.data_r_2026_sv2v_reg ;
  assign \piso.data_r [2025] = \piso.data_r_2025_sv2v_reg ;
  assign \piso.data_r [2024] = \piso.data_r_2024_sv2v_reg ;
  assign \piso.data_r [2023] = \piso.data_r_2023_sv2v_reg ;
  assign \piso.data_r [2022] = \piso.data_r_2022_sv2v_reg ;
  assign \piso.data_r [2021] = \piso.data_r_2021_sv2v_reg ;
  assign \piso.data_r [2020] = \piso.data_r_2020_sv2v_reg ;
  assign \piso.data_r [2019] = \piso.data_r_2019_sv2v_reg ;
  assign \piso.data_r [2018] = \piso.data_r_2018_sv2v_reg ;
  assign \piso.data_r [2017] = \piso.data_r_2017_sv2v_reg ;
  assign \piso.data_r [2016] = \piso.data_r_2016_sv2v_reg ;
  assign \piso.data_r [2015] = \piso.data_r_2015_sv2v_reg ;
  assign \piso.data_r [2014] = \piso.data_r_2014_sv2v_reg ;
  assign \piso.data_r [2013] = \piso.data_r_2013_sv2v_reg ;
  assign \piso.data_r [2012] = \piso.data_r_2012_sv2v_reg ;
  assign \piso.data_r [2011] = \piso.data_r_2011_sv2v_reg ;
  assign \piso.data_r [2010] = \piso.data_r_2010_sv2v_reg ;
  assign \piso.data_r [2009] = \piso.data_r_2009_sv2v_reg ;
  assign \piso.data_r [2008] = \piso.data_r_2008_sv2v_reg ;
  assign \piso.data_r [2007] = \piso.data_r_2007_sv2v_reg ;
  assign \piso.data_r [2006] = \piso.data_r_2006_sv2v_reg ;
  assign \piso.data_r [2005] = \piso.data_r_2005_sv2v_reg ;
  assign \piso.data_r [2004] = \piso.data_r_2004_sv2v_reg ;
  assign \piso.data_r [2003] = \piso.data_r_2003_sv2v_reg ;
  assign \piso.data_r [2002] = \piso.data_r_2002_sv2v_reg ;
  assign \piso.data_r [2001] = \piso.data_r_2001_sv2v_reg ;
  assign \piso.data_r [2000] = \piso.data_r_2000_sv2v_reg ;
  assign \piso.data_r [1999] = \piso.data_r_1999_sv2v_reg ;
  assign \piso.data_r [1998] = \piso.data_r_1998_sv2v_reg ;
  assign \piso.data_r [1997] = \piso.data_r_1997_sv2v_reg ;
  assign \piso.data_r [1996] = \piso.data_r_1996_sv2v_reg ;
  assign \piso.data_r [1995] = \piso.data_r_1995_sv2v_reg ;
  assign \piso.data_r [1994] = \piso.data_r_1994_sv2v_reg ;
  assign \piso.data_r [1993] = \piso.data_r_1993_sv2v_reg ;
  assign \piso.data_r [1992] = \piso.data_r_1992_sv2v_reg ;
  assign \piso.data_r [1991] = \piso.data_r_1991_sv2v_reg ;
  assign \piso.data_r [1990] = \piso.data_r_1990_sv2v_reg ;
  assign \piso.data_r [1989] = \piso.data_r_1989_sv2v_reg ;
  assign \piso.data_r [1988] = \piso.data_r_1988_sv2v_reg ;
  assign \piso.data_r [1987] = \piso.data_r_1987_sv2v_reg ;
  assign \piso.data_r [1986] = \piso.data_r_1986_sv2v_reg ;
  assign \piso.data_r [1985] = \piso.data_r_1985_sv2v_reg ;
  assign \piso.data_r [1984] = \piso.data_r_1984_sv2v_reg ;
  assign \piso.data_r [1983] = \piso.data_r_1983_sv2v_reg ;
  assign \piso.data_r [1982] = \piso.data_r_1982_sv2v_reg ;
  assign \piso.data_r [1981] = \piso.data_r_1981_sv2v_reg ;
  assign \piso.data_r [1980] = \piso.data_r_1980_sv2v_reg ;
  assign \piso.data_r [1979] = \piso.data_r_1979_sv2v_reg ;
  assign \piso.data_r [1978] = \piso.data_r_1978_sv2v_reg ;
  assign \piso.data_r [1977] = \piso.data_r_1977_sv2v_reg ;
  assign \piso.data_r [1976] = \piso.data_r_1976_sv2v_reg ;
  assign \piso.data_r [1975] = \piso.data_r_1975_sv2v_reg ;
  assign \piso.data_r [1974] = \piso.data_r_1974_sv2v_reg ;
  assign \piso.data_r [1973] = \piso.data_r_1973_sv2v_reg ;
  assign \piso.data_r [1972] = \piso.data_r_1972_sv2v_reg ;
  assign \piso.data_r [1971] = \piso.data_r_1971_sv2v_reg ;
  assign \piso.data_r [1970] = \piso.data_r_1970_sv2v_reg ;
  assign \piso.data_r [1969] = \piso.data_r_1969_sv2v_reg ;
  assign \piso.data_r [1968] = \piso.data_r_1968_sv2v_reg ;
  assign \piso.data_r [1967] = \piso.data_r_1967_sv2v_reg ;
  assign \piso.data_r [1966] = \piso.data_r_1966_sv2v_reg ;
  assign \piso.data_r [1965] = \piso.data_r_1965_sv2v_reg ;
  assign \piso.data_r [1964] = \piso.data_r_1964_sv2v_reg ;
  assign \piso.data_r [1963] = \piso.data_r_1963_sv2v_reg ;
  assign \piso.data_r [1962] = \piso.data_r_1962_sv2v_reg ;
  assign \piso.data_r [1961] = \piso.data_r_1961_sv2v_reg ;
  assign \piso.data_r [1960] = \piso.data_r_1960_sv2v_reg ;
  assign \piso.data_r [1959] = \piso.data_r_1959_sv2v_reg ;
  assign \piso.data_r [1958] = \piso.data_r_1958_sv2v_reg ;
  assign \piso.data_r [1957] = \piso.data_r_1957_sv2v_reg ;
  assign \piso.data_r [1956] = \piso.data_r_1956_sv2v_reg ;
  assign \piso.data_r [1955] = \piso.data_r_1955_sv2v_reg ;
  assign \piso.data_r [1954] = \piso.data_r_1954_sv2v_reg ;
  assign \piso.data_r [1953] = \piso.data_r_1953_sv2v_reg ;
  assign \piso.data_r [1952] = \piso.data_r_1952_sv2v_reg ;
  assign \piso.data_r [1951] = \piso.data_r_1951_sv2v_reg ;
  assign \piso.data_r [1950] = \piso.data_r_1950_sv2v_reg ;
  assign \piso.data_r [1949] = \piso.data_r_1949_sv2v_reg ;
  assign \piso.data_r [1948] = \piso.data_r_1948_sv2v_reg ;
  assign \piso.data_r [1947] = \piso.data_r_1947_sv2v_reg ;
  assign \piso.data_r [1946] = \piso.data_r_1946_sv2v_reg ;
  assign \piso.data_r [1945] = \piso.data_r_1945_sv2v_reg ;
  assign \piso.data_r [1944] = \piso.data_r_1944_sv2v_reg ;
  assign \piso.data_r [1943] = \piso.data_r_1943_sv2v_reg ;
  assign \piso.data_r [1942] = \piso.data_r_1942_sv2v_reg ;
  assign \piso.data_r [1941] = \piso.data_r_1941_sv2v_reg ;
  assign \piso.data_r [1940] = \piso.data_r_1940_sv2v_reg ;
  assign \piso.data_r [1939] = \piso.data_r_1939_sv2v_reg ;
  assign \piso.data_r [1938] = \piso.data_r_1938_sv2v_reg ;
  assign \piso.data_r [1937] = \piso.data_r_1937_sv2v_reg ;
  assign \piso.data_r [1936] = \piso.data_r_1936_sv2v_reg ;
  assign \piso.data_r [1935] = \piso.data_r_1935_sv2v_reg ;
  assign \piso.data_r [1934] = \piso.data_r_1934_sv2v_reg ;
  assign \piso.data_r [1933] = \piso.data_r_1933_sv2v_reg ;
  assign \piso.data_r [1932] = \piso.data_r_1932_sv2v_reg ;
  assign \piso.data_r [1931] = \piso.data_r_1931_sv2v_reg ;
  assign \piso.data_r [1930] = \piso.data_r_1930_sv2v_reg ;
  assign \piso.data_r [1929] = \piso.data_r_1929_sv2v_reg ;
  assign \piso.data_r [1928] = \piso.data_r_1928_sv2v_reg ;
  assign \piso.data_r [1927] = \piso.data_r_1927_sv2v_reg ;
  assign \piso.data_r [1926] = \piso.data_r_1926_sv2v_reg ;
  assign \piso.data_r [1925] = \piso.data_r_1925_sv2v_reg ;
  assign \piso.data_r [1924] = \piso.data_r_1924_sv2v_reg ;
  assign \piso.data_r [1923] = \piso.data_r_1923_sv2v_reg ;
  assign \piso.data_r [1922] = \piso.data_r_1922_sv2v_reg ;
  assign \piso.data_r [1921] = \piso.data_r_1921_sv2v_reg ;
  assign \piso.data_r [1920] = \piso.data_r_1920_sv2v_reg ;
  assign \piso.data_r [1919] = \piso.data_r_1919_sv2v_reg ;
  assign \piso.data_r [1918] = \piso.data_r_1918_sv2v_reg ;
  assign \piso.data_r [1917] = \piso.data_r_1917_sv2v_reg ;
  assign \piso.data_r [1916] = \piso.data_r_1916_sv2v_reg ;
  assign \piso.data_r [1915] = \piso.data_r_1915_sv2v_reg ;
  assign \piso.data_r [1914] = \piso.data_r_1914_sv2v_reg ;
  assign \piso.data_r [1913] = \piso.data_r_1913_sv2v_reg ;
  assign \piso.data_r [1912] = \piso.data_r_1912_sv2v_reg ;
  assign \piso.data_r [1911] = \piso.data_r_1911_sv2v_reg ;
  assign \piso.data_r [1910] = \piso.data_r_1910_sv2v_reg ;
  assign \piso.data_r [1909] = \piso.data_r_1909_sv2v_reg ;
  assign \piso.data_r [1908] = \piso.data_r_1908_sv2v_reg ;
  assign \piso.data_r [1907] = \piso.data_r_1907_sv2v_reg ;
  assign \piso.data_r [1906] = \piso.data_r_1906_sv2v_reg ;
  assign \piso.data_r [1905] = \piso.data_r_1905_sv2v_reg ;
  assign \piso.data_r [1904] = \piso.data_r_1904_sv2v_reg ;
  assign \piso.data_r [1903] = \piso.data_r_1903_sv2v_reg ;
  assign \piso.data_r [1902] = \piso.data_r_1902_sv2v_reg ;
  assign \piso.data_r [1901] = \piso.data_r_1901_sv2v_reg ;
  assign \piso.data_r [1900] = \piso.data_r_1900_sv2v_reg ;
  assign \piso.data_r [1899] = \piso.data_r_1899_sv2v_reg ;
  assign \piso.data_r [1898] = \piso.data_r_1898_sv2v_reg ;
  assign \piso.data_r [1897] = \piso.data_r_1897_sv2v_reg ;
  assign \piso.data_r [1896] = \piso.data_r_1896_sv2v_reg ;
  assign \piso.data_r [1895] = \piso.data_r_1895_sv2v_reg ;
  assign \piso.data_r [1894] = \piso.data_r_1894_sv2v_reg ;
  assign \piso.data_r [1893] = \piso.data_r_1893_sv2v_reg ;
  assign \piso.data_r [1892] = \piso.data_r_1892_sv2v_reg ;
  assign \piso.data_r [1891] = \piso.data_r_1891_sv2v_reg ;
  assign \piso.data_r [1890] = \piso.data_r_1890_sv2v_reg ;
  assign \piso.data_r [1889] = \piso.data_r_1889_sv2v_reg ;
  assign \piso.data_r [1888] = \piso.data_r_1888_sv2v_reg ;
  assign \piso.data_r [1887] = \piso.data_r_1887_sv2v_reg ;
  assign \piso.data_r [1886] = \piso.data_r_1886_sv2v_reg ;
  assign \piso.data_r [1885] = \piso.data_r_1885_sv2v_reg ;
  assign \piso.data_r [1884] = \piso.data_r_1884_sv2v_reg ;
  assign \piso.data_r [1883] = \piso.data_r_1883_sv2v_reg ;
  assign \piso.data_r [1882] = \piso.data_r_1882_sv2v_reg ;
  assign \piso.data_r [1881] = \piso.data_r_1881_sv2v_reg ;
  assign \piso.data_r [1880] = \piso.data_r_1880_sv2v_reg ;
  assign \piso.data_r [1879] = \piso.data_r_1879_sv2v_reg ;
  assign \piso.data_r [1878] = \piso.data_r_1878_sv2v_reg ;
  assign \piso.data_r [1877] = \piso.data_r_1877_sv2v_reg ;
  assign \piso.data_r [1876] = \piso.data_r_1876_sv2v_reg ;
  assign \piso.data_r [1875] = \piso.data_r_1875_sv2v_reg ;
  assign \piso.data_r [1874] = \piso.data_r_1874_sv2v_reg ;
  assign \piso.data_r [1873] = \piso.data_r_1873_sv2v_reg ;
  assign \piso.data_r [1872] = \piso.data_r_1872_sv2v_reg ;
  assign \piso.data_r [1871] = \piso.data_r_1871_sv2v_reg ;
  assign \piso.data_r [1870] = \piso.data_r_1870_sv2v_reg ;
  assign \piso.data_r [1869] = \piso.data_r_1869_sv2v_reg ;
  assign \piso.data_r [1868] = \piso.data_r_1868_sv2v_reg ;
  assign \piso.data_r [1867] = \piso.data_r_1867_sv2v_reg ;
  assign \piso.data_r [1866] = \piso.data_r_1866_sv2v_reg ;
  assign \piso.data_r [1865] = \piso.data_r_1865_sv2v_reg ;
  assign \piso.data_r [1864] = \piso.data_r_1864_sv2v_reg ;
  assign \piso.data_r [1863] = \piso.data_r_1863_sv2v_reg ;
  assign \piso.data_r [1862] = \piso.data_r_1862_sv2v_reg ;
  assign \piso.data_r [1861] = \piso.data_r_1861_sv2v_reg ;
  assign \piso.data_r [1860] = \piso.data_r_1860_sv2v_reg ;
  assign \piso.data_r [1859] = \piso.data_r_1859_sv2v_reg ;
  assign \piso.data_r [1858] = \piso.data_r_1858_sv2v_reg ;
  assign \piso.data_r [1857] = \piso.data_r_1857_sv2v_reg ;
  assign \piso.data_r [1856] = \piso.data_r_1856_sv2v_reg ;
  assign \piso.data_r [1855] = \piso.data_r_1855_sv2v_reg ;
  assign \piso.data_r [1854] = \piso.data_r_1854_sv2v_reg ;
  assign \piso.data_r [1853] = \piso.data_r_1853_sv2v_reg ;
  assign \piso.data_r [1852] = \piso.data_r_1852_sv2v_reg ;
  assign \piso.data_r [1851] = \piso.data_r_1851_sv2v_reg ;
  assign \piso.data_r [1850] = \piso.data_r_1850_sv2v_reg ;
  assign \piso.data_r [1849] = \piso.data_r_1849_sv2v_reg ;
  assign \piso.data_r [1848] = \piso.data_r_1848_sv2v_reg ;
  assign \piso.data_r [1847] = \piso.data_r_1847_sv2v_reg ;
  assign \piso.data_r [1846] = \piso.data_r_1846_sv2v_reg ;
  assign \piso.data_r [1845] = \piso.data_r_1845_sv2v_reg ;
  assign \piso.data_r [1844] = \piso.data_r_1844_sv2v_reg ;
  assign \piso.data_r [1843] = \piso.data_r_1843_sv2v_reg ;
  assign \piso.data_r [1842] = \piso.data_r_1842_sv2v_reg ;
  assign \piso.data_r [1841] = \piso.data_r_1841_sv2v_reg ;
  assign \piso.data_r [1840] = \piso.data_r_1840_sv2v_reg ;
  assign \piso.data_r [1839] = \piso.data_r_1839_sv2v_reg ;
  assign \piso.data_r [1838] = \piso.data_r_1838_sv2v_reg ;
  assign \piso.data_r [1837] = \piso.data_r_1837_sv2v_reg ;
  assign \piso.data_r [1836] = \piso.data_r_1836_sv2v_reg ;
  assign \piso.data_r [1835] = \piso.data_r_1835_sv2v_reg ;
  assign \piso.data_r [1834] = \piso.data_r_1834_sv2v_reg ;
  assign \piso.data_r [1833] = \piso.data_r_1833_sv2v_reg ;
  assign \piso.data_r [1832] = \piso.data_r_1832_sv2v_reg ;
  assign \piso.data_r [1831] = \piso.data_r_1831_sv2v_reg ;
  assign \piso.data_r [1830] = \piso.data_r_1830_sv2v_reg ;
  assign \piso.data_r [1829] = \piso.data_r_1829_sv2v_reg ;
  assign \piso.data_r [1828] = \piso.data_r_1828_sv2v_reg ;
  assign \piso.data_r [1827] = \piso.data_r_1827_sv2v_reg ;
  assign \piso.data_r [1826] = \piso.data_r_1826_sv2v_reg ;
  assign \piso.data_r [1825] = \piso.data_r_1825_sv2v_reg ;
  assign \piso.data_r [1824] = \piso.data_r_1824_sv2v_reg ;
  assign \piso.data_r [1823] = \piso.data_r_1823_sv2v_reg ;
  assign \piso.data_r [1822] = \piso.data_r_1822_sv2v_reg ;
  assign \piso.data_r [1821] = \piso.data_r_1821_sv2v_reg ;
  assign \piso.data_r [1820] = \piso.data_r_1820_sv2v_reg ;
  assign \piso.data_r [1819] = \piso.data_r_1819_sv2v_reg ;
  assign \piso.data_r [1818] = \piso.data_r_1818_sv2v_reg ;
  assign \piso.data_r [1817] = \piso.data_r_1817_sv2v_reg ;
  assign \piso.data_r [1816] = \piso.data_r_1816_sv2v_reg ;
  assign \piso.data_r [1815] = \piso.data_r_1815_sv2v_reg ;
  assign \piso.data_r [1814] = \piso.data_r_1814_sv2v_reg ;
  assign \piso.data_r [1813] = \piso.data_r_1813_sv2v_reg ;
  assign \piso.data_r [1812] = \piso.data_r_1812_sv2v_reg ;
  assign \piso.data_r [1811] = \piso.data_r_1811_sv2v_reg ;
  assign \piso.data_r [1810] = \piso.data_r_1810_sv2v_reg ;
  assign \piso.data_r [1809] = \piso.data_r_1809_sv2v_reg ;
  assign \piso.data_r [1808] = \piso.data_r_1808_sv2v_reg ;
  assign \piso.data_r [1807] = \piso.data_r_1807_sv2v_reg ;
  assign \piso.data_r [1806] = \piso.data_r_1806_sv2v_reg ;
  assign \piso.data_r [1805] = \piso.data_r_1805_sv2v_reg ;
  assign \piso.data_r [1804] = \piso.data_r_1804_sv2v_reg ;
  assign \piso.data_r [1803] = \piso.data_r_1803_sv2v_reg ;
  assign \piso.data_r [1802] = \piso.data_r_1802_sv2v_reg ;
  assign \piso.data_r [1801] = \piso.data_r_1801_sv2v_reg ;
  assign \piso.data_r [1800] = \piso.data_r_1800_sv2v_reg ;
  assign \piso.data_r [1799] = \piso.data_r_1799_sv2v_reg ;
  assign \piso.data_r [1798] = \piso.data_r_1798_sv2v_reg ;
  assign \piso.data_r [1797] = \piso.data_r_1797_sv2v_reg ;
  assign \piso.data_r [1796] = \piso.data_r_1796_sv2v_reg ;
  assign \piso.data_r [1795] = \piso.data_r_1795_sv2v_reg ;
  assign \piso.data_r [1794] = \piso.data_r_1794_sv2v_reg ;
  assign \piso.data_r [1793] = \piso.data_r_1793_sv2v_reg ;
  assign \piso.data_r [1792] = \piso.data_r_1792_sv2v_reg ;
  assign \piso.data_r [1791] = \piso.data_r_1791_sv2v_reg ;
  assign \piso.data_r [1790] = \piso.data_r_1790_sv2v_reg ;
  assign \piso.data_r [1789] = \piso.data_r_1789_sv2v_reg ;
  assign \piso.data_r [1788] = \piso.data_r_1788_sv2v_reg ;
  assign \piso.data_r [1787] = \piso.data_r_1787_sv2v_reg ;
  assign \piso.data_r [1786] = \piso.data_r_1786_sv2v_reg ;
  assign \piso.data_r [1785] = \piso.data_r_1785_sv2v_reg ;
  assign \piso.data_r [1784] = \piso.data_r_1784_sv2v_reg ;
  assign \piso.data_r [1783] = \piso.data_r_1783_sv2v_reg ;
  assign \piso.data_r [1782] = \piso.data_r_1782_sv2v_reg ;
  assign \piso.data_r [1781] = \piso.data_r_1781_sv2v_reg ;
  assign \piso.data_r [1780] = \piso.data_r_1780_sv2v_reg ;
  assign \piso.data_r [1779] = \piso.data_r_1779_sv2v_reg ;
  assign \piso.data_r [1778] = \piso.data_r_1778_sv2v_reg ;
  assign \piso.data_r [1777] = \piso.data_r_1777_sv2v_reg ;
  assign \piso.data_r [1776] = \piso.data_r_1776_sv2v_reg ;
  assign \piso.data_r [1775] = \piso.data_r_1775_sv2v_reg ;
  assign \piso.data_r [1774] = \piso.data_r_1774_sv2v_reg ;
  assign \piso.data_r [1773] = \piso.data_r_1773_sv2v_reg ;
  assign \piso.data_r [1772] = \piso.data_r_1772_sv2v_reg ;
  assign \piso.data_r [1771] = \piso.data_r_1771_sv2v_reg ;
  assign \piso.data_r [1770] = \piso.data_r_1770_sv2v_reg ;
  assign \piso.data_r [1769] = \piso.data_r_1769_sv2v_reg ;
  assign \piso.data_r [1768] = \piso.data_r_1768_sv2v_reg ;
  assign \piso.data_r [1767] = \piso.data_r_1767_sv2v_reg ;
  assign \piso.data_r [1766] = \piso.data_r_1766_sv2v_reg ;
  assign \piso.data_r [1765] = \piso.data_r_1765_sv2v_reg ;
  assign \piso.data_r [1764] = \piso.data_r_1764_sv2v_reg ;
  assign \piso.data_r [1763] = \piso.data_r_1763_sv2v_reg ;
  assign \piso.data_r [1762] = \piso.data_r_1762_sv2v_reg ;
  assign \piso.data_r [1761] = \piso.data_r_1761_sv2v_reg ;
  assign \piso.data_r [1760] = \piso.data_r_1760_sv2v_reg ;
  assign \piso.data_r [1759] = \piso.data_r_1759_sv2v_reg ;
  assign \piso.data_r [1758] = \piso.data_r_1758_sv2v_reg ;
  assign \piso.data_r [1757] = \piso.data_r_1757_sv2v_reg ;
  assign \piso.data_r [1756] = \piso.data_r_1756_sv2v_reg ;
  assign \piso.data_r [1755] = \piso.data_r_1755_sv2v_reg ;
  assign \piso.data_r [1754] = \piso.data_r_1754_sv2v_reg ;
  assign \piso.data_r [1753] = \piso.data_r_1753_sv2v_reg ;
  assign \piso.data_r [1752] = \piso.data_r_1752_sv2v_reg ;
  assign \piso.data_r [1751] = \piso.data_r_1751_sv2v_reg ;
  assign \piso.data_r [1750] = \piso.data_r_1750_sv2v_reg ;
  assign \piso.data_r [1749] = \piso.data_r_1749_sv2v_reg ;
  assign \piso.data_r [1748] = \piso.data_r_1748_sv2v_reg ;
  assign \piso.data_r [1747] = \piso.data_r_1747_sv2v_reg ;
  assign \piso.data_r [1746] = \piso.data_r_1746_sv2v_reg ;
  assign \piso.data_r [1745] = \piso.data_r_1745_sv2v_reg ;
  assign \piso.data_r [1744] = \piso.data_r_1744_sv2v_reg ;
  assign \piso.data_r [1743] = \piso.data_r_1743_sv2v_reg ;
  assign \piso.data_r [1742] = \piso.data_r_1742_sv2v_reg ;
  assign \piso.data_r [1741] = \piso.data_r_1741_sv2v_reg ;
  assign \piso.data_r [1740] = \piso.data_r_1740_sv2v_reg ;
  assign \piso.data_r [1739] = \piso.data_r_1739_sv2v_reg ;
  assign \piso.data_r [1738] = \piso.data_r_1738_sv2v_reg ;
  assign \piso.data_r [1737] = \piso.data_r_1737_sv2v_reg ;
  assign \piso.data_r [1736] = \piso.data_r_1736_sv2v_reg ;
  assign \piso.data_r [1735] = \piso.data_r_1735_sv2v_reg ;
  assign \piso.data_r [1734] = \piso.data_r_1734_sv2v_reg ;
  assign \piso.data_r [1733] = \piso.data_r_1733_sv2v_reg ;
  assign \piso.data_r [1732] = \piso.data_r_1732_sv2v_reg ;
  assign \piso.data_r [1731] = \piso.data_r_1731_sv2v_reg ;
  assign \piso.data_r [1730] = \piso.data_r_1730_sv2v_reg ;
  assign \piso.data_r [1729] = \piso.data_r_1729_sv2v_reg ;
  assign \piso.data_r [1728] = \piso.data_r_1728_sv2v_reg ;
  assign \piso.data_r [1727] = \piso.data_r_1727_sv2v_reg ;
  assign \piso.data_r [1726] = \piso.data_r_1726_sv2v_reg ;
  assign \piso.data_r [1725] = \piso.data_r_1725_sv2v_reg ;
  assign \piso.data_r [1724] = \piso.data_r_1724_sv2v_reg ;
  assign \piso.data_r [1723] = \piso.data_r_1723_sv2v_reg ;
  assign \piso.data_r [1722] = \piso.data_r_1722_sv2v_reg ;
  assign \piso.data_r [1721] = \piso.data_r_1721_sv2v_reg ;
  assign \piso.data_r [1720] = \piso.data_r_1720_sv2v_reg ;
  assign \piso.data_r [1719] = \piso.data_r_1719_sv2v_reg ;
  assign \piso.data_r [1718] = \piso.data_r_1718_sv2v_reg ;
  assign \piso.data_r [1717] = \piso.data_r_1717_sv2v_reg ;
  assign \piso.data_r [1716] = \piso.data_r_1716_sv2v_reg ;
  assign \piso.data_r [1715] = \piso.data_r_1715_sv2v_reg ;
  assign \piso.data_r [1714] = \piso.data_r_1714_sv2v_reg ;
  assign \piso.data_r [1713] = \piso.data_r_1713_sv2v_reg ;
  assign \piso.data_r [1712] = \piso.data_r_1712_sv2v_reg ;
  assign \piso.data_r [1711] = \piso.data_r_1711_sv2v_reg ;
  assign \piso.data_r [1710] = \piso.data_r_1710_sv2v_reg ;
  assign \piso.data_r [1709] = \piso.data_r_1709_sv2v_reg ;
  assign \piso.data_r [1708] = \piso.data_r_1708_sv2v_reg ;
  assign \piso.data_r [1707] = \piso.data_r_1707_sv2v_reg ;
  assign \piso.data_r [1706] = \piso.data_r_1706_sv2v_reg ;
  assign \piso.data_r [1705] = \piso.data_r_1705_sv2v_reg ;
  assign \piso.data_r [1704] = \piso.data_r_1704_sv2v_reg ;
  assign \piso.data_r [1703] = \piso.data_r_1703_sv2v_reg ;
  assign \piso.data_r [1702] = \piso.data_r_1702_sv2v_reg ;
  assign \piso.data_r [1701] = \piso.data_r_1701_sv2v_reg ;
  assign \piso.data_r [1700] = \piso.data_r_1700_sv2v_reg ;
  assign \piso.data_r [1699] = \piso.data_r_1699_sv2v_reg ;
  assign \piso.data_r [1698] = \piso.data_r_1698_sv2v_reg ;
  assign \piso.data_r [1697] = \piso.data_r_1697_sv2v_reg ;
  assign \piso.data_r [1696] = \piso.data_r_1696_sv2v_reg ;
  assign \piso.data_r [1695] = \piso.data_r_1695_sv2v_reg ;
  assign \piso.data_r [1694] = \piso.data_r_1694_sv2v_reg ;
  assign \piso.data_r [1693] = \piso.data_r_1693_sv2v_reg ;
  assign \piso.data_r [1692] = \piso.data_r_1692_sv2v_reg ;
  assign \piso.data_r [1691] = \piso.data_r_1691_sv2v_reg ;
  assign \piso.data_r [1690] = \piso.data_r_1690_sv2v_reg ;
  assign \piso.data_r [1689] = \piso.data_r_1689_sv2v_reg ;
  assign \piso.data_r [1688] = \piso.data_r_1688_sv2v_reg ;
  assign \piso.data_r [1687] = \piso.data_r_1687_sv2v_reg ;
  assign \piso.data_r [1686] = \piso.data_r_1686_sv2v_reg ;
  assign \piso.data_r [1685] = \piso.data_r_1685_sv2v_reg ;
  assign \piso.data_r [1684] = \piso.data_r_1684_sv2v_reg ;
  assign \piso.data_r [1683] = \piso.data_r_1683_sv2v_reg ;
  assign \piso.data_r [1682] = \piso.data_r_1682_sv2v_reg ;
  assign \piso.data_r [1681] = \piso.data_r_1681_sv2v_reg ;
  assign \piso.data_r [1680] = \piso.data_r_1680_sv2v_reg ;
  assign \piso.data_r [1679] = \piso.data_r_1679_sv2v_reg ;
  assign \piso.data_r [1678] = \piso.data_r_1678_sv2v_reg ;
  assign \piso.data_r [1677] = \piso.data_r_1677_sv2v_reg ;
  assign \piso.data_r [1676] = \piso.data_r_1676_sv2v_reg ;
  assign \piso.data_r [1675] = \piso.data_r_1675_sv2v_reg ;
  assign \piso.data_r [1674] = \piso.data_r_1674_sv2v_reg ;
  assign \piso.data_r [1673] = \piso.data_r_1673_sv2v_reg ;
  assign \piso.data_r [1672] = \piso.data_r_1672_sv2v_reg ;
  assign \piso.data_r [1671] = \piso.data_r_1671_sv2v_reg ;
  assign \piso.data_r [1670] = \piso.data_r_1670_sv2v_reg ;
  assign \piso.data_r [1669] = \piso.data_r_1669_sv2v_reg ;
  assign \piso.data_r [1668] = \piso.data_r_1668_sv2v_reg ;
  assign \piso.data_r [1667] = \piso.data_r_1667_sv2v_reg ;
  assign \piso.data_r [1666] = \piso.data_r_1666_sv2v_reg ;
  assign \piso.data_r [1665] = \piso.data_r_1665_sv2v_reg ;
  assign \piso.data_r [1664] = \piso.data_r_1664_sv2v_reg ;
  assign \piso.data_r [1663] = \piso.data_r_1663_sv2v_reg ;
  assign \piso.data_r [1662] = \piso.data_r_1662_sv2v_reg ;
  assign \piso.data_r [1661] = \piso.data_r_1661_sv2v_reg ;
  assign \piso.data_r [1660] = \piso.data_r_1660_sv2v_reg ;
  assign \piso.data_r [1659] = \piso.data_r_1659_sv2v_reg ;
  assign \piso.data_r [1658] = \piso.data_r_1658_sv2v_reg ;
  assign \piso.data_r [1657] = \piso.data_r_1657_sv2v_reg ;
  assign \piso.data_r [1656] = \piso.data_r_1656_sv2v_reg ;
  assign \piso.data_r [1655] = \piso.data_r_1655_sv2v_reg ;
  assign \piso.data_r [1654] = \piso.data_r_1654_sv2v_reg ;
  assign \piso.data_r [1653] = \piso.data_r_1653_sv2v_reg ;
  assign \piso.data_r [1652] = \piso.data_r_1652_sv2v_reg ;
  assign \piso.data_r [1651] = \piso.data_r_1651_sv2v_reg ;
  assign \piso.data_r [1650] = \piso.data_r_1650_sv2v_reg ;
  assign \piso.data_r [1649] = \piso.data_r_1649_sv2v_reg ;
  assign \piso.data_r [1648] = \piso.data_r_1648_sv2v_reg ;
  assign \piso.data_r [1647] = \piso.data_r_1647_sv2v_reg ;
  assign \piso.data_r [1646] = \piso.data_r_1646_sv2v_reg ;
  assign \piso.data_r [1645] = \piso.data_r_1645_sv2v_reg ;
  assign \piso.data_r [1644] = \piso.data_r_1644_sv2v_reg ;
  assign \piso.data_r [1643] = \piso.data_r_1643_sv2v_reg ;
  assign \piso.data_r [1642] = \piso.data_r_1642_sv2v_reg ;
  assign \piso.data_r [1641] = \piso.data_r_1641_sv2v_reg ;
  assign \piso.data_r [1640] = \piso.data_r_1640_sv2v_reg ;
  assign \piso.data_r [1639] = \piso.data_r_1639_sv2v_reg ;
  assign \piso.data_r [1638] = \piso.data_r_1638_sv2v_reg ;
  assign \piso.data_r [1637] = \piso.data_r_1637_sv2v_reg ;
  assign \piso.data_r [1636] = \piso.data_r_1636_sv2v_reg ;
  assign \piso.data_r [1635] = \piso.data_r_1635_sv2v_reg ;
  assign \piso.data_r [1634] = \piso.data_r_1634_sv2v_reg ;
  assign \piso.data_r [1633] = \piso.data_r_1633_sv2v_reg ;
  assign \piso.data_r [1632] = \piso.data_r_1632_sv2v_reg ;
  assign \piso.data_r [1631] = \piso.data_r_1631_sv2v_reg ;
  assign \piso.data_r [1630] = \piso.data_r_1630_sv2v_reg ;
  assign \piso.data_r [1629] = \piso.data_r_1629_sv2v_reg ;
  assign \piso.data_r [1628] = \piso.data_r_1628_sv2v_reg ;
  assign \piso.data_r [1627] = \piso.data_r_1627_sv2v_reg ;
  assign \piso.data_r [1626] = \piso.data_r_1626_sv2v_reg ;
  assign \piso.data_r [1625] = \piso.data_r_1625_sv2v_reg ;
  assign \piso.data_r [1624] = \piso.data_r_1624_sv2v_reg ;
  assign \piso.data_r [1623] = \piso.data_r_1623_sv2v_reg ;
  assign \piso.data_r [1622] = \piso.data_r_1622_sv2v_reg ;
  assign \piso.data_r [1621] = \piso.data_r_1621_sv2v_reg ;
  assign \piso.data_r [1620] = \piso.data_r_1620_sv2v_reg ;
  assign \piso.data_r [1619] = \piso.data_r_1619_sv2v_reg ;
  assign \piso.data_r [1618] = \piso.data_r_1618_sv2v_reg ;
  assign \piso.data_r [1617] = \piso.data_r_1617_sv2v_reg ;
  assign \piso.data_r [1616] = \piso.data_r_1616_sv2v_reg ;
  assign \piso.data_r [1615] = \piso.data_r_1615_sv2v_reg ;
  assign \piso.data_r [1614] = \piso.data_r_1614_sv2v_reg ;
  assign \piso.data_r [1613] = \piso.data_r_1613_sv2v_reg ;
  assign \piso.data_r [1612] = \piso.data_r_1612_sv2v_reg ;
  assign \piso.data_r [1611] = \piso.data_r_1611_sv2v_reg ;
  assign \piso.data_r [1610] = \piso.data_r_1610_sv2v_reg ;
  assign \piso.data_r [1609] = \piso.data_r_1609_sv2v_reg ;
  assign \piso.data_r [1608] = \piso.data_r_1608_sv2v_reg ;
  assign \piso.data_r [1607] = \piso.data_r_1607_sv2v_reg ;
  assign \piso.data_r [1606] = \piso.data_r_1606_sv2v_reg ;
  assign \piso.data_r [1605] = \piso.data_r_1605_sv2v_reg ;
  assign \piso.data_r [1604] = \piso.data_r_1604_sv2v_reg ;
  assign \piso.data_r [1603] = \piso.data_r_1603_sv2v_reg ;
  assign \piso.data_r [1602] = \piso.data_r_1602_sv2v_reg ;
  assign \piso.data_r [1601] = \piso.data_r_1601_sv2v_reg ;
  assign \piso.data_r [1600] = \piso.data_r_1600_sv2v_reg ;
  assign \piso.data_r [1599] = \piso.data_r_1599_sv2v_reg ;
  assign \piso.data_r [1598] = \piso.data_r_1598_sv2v_reg ;
  assign \piso.data_r [1597] = \piso.data_r_1597_sv2v_reg ;
  assign \piso.data_r [1596] = \piso.data_r_1596_sv2v_reg ;
  assign \piso.data_r [1595] = \piso.data_r_1595_sv2v_reg ;
  assign \piso.data_r [1594] = \piso.data_r_1594_sv2v_reg ;
  assign \piso.data_r [1593] = \piso.data_r_1593_sv2v_reg ;
  assign \piso.data_r [1592] = \piso.data_r_1592_sv2v_reg ;
  assign \piso.data_r [1591] = \piso.data_r_1591_sv2v_reg ;
  assign \piso.data_r [1590] = \piso.data_r_1590_sv2v_reg ;
  assign \piso.data_r [1589] = \piso.data_r_1589_sv2v_reg ;
  assign \piso.data_r [1588] = \piso.data_r_1588_sv2v_reg ;
  assign \piso.data_r [1587] = \piso.data_r_1587_sv2v_reg ;
  assign \piso.data_r [1586] = \piso.data_r_1586_sv2v_reg ;
  assign \piso.data_r [1585] = \piso.data_r_1585_sv2v_reg ;
  assign \piso.data_r [1584] = \piso.data_r_1584_sv2v_reg ;
  assign \piso.data_r [1583] = \piso.data_r_1583_sv2v_reg ;
  assign \piso.data_r [1582] = \piso.data_r_1582_sv2v_reg ;
  assign \piso.data_r [1581] = \piso.data_r_1581_sv2v_reg ;
  assign \piso.data_r [1580] = \piso.data_r_1580_sv2v_reg ;
  assign \piso.data_r [1579] = \piso.data_r_1579_sv2v_reg ;
  assign \piso.data_r [1578] = \piso.data_r_1578_sv2v_reg ;
  assign \piso.data_r [1577] = \piso.data_r_1577_sv2v_reg ;
  assign \piso.data_r [1576] = \piso.data_r_1576_sv2v_reg ;
  assign \piso.data_r [1575] = \piso.data_r_1575_sv2v_reg ;
  assign \piso.data_r [1574] = \piso.data_r_1574_sv2v_reg ;
  assign \piso.data_r [1573] = \piso.data_r_1573_sv2v_reg ;
  assign \piso.data_r [1572] = \piso.data_r_1572_sv2v_reg ;
  assign \piso.data_r [1571] = \piso.data_r_1571_sv2v_reg ;
  assign \piso.data_r [1570] = \piso.data_r_1570_sv2v_reg ;
  assign \piso.data_r [1569] = \piso.data_r_1569_sv2v_reg ;
  assign \piso.data_r [1568] = \piso.data_r_1568_sv2v_reg ;
  assign \piso.data_r [1567] = \piso.data_r_1567_sv2v_reg ;
  assign \piso.data_r [1566] = \piso.data_r_1566_sv2v_reg ;
  assign \piso.data_r [1565] = \piso.data_r_1565_sv2v_reg ;
  assign \piso.data_r [1564] = \piso.data_r_1564_sv2v_reg ;
  assign \piso.data_r [1563] = \piso.data_r_1563_sv2v_reg ;
  assign \piso.data_r [1562] = \piso.data_r_1562_sv2v_reg ;
  assign \piso.data_r [1561] = \piso.data_r_1561_sv2v_reg ;
  assign \piso.data_r [1560] = \piso.data_r_1560_sv2v_reg ;
  assign \piso.data_r [1559] = \piso.data_r_1559_sv2v_reg ;
  assign \piso.data_r [1558] = \piso.data_r_1558_sv2v_reg ;
  assign \piso.data_r [1557] = \piso.data_r_1557_sv2v_reg ;
  assign \piso.data_r [1556] = \piso.data_r_1556_sv2v_reg ;
  assign \piso.data_r [1555] = \piso.data_r_1555_sv2v_reg ;
  assign \piso.data_r [1554] = \piso.data_r_1554_sv2v_reg ;
  assign \piso.data_r [1553] = \piso.data_r_1553_sv2v_reg ;
  assign \piso.data_r [1552] = \piso.data_r_1552_sv2v_reg ;
  assign \piso.data_r [1551] = \piso.data_r_1551_sv2v_reg ;
  assign \piso.data_r [1550] = \piso.data_r_1550_sv2v_reg ;
  assign \piso.data_r [1549] = \piso.data_r_1549_sv2v_reg ;
  assign \piso.data_r [1548] = \piso.data_r_1548_sv2v_reg ;
  assign \piso.data_r [1547] = \piso.data_r_1547_sv2v_reg ;
  assign \piso.data_r [1546] = \piso.data_r_1546_sv2v_reg ;
  assign \piso.data_r [1545] = \piso.data_r_1545_sv2v_reg ;
  assign \piso.data_r [1544] = \piso.data_r_1544_sv2v_reg ;
  assign \piso.data_r [1543] = \piso.data_r_1543_sv2v_reg ;
  assign \piso.data_r [1542] = \piso.data_r_1542_sv2v_reg ;
  assign \piso.data_r [1541] = \piso.data_r_1541_sv2v_reg ;
  assign \piso.data_r [1540] = \piso.data_r_1540_sv2v_reg ;
  assign \piso.data_r [1539] = \piso.data_r_1539_sv2v_reg ;
  assign \piso.data_r [1538] = \piso.data_r_1538_sv2v_reg ;
  assign \piso.data_r [1537] = \piso.data_r_1537_sv2v_reg ;
  assign \piso.data_r [1536] = \piso.data_r_1536_sv2v_reg ;
  assign \piso.data_r [1535] = \piso.data_r_1535_sv2v_reg ;
  assign \piso.data_r [1534] = \piso.data_r_1534_sv2v_reg ;
  assign \piso.data_r [1533] = \piso.data_r_1533_sv2v_reg ;
  assign \piso.data_r [1532] = \piso.data_r_1532_sv2v_reg ;
  assign \piso.data_r [1531] = \piso.data_r_1531_sv2v_reg ;
  assign \piso.data_r [1530] = \piso.data_r_1530_sv2v_reg ;
  assign \piso.data_r [1529] = \piso.data_r_1529_sv2v_reg ;
  assign \piso.data_r [1528] = \piso.data_r_1528_sv2v_reg ;
  assign \piso.data_r [1527] = \piso.data_r_1527_sv2v_reg ;
  assign \piso.data_r [1526] = \piso.data_r_1526_sv2v_reg ;
  assign \piso.data_r [1525] = \piso.data_r_1525_sv2v_reg ;
  assign \piso.data_r [1524] = \piso.data_r_1524_sv2v_reg ;
  assign \piso.data_r [1523] = \piso.data_r_1523_sv2v_reg ;
  assign \piso.data_r [1522] = \piso.data_r_1522_sv2v_reg ;
  assign \piso.data_r [1521] = \piso.data_r_1521_sv2v_reg ;
  assign \piso.data_r [1520] = \piso.data_r_1520_sv2v_reg ;
  assign \piso.data_r [1519] = \piso.data_r_1519_sv2v_reg ;
  assign \piso.data_r [1518] = \piso.data_r_1518_sv2v_reg ;
  assign \piso.data_r [1517] = \piso.data_r_1517_sv2v_reg ;
  assign \piso.data_r [1516] = \piso.data_r_1516_sv2v_reg ;
  assign \piso.data_r [1515] = \piso.data_r_1515_sv2v_reg ;
  assign \piso.data_r [1514] = \piso.data_r_1514_sv2v_reg ;
  assign \piso.data_r [1513] = \piso.data_r_1513_sv2v_reg ;
  assign \piso.data_r [1512] = \piso.data_r_1512_sv2v_reg ;
  assign \piso.data_r [1511] = \piso.data_r_1511_sv2v_reg ;
  assign \piso.data_r [1510] = \piso.data_r_1510_sv2v_reg ;
  assign \piso.data_r [1509] = \piso.data_r_1509_sv2v_reg ;
  assign \piso.data_r [1508] = \piso.data_r_1508_sv2v_reg ;
  assign \piso.data_r [1507] = \piso.data_r_1507_sv2v_reg ;
  assign \piso.data_r [1506] = \piso.data_r_1506_sv2v_reg ;
  assign \piso.data_r [1505] = \piso.data_r_1505_sv2v_reg ;
  assign \piso.data_r [1504] = \piso.data_r_1504_sv2v_reg ;
  assign \piso.data_r [1503] = \piso.data_r_1503_sv2v_reg ;
  assign \piso.data_r [1502] = \piso.data_r_1502_sv2v_reg ;
  assign \piso.data_r [1501] = \piso.data_r_1501_sv2v_reg ;
  assign \piso.data_r [1500] = \piso.data_r_1500_sv2v_reg ;
  assign \piso.data_r [1499] = \piso.data_r_1499_sv2v_reg ;
  assign \piso.data_r [1498] = \piso.data_r_1498_sv2v_reg ;
  assign \piso.data_r [1497] = \piso.data_r_1497_sv2v_reg ;
  assign \piso.data_r [1496] = \piso.data_r_1496_sv2v_reg ;
  assign \piso.data_r [1495] = \piso.data_r_1495_sv2v_reg ;
  assign \piso.data_r [1494] = \piso.data_r_1494_sv2v_reg ;
  assign \piso.data_r [1493] = \piso.data_r_1493_sv2v_reg ;
  assign \piso.data_r [1492] = \piso.data_r_1492_sv2v_reg ;
  assign \piso.data_r [1491] = \piso.data_r_1491_sv2v_reg ;
  assign \piso.data_r [1490] = \piso.data_r_1490_sv2v_reg ;
  assign \piso.data_r [1489] = \piso.data_r_1489_sv2v_reg ;
  assign \piso.data_r [1488] = \piso.data_r_1488_sv2v_reg ;
  assign \piso.data_r [1487] = \piso.data_r_1487_sv2v_reg ;
  assign \piso.data_r [1486] = \piso.data_r_1486_sv2v_reg ;
  assign \piso.data_r [1485] = \piso.data_r_1485_sv2v_reg ;
  assign \piso.data_r [1484] = \piso.data_r_1484_sv2v_reg ;
  assign \piso.data_r [1483] = \piso.data_r_1483_sv2v_reg ;
  assign \piso.data_r [1482] = \piso.data_r_1482_sv2v_reg ;
  assign \piso.data_r [1481] = \piso.data_r_1481_sv2v_reg ;
  assign \piso.data_r [1480] = \piso.data_r_1480_sv2v_reg ;
  assign \piso.data_r [1479] = \piso.data_r_1479_sv2v_reg ;
  assign \piso.data_r [1478] = \piso.data_r_1478_sv2v_reg ;
  assign \piso.data_r [1477] = \piso.data_r_1477_sv2v_reg ;
  assign \piso.data_r [1476] = \piso.data_r_1476_sv2v_reg ;
  assign \piso.data_r [1475] = \piso.data_r_1475_sv2v_reg ;
  assign \piso.data_r [1474] = \piso.data_r_1474_sv2v_reg ;
  assign \piso.data_r [1473] = \piso.data_r_1473_sv2v_reg ;
  assign \piso.data_r [1472] = \piso.data_r_1472_sv2v_reg ;
  assign \piso.data_r [1471] = \piso.data_r_1471_sv2v_reg ;
  assign \piso.data_r [1470] = \piso.data_r_1470_sv2v_reg ;
  assign \piso.data_r [1469] = \piso.data_r_1469_sv2v_reg ;
  assign \piso.data_r [1468] = \piso.data_r_1468_sv2v_reg ;
  assign \piso.data_r [1467] = \piso.data_r_1467_sv2v_reg ;
  assign \piso.data_r [1466] = \piso.data_r_1466_sv2v_reg ;
  assign \piso.data_r [1465] = \piso.data_r_1465_sv2v_reg ;
  assign \piso.data_r [1464] = \piso.data_r_1464_sv2v_reg ;
  assign \piso.data_r [1463] = \piso.data_r_1463_sv2v_reg ;
  assign \piso.data_r [1462] = \piso.data_r_1462_sv2v_reg ;
  assign \piso.data_r [1461] = \piso.data_r_1461_sv2v_reg ;
  assign \piso.data_r [1460] = \piso.data_r_1460_sv2v_reg ;
  assign \piso.data_r [1459] = \piso.data_r_1459_sv2v_reg ;
  assign \piso.data_r [1458] = \piso.data_r_1458_sv2v_reg ;
  assign \piso.data_r [1457] = \piso.data_r_1457_sv2v_reg ;
  assign \piso.data_r [1456] = \piso.data_r_1456_sv2v_reg ;
  assign \piso.data_r [1455] = \piso.data_r_1455_sv2v_reg ;
  assign \piso.data_r [1454] = \piso.data_r_1454_sv2v_reg ;
  assign \piso.data_r [1453] = \piso.data_r_1453_sv2v_reg ;
  assign \piso.data_r [1452] = \piso.data_r_1452_sv2v_reg ;
  assign \piso.data_r [1451] = \piso.data_r_1451_sv2v_reg ;
  assign \piso.data_r [1450] = \piso.data_r_1450_sv2v_reg ;
  assign \piso.data_r [1449] = \piso.data_r_1449_sv2v_reg ;
  assign \piso.data_r [1448] = \piso.data_r_1448_sv2v_reg ;
  assign \piso.data_r [1447] = \piso.data_r_1447_sv2v_reg ;
  assign \piso.data_r [1446] = \piso.data_r_1446_sv2v_reg ;
  assign \piso.data_r [1445] = \piso.data_r_1445_sv2v_reg ;
  assign \piso.data_r [1444] = \piso.data_r_1444_sv2v_reg ;
  assign \piso.data_r [1443] = \piso.data_r_1443_sv2v_reg ;
  assign \piso.data_r [1442] = \piso.data_r_1442_sv2v_reg ;
  assign \piso.data_r [1441] = \piso.data_r_1441_sv2v_reg ;
  assign \piso.data_r [1440] = \piso.data_r_1440_sv2v_reg ;
  assign \piso.data_r [1439] = \piso.data_r_1439_sv2v_reg ;
  assign \piso.data_r [1438] = \piso.data_r_1438_sv2v_reg ;
  assign \piso.data_r [1437] = \piso.data_r_1437_sv2v_reg ;
  assign \piso.data_r [1436] = \piso.data_r_1436_sv2v_reg ;
  assign \piso.data_r [1435] = \piso.data_r_1435_sv2v_reg ;
  assign \piso.data_r [1434] = \piso.data_r_1434_sv2v_reg ;
  assign \piso.data_r [1433] = \piso.data_r_1433_sv2v_reg ;
  assign \piso.data_r [1432] = \piso.data_r_1432_sv2v_reg ;
  assign \piso.data_r [1431] = \piso.data_r_1431_sv2v_reg ;
  assign \piso.data_r [1430] = \piso.data_r_1430_sv2v_reg ;
  assign \piso.data_r [1429] = \piso.data_r_1429_sv2v_reg ;
  assign \piso.data_r [1428] = \piso.data_r_1428_sv2v_reg ;
  assign \piso.data_r [1427] = \piso.data_r_1427_sv2v_reg ;
  assign \piso.data_r [1426] = \piso.data_r_1426_sv2v_reg ;
  assign \piso.data_r [1425] = \piso.data_r_1425_sv2v_reg ;
  assign \piso.data_r [1424] = \piso.data_r_1424_sv2v_reg ;
  assign \piso.data_r [1423] = \piso.data_r_1423_sv2v_reg ;
  assign \piso.data_r [1422] = \piso.data_r_1422_sv2v_reg ;
  assign \piso.data_r [1421] = \piso.data_r_1421_sv2v_reg ;
  assign \piso.data_r [1420] = \piso.data_r_1420_sv2v_reg ;
  assign \piso.data_r [1419] = \piso.data_r_1419_sv2v_reg ;
  assign \piso.data_r [1418] = \piso.data_r_1418_sv2v_reg ;
  assign \piso.data_r [1417] = \piso.data_r_1417_sv2v_reg ;
  assign \piso.data_r [1416] = \piso.data_r_1416_sv2v_reg ;
  assign \piso.data_r [1415] = \piso.data_r_1415_sv2v_reg ;
  assign \piso.data_r [1414] = \piso.data_r_1414_sv2v_reg ;
  assign \piso.data_r [1413] = \piso.data_r_1413_sv2v_reg ;
  assign \piso.data_r [1412] = \piso.data_r_1412_sv2v_reg ;
  assign \piso.data_r [1411] = \piso.data_r_1411_sv2v_reg ;
  assign \piso.data_r [1410] = \piso.data_r_1410_sv2v_reg ;
  assign \piso.data_r [1409] = \piso.data_r_1409_sv2v_reg ;
  assign \piso.data_r [1408] = \piso.data_r_1408_sv2v_reg ;
  assign \piso.data_r [1407] = \piso.data_r_1407_sv2v_reg ;
  assign \piso.data_r [1406] = \piso.data_r_1406_sv2v_reg ;
  assign \piso.data_r [1405] = \piso.data_r_1405_sv2v_reg ;
  assign \piso.data_r [1404] = \piso.data_r_1404_sv2v_reg ;
  assign \piso.data_r [1403] = \piso.data_r_1403_sv2v_reg ;
  assign \piso.data_r [1402] = \piso.data_r_1402_sv2v_reg ;
  assign \piso.data_r [1401] = \piso.data_r_1401_sv2v_reg ;
  assign \piso.data_r [1400] = \piso.data_r_1400_sv2v_reg ;
  assign \piso.data_r [1399] = \piso.data_r_1399_sv2v_reg ;
  assign \piso.data_r [1398] = \piso.data_r_1398_sv2v_reg ;
  assign \piso.data_r [1397] = \piso.data_r_1397_sv2v_reg ;
  assign \piso.data_r [1396] = \piso.data_r_1396_sv2v_reg ;
  assign \piso.data_r [1395] = \piso.data_r_1395_sv2v_reg ;
  assign \piso.data_r [1394] = \piso.data_r_1394_sv2v_reg ;
  assign \piso.data_r [1393] = \piso.data_r_1393_sv2v_reg ;
  assign \piso.data_r [1392] = \piso.data_r_1392_sv2v_reg ;
  assign \piso.data_r [1391] = \piso.data_r_1391_sv2v_reg ;
  assign \piso.data_r [1390] = \piso.data_r_1390_sv2v_reg ;
  assign \piso.data_r [1389] = \piso.data_r_1389_sv2v_reg ;
  assign \piso.data_r [1388] = \piso.data_r_1388_sv2v_reg ;
  assign \piso.data_r [1387] = \piso.data_r_1387_sv2v_reg ;
  assign \piso.data_r [1386] = \piso.data_r_1386_sv2v_reg ;
  assign \piso.data_r [1385] = \piso.data_r_1385_sv2v_reg ;
  assign \piso.data_r [1384] = \piso.data_r_1384_sv2v_reg ;
  assign \piso.data_r [1383] = \piso.data_r_1383_sv2v_reg ;
  assign \piso.data_r [1382] = \piso.data_r_1382_sv2v_reg ;
  assign \piso.data_r [1381] = \piso.data_r_1381_sv2v_reg ;
  assign \piso.data_r [1380] = \piso.data_r_1380_sv2v_reg ;
  assign \piso.data_r [1379] = \piso.data_r_1379_sv2v_reg ;
  assign \piso.data_r [1378] = \piso.data_r_1378_sv2v_reg ;
  assign \piso.data_r [1377] = \piso.data_r_1377_sv2v_reg ;
  assign \piso.data_r [1376] = \piso.data_r_1376_sv2v_reg ;
  assign \piso.data_r [1375] = \piso.data_r_1375_sv2v_reg ;
  assign \piso.data_r [1374] = \piso.data_r_1374_sv2v_reg ;
  assign \piso.data_r [1373] = \piso.data_r_1373_sv2v_reg ;
  assign \piso.data_r [1372] = \piso.data_r_1372_sv2v_reg ;
  assign \piso.data_r [1371] = \piso.data_r_1371_sv2v_reg ;
  assign \piso.data_r [1370] = \piso.data_r_1370_sv2v_reg ;
  assign \piso.data_r [1369] = \piso.data_r_1369_sv2v_reg ;
  assign \piso.data_r [1368] = \piso.data_r_1368_sv2v_reg ;
  assign \piso.data_r [1367] = \piso.data_r_1367_sv2v_reg ;
  assign \piso.data_r [1366] = \piso.data_r_1366_sv2v_reg ;
  assign \piso.data_r [1365] = \piso.data_r_1365_sv2v_reg ;
  assign \piso.data_r [1364] = \piso.data_r_1364_sv2v_reg ;
  assign \piso.data_r [1363] = \piso.data_r_1363_sv2v_reg ;
  assign \piso.data_r [1362] = \piso.data_r_1362_sv2v_reg ;
  assign \piso.data_r [1361] = \piso.data_r_1361_sv2v_reg ;
  assign \piso.data_r [1360] = \piso.data_r_1360_sv2v_reg ;
  assign \piso.data_r [1359] = \piso.data_r_1359_sv2v_reg ;
  assign \piso.data_r [1358] = \piso.data_r_1358_sv2v_reg ;
  assign \piso.data_r [1357] = \piso.data_r_1357_sv2v_reg ;
  assign \piso.data_r [1356] = \piso.data_r_1356_sv2v_reg ;
  assign \piso.data_r [1355] = \piso.data_r_1355_sv2v_reg ;
  assign \piso.data_r [1354] = \piso.data_r_1354_sv2v_reg ;
  assign \piso.data_r [1353] = \piso.data_r_1353_sv2v_reg ;
  assign \piso.data_r [1352] = \piso.data_r_1352_sv2v_reg ;
  assign \piso.data_r [1351] = \piso.data_r_1351_sv2v_reg ;
  assign \piso.data_r [1350] = \piso.data_r_1350_sv2v_reg ;
  assign \piso.data_r [1349] = \piso.data_r_1349_sv2v_reg ;
  assign \piso.data_r [1348] = \piso.data_r_1348_sv2v_reg ;
  assign \piso.data_r [1347] = \piso.data_r_1347_sv2v_reg ;
  assign \piso.data_r [1346] = \piso.data_r_1346_sv2v_reg ;
  assign \piso.data_r [1345] = \piso.data_r_1345_sv2v_reg ;
  assign \piso.data_r [1344] = \piso.data_r_1344_sv2v_reg ;
  assign \piso.data_r [1343] = \piso.data_r_1343_sv2v_reg ;
  assign \piso.data_r [1342] = \piso.data_r_1342_sv2v_reg ;
  assign \piso.data_r [1341] = \piso.data_r_1341_sv2v_reg ;
  assign \piso.data_r [1340] = \piso.data_r_1340_sv2v_reg ;
  assign \piso.data_r [1339] = \piso.data_r_1339_sv2v_reg ;
  assign \piso.data_r [1338] = \piso.data_r_1338_sv2v_reg ;
  assign \piso.data_r [1337] = \piso.data_r_1337_sv2v_reg ;
  assign \piso.data_r [1336] = \piso.data_r_1336_sv2v_reg ;
  assign \piso.data_r [1335] = \piso.data_r_1335_sv2v_reg ;
  assign \piso.data_r [1334] = \piso.data_r_1334_sv2v_reg ;
  assign \piso.data_r [1333] = \piso.data_r_1333_sv2v_reg ;
  assign \piso.data_r [1332] = \piso.data_r_1332_sv2v_reg ;
  assign \piso.data_r [1331] = \piso.data_r_1331_sv2v_reg ;
  assign \piso.data_r [1330] = \piso.data_r_1330_sv2v_reg ;
  assign \piso.data_r [1329] = \piso.data_r_1329_sv2v_reg ;
  assign \piso.data_r [1328] = \piso.data_r_1328_sv2v_reg ;
  assign \piso.data_r [1327] = \piso.data_r_1327_sv2v_reg ;
  assign \piso.data_r [1326] = \piso.data_r_1326_sv2v_reg ;
  assign \piso.data_r [1325] = \piso.data_r_1325_sv2v_reg ;
  assign \piso.data_r [1324] = \piso.data_r_1324_sv2v_reg ;
  assign \piso.data_r [1323] = \piso.data_r_1323_sv2v_reg ;
  assign \piso.data_r [1322] = \piso.data_r_1322_sv2v_reg ;
  assign \piso.data_r [1321] = \piso.data_r_1321_sv2v_reg ;
  assign \piso.data_r [1320] = \piso.data_r_1320_sv2v_reg ;
  assign \piso.data_r [1319] = \piso.data_r_1319_sv2v_reg ;
  assign \piso.data_r [1318] = \piso.data_r_1318_sv2v_reg ;
  assign \piso.data_r [1317] = \piso.data_r_1317_sv2v_reg ;
  assign \piso.data_r [1316] = \piso.data_r_1316_sv2v_reg ;
  assign \piso.data_r [1315] = \piso.data_r_1315_sv2v_reg ;
  assign \piso.data_r [1314] = \piso.data_r_1314_sv2v_reg ;
  assign \piso.data_r [1313] = \piso.data_r_1313_sv2v_reg ;
  assign \piso.data_r [1312] = \piso.data_r_1312_sv2v_reg ;
  assign \piso.data_r [1311] = \piso.data_r_1311_sv2v_reg ;
  assign \piso.data_r [1310] = \piso.data_r_1310_sv2v_reg ;
  assign \piso.data_r [1309] = \piso.data_r_1309_sv2v_reg ;
  assign \piso.data_r [1308] = \piso.data_r_1308_sv2v_reg ;
  assign \piso.data_r [1307] = \piso.data_r_1307_sv2v_reg ;
  assign \piso.data_r [1306] = \piso.data_r_1306_sv2v_reg ;
  assign \piso.data_r [1305] = \piso.data_r_1305_sv2v_reg ;
  assign \piso.data_r [1304] = \piso.data_r_1304_sv2v_reg ;
  assign \piso.data_r [1303] = \piso.data_r_1303_sv2v_reg ;
  assign \piso.data_r [1302] = \piso.data_r_1302_sv2v_reg ;
  assign \piso.data_r [1301] = \piso.data_r_1301_sv2v_reg ;
  assign \piso.data_r [1300] = \piso.data_r_1300_sv2v_reg ;
  assign \piso.data_r [1299] = \piso.data_r_1299_sv2v_reg ;
  assign \piso.data_r [1298] = \piso.data_r_1298_sv2v_reg ;
  assign \piso.data_r [1297] = \piso.data_r_1297_sv2v_reg ;
  assign \piso.data_r [1296] = \piso.data_r_1296_sv2v_reg ;
  assign \piso.data_r [1295] = \piso.data_r_1295_sv2v_reg ;
  assign \piso.data_r [1294] = \piso.data_r_1294_sv2v_reg ;
  assign \piso.data_r [1293] = \piso.data_r_1293_sv2v_reg ;
  assign \piso.data_r [1292] = \piso.data_r_1292_sv2v_reg ;
  assign \piso.data_r [1291] = \piso.data_r_1291_sv2v_reg ;
  assign \piso.data_r [1290] = \piso.data_r_1290_sv2v_reg ;
  assign \piso.data_r [1289] = \piso.data_r_1289_sv2v_reg ;
  assign \piso.data_r [1288] = \piso.data_r_1288_sv2v_reg ;
  assign \piso.data_r [1287] = \piso.data_r_1287_sv2v_reg ;
  assign \piso.data_r [1286] = \piso.data_r_1286_sv2v_reg ;
  assign \piso.data_r [1285] = \piso.data_r_1285_sv2v_reg ;
  assign \piso.data_r [1284] = \piso.data_r_1284_sv2v_reg ;
  assign \piso.data_r [1283] = \piso.data_r_1283_sv2v_reg ;
  assign \piso.data_r [1282] = \piso.data_r_1282_sv2v_reg ;
  assign \piso.data_r [1281] = \piso.data_r_1281_sv2v_reg ;
  assign \piso.data_r [1280] = \piso.data_r_1280_sv2v_reg ;
  assign \piso.data_r [1279] = \piso.data_r_1279_sv2v_reg ;
  assign \piso.data_r [1278] = \piso.data_r_1278_sv2v_reg ;
  assign \piso.data_r [1277] = \piso.data_r_1277_sv2v_reg ;
  assign \piso.data_r [1276] = \piso.data_r_1276_sv2v_reg ;
  assign \piso.data_r [1275] = \piso.data_r_1275_sv2v_reg ;
  assign \piso.data_r [1274] = \piso.data_r_1274_sv2v_reg ;
  assign \piso.data_r [1273] = \piso.data_r_1273_sv2v_reg ;
  assign \piso.data_r [1272] = \piso.data_r_1272_sv2v_reg ;
  assign \piso.data_r [1271] = \piso.data_r_1271_sv2v_reg ;
  assign \piso.data_r [1270] = \piso.data_r_1270_sv2v_reg ;
  assign \piso.data_r [1269] = \piso.data_r_1269_sv2v_reg ;
  assign \piso.data_r [1268] = \piso.data_r_1268_sv2v_reg ;
  assign \piso.data_r [1267] = \piso.data_r_1267_sv2v_reg ;
  assign \piso.data_r [1266] = \piso.data_r_1266_sv2v_reg ;
  assign \piso.data_r [1265] = \piso.data_r_1265_sv2v_reg ;
  assign \piso.data_r [1264] = \piso.data_r_1264_sv2v_reg ;
  assign \piso.data_r [1263] = \piso.data_r_1263_sv2v_reg ;
  assign \piso.data_r [1262] = \piso.data_r_1262_sv2v_reg ;
  assign \piso.data_r [1261] = \piso.data_r_1261_sv2v_reg ;
  assign \piso.data_r [1260] = \piso.data_r_1260_sv2v_reg ;
  assign \piso.data_r [1259] = \piso.data_r_1259_sv2v_reg ;
  assign \piso.data_r [1258] = \piso.data_r_1258_sv2v_reg ;
  assign \piso.data_r [1257] = \piso.data_r_1257_sv2v_reg ;
  assign \piso.data_r [1256] = \piso.data_r_1256_sv2v_reg ;
  assign \piso.data_r [1255] = \piso.data_r_1255_sv2v_reg ;
  assign \piso.data_r [1254] = \piso.data_r_1254_sv2v_reg ;
  assign \piso.data_r [1253] = \piso.data_r_1253_sv2v_reg ;
  assign \piso.data_r [1252] = \piso.data_r_1252_sv2v_reg ;
  assign \piso.data_r [1251] = \piso.data_r_1251_sv2v_reg ;
  assign \piso.data_r [1250] = \piso.data_r_1250_sv2v_reg ;
  assign \piso.data_r [1249] = \piso.data_r_1249_sv2v_reg ;
  assign \piso.data_r [1248] = \piso.data_r_1248_sv2v_reg ;
  assign \piso.data_r [1247] = \piso.data_r_1247_sv2v_reg ;
  assign \piso.data_r [1246] = \piso.data_r_1246_sv2v_reg ;
  assign \piso.data_r [1245] = \piso.data_r_1245_sv2v_reg ;
  assign \piso.data_r [1244] = \piso.data_r_1244_sv2v_reg ;
  assign \piso.data_r [1243] = \piso.data_r_1243_sv2v_reg ;
  assign \piso.data_r [1242] = \piso.data_r_1242_sv2v_reg ;
  assign \piso.data_r [1241] = \piso.data_r_1241_sv2v_reg ;
  assign \piso.data_r [1240] = \piso.data_r_1240_sv2v_reg ;
  assign \piso.data_r [1239] = \piso.data_r_1239_sv2v_reg ;
  assign \piso.data_r [1238] = \piso.data_r_1238_sv2v_reg ;
  assign \piso.data_r [1237] = \piso.data_r_1237_sv2v_reg ;
  assign \piso.data_r [1236] = \piso.data_r_1236_sv2v_reg ;
  assign \piso.data_r [1235] = \piso.data_r_1235_sv2v_reg ;
  assign \piso.data_r [1234] = \piso.data_r_1234_sv2v_reg ;
  assign \piso.data_r [1233] = \piso.data_r_1233_sv2v_reg ;
  assign \piso.data_r [1232] = \piso.data_r_1232_sv2v_reg ;
  assign \piso.data_r [1231] = \piso.data_r_1231_sv2v_reg ;
  assign \piso.data_r [1230] = \piso.data_r_1230_sv2v_reg ;
  assign \piso.data_r [1229] = \piso.data_r_1229_sv2v_reg ;
  assign \piso.data_r [1228] = \piso.data_r_1228_sv2v_reg ;
  assign \piso.data_r [1227] = \piso.data_r_1227_sv2v_reg ;
  assign \piso.data_r [1226] = \piso.data_r_1226_sv2v_reg ;
  assign \piso.data_r [1225] = \piso.data_r_1225_sv2v_reg ;
  assign \piso.data_r [1224] = \piso.data_r_1224_sv2v_reg ;
  assign \piso.data_r [1223] = \piso.data_r_1223_sv2v_reg ;
  assign \piso.data_r [1222] = \piso.data_r_1222_sv2v_reg ;
  assign \piso.data_r [1221] = \piso.data_r_1221_sv2v_reg ;
  assign \piso.data_r [1220] = \piso.data_r_1220_sv2v_reg ;
  assign \piso.data_r [1219] = \piso.data_r_1219_sv2v_reg ;
  assign \piso.data_r [1218] = \piso.data_r_1218_sv2v_reg ;
  assign \piso.data_r [1217] = \piso.data_r_1217_sv2v_reg ;
  assign \piso.data_r [1216] = \piso.data_r_1216_sv2v_reg ;
  assign \piso.data_r [1215] = \piso.data_r_1215_sv2v_reg ;
  assign \piso.data_r [1214] = \piso.data_r_1214_sv2v_reg ;
  assign \piso.data_r [1213] = \piso.data_r_1213_sv2v_reg ;
  assign \piso.data_r [1212] = \piso.data_r_1212_sv2v_reg ;
  assign \piso.data_r [1211] = \piso.data_r_1211_sv2v_reg ;
  assign \piso.data_r [1210] = \piso.data_r_1210_sv2v_reg ;
  assign \piso.data_r [1209] = \piso.data_r_1209_sv2v_reg ;
  assign \piso.data_r [1208] = \piso.data_r_1208_sv2v_reg ;
  assign \piso.data_r [1207] = \piso.data_r_1207_sv2v_reg ;
  assign \piso.data_r [1206] = \piso.data_r_1206_sv2v_reg ;
  assign \piso.data_r [1205] = \piso.data_r_1205_sv2v_reg ;
  assign \piso.data_r [1204] = \piso.data_r_1204_sv2v_reg ;
  assign \piso.data_r [1203] = \piso.data_r_1203_sv2v_reg ;
  assign \piso.data_r [1202] = \piso.data_r_1202_sv2v_reg ;
  assign \piso.data_r [1201] = \piso.data_r_1201_sv2v_reg ;
  assign \piso.data_r [1200] = \piso.data_r_1200_sv2v_reg ;
  assign \piso.data_r [1199] = \piso.data_r_1199_sv2v_reg ;
  assign \piso.data_r [1198] = \piso.data_r_1198_sv2v_reg ;
  assign \piso.data_r [1197] = \piso.data_r_1197_sv2v_reg ;
  assign \piso.data_r [1196] = \piso.data_r_1196_sv2v_reg ;
  assign \piso.data_r [1195] = \piso.data_r_1195_sv2v_reg ;
  assign \piso.data_r [1194] = \piso.data_r_1194_sv2v_reg ;
  assign \piso.data_r [1193] = \piso.data_r_1193_sv2v_reg ;
  assign \piso.data_r [1192] = \piso.data_r_1192_sv2v_reg ;
  assign \piso.data_r [1191] = \piso.data_r_1191_sv2v_reg ;
  assign \piso.data_r [1190] = \piso.data_r_1190_sv2v_reg ;
  assign \piso.data_r [1189] = \piso.data_r_1189_sv2v_reg ;
  assign \piso.data_r [1188] = \piso.data_r_1188_sv2v_reg ;
  assign \piso.data_r [1187] = \piso.data_r_1187_sv2v_reg ;
  assign \piso.data_r [1186] = \piso.data_r_1186_sv2v_reg ;
  assign \piso.data_r [1185] = \piso.data_r_1185_sv2v_reg ;
  assign \piso.data_r [1184] = \piso.data_r_1184_sv2v_reg ;
  assign \piso.data_r [1183] = \piso.data_r_1183_sv2v_reg ;
  assign \piso.data_r [1182] = \piso.data_r_1182_sv2v_reg ;
  assign \piso.data_r [1181] = \piso.data_r_1181_sv2v_reg ;
  assign \piso.data_r [1180] = \piso.data_r_1180_sv2v_reg ;
  assign \piso.data_r [1179] = \piso.data_r_1179_sv2v_reg ;
  assign \piso.data_r [1178] = \piso.data_r_1178_sv2v_reg ;
  assign \piso.data_r [1177] = \piso.data_r_1177_sv2v_reg ;
  assign \piso.data_r [1176] = \piso.data_r_1176_sv2v_reg ;
  assign \piso.data_r [1175] = \piso.data_r_1175_sv2v_reg ;
  assign \piso.data_r [1174] = \piso.data_r_1174_sv2v_reg ;
  assign \piso.data_r [1173] = \piso.data_r_1173_sv2v_reg ;
  assign \piso.data_r [1172] = \piso.data_r_1172_sv2v_reg ;
  assign \piso.data_r [1171] = \piso.data_r_1171_sv2v_reg ;
  assign \piso.data_r [1170] = \piso.data_r_1170_sv2v_reg ;
  assign \piso.data_r [1169] = \piso.data_r_1169_sv2v_reg ;
  assign \piso.data_r [1168] = \piso.data_r_1168_sv2v_reg ;
  assign \piso.data_r [1167] = \piso.data_r_1167_sv2v_reg ;
  assign \piso.data_r [1166] = \piso.data_r_1166_sv2v_reg ;
  assign \piso.data_r [1165] = \piso.data_r_1165_sv2v_reg ;
  assign \piso.data_r [1164] = \piso.data_r_1164_sv2v_reg ;
  assign \piso.data_r [1163] = \piso.data_r_1163_sv2v_reg ;
  assign \piso.data_r [1162] = \piso.data_r_1162_sv2v_reg ;
  assign \piso.data_r [1161] = \piso.data_r_1161_sv2v_reg ;
  assign \piso.data_r [1160] = \piso.data_r_1160_sv2v_reg ;
  assign \piso.data_r [1159] = \piso.data_r_1159_sv2v_reg ;
  assign \piso.data_r [1158] = \piso.data_r_1158_sv2v_reg ;
  assign \piso.data_r [1157] = \piso.data_r_1157_sv2v_reg ;
  assign \piso.data_r [1156] = \piso.data_r_1156_sv2v_reg ;
  assign \piso.data_r [1155] = \piso.data_r_1155_sv2v_reg ;
  assign \piso.data_r [1154] = \piso.data_r_1154_sv2v_reg ;
  assign \piso.data_r [1153] = \piso.data_r_1153_sv2v_reg ;
  assign \piso.data_r [1152] = \piso.data_r_1152_sv2v_reg ;
  assign \piso.data_r [1151] = \piso.data_r_1151_sv2v_reg ;
  assign \piso.data_r [1150] = \piso.data_r_1150_sv2v_reg ;
  assign \piso.data_r [1149] = \piso.data_r_1149_sv2v_reg ;
  assign \piso.data_r [1148] = \piso.data_r_1148_sv2v_reg ;
  assign \piso.data_r [1147] = \piso.data_r_1147_sv2v_reg ;
  assign \piso.data_r [1146] = \piso.data_r_1146_sv2v_reg ;
  assign \piso.data_r [1145] = \piso.data_r_1145_sv2v_reg ;
  assign \piso.data_r [1144] = \piso.data_r_1144_sv2v_reg ;
  assign \piso.data_r [1143] = \piso.data_r_1143_sv2v_reg ;
  assign \piso.data_r [1142] = \piso.data_r_1142_sv2v_reg ;
  assign \piso.data_r [1141] = \piso.data_r_1141_sv2v_reg ;
  assign \piso.data_r [1140] = \piso.data_r_1140_sv2v_reg ;
  assign \piso.data_r [1139] = \piso.data_r_1139_sv2v_reg ;
  assign \piso.data_r [1138] = \piso.data_r_1138_sv2v_reg ;
  assign \piso.data_r [1137] = \piso.data_r_1137_sv2v_reg ;
  assign \piso.data_r [1136] = \piso.data_r_1136_sv2v_reg ;
  assign \piso.data_r [1135] = \piso.data_r_1135_sv2v_reg ;
  assign \piso.data_r [1134] = \piso.data_r_1134_sv2v_reg ;
  assign \piso.data_r [1133] = \piso.data_r_1133_sv2v_reg ;
  assign \piso.data_r [1132] = \piso.data_r_1132_sv2v_reg ;
  assign \piso.data_r [1131] = \piso.data_r_1131_sv2v_reg ;
  assign \piso.data_r [1130] = \piso.data_r_1130_sv2v_reg ;
  assign \piso.data_r [1129] = \piso.data_r_1129_sv2v_reg ;
  assign \piso.data_r [1128] = \piso.data_r_1128_sv2v_reg ;
  assign \piso.data_r [1127] = \piso.data_r_1127_sv2v_reg ;
  assign \piso.data_r [1126] = \piso.data_r_1126_sv2v_reg ;
  assign \piso.data_r [1125] = \piso.data_r_1125_sv2v_reg ;
  assign \piso.data_r [1124] = \piso.data_r_1124_sv2v_reg ;
  assign \piso.data_r [1123] = \piso.data_r_1123_sv2v_reg ;
  assign \piso.data_r [1122] = \piso.data_r_1122_sv2v_reg ;
  assign \piso.data_r [1121] = \piso.data_r_1121_sv2v_reg ;
  assign \piso.data_r [1120] = \piso.data_r_1120_sv2v_reg ;
  assign \piso.data_r [1119] = \piso.data_r_1119_sv2v_reg ;
  assign \piso.data_r [1118] = \piso.data_r_1118_sv2v_reg ;
  assign \piso.data_r [1117] = \piso.data_r_1117_sv2v_reg ;
  assign \piso.data_r [1116] = \piso.data_r_1116_sv2v_reg ;
  assign \piso.data_r [1115] = \piso.data_r_1115_sv2v_reg ;
  assign \piso.data_r [1114] = \piso.data_r_1114_sv2v_reg ;
  assign \piso.data_r [1113] = \piso.data_r_1113_sv2v_reg ;
  assign \piso.data_r [1112] = \piso.data_r_1112_sv2v_reg ;
  assign \piso.data_r [1111] = \piso.data_r_1111_sv2v_reg ;
  assign \piso.data_r [1110] = \piso.data_r_1110_sv2v_reg ;
  assign \piso.data_r [1109] = \piso.data_r_1109_sv2v_reg ;
  assign \piso.data_r [1108] = \piso.data_r_1108_sv2v_reg ;
  assign \piso.data_r [1107] = \piso.data_r_1107_sv2v_reg ;
  assign \piso.data_r [1106] = \piso.data_r_1106_sv2v_reg ;
  assign \piso.data_r [1105] = \piso.data_r_1105_sv2v_reg ;
  assign \piso.data_r [1104] = \piso.data_r_1104_sv2v_reg ;
  assign \piso.data_r [1103] = \piso.data_r_1103_sv2v_reg ;
  assign \piso.data_r [1102] = \piso.data_r_1102_sv2v_reg ;
  assign \piso.data_r [1101] = \piso.data_r_1101_sv2v_reg ;
  assign \piso.data_r [1100] = \piso.data_r_1100_sv2v_reg ;
  assign \piso.data_r [1099] = \piso.data_r_1099_sv2v_reg ;
  assign \piso.data_r [1098] = \piso.data_r_1098_sv2v_reg ;
  assign \piso.data_r [1097] = \piso.data_r_1097_sv2v_reg ;
  assign \piso.data_r [1096] = \piso.data_r_1096_sv2v_reg ;
  assign \piso.data_r [1095] = \piso.data_r_1095_sv2v_reg ;
  assign \piso.data_r [1094] = \piso.data_r_1094_sv2v_reg ;
  assign \piso.data_r [1093] = \piso.data_r_1093_sv2v_reg ;
  assign \piso.data_r [1092] = \piso.data_r_1092_sv2v_reg ;
  assign \piso.data_r [1091] = \piso.data_r_1091_sv2v_reg ;
  assign \piso.data_r [1090] = \piso.data_r_1090_sv2v_reg ;
  assign \piso.data_r [1089] = \piso.data_r_1089_sv2v_reg ;
  assign \piso.data_r [1088] = \piso.data_r_1088_sv2v_reg ;
  assign \piso.data_r [1087] = \piso.data_r_1087_sv2v_reg ;
  assign \piso.data_r [1086] = \piso.data_r_1086_sv2v_reg ;
  assign \piso.data_r [1085] = \piso.data_r_1085_sv2v_reg ;
  assign \piso.data_r [1084] = \piso.data_r_1084_sv2v_reg ;
  assign \piso.data_r [1083] = \piso.data_r_1083_sv2v_reg ;
  assign \piso.data_r [1082] = \piso.data_r_1082_sv2v_reg ;
  assign \piso.data_r [1081] = \piso.data_r_1081_sv2v_reg ;
  assign \piso.data_r [1080] = \piso.data_r_1080_sv2v_reg ;
  assign \piso.data_r [1079] = \piso.data_r_1079_sv2v_reg ;
  assign \piso.data_r [1078] = \piso.data_r_1078_sv2v_reg ;
  assign \piso.data_r [1077] = \piso.data_r_1077_sv2v_reg ;
  assign \piso.data_r [1076] = \piso.data_r_1076_sv2v_reg ;
  assign \piso.data_r [1075] = \piso.data_r_1075_sv2v_reg ;
  assign \piso.data_r [1074] = \piso.data_r_1074_sv2v_reg ;
  assign \piso.data_r [1073] = \piso.data_r_1073_sv2v_reg ;
  assign \piso.data_r [1072] = \piso.data_r_1072_sv2v_reg ;
  assign \piso.data_r [1071] = \piso.data_r_1071_sv2v_reg ;
  assign \piso.data_r [1070] = \piso.data_r_1070_sv2v_reg ;
  assign \piso.data_r [1069] = \piso.data_r_1069_sv2v_reg ;
  assign \piso.data_r [1068] = \piso.data_r_1068_sv2v_reg ;
  assign \piso.data_r [1067] = \piso.data_r_1067_sv2v_reg ;
  assign \piso.data_r [1066] = \piso.data_r_1066_sv2v_reg ;
  assign \piso.data_r [1065] = \piso.data_r_1065_sv2v_reg ;
  assign \piso.data_r [1064] = \piso.data_r_1064_sv2v_reg ;
  assign \piso.data_r [1063] = \piso.data_r_1063_sv2v_reg ;
  assign \piso.data_r [1062] = \piso.data_r_1062_sv2v_reg ;
  assign \piso.data_r [1061] = \piso.data_r_1061_sv2v_reg ;
  assign \piso.data_r [1060] = \piso.data_r_1060_sv2v_reg ;
  assign \piso.data_r [1059] = \piso.data_r_1059_sv2v_reg ;
  assign \piso.data_r [1058] = \piso.data_r_1058_sv2v_reg ;
  assign \piso.data_r [1057] = \piso.data_r_1057_sv2v_reg ;
  assign \piso.data_r [1056] = \piso.data_r_1056_sv2v_reg ;
  assign \piso.data_r [1055] = \piso.data_r_1055_sv2v_reg ;
  assign \piso.data_r [1054] = \piso.data_r_1054_sv2v_reg ;
  assign \piso.data_r [1053] = \piso.data_r_1053_sv2v_reg ;
  assign \piso.data_r [1052] = \piso.data_r_1052_sv2v_reg ;
  assign \piso.data_r [1051] = \piso.data_r_1051_sv2v_reg ;
  assign \piso.data_r [1050] = \piso.data_r_1050_sv2v_reg ;
  assign \piso.data_r [1049] = \piso.data_r_1049_sv2v_reg ;
  assign \piso.data_r [1048] = \piso.data_r_1048_sv2v_reg ;
  assign \piso.data_r [1047] = \piso.data_r_1047_sv2v_reg ;
  assign \piso.data_r [1046] = \piso.data_r_1046_sv2v_reg ;
  assign \piso.data_r [1045] = \piso.data_r_1045_sv2v_reg ;
  assign \piso.data_r [1044] = \piso.data_r_1044_sv2v_reg ;
  assign \piso.data_r [1043] = \piso.data_r_1043_sv2v_reg ;
  assign \piso.data_r [1042] = \piso.data_r_1042_sv2v_reg ;
  assign \piso.data_r [1041] = \piso.data_r_1041_sv2v_reg ;
  assign \piso.data_r [1040] = \piso.data_r_1040_sv2v_reg ;
  assign \piso.data_r [1039] = \piso.data_r_1039_sv2v_reg ;
  assign \piso.data_r [1038] = \piso.data_r_1038_sv2v_reg ;
  assign \piso.data_r [1037] = \piso.data_r_1037_sv2v_reg ;
  assign \piso.data_r [1036] = \piso.data_r_1036_sv2v_reg ;
  assign \piso.data_r [1035] = \piso.data_r_1035_sv2v_reg ;
  assign \piso.data_r [1034] = \piso.data_r_1034_sv2v_reg ;
  assign \piso.data_r [1033] = \piso.data_r_1033_sv2v_reg ;
  assign \piso.data_r [1032] = \piso.data_r_1032_sv2v_reg ;
  assign \piso.data_r [1031] = \piso.data_r_1031_sv2v_reg ;
  assign \piso.data_r [1030] = \piso.data_r_1030_sv2v_reg ;
  assign \piso.data_r [1029] = \piso.data_r_1029_sv2v_reg ;
  assign \piso.data_r [1028] = \piso.data_r_1028_sv2v_reg ;
  assign \piso.data_r [1027] = \piso.data_r_1027_sv2v_reg ;
  assign \piso.data_r [1026] = \piso.data_r_1026_sv2v_reg ;
  assign \piso.data_r [1025] = \piso.data_r_1025_sv2v_reg ;
  assign \piso.data_r [1024] = \piso.data_r_1024_sv2v_reg ;
  assign \piso.data_r [1023] = \piso.data_r_1023_sv2v_reg ;
  assign \piso.data_r [1022] = \piso.data_r_1022_sv2v_reg ;
  assign \piso.data_r [1021] = \piso.data_r_1021_sv2v_reg ;
  assign \piso.data_r [1020] = \piso.data_r_1020_sv2v_reg ;
  assign \piso.data_r [1019] = \piso.data_r_1019_sv2v_reg ;
  assign \piso.data_r [1018] = \piso.data_r_1018_sv2v_reg ;
  assign \piso.data_r [1017] = \piso.data_r_1017_sv2v_reg ;
  assign \piso.data_r [1016] = \piso.data_r_1016_sv2v_reg ;
  assign \piso.data_r [1015] = \piso.data_r_1015_sv2v_reg ;
  assign \piso.data_r [1014] = \piso.data_r_1014_sv2v_reg ;
  assign \piso.data_r [1013] = \piso.data_r_1013_sv2v_reg ;
  assign \piso.data_r [1012] = \piso.data_r_1012_sv2v_reg ;
  assign \piso.data_r [1011] = \piso.data_r_1011_sv2v_reg ;
  assign \piso.data_r [1010] = \piso.data_r_1010_sv2v_reg ;
  assign \piso.data_r [1009] = \piso.data_r_1009_sv2v_reg ;
  assign \piso.data_r [1008] = \piso.data_r_1008_sv2v_reg ;
  assign \piso.data_r [1007] = \piso.data_r_1007_sv2v_reg ;
  assign \piso.data_r [1006] = \piso.data_r_1006_sv2v_reg ;
  assign \piso.data_r [1005] = \piso.data_r_1005_sv2v_reg ;
  assign \piso.data_r [1004] = \piso.data_r_1004_sv2v_reg ;
  assign \piso.data_r [1003] = \piso.data_r_1003_sv2v_reg ;
  assign \piso.data_r [1002] = \piso.data_r_1002_sv2v_reg ;
  assign \piso.data_r [1001] = \piso.data_r_1001_sv2v_reg ;
  assign \piso.data_r [1000] = \piso.data_r_1000_sv2v_reg ;
  assign \piso.data_r [999] = \piso.data_r_999_sv2v_reg ;
  assign \piso.data_r [998] = \piso.data_r_998_sv2v_reg ;
  assign \piso.data_r [997] = \piso.data_r_997_sv2v_reg ;
  assign \piso.data_r [996] = \piso.data_r_996_sv2v_reg ;
  assign \piso.data_r [995] = \piso.data_r_995_sv2v_reg ;
  assign \piso.data_r [994] = \piso.data_r_994_sv2v_reg ;
  assign \piso.data_r [993] = \piso.data_r_993_sv2v_reg ;
  assign \piso.data_r [992] = \piso.data_r_992_sv2v_reg ;
  assign \piso.data_r [991] = \piso.data_r_991_sv2v_reg ;
  assign \piso.data_r [990] = \piso.data_r_990_sv2v_reg ;
  assign \piso.data_r [989] = \piso.data_r_989_sv2v_reg ;
  assign \piso.data_r [988] = \piso.data_r_988_sv2v_reg ;
  assign \piso.data_r [987] = \piso.data_r_987_sv2v_reg ;
  assign \piso.data_r [986] = \piso.data_r_986_sv2v_reg ;
  assign \piso.data_r [985] = \piso.data_r_985_sv2v_reg ;
  assign \piso.data_r [984] = \piso.data_r_984_sv2v_reg ;
  assign \piso.data_r [983] = \piso.data_r_983_sv2v_reg ;
  assign \piso.data_r [982] = \piso.data_r_982_sv2v_reg ;
  assign \piso.data_r [981] = \piso.data_r_981_sv2v_reg ;
  assign \piso.data_r [980] = \piso.data_r_980_sv2v_reg ;
  assign \piso.data_r [979] = \piso.data_r_979_sv2v_reg ;
  assign \piso.data_r [978] = \piso.data_r_978_sv2v_reg ;
  assign \piso.data_r [977] = \piso.data_r_977_sv2v_reg ;
  assign \piso.data_r [976] = \piso.data_r_976_sv2v_reg ;
  assign \piso.data_r [975] = \piso.data_r_975_sv2v_reg ;
  assign \piso.data_r [974] = \piso.data_r_974_sv2v_reg ;
  assign \piso.data_r [973] = \piso.data_r_973_sv2v_reg ;
  assign \piso.data_r [972] = \piso.data_r_972_sv2v_reg ;
  assign \piso.data_r [971] = \piso.data_r_971_sv2v_reg ;
  assign \piso.data_r [970] = \piso.data_r_970_sv2v_reg ;
  assign \piso.data_r [969] = \piso.data_r_969_sv2v_reg ;
  assign \piso.data_r [968] = \piso.data_r_968_sv2v_reg ;
  assign \piso.data_r [967] = \piso.data_r_967_sv2v_reg ;
  assign \piso.data_r [966] = \piso.data_r_966_sv2v_reg ;
  assign \piso.data_r [965] = \piso.data_r_965_sv2v_reg ;
  assign \piso.data_r [964] = \piso.data_r_964_sv2v_reg ;
  assign \piso.data_r [963] = \piso.data_r_963_sv2v_reg ;
  assign \piso.data_r [962] = \piso.data_r_962_sv2v_reg ;
  assign \piso.data_r [961] = \piso.data_r_961_sv2v_reg ;
  assign \piso.data_r [960] = \piso.data_r_960_sv2v_reg ;
  assign \piso.data_r [959] = \piso.data_r_959_sv2v_reg ;
  assign \piso.data_r [958] = \piso.data_r_958_sv2v_reg ;
  assign \piso.data_r [957] = \piso.data_r_957_sv2v_reg ;
  assign \piso.data_r [956] = \piso.data_r_956_sv2v_reg ;
  assign \piso.data_r [955] = \piso.data_r_955_sv2v_reg ;
  assign \piso.data_r [954] = \piso.data_r_954_sv2v_reg ;
  assign \piso.data_r [953] = \piso.data_r_953_sv2v_reg ;
  assign \piso.data_r [952] = \piso.data_r_952_sv2v_reg ;
  assign \piso.data_r [951] = \piso.data_r_951_sv2v_reg ;
  assign \piso.data_r [950] = \piso.data_r_950_sv2v_reg ;
  assign \piso.data_r [949] = \piso.data_r_949_sv2v_reg ;
  assign \piso.data_r [948] = \piso.data_r_948_sv2v_reg ;
  assign \piso.data_r [947] = \piso.data_r_947_sv2v_reg ;
  assign \piso.data_r [946] = \piso.data_r_946_sv2v_reg ;
  assign \piso.data_r [945] = \piso.data_r_945_sv2v_reg ;
  assign \piso.data_r [944] = \piso.data_r_944_sv2v_reg ;
  assign \piso.data_r [943] = \piso.data_r_943_sv2v_reg ;
  assign \piso.data_r [942] = \piso.data_r_942_sv2v_reg ;
  assign \piso.data_r [941] = \piso.data_r_941_sv2v_reg ;
  assign \piso.data_r [940] = \piso.data_r_940_sv2v_reg ;
  assign \piso.data_r [939] = \piso.data_r_939_sv2v_reg ;
  assign \piso.data_r [938] = \piso.data_r_938_sv2v_reg ;
  assign \piso.data_r [937] = \piso.data_r_937_sv2v_reg ;
  assign \piso.data_r [936] = \piso.data_r_936_sv2v_reg ;
  assign \piso.data_r [935] = \piso.data_r_935_sv2v_reg ;
  assign \piso.data_r [934] = \piso.data_r_934_sv2v_reg ;
  assign \piso.data_r [933] = \piso.data_r_933_sv2v_reg ;
  assign \piso.data_r [932] = \piso.data_r_932_sv2v_reg ;
  assign \piso.data_r [931] = \piso.data_r_931_sv2v_reg ;
  assign \piso.data_r [930] = \piso.data_r_930_sv2v_reg ;
  assign \piso.data_r [929] = \piso.data_r_929_sv2v_reg ;
  assign \piso.data_r [928] = \piso.data_r_928_sv2v_reg ;
  assign \piso.data_r [927] = \piso.data_r_927_sv2v_reg ;
  assign \piso.data_r [926] = \piso.data_r_926_sv2v_reg ;
  assign \piso.data_r [925] = \piso.data_r_925_sv2v_reg ;
  assign \piso.data_r [924] = \piso.data_r_924_sv2v_reg ;
  assign \piso.data_r [923] = \piso.data_r_923_sv2v_reg ;
  assign \piso.data_r [922] = \piso.data_r_922_sv2v_reg ;
  assign \piso.data_r [921] = \piso.data_r_921_sv2v_reg ;
  assign \piso.data_r [920] = \piso.data_r_920_sv2v_reg ;
  assign \piso.data_r [919] = \piso.data_r_919_sv2v_reg ;
  assign \piso.data_r [918] = \piso.data_r_918_sv2v_reg ;
  assign \piso.data_r [917] = \piso.data_r_917_sv2v_reg ;
  assign \piso.data_r [916] = \piso.data_r_916_sv2v_reg ;
  assign \piso.data_r [915] = \piso.data_r_915_sv2v_reg ;
  assign \piso.data_r [914] = \piso.data_r_914_sv2v_reg ;
  assign \piso.data_r [913] = \piso.data_r_913_sv2v_reg ;
  assign \piso.data_r [912] = \piso.data_r_912_sv2v_reg ;
  assign \piso.data_r [911] = \piso.data_r_911_sv2v_reg ;
  assign \piso.data_r [910] = \piso.data_r_910_sv2v_reg ;
  assign \piso.data_r [909] = \piso.data_r_909_sv2v_reg ;
  assign \piso.data_r [908] = \piso.data_r_908_sv2v_reg ;
  assign \piso.data_r [907] = \piso.data_r_907_sv2v_reg ;
  assign \piso.data_r [906] = \piso.data_r_906_sv2v_reg ;
  assign \piso.data_r [905] = \piso.data_r_905_sv2v_reg ;
  assign \piso.data_r [904] = \piso.data_r_904_sv2v_reg ;
  assign \piso.data_r [903] = \piso.data_r_903_sv2v_reg ;
  assign \piso.data_r [902] = \piso.data_r_902_sv2v_reg ;
  assign \piso.data_r [901] = \piso.data_r_901_sv2v_reg ;
  assign \piso.data_r [900] = \piso.data_r_900_sv2v_reg ;
  assign \piso.data_r [899] = \piso.data_r_899_sv2v_reg ;
  assign \piso.data_r [898] = \piso.data_r_898_sv2v_reg ;
  assign \piso.data_r [897] = \piso.data_r_897_sv2v_reg ;
  assign \piso.data_r [896] = \piso.data_r_896_sv2v_reg ;
  assign \piso.data_r [895] = \piso.data_r_895_sv2v_reg ;
  assign \piso.data_r [894] = \piso.data_r_894_sv2v_reg ;
  assign \piso.data_r [893] = \piso.data_r_893_sv2v_reg ;
  assign \piso.data_r [892] = \piso.data_r_892_sv2v_reg ;
  assign \piso.data_r [891] = \piso.data_r_891_sv2v_reg ;
  assign \piso.data_r [890] = \piso.data_r_890_sv2v_reg ;
  assign \piso.data_r [889] = \piso.data_r_889_sv2v_reg ;
  assign \piso.data_r [888] = \piso.data_r_888_sv2v_reg ;
  assign \piso.data_r [887] = \piso.data_r_887_sv2v_reg ;
  assign \piso.data_r [886] = \piso.data_r_886_sv2v_reg ;
  assign \piso.data_r [885] = \piso.data_r_885_sv2v_reg ;
  assign \piso.data_r [884] = \piso.data_r_884_sv2v_reg ;
  assign \piso.data_r [883] = \piso.data_r_883_sv2v_reg ;
  assign \piso.data_r [882] = \piso.data_r_882_sv2v_reg ;
  assign \piso.data_r [881] = \piso.data_r_881_sv2v_reg ;
  assign \piso.data_r [880] = \piso.data_r_880_sv2v_reg ;
  assign \piso.data_r [879] = \piso.data_r_879_sv2v_reg ;
  assign \piso.data_r [878] = \piso.data_r_878_sv2v_reg ;
  assign \piso.data_r [877] = \piso.data_r_877_sv2v_reg ;
  assign \piso.data_r [876] = \piso.data_r_876_sv2v_reg ;
  assign \piso.data_r [875] = \piso.data_r_875_sv2v_reg ;
  assign \piso.data_r [874] = \piso.data_r_874_sv2v_reg ;
  assign \piso.data_r [873] = \piso.data_r_873_sv2v_reg ;
  assign \piso.data_r [872] = \piso.data_r_872_sv2v_reg ;
  assign \piso.data_r [871] = \piso.data_r_871_sv2v_reg ;
  assign \piso.data_r [870] = \piso.data_r_870_sv2v_reg ;
  assign \piso.data_r [869] = \piso.data_r_869_sv2v_reg ;
  assign \piso.data_r [868] = \piso.data_r_868_sv2v_reg ;
  assign \piso.data_r [867] = \piso.data_r_867_sv2v_reg ;
  assign \piso.data_r [866] = \piso.data_r_866_sv2v_reg ;
  assign \piso.data_r [865] = \piso.data_r_865_sv2v_reg ;
  assign \piso.data_r [864] = \piso.data_r_864_sv2v_reg ;
  assign \piso.data_r [863] = \piso.data_r_863_sv2v_reg ;
  assign \piso.data_r [862] = \piso.data_r_862_sv2v_reg ;
  assign \piso.data_r [861] = \piso.data_r_861_sv2v_reg ;
  assign \piso.data_r [860] = \piso.data_r_860_sv2v_reg ;
  assign \piso.data_r [859] = \piso.data_r_859_sv2v_reg ;
  assign \piso.data_r [858] = \piso.data_r_858_sv2v_reg ;
  assign \piso.data_r [857] = \piso.data_r_857_sv2v_reg ;
  assign \piso.data_r [856] = \piso.data_r_856_sv2v_reg ;
  assign \piso.data_r [855] = \piso.data_r_855_sv2v_reg ;
  assign \piso.data_r [854] = \piso.data_r_854_sv2v_reg ;
  assign \piso.data_r [853] = \piso.data_r_853_sv2v_reg ;
  assign \piso.data_r [852] = \piso.data_r_852_sv2v_reg ;
  assign \piso.data_r [851] = \piso.data_r_851_sv2v_reg ;
  assign \piso.data_r [850] = \piso.data_r_850_sv2v_reg ;
  assign \piso.data_r [849] = \piso.data_r_849_sv2v_reg ;
  assign \piso.data_r [848] = \piso.data_r_848_sv2v_reg ;
  assign \piso.data_r [847] = \piso.data_r_847_sv2v_reg ;
  assign \piso.data_r [846] = \piso.data_r_846_sv2v_reg ;
  assign \piso.data_r [845] = \piso.data_r_845_sv2v_reg ;
  assign \piso.data_r [844] = \piso.data_r_844_sv2v_reg ;
  assign \piso.data_r [843] = \piso.data_r_843_sv2v_reg ;
  assign \piso.data_r [842] = \piso.data_r_842_sv2v_reg ;
  assign \piso.data_r [841] = \piso.data_r_841_sv2v_reg ;
  assign \piso.data_r [840] = \piso.data_r_840_sv2v_reg ;
  assign \piso.data_r [839] = \piso.data_r_839_sv2v_reg ;
  assign \piso.data_r [838] = \piso.data_r_838_sv2v_reg ;
  assign \piso.data_r [837] = \piso.data_r_837_sv2v_reg ;
  assign \piso.data_r [836] = \piso.data_r_836_sv2v_reg ;
  assign \piso.data_r [835] = \piso.data_r_835_sv2v_reg ;
  assign \piso.data_r [834] = \piso.data_r_834_sv2v_reg ;
  assign \piso.data_r [833] = \piso.data_r_833_sv2v_reg ;
  assign \piso.data_r [832] = \piso.data_r_832_sv2v_reg ;
  assign \piso.data_r [831] = \piso.data_r_831_sv2v_reg ;
  assign \piso.data_r [830] = \piso.data_r_830_sv2v_reg ;
  assign \piso.data_r [829] = \piso.data_r_829_sv2v_reg ;
  assign \piso.data_r [828] = \piso.data_r_828_sv2v_reg ;
  assign \piso.data_r [827] = \piso.data_r_827_sv2v_reg ;
  assign \piso.data_r [826] = \piso.data_r_826_sv2v_reg ;
  assign \piso.data_r [825] = \piso.data_r_825_sv2v_reg ;
  assign \piso.data_r [824] = \piso.data_r_824_sv2v_reg ;
  assign \piso.data_r [823] = \piso.data_r_823_sv2v_reg ;
  assign \piso.data_r [822] = \piso.data_r_822_sv2v_reg ;
  assign \piso.data_r [821] = \piso.data_r_821_sv2v_reg ;
  assign \piso.data_r [820] = \piso.data_r_820_sv2v_reg ;
  assign \piso.data_r [819] = \piso.data_r_819_sv2v_reg ;
  assign \piso.data_r [818] = \piso.data_r_818_sv2v_reg ;
  assign \piso.data_r [817] = \piso.data_r_817_sv2v_reg ;
  assign \piso.data_r [816] = \piso.data_r_816_sv2v_reg ;
  assign \piso.data_r [815] = \piso.data_r_815_sv2v_reg ;
  assign \piso.data_r [814] = \piso.data_r_814_sv2v_reg ;
  assign \piso.data_r [813] = \piso.data_r_813_sv2v_reg ;
  assign \piso.data_r [812] = \piso.data_r_812_sv2v_reg ;
  assign \piso.data_r [811] = \piso.data_r_811_sv2v_reg ;
  assign \piso.data_r [810] = \piso.data_r_810_sv2v_reg ;
  assign \piso.data_r [809] = \piso.data_r_809_sv2v_reg ;
  assign \piso.data_r [808] = \piso.data_r_808_sv2v_reg ;
  assign \piso.data_r [807] = \piso.data_r_807_sv2v_reg ;
  assign \piso.data_r [806] = \piso.data_r_806_sv2v_reg ;
  assign \piso.data_r [805] = \piso.data_r_805_sv2v_reg ;
  assign \piso.data_r [804] = \piso.data_r_804_sv2v_reg ;
  assign \piso.data_r [803] = \piso.data_r_803_sv2v_reg ;
  assign \piso.data_r [802] = \piso.data_r_802_sv2v_reg ;
  assign \piso.data_r [801] = \piso.data_r_801_sv2v_reg ;
  assign \piso.data_r [800] = \piso.data_r_800_sv2v_reg ;
  assign \piso.data_r [799] = \piso.data_r_799_sv2v_reg ;
  assign \piso.data_r [798] = \piso.data_r_798_sv2v_reg ;
  assign \piso.data_r [797] = \piso.data_r_797_sv2v_reg ;
  assign \piso.data_r [796] = \piso.data_r_796_sv2v_reg ;
  assign \piso.data_r [795] = \piso.data_r_795_sv2v_reg ;
  assign \piso.data_r [794] = \piso.data_r_794_sv2v_reg ;
  assign \piso.data_r [793] = \piso.data_r_793_sv2v_reg ;
  assign \piso.data_r [792] = \piso.data_r_792_sv2v_reg ;
  assign \piso.data_r [791] = \piso.data_r_791_sv2v_reg ;
  assign \piso.data_r [790] = \piso.data_r_790_sv2v_reg ;
  assign \piso.data_r [789] = \piso.data_r_789_sv2v_reg ;
  assign \piso.data_r [788] = \piso.data_r_788_sv2v_reg ;
  assign \piso.data_r [787] = \piso.data_r_787_sv2v_reg ;
  assign \piso.data_r [786] = \piso.data_r_786_sv2v_reg ;
  assign \piso.data_r [785] = \piso.data_r_785_sv2v_reg ;
  assign \piso.data_r [784] = \piso.data_r_784_sv2v_reg ;
  assign \piso.data_r [783] = \piso.data_r_783_sv2v_reg ;
  assign \piso.data_r [782] = \piso.data_r_782_sv2v_reg ;
  assign \piso.data_r [781] = \piso.data_r_781_sv2v_reg ;
  assign \piso.data_r [780] = \piso.data_r_780_sv2v_reg ;
  assign \piso.data_r [779] = \piso.data_r_779_sv2v_reg ;
  assign \piso.data_r [778] = \piso.data_r_778_sv2v_reg ;
  assign \piso.data_r [777] = \piso.data_r_777_sv2v_reg ;
  assign \piso.data_r [776] = \piso.data_r_776_sv2v_reg ;
  assign \piso.data_r [775] = \piso.data_r_775_sv2v_reg ;
  assign \piso.data_r [774] = \piso.data_r_774_sv2v_reg ;
  assign \piso.data_r [773] = \piso.data_r_773_sv2v_reg ;
  assign \piso.data_r [772] = \piso.data_r_772_sv2v_reg ;
  assign \piso.data_r [771] = \piso.data_r_771_sv2v_reg ;
  assign \piso.data_r [770] = \piso.data_r_770_sv2v_reg ;
  assign \piso.data_r [769] = \piso.data_r_769_sv2v_reg ;
  assign \piso.data_r [768] = \piso.data_r_768_sv2v_reg ;
  assign \piso.data_r [767] = \piso.data_r_767_sv2v_reg ;
  assign \piso.data_r [766] = \piso.data_r_766_sv2v_reg ;
  assign \piso.data_r [765] = \piso.data_r_765_sv2v_reg ;
  assign \piso.data_r [764] = \piso.data_r_764_sv2v_reg ;
  assign \piso.data_r [763] = \piso.data_r_763_sv2v_reg ;
  assign \piso.data_r [762] = \piso.data_r_762_sv2v_reg ;
  assign \piso.data_r [761] = \piso.data_r_761_sv2v_reg ;
  assign \piso.data_r [760] = \piso.data_r_760_sv2v_reg ;
  assign \piso.data_r [759] = \piso.data_r_759_sv2v_reg ;
  assign \piso.data_r [758] = \piso.data_r_758_sv2v_reg ;
  assign \piso.data_r [757] = \piso.data_r_757_sv2v_reg ;
  assign \piso.data_r [756] = \piso.data_r_756_sv2v_reg ;
  assign \piso.data_r [755] = \piso.data_r_755_sv2v_reg ;
  assign \piso.data_r [754] = \piso.data_r_754_sv2v_reg ;
  assign \piso.data_r [753] = \piso.data_r_753_sv2v_reg ;
  assign \piso.data_r [752] = \piso.data_r_752_sv2v_reg ;
  assign \piso.data_r [751] = \piso.data_r_751_sv2v_reg ;
  assign \piso.data_r [750] = \piso.data_r_750_sv2v_reg ;
  assign \piso.data_r [749] = \piso.data_r_749_sv2v_reg ;
  assign \piso.data_r [748] = \piso.data_r_748_sv2v_reg ;
  assign \piso.data_r [747] = \piso.data_r_747_sv2v_reg ;
  assign \piso.data_r [746] = \piso.data_r_746_sv2v_reg ;
  assign \piso.data_r [745] = \piso.data_r_745_sv2v_reg ;
  assign \piso.data_r [744] = \piso.data_r_744_sv2v_reg ;
  assign \piso.data_r [743] = \piso.data_r_743_sv2v_reg ;
  assign \piso.data_r [742] = \piso.data_r_742_sv2v_reg ;
  assign \piso.data_r [741] = \piso.data_r_741_sv2v_reg ;
  assign \piso.data_r [740] = \piso.data_r_740_sv2v_reg ;
  assign \piso.data_r [739] = \piso.data_r_739_sv2v_reg ;
  assign \piso.data_r [738] = \piso.data_r_738_sv2v_reg ;
  assign \piso.data_r [737] = \piso.data_r_737_sv2v_reg ;
  assign \piso.data_r [736] = \piso.data_r_736_sv2v_reg ;
  assign \piso.data_r [735] = \piso.data_r_735_sv2v_reg ;
  assign \piso.data_r [734] = \piso.data_r_734_sv2v_reg ;
  assign \piso.data_r [733] = \piso.data_r_733_sv2v_reg ;
  assign \piso.data_r [732] = \piso.data_r_732_sv2v_reg ;
  assign \piso.data_r [731] = \piso.data_r_731_sv2v_reg ;
  assign \piso.data_r [730] = \piso.data_r_730_sv2v_reg ;
  assign \piso.data_r [729] = \piso.data_r_729_sv2v_reg ;
  assign \piso.data_r [728] = \piso.data_r_728_sv2v_reg ;
  assign \piso.data_r [727] = \piso.data_r_727_sv2v_reg ;
  assign \piso.data_r [726] = \piso.data_r_726_sv2v_reg ;
  assign \piso.data_r [725] = \piso.data_r_725_sv2v_reg ;
  assign \piso.data_r [724] = \piso.data_r_724_sv2v_reg ;
  assign \piso.data_r [723] = \piso.data_r_723_sv2v_reg ;
  assign \piso.data_r [722] = \piso.data_r_722_sv2v_reg ;
  assign \piso.data_r [721] = \piso.data_r_721_sv2v_reg ;
  assign \piso.data_r [720] = \piso.data_r_720_sv2v_reg ;
  assign \piso.data_r [719] = \piso.data_r_719_sv2v_reg ;
  assign \piso.data_r [718] = \piso.data_r_718_sv2v_reg ;
  assign \piso.data_r [717] = \piso.data_r_717_sv2v_reg ;
  assign \piso.data_r [716] = \piso.data_r_716_sv2v_reg ;
  assign \piso.data_r [715] = \piso.data_r_715_sv2v_reg ;
  assign \piso.data_r [714] = \piso.data_r_714_sv2v_reg ;
  assign \piso.data_r [713] = \piso.data_r_713_sv2v_reg ;
  assign \piso.data_r [712] = \piso.data_r_712_sv2v_reg ;
  assign \piso.data_r [711] = \piso.data_r_711_sv2v_reg ;
  assign \piso.data_r [710] = \piso.data_r_710_sv2v_reg ;
  assign \piso.data_r [709] = \piso.data_r_709_sv2v_reg ;
  assign \piso.data_r [708] = \piso.data_r_708_sv2v_reg ;
  assign \piso.data_r [707] = \piso.data_r_707_sv2v_reg ;
  assign \piso.data_r [706] = \piso.data_r_706_sv2v_reg ;
  assign \piso.data_r [705] = \piso.data_r_705_sv2v_reg ;
  assign \piso.data_r [704] = \piso.data_r_704_sv2v_reg ;
  assign \piso.data_r [703] = \piso.data_r_703_sv2v_reg ;
  assign \piso.data_r [702] = \piso.data_r_702_sv2v_reg ;
  assign \piso.data_r [701] = \piso.data_r_701_sv2v_reg ;
  assign \piso.data_r [700] = \piso.data_r_700_sv2v_reg ;
  assign \piso.data_r [699] = \piso.data_r_699_sv2v_reg ;
  assign \piso.data_r [698] = \piso.data_r_698_sv2v_reg ;
  assign \piso.data_r [697] = \piso.data_r_697_sv2v_reg ;
  assign \piso.data_r [696] = \piso.data_r_696_sv2v_reg ;
  assign \piso.data_r [695] = \piso.data_r_695_sv2v_reg ;
  assign \piso.data_r [694] = \piso.data_r_694_sv2v_reg ;
  assign \piso.data_r [693] = \piso.data_r_693_sv2v_reg ;
  assign \piso.data_r [692] = \piso.data_r_692_sv2v_reg ;
  assign \piso.data_r [691] = \piso.data_r_691_sv2v_reg ;
  assign \piso.data_r [690] = \piso.data_r_690_sv2v_reg ;
  assign \piso.data_r [689] = \piso.data_r_689_sv2v_reg ;
  assign \piso.data_r [688] = \piso.data_r_688_sv2v_reg ;
  assign \piso.data_r [687] = \piso.data_r_687_sv2v_reg ;
  assign \piso.data_r [686] = \piso.data_r_686_sv2v_reg ;
  assign \piso.data_r [685] = \piso.data_r_685_sv2v_reg ;
  assign \piso.data_r [684] = \piso.data_r_684_sv2v_reg ;
  assign \piso.data_r [683] = \piso.data_r_683_sv2v_reg ;
  assign \piso.data_r [682] = \piso.data_r_682_sv2v_reg ;
  assign \piso.data_r [681] = \piso.data_r_681_sv2v_reg ;
  assign \piso.data_r [680] = \piso.data_r_680_sv2v_reg ;
  assign \piso.data_r [679] = \piso.data_r_679_sv2v_reg ;
  assign \piso.data_r [678] = \piso.data_r_678_sv2v_reg ;
  assign \piso.data_r [677] = \piso.data_r_677_sv2v_reg ;
  assign \piso.data_r [676] = \piso.data_r_676_sv2v_reg ;
  assign \piso.data_r [675] = \piso.data_r_675_sv2v_reg ;
  assign \piso.data_r [674] = \piso.data_r_674_sv2v_reg ;
  assign \piso.data_r [673] = \piso.data_r_673_sv2v_reg ;
  assign \piso.data_r [672] = \piso.data_r_672_sv2v_reg ;
  assign \piso.data_r [671] = \piso.data_r_671_sv2v_reg ;
  assign \piso.data_r [670] = \piso.data_r_670_sv2v_reg ;
  assign \piso.data_r [669] = \piso.data_r_669_sv2v_reg ;
  assign \piso.data_r [668] = \piso.data_r_668_sv2v_reg ;
  assign \piso.data_r [667] = \piso.data_r_667_sv2v_reg ;
  assign \piso.data_r [666] = \piso.data_r_666_sv2v_reg ;
  assign \piso.data_r [665] = \piso.data_r_665_sv2v_reg ;
  assign \piso.data_r [664] = \piso.data_r_664_sv2v_reg ;
  assign \piso.data_r [663] = \piso.data_r_663_sv2v_reg ;
  assign \piso.data_r [662] = \piso.data_r_662_sv2v_reg ;
  assign \piso.data_r [661] = \piso.data_r_661_sv2v_reg ;
  assign \piso.data_r [660] = \piso.data_r_660_sv2v_reg ;
  assign \piso.data_r [659] = \piso.data_r_659_sv2v_reg ;
  assign \piso.data_r [658] = \piso.data_r_658_sv2v_reg ;
  assign \piso.data_r [657] = \piso.data_r_657_sv2v_reg ;
  assign \piso.data_r [656] = \piso.data_r_656_sv2v_reg ;
  assign \piso.data_r [655] = \piso.data_r_655_sv2v_reg ;
  assign \piso.data_r [654] = \piso.data_r_654_sv2v_reg ;
  assign \piso.data_r [653] = \piso.data_r_653_sv2v_reg ;
  assign \piso.data_r [652] = \piso.data_r_652_sv2v_reg ;
  assign \piso.data_r [651] = \piso.data_r_651_sv2v_reg ;
  assign \piso.data_r [650] = \piso.data_r_650_sv2v_reg ;
  assign \piso.data_r [649] = \piso.data_r_649_sv2v_reg ;
  assign \piso.data_r [648] = \piso.data_r_648_sv2v_reg ;
  assign \piso.data_r [647] = \piso.data_r_647_sv2v_reg ;
  assign \piso.data_r [646] = \piso.data_r_646_sv2v_reg ;
  assign \piso.data_r [645] = \piso.data_r_645_sv2v_reg ;
  assign \piso.data_r [644] = \piso.data_r_644_sv2v_reg ;
  assign \piso.data_r [643] = \piso.data_r_643_sv2v_reg ;
  assign \piso.data_r [642] = \piso.data_r_642_sv2v_reg ;
  assign \piso.data_r [641] = \piso.data_r_641_sv2v_reg ;
  assign \piso.data_r [640] = \piso.data_r_640_sv2v_reg ;
  assign \piso.data_r [639] = \piso.data_r_639_sv2v_reg ;
  assign \piso.data_r [638] = \piso.data_r_638_sv2v_reg ;
  assign \piso.data_r [637] = \piso.data_r_637_sv2v_reg ;
  assign \piso.data_r [636] = \piso.data_r_636_sv2v_reg ;
  assign \piso.data_r [635] = \piso.data_r_635_sv2v_reg ;
  assign \piso.data_r [634] = \piso.data_r_634_sv2v_reg ;
  assign \piso.data_r [633] = \piso.data_r_633_sv2v_reg ;
  assign \piso.data_r [632] = \piso.data_r_632_sv2v_reg ;
  assign \piso.data_r [631] = \piso.data_r_631_sv2v_reg ;
  assign \piso.data_r [630] = \piso.data_r_630_sv2v_reg ;
  assign \piso.data_r [629] = \piso.data_r_629_sv2v_reg ;
  assign \piso.data_r [628] = \piso.data_r_628_sv2v_reg ;
  assign \piso.data_r [627] = \piso.data_r_627_sv2v_reg ;
  assign \piso.data_r [626] = \piso.data_r_626_sv2v_reg ;
  assign \piso.data_r [625] = \piso.data_r_625_sv2v_reg ;
  assign \piso.data_r [624] = \piso.data_r_624_sv2v_reg ;
  assign \piso.data_r [623] = \piso.data_r_623_sv2v_reg ;
  assign \piso.data_r [622] = \piso.data_r_622_sv2v_reg ;
  assign \piso.data_r [621] = \piso.data_r_621_sv2v_reg ;
  assign \piso.data_r [620] = \piso.data_r_620_sv2v_reg ;
  assign \piso.data_r [619] = \piso.data_r_619_sv2v_reg ;
  assign \piso.data_r [618] = \piso.data_r_618_sv2v_reg ;
  assign \piso.data_r [617] = \piso.data_r_617_sv2v_reg ;
  assign \piso.data_r [616] = \piso.data_r_616_sv2v_reg ;
  assign \piso.data_r [615] = \piso.data_r_615_sv2v_reg ;
  assign \piso.data_r [614] = \piso.data_r_614_sv2v_reg ;
  assign \piso.data_r [613] = \piso.data_r_613_sv2v_reg ;
  assign \piso.data_r [612] = \piso.data_r_612_sv2v_reg ;
  assign \piso.data_r [611] = \piso.data_r_611_sv2v_reg ;
  assign \piso.data_r [610] = \piso.data_r_610_sv2v_reg ;
  assign \piso.data_r [609] = \piso.data_r_609_sv2v_reg ;
  assign \piso.data_r [608] = \piso.data_r_608_sv2v_reg ;
  assign \piso.data_r [607] = \piso.data_r_607_sv2v_reg ;
  assign \piso.data_r [606] = \piso.data_r_606_sv2v_reg ;
  assign \piso.data_r [605] = \piso.data_r_605_sv2v_reg ;
  assign \piso.data_r [604] = \piso.data_r_604_sv2v_reg ;
  assign \piso.data_r [603] = \piso.data_r_603_sv2v_reg ;
  assign \piso.data_r [602] = \piso.data_r_602_sv2v_reg ;
  assign \piso.data_r [601] = \piso.data_r_601_sv2v_reg ;
  assign \piso.data_r [600] = \piso.data_r_600_sv2v_reg ;
  assign \piso.data_r [599] = \piso.data_r_599_sv2v_reg ;
  assign \piso.data_r [598] = \piso.data_r_598_sv2v_reg ;
  assign \piso.data_r [597] = \piso.data_r_597_sv2v_reg ;
  assign \piso.data_r [596] = \piso.data_r_596_sv2v_reg ;
  assign \piso.data_r [595] = \piso.data_r_595_sv2v_reg ;
  assign \piso.data_r [594] = \piso.data_r_594_sv2v_reg ;
  assign \piso.data_r [593] = \piso.data_r_593_sv2v_reg ;
  assign \piso.data_r [592] = \piso.data_r_592_sv2v_reg ;
  assign \piso.data_r [591] = \piso.data_r_591_sv2v_reg ;
  assign \piso.data_r [590] = \piso.data_r_590_sv2v_reg ;
  assign \piso.data_r [589] = \piso.data_r_589_sv2v_reg ;
  assign \piso.data_r [588] = \piso.data_r_588_sv2v_reg ;
  assign \piso.data_r [587] = \piso.data_r_587_sv2v_reg ;
  assign \piso.data_r [586] = \piso.data_r_586_sv2v_reg ;
  assign \piso.data_r [585] = \piso.data_r_585_sv2v_reg ;
  assign \piso.data_r [584] = \piso.data_r_584_sv2v_reg ;
  assign \piso.data_r [583] = \piso.data_r_583_sv2v_reg ;
  assign \piso.data_r [582] = \piso.data_r_582_sv2v_reg ;
  assign \piso.data_r [581] = \piso.data_r_581_sv2v_reg ;
  assign \piso.data_r [580] = \piso.data_r_580_sv2v_reg ;
  assign \piso.data_r [579] = \piso.data_r_579_sv2v_reg ;
  assign \piso.data_r [578] = \piso.data_r_578_sv2v_reg ;
  assign \piso.data_r [577] = \piso.data_r_577_sv2v_reg ;
  assign \piso.data_r [576] = \piso.data_r_576_sv2v_reg ;
  assign \piso.data_r [575] = \piso.data_r_575_sv2v_reg ;
  assign \piso.data_r [574] = \piso.data_r_574_sv2v_reg ;
  assign \piso.data_r [573] = \piso.data_r_573_sv2v_reg ;
  assign \piso.data_r [572] = \piso.data_r_572_sv2v_reg ;
  assign \piso.data_r [571] = \piso.data_r_571_sv2v_reg ;
  assign \piso.data_r [570] = \piso.data_r_570_sv2v_reg ;
  assign \piso.data_r [569] = \piso.data_r_569_sv2v_reg ;
  assign \piso.data_r [568] = \piso.data_r_568_sv2v_reg ;
  assign \piso.data_r [567] = \piso.data_r_567_sv2v_reg ;
  assign \piso.data_r [566] = \piso.data_r_566_sv2v_reg ;
  assign \piso.data_r [565] = \piso.data_r_565_sv2v_reg ;
  assign \piso.data_r [564] = \piso.data_r_564_sv2v_reg ;
  assign \piso.data_r [563] = \piso.data_r_563_sv2v_reg ;
  assign \piso.data_r [562] = \piso.data_r_562_sv2v_reg ;
  assign \piso.data_r [561] = \piso.data_r_561_sv2v_reg ;
  assign \piso.data_r [560] = \piso.data_r_560_sv2v_reg ;
  assign \piso.data_r [559] = \piso.data_r_559_sv2v_reg ;
  assign \piso.data_r [558] = \piso.data_r_558_sv2v_reg ;
  assign \piso.data_r [557] = \piso.data_r_557_sv2v_reg ;
  assign \piso.data_r [556] = \piso.data_r_556_sv2v_reg ;
  assign \piso.data_r [555] = \piso.data_r_555_sv2v_reg ;
  assign \piso.data_r [554] = \piso.data_r_554_sv2v_reg ;
  assign \piso.data_r [553] = \piso.data_r_553_sv2v_reg ;
  assign \piso.data_r [552] = \piso.data_r_552_sv2v_reg ;
  assign \piso.data_r [551] = \piso.data_r_551_sv2v_reg ;
  assign \piso.data_r [550] = \piso.data_r_550_sv2v_reg ;
  assign \piso.data_r [549] = \piso.data_r_549_sv2v_reg ;
  assign \piso.data_r [548] = \piso.data_r_548_sv2v_reg ;
  assign \piso.data_r [547] = \piso.data_r_547_sv2v_reg ;
  assign \piso.data_r [546] = \piso.data_r_546_sv2v_reg ;
  assign \piso.data_r [545] = \piso.data_r_545_sv2v_reg ;
  assign \piso.data_r [544] = \piso.data_r_544_sv2v_reg ;
  assign \piso.data_r [543] = \piso.data_r_543_sv2v_reg ;
  assign \piso.data_r [542] = \piso.data_r_542_sv2v_reg ;
  assign \piso.data_r [541] = \piso.data_r_541_sv2v_reg ;
  assign \piso.data_r [540] = \piso.data_r_540_sv2v_reg ;
  assign \piso.data_r [539] = \piso.data_r_539_sv2v_reg ;
  assign \piso.data_r [538] = \piso.data_r_538_sv2v_reg ;
  assign \piso.data_r [537] = \piso.data_r_537_sv2v_reg ;
  assign \piso.data_r [536] = \piso.data_r_536_sv2v_reg ;
  assign \piso.data_r [535] = \piso.data_r_535_sv2v_reg ;
  assign \piso.data_r [534] = \piso.data_r_534_sv2v_reg ;
  assign \piso.data_r [533] = \piso.data_r_533_sv2v_reg ;
  assign \piso.data_r [532] = \piso.data_r_532_sv2v_reg ;
  assign \piso.data_r [531] = \piso.data_r_531_sv2v_reg ;
  assign \piso.data_r [530] = \piso.data_r_530_sv2v_reg ;
  assign \piso.data_r [529] = \piso.data_r_529_sv2v_reg ;
  assign \piso.data_r [528] = \piso.data_r_528_sv2v_reg ;
  assign \piso.data_r [527] = \piso.data_r_527_sv2v_reg ;
  assign \piso.data_r [526] = \piso.data_r_526_sv2v_reg ;
  assign \piso.data_r [525] = \piso.data_r_525_sv2v_reg ;
  assign \piso.data_r [524] = \piso.data_r_524_sv2v_reg ;
  assign \piso.data_r [523] = \piso.data_r_523_sv2v_reg ;
  assign \piso.data_r [522] = \piso.data_r_522_sv2v_reg ;
  assign \piso.data_r [521] = \piso.data_r_521_sv2v_reg ;
  assign \piso.data_r [520] = \piso.data_r_520_sv2v_reg ;
  assign \piso.data_r [519] = \piso.data_r_519_sv2v_reg ;
  assign \piso.data_r [518] = \piso.data_r_518_sv2v_reg ;
  assign \piso.data_r [517] = \piso.data_r_517_sv2v_reg ;
  assign \piso.data_r [516] = \piso.data_r_516_sv2v_reg ;
  assign \piso.data_r [515] = \piso.data_r_515_sv2v_reg ;
  assign \piso.data_r [514] = \piso.data_r_514_sv2v_reg ;
  assign \piso.data_r [513] = \piso.data_r_513_sv2v_reg ;
  assign \piso.data_r [512] = \piso.data_r_512_sv2v_reg ;
  assign \piso.data_r [511] = \piso.data_r_511_sv2v_reg ;
  assign \piso.data_r [510] = \piso.data_r_510_sv2v_reg ;
  assign \piso.data_r [509] = \piso.data_r_509_sv2v_reg ;
  assign \piso.data_r [508] = \piso.data_r_508_sv2v_reg ;
  assign \piso.data_r [507] = \piso.data_r_507_sv2v_reg ;
  assign \piso.data_r [506] = \piso.data_r_506_sv2v_reg ;
  assign \piso.data_r [505] = \piso.data_r_505_sv2v_reg ;
  assign \piso.data_r [504] = \piso.data_r_504_sv2v_reg ;
  assign \piso.data_r [503] = \piso.data_r_503_sv2v_reg ;
  assign \piso.data_r [502] = \piso.data_r_502_sv2v_reg ;
  assign \piso.data_r [501] = \piso.data_r_501_sv2v_reg ;
  assign \piso.data_r [500] = \piso.data_r_500_sv2v_reg ;
  assign \piso.data_r [499] = \piso.data_r_499_sv2v_reg ;
  assign \piso.data_r [498] = \piso.data_r_498_sv2v_reg ;
  assign \piso.data_r [497] = \piso.data_r_497_sv2v_reg ;
  assign \piso.data_r [496] = \piso.data_r_496_sv2v_reg ;
  assign \piso.data_r [495] = \piso.data_r_495_sv2v_reg ;
  assign \piso.data_r [494] = \piso.data_r_494_sv2v_reg ;
  assign \piso.data_r [493] = \piso.data_r_493_sv2v_reg ;
  assign \piso.data_r [492] = \piso.data_r_492_sv2v_reg ;
  assign \piso.data_r [491] = \piso.data_r_491_sv2v_reg ;
  assign \piso.data_r [490] = \piso.data_r_490_sv2v_reg ;
  assign \piso.data_r [489] = \piso.data_r_489_sv2v_reg ;
  assign \piso.data_r [488] = \piso.data_r_488_sv2v_reg ;
  assign \piso.data_r [487] = \piso.data_r_487_sv2v_reg ;
  assign \piso.data_r [486] = \piso.data_r_486_sv2v_reg ;
  assign \piso.data_r [485] = \piso.data_r_485_sv2v_reg ;
  assign \piso.data_r [484] = \piso.data_r_484_sv2v_reg ;
  assign \piso.data_r [483] = \piso.data_r_483_sv2v_reg ;
  assign \piso.data_r [482] = \piso.data_r_482_sv2v_reg ;
  assign \piso.data_r [481] = \piso.data_r_481_sv2v_reg ;
  assign \piso.data_r [480] = \piso.data_r_480_sv2v_reg ;
  assign \piso.data_r [479] = \piso.data_r_479_sv2v_reg ;
  assign \piso.data_r [478] = \piso.data_r_478_sv2v_reg ;
  assign \piso.data_r [477] = \piso.data_r_477_sv2v_reg ;
  assign \piso.data_r [476] = \piso.data_r_476_sv2v_reg ;
  assign \piso.data_r [475] = \piso.data_r_475_sv2v_reg ;
  assign \piso.data_r [474] = \piso.data_r_474_sv2v_reg ;
  assign \piso.data_r [473] = \piso.data_r_473_sv2v_reg ;
  assign \piso.data_r [472] = \piso.data_r_472_sv2v_reg ;
  assign \piso.data_r [471] = \piso.data_r_471_sv2v_reg ;
  assign \piso.data_r [470] = \piso.data_r_470_sv2v_reg ;
  assign \piso.data_r [469] = \piso.data_r_469_sv2v_reg ;
  assign \piso.data_r [468] = \piso.data_r_468_sv2v_reg ;
  assign \piso.data_r [467] = \piso.data_r_467_sv2v_reg ;
  assign \piso.data_r [466] = \piso.data_r_466_sv2v_reg ;
  assign \piso.data_r [465] = \piso.data_r_465_sv2v_reg ;
  assign \piso.data_r [464] = \piso.data_r_464_sv2v_reg ;
  assign \piso.data_r [463] = \piso.data_r_463_sv2v_reg ;
  assign \piso.data_r [462] = \piso.data_r_462_sv2v_reg ;
  assign \piso.data_r [461] = \piso.data_r_461_sv2v_reg ;
  assign \piso.data_r [460] = \piso.data_r_460_sv2v_reg ;
  assign \piso.data_r [459] = \piso.data_r_459_sv2v_reg ;
  assign \piso.data_r [458] = \piso.data_r_458_sv2v_reg ;
  assign \piso.data_r [457] = \piso.data_r_457_sv2v_reg ;
  assign \piso.data_r [456] = \piso.data_r_456_sv2v_reg ;
  assign \piso.data_r [455] = \piso.data_r_455_sv2v_reg ;
  assign \piso.data_r [454] = \piso.data_r_454_sv2v_reg ;
  assign \piso.data_r [453] = \piso.data_r_453_sv2v_reg ;
  assign \piso.data_r [452] = \piso.data_r_452_sv2v_reg ;
  assign \piso.data_r [451] = \piso.data_r_451_sv2v_reg ;
  assign \piso.data_r [450] = \piso.data_r_450_sv2v_reg ;
  assign \piso.data_r [449] = \piso.data_r_449_sv2v_reg ;
  assign \piso.data_r [448] = \piso.data_r_448_sv2v_reg ;
  assign \piso.data_r [447] = \piso.data_r_447_sv2v_reg ;
  assign \piso.data_r [446] = \piso.data_r_446_sv2v_reg ;
  assign \piso.data_r [445] = \piso.data_r_445_sv2v_reg ;
  assign \piso.data_r [444] = \piso.data_r_444_sv2v_reg ;
  assign \piso.data_r [443] = \piso.data_r_443_sv2v_reg ;
  assign \piso.data_r [442] = \piso.data_r_442_sv2v_reg ;
  assign \piso.data_r [441] = \piso.data_r_441_sv2v_reg ;
  assign \piso.data_r [440] = \piso.data_r_440_sv2v_reg ;
  assign \piso.data_r [439] = \piso.data_r_439_sv2v_reg ;
  assign \piso.data_r [438] = \piso.data_r_438_sv2v_reg ;
  assign \piso.data_r [437] = \piso.data_r_437_sv2v_reg ;
  assign \piso.data_r [436] = \piso.data_r_436_sv2v_reg ;
  assign \piso.data_r [435] = \piso.data_r_435_sv2v_reg ;
  assign \piso.data_r [434] = \piso.data_r_434_sv2v_reg ;
  assign \piso.data_r [433] = \piso.data_r_433_sv2v_reg ;
  assign \piso.data_r [432] = \piso.data_r_432_sv2v_reg ;
  assign \piso.data_r [431] = \piso.data_r_431_sv2v_reg ;
  assign \piso.data_r [430] = \piso.data_r_430_sv2v_reg ;
  assign \piso.data_r [429] = \piso.data_r_429_sv2v_reg ;
  assign \piso.data_r [428] = \piso.data_r_428_sv2v_reg ;
  assign \piso.data_r [427] = \piso.data_r_427_sv2v_reg ;
  assign \piso.data_r [426] = \piso.data_r_426_sv2v_reg ;
  assign \piso.data_r [425] = \piso.data_r_425_sv2v_reg ;
  assign \piso.data_r [424] = \piso.data_r_424_sv2v_reg ;
  assign \piso.data_r [423] = \piso.data_r_423_sv2v_reg ;
  assign \piso.data_r [422] = \piso.data_r_422_sv2v_reg ;
  assign \piso.data_r [421] = \piso.data_r_421_sv2v_reg ;
  assign \piso.data_r [420] = \piso.data_r_420_sv2v_reg ;
  assign \piso.data_r [419] = \piso.data_r_419_sv2v_reg ;
  assign \piso.data_r [418] = \piso.data_r_418_sv2v_reg ;
  assign \piso.data_r [417] = \piso.data_r_417_sv2v_reg ;
  assign \piso.data_r [416] = \piso.data_r_416_sv2v_reg ;
  assign \piso.data_r [415] = \piso.data_r_415_sv2v_reg ;
  assign \piso.data_r [414] = \piso.data_r_414_sv2v_reg ;
  assign \piso.data_r [413] = \piso.data_r_413_sv2v_reg ;
  assign \piso.data_r [412] = \piso.data_r_412_sv2v_reg ;
  assign \piso.data_r [411] = \piso.data_r_411_sv2v_reg ;
  assign \piso.data_r [410] = \piso.data_r_410_sv2v_reg ;
  assign \piso.data_r [409] = \piso.data_r_409_sv2v_reg ;
  assign \piso.data_r [408] = \piso.data_r_408_sv2v_reg ;
  assign \piso.data_r [407] = \piso.data_r_407_sv2v_reg ;
  assign \piso.data_r [406] = \piso.data_r_406_sv2v_reg ;
  assign \piso.data_r [405] = \piso.data_r_405_sv2v_reg ;
  assign \piso.data_r [404] = \piso.data_r_404_sv2v_reg ;
  assign \piso.data_r [403] = \piso.data_r_403_sv2v_reg ;
  assign \piso.data_r [402] = \piso.data_r_402_sv2v_reg ;
  assign \piso.data_r [401] = \piso.data_r_401_sv2v_reg ;
  assign \piso.data_r [400] = \piso.data_r_400_sv2v_reg ;
  assign \piso.data_r [399] = \piso.data_r_399_sv2v_reg ;
  assign \piso.data_r [398] = \piso.data_r_398_sv2v_reg ;
  assign \piso.data_r [397] = \piso.data_r_397_sv2v_reg ;
  assign \piso.data_r [396] = \piso.data_r_396_sv2v_reg ;
  assign \piso.data_r [395] = \piso.data_r_395_sv2v_reg ;
  assign \piso.data_r [394] = \piso.data_r_394_sv2v_reg ;
  assign \piso.data_r [393] = \piso.data_r_393_sv2v_reg ;
  assign \piso.data_r [392] = \piso.data_r_392_sv2v_reg ;
  assign \piso.data_r [391] = \piso.data_r_391_sv2v_reg ;
  assign \piso.data_r [390] = \piso.data_r_390_sv2v_reg ;
  assign \piso.data_r [389] = \piso.data_r_389_sv2v_reg ;
  assign \piso.data_r [388] = \piso.data_r_388_sv2v_reg ;
  assign \piso.data_r [387] = \piso.data_r_387_sv2v_reg ;
  assign \piso.data_r [386] = \piso.data_r_386_sv2v_reg ;
  assign \piso.data_r [385] = \piso.data_r_385_sv2v_reg ;
  assign \piso.data_r [384] = \piso.data_r_384_sv2v_reg ;
  assign \piso.data_r [383] = \piso.data_r_383_sv2v_reg ;
  assign \piso.data_r [382] = \piso.data_r_382_sv2v_reg ;
  assign \piso.data_r [381] = \piso.data_r_381_sv2v_reg ;
  assign \piso.data_r [380] = \piso.data_r_380_sv2v_reg ;
  assign \piso.data_r [379] = \piso.data_r_379_sv2v_reg ;
  assign \piso.data_r [378] = \piso.data_r_378_sv2v_reg ;
  assign \piso.data_r [377] = \piso.data_r_377_sv2v_reg ;
  assign \piso.data_r [376] = \piso.data_r_376_sv2v_reg ;
  assign \piso.data_r [375] = \piso.data_r_375_sv2v_reg ;
  assign \piso.data_r [374] = \piso.data_r_374_sv2v_reg ;
  assign \piso.data_r [373] = \piso.data_r_373_sv2v_reg ;
  assign \piso.data_r [372] = \piso.data_r_372_sv2v_reg ;
  assign \piso.data_r [371] = \piso.data_r_371_sv2v_reg ;
  assign \piso.data_r [370] = \piso.data_r_370_sv2v_reg ;
  assign \piso.data_r [369] = \piso.data_r_369_sv2v_reg ;
  assign \piso.data_r [368] = \piso.data_r_368_sv2v_reg ;
  assign \piso.data_r [367] = \piso.data_r_367_sv2v_reg ;
  assign \piso.data_r [366] = \piso.data_r_366_sv2v_reg ;
  assign \piso.data_r [365] = \piso.data_r_365_sv2v_reg ;
  assign \piso.data_r [364] = \piso.data_r_364_sv2v_reg ;
  assign \piso.data_r [363] = \piso.data_r_363_sv2v_reg ;
  assign \piso.data_r [362] = \piso.data_r_362_sv2v_reg ;
  assign \piso.data_r [361] = \piso.data_r_361_sv2v_reg ;
  assign \piso.data_r [360] = \piso.data_r_360_sv2v_reg ;
  assign \piso.data_r [359] = \piso.data_r_359_sv2v_reg ;
  assign \piso.data_r [358] = \piso.data_r_358_sv2v_reg ;
  assign \piso.data_r [357] = \piso.data_r_357_sv2v_reg ;
  assign \piso.data_r [356] = \piso.data_r_356_sv2v_reg ;
  assign \piso.data_r [355] = \piso.data_r_355_sv2v_reg ;
  assign \piso.data_r [354] = \piso.data_r_354_sv2v_reg ;
  assign \piso.data_r [353] = \piso.data_r_353_sv2v_reg ;
  assign \piso.data_r [352] = \piso.data_r_352_sv2v_reg ;
  assign \piso.data_r [351] = \piso.data_r_351_sv2v_reg ;
  assign \piso.data_r [350] = \piso.data_r_350_sv2v_reg ;
  assign \piso.data_r [349] = \piso.data_r_349_sv2v_reg ;
  assign \piso.data_r [348] = \piso.data_r_348_sv2v_reg ;
  assign \piso.data_r [347] = \piso.data_r_347_sv2v_reg ;
  assign \piso.data_r [346] = \piso.data_r_346_sv2v_reg ;
  assign \piso.data_r [345] = \piso.data_r_345_sv2v_reg ;
  assign \piso.data_r [344] = \piso.data_r_344_sv2v_reg ;
  assign \piso.data_r [343] = \piso.data_r_343_sv2v_reg ;
  assign \piso.data_r [342] = \piso.data_r_342_sv2v_reg ;
  assign \piso.data_r [341] = \piso.data_r_341_sv2v_reg ;
  assign \piso.data_r [340] = \piso.data_r_340_sv2v_reg ;
  assign \piso.data_r [339] = \piso.data_r_339_sv2v_reg ;
  assign \piso.data_r [338] = \piso.data_r_338_sv2v_reg ;
  assign \piso.data_r [337] = \piso.data_r_337_sv2v_reg ;
  assign \piso.data_r [336] = \piso.data_r_336_sv2v_reg ;
  assign \piso.data_r [335] = \piso.data_r_335_sv2v_reg ;
  assign \piso.data_r [334] = \piso.data_r_334_sv2v_reg ;
  assign \piso.data_r [333] = \piso.data_r_333_sv2v_reg ;
  assign \piso.data_r [332] = \piso.data_r_332_sv2v_reg ;
  assign \piso.data_r [331] = \piso.data_r_331_sv2v_reg ;
  assign \piso.data_r [330] = \piso.data_r_330_sv2v_reg ;
  assign \piso.data_r [329] = \piso.data_r_329_sv2v_reg ;
  assign \piso.data_r [328] = \piso.data_r_328_sv2v_reg ;
  assign \piso.data_r [327] = \piso.data_r_327_sv2v_reg ;
  assign \piso.data_r [326] = \piso.data_r_326_sv2v_reg ;
  assign \piso.data_r [325] = \piso.data_r_325_sv2v_reg ;
  assign \piso.data_r [324] = \piso.data_r_324_sv2v_reg ;
  assign \piso.data_r [323] = \piso.data_r_323_sv2v_reg ;
  assign \piso.data_r [322] = \piso.data_r_322_sv2v_reg ;
  assign \piso.data_r [321] = \piso.data_r_321_sv2v_reg ;
  assign \piso.data_r [320] = \piso.data_r_320_sv2v_reg ;
  assign \piso.data_r [319] = \piso.data_r_319_sv2v_reg ;
  assign \piso.data_r [318] = \piso.data_r_318_sv2v_reg ;
  assign \piso.data_r [317] = \piso.data_r_317_sv2v_reg ;
  assign \piso.data_r [316] = \piso.data_r_316_sv2v_reg ;
  assign \piso.data_r [315] = \piso.data_r_315_sv2v_reg ;
  assign \piso.data_r [314] = \piso.data_r_314_sv2v_reg ;
  assign \piso.data_r [313] = \piso.data_r_313_sv2v_reg ;
  assign \piso.data_r [312] = \piso.data_r_312_sv2v_reg ;
  assign \piso.data_r [311] = \piso.data_r_311_sv2v_reg ;
  assign \piso.data_r [310] = \piso.data_r_310_sv2v_reg ;
  assign \piso.data_r [309] = \piso.data_r_309_sv2v_reg ;
  assign \piso.data_r [308] = \piso.data_r_308_sv2v_reg ;
  assign \piso.data_r [307] = \piso.data_r_307_sv2v_reg ;
  assign \piso.data_r [306] = \piso.data_r_306_sv2v_reg ;
  assign \piso.data_r [305] = \piso.data_r_305_sv2v_reg ;
  assign \piso.data_r [304] = \piso.data_r_304_sv2v_reg ;
  assign \piso.data_r [303] = \piso.data_r_303_sv2v_reg ;
  assign \piso.data_r [302] = \piso.data_r_302_sv2v_reg ;
  assign \piso.data_r [301] = \piso.data_r_301_sv2v_reg ;
  assign \piso.data_r [300] = \piso.data_r_300_sv2v_reg ;
  assign \piso.data_r [299] = \piso.data_r_299_sv2v_reg ;
  assign \piso.data_r [298] = \piso.data_r_298_sv2v_reg ;
  assign \piso.data_r [297] = \piso.data_r_297_sv2v_reg ;
  assign \piso.data_r [296] = \piso.data_r_296_sv2v_reg ;
  assign \piso.data_r [295] = \piso.data_r_295_sv2v_reg ;
  assign \piso.data_r [294] = \piso.data_r_294_sv2v_reg ;
  assign \piso.data_r [293] = \piso.data_r_293_sv2v_reg ;
  assign \piso.data_r [292] = \piso.data_r_292_sv2v_reg ;
  assign \piso.data_r [291] = \piso.data_r_291_sv2v_reg ;
  assign \piso.data_r [290] = \piso.data_r_290_sv2v_reg ;
  assign \piso.data_r [289] = \piso.data_r_289_sv2v_reg ;
  assign \piso.data_r [288] = \piso.data_r_288_sv2v_reg ;
  assign \piso.data_r [287] = \piso.data_r_287_sv2v_reg ;
  assign \piso.data_r [286] = \piso.data_r_286_sv2v_reg ;
  assign \piso.data_r [285] = \piso.data_r_285_sv2v_reg ;
  assign \piso.data_r [284] = \piso.data_r_284_sv2v_reg ;
  assign \piso.data_r [283] = \piso.data_r_283_sv2v_reg ;
  assign \piso.data_r [282] = \piso.data_r_282_sv2v_reg ;
  assign \piso.data_r [281] = \piso.data_r_281_sv2v_reg ;
  assign \piso.data_r [280] = \piso.data_r_280_sv2v_reg ;
  assign \piso.data_r [279] = \piso.data_r_279_sv2v_reg ;
  assign \piso.data_r [278] = \piso.data_r_278_sv2v_reg ;
  assign \piso.data_r [277] = \piso.data_r_277_sv2v_reg ;
  assign \piso.data_r [276] = \piso.data_r_276_sv2v_reg ;
  assign \piso.data_r [275] = \piso.data_r_275_sv2v_reg ;
  assign \piso.data_r [274] = \piso.data_r_274_sv2v_reg ;
  assign \piso.data_r [273] = \piso.data_r_273_sv2v_reg ;
  assign \piso.data_r [272] = \piso.data_r_272_sv2v_reg ;
  assign \piso.data_r [271] = \piso.data_r_271_sv2v_reg ;
  assign \piso.data_r [270] = \piso.data_r_270_sv2v_reg ;
  assign \piso.data_r [269] = \piso.data_r_269_sv2v_reg ;
  assign \piso.data_r [268] = \piso.data_r_268_sv2v_reg ;
  assign \piso.data_r [267] = \piso.data_r_267_sv2v_reg ;
  assign \piso.data_r [266] = \piso.data_r_266_sv2v_reg ;
  assign \piso.data_r [265] = \piso.data_r_265_sv2v_reg ;
  assign \piso.data_r [264] = \piso.data_r_264_sv2v_reg ;
  assign \piso.data_r [263] = \piso.data_r_263_sv2v_reg ;
  assign \piso.data_r [262] = \piso.data_r_262_sv2v_reg ;
  assign \piso.data_r [261] = \piso.data_r_261_sv2v_reg ;
  assign \piso.data_r [260] = \piso.data_r_260_sv2v_reg ;
  assign \piso.data_r [259] = \piso.data_r_259_sv2v_reg ;
  assign \piso.data_r [258] = \piso.data_r_258_sv2v_reg ;
  assign \piso.data_r [257] = \piso.data_r_257_sv2v_reg ;
  assign \piso.data_r [256] = \piso.data_r_256_sv2v_reg ;
  assign \piso.data_r [255] = \piso.data_r_255_sv2v_reg ;
  assign \piso.data_r [254] = \piso.data_r_254_sv2v_reg ;
  assign \piso.data_r [253] = \piso.data_r_253_sv2v_reg ;
  assign \piso.data_r [252] = \piso.data_r_252_sv2v_reg ;
  assign \piso.data_r [251] = \piso.data_r_251_sv2v_reg ;
  assign \piso.data_r [250] = \piso.data_r_250_sv2v_reg ;
  assign \piso.data_r [249] = \piso.data_r_249_sv2v_reg ;
  assign \piso.data_r [248] = \piso.data_r_248_sv2v_reg ;
  assign \piso.data_r [247] = \piso.data_r_247_sv2v_reg ;
  assign \piso.data_r [246] = \piso.data_r_246_sv2v_reg ;
  assign \piso.data_r [245] = \piso.data_r_245_sv2v_reg ;
  assign \piso.data_r [244] = \piso.data_r_244_sv2v_reg ;
  assign \piso.data_r [243] = \piso.data_r_243_sv2v_reg ;
  assign \piso.data_r [242] = \piso.data_r_242_sv2v_reg ;
  assign \piso.data_r [241] = \piso.data_r_241_sv2v_reg ;
  assign \piso.data_r [240] = \piso.data_r_240_sv2v_reg ;
  assign \piso.data_r [239] = \piso.data_r_239_sv2v_reg ;
  assign \piso.data_r [238] = \piso.data_r_238_sv2v_reg ;
  assign \piso.data_r [237] = \piso.data_r_237_sv2v_reg ;
  assign \piso.data_r [236] = \piso.data_r_236_sv2v_reg ;
  assign \piso.data_r [235] = \piso.data_r_235_sv2v_reg ;
  assign \piso.data_r [234] = \piso.data_r_234_sv2v_reg ;
  assign \piso.data_r [233] = \piso.data_r_233_sv2v_reg ;
  assign \piso.data_r [232] = \piso.data_r_232_sv2v_reg ;
  assign \piso.data_r [231] = \piso.data_r_231_sv2v_reg ;
  assign \piso.data_r [230] = \piso.data_r_230_sv2v_reg ;
  assign \piso.data_r [229] = \piso.data_r_229_sv2v_reg ;
  assign \piso.data_r [228] = \piso.data_r_228_sv2v_reg ;
  assign \piso.data_r [227] = \piso.data_r_227_sv2v_reg ;
  assign \piso.data_r [226] = \piso.data_r_226_sv2v_reg ;
  assign \piso.data_r [225] = \piso.data_r_225_sv2v_reg ;
  assign \piso.data_r [224] = \piso.data_r_224_sv2v_reg ;
  assign \piso.data_r [223] = \piso.data_r_223_sv2v_reg ;
  assign \piso.data_r [222] = \piso.data_r_222_sv2v_reg ;
  assign \piso.data_r [221] = \piso.data_r_221_sv2v_reg ;
  assign \piso.data_r [220] = \piso.data_r_220_sv2v_reg ;
  assign \piso.data_r [219] = \piso.data_r_219_sv2v_reg ;
  assign \piso.data_r [218] = \piso.data_r_218_sv2v_reg ;
  assign \piso.data_r [217] = \piso.data_r_217_sv2v_reg ;
  assign \piso.data_r [216] = \piso.data_r_216_sv2v_reg ;
  assign \piso.data_r [215] = \piso.data_r_215_sv2v_reg ;
  assign \piso.data_r [214] = \piso.data_r_214_sv2v_reg ;
  assign \piso.data_r [213] = \piso.data_r_213_sv2v_reg ;
  assign \piso.data_r [212] = \piso.data_r_212_sv2v_reg ;
  assign \piso.data_r [211] = \piso.data_r_211_sv2v_reg ;
  assign \piso.data_r [210] = \piso.data_r_210_sv2v_reg ;
  assign \piso.data_r [209] = \piso.data_r_209_sv2v_reg ;
  assign \piso.data_r [208] = \piso.data_r_208_sv2v_reg ;
  assign \piso.data_r [207] = \piso.data_r_207_sv2v_reg ;
  assign \piso.data_r [206] = \piso.data_r_206_sv2v_reg ;
  assign \piso.data_r [205] = \piso.data_r_205_sv2v_reg ;
  assign \piso.data_r [204] = \piso.data_r_204_sv2v_reg ;
  assign \piso.data_r [203] = \piso.data_r_203_sv2v_reg ;
  assign \piso.data_r [202] = \piso.data_r_202_sv2v_reg ;
  assign \piso.data_r [201] = \piso.data_r_201_sv2v_reg ;
  assign \piso.data_r [200] = \piso.data_r_200_sv2v_reg ;
  assign \piso.data_r [199] = \piso.data_r_199_sv2v_reg ;
  assign \piso.data_r [198] = \piso.data_r_198_sv2v_reg ;
  assign \piso.data_r [197] = \piso.data_r_197_sv2v_reg ;
  assign \piso.data_r [196] = \piso.data_r_196_sv2v_reg ;
  assign \piso.data_r [195] = \piso.data_r_195_sv2v_reg ;
  assign \piso.data_r [194] = \piso.data_r_194_sv2v_reg ;
  assign \piso.data_r [193] = \piso.data_r_193_sv2v_reg ;
  assign \piso.data_r [192] = \piso.data_r_192_sv2v_reg ;
  assign \piso.data_r [191] = \piso.data_r_191_sv2v_reg ;
  assign \piso.data_r [190] = \piso.data_r_190_sv2v_reg ;
  assign \piso.data_r [189] = \piso.data_r_189_sv2v_reg ;
  assign \piso.data_r [188] = \piso.data_r_188_sv2v_reg ;
  assign \piso.data_r [187] = \piso.data_r_187_sv2v_reg ;
  assign \piso.data_r [186] = \piso.data_r_186_sv2v_reg ;
  assign \piso.data_r [185] = \piso.data_r_185_sv2v_reg ;
  assign \piso.data_r [184] = \piso.data_r_184_sv2v_reg ;
  assign \piso.data_r [183] = \piso.data_r_183_sv2v_reg ;
  assign \piso.data_r [182] = \piso.data_r_182_sv2v_reg ;
  assign \piso.data_r [181] = \piso.data_r_181_sv2v_reg ;
  assign \piso.data_r [180] = \piso.data_r_180_sv2v_reg ;
  assign \piso.data_r [179] = \piso.data_r_179_sv2v_reg ;
  assign \piso.data_r [178] = \piso.data_r_178_sv2v_reg ;
  assign \piso.data_r [177] = \piso.data_r_177_sv2v_reg ;
  assign \piso.data_r [176] = \piso.data_r_176_sv2v_reg ;
  assign \piso.data_r [175] = \piso.data_r_175_sv2v_reg ;
  assign \piso.data_r [174] = \piso.data_r_174_sv2v_reg ;
  assign \piso.data_r [173] = \piso.data_r_173_sv2v_reg ;
  assign \piso.data_r [172] = \piso.data_r_172_sv2v_reg ;
  assign \piso.data_r [171] = \piso.data_r_171_sv2v_reg ;
  assign \piso.data_r [170] = \piso.data_r_170_sv2v_reg ;
  assign \piso.data_r [169] = \piso.data_r_169_sv2v_reg ;
  assign \piso.data_r [168] = \piso.data_r_168_sv2v_reg ;
  assign \piso.data_r [167] = \piso.data_r_167_sv2v_reg ;
  assign \piso.data_r [166] = \piso.data_r_166_sv2v_reg ;
  assign \piso.data_r [165] = \piso.data_r_165_sv2v_reg ;
  assign \piso.data_r [164] = \piso.data_r_164_sv2v_reg ;
  assign \piso.data_r [163] = \piso.data_r_163_sv2v_reg ;
  assign \piso.data_r [162] = \piso.data_r_162_sv2v_reg ;
  assign \piso.data_r [161] = \piso.data_r_161_sv2v_reg ;
  assign \piso.data_r [160] = \piso.data_r_160_sv2v_reg ;
  assign \piso.data_r [159] = \piso.data_r_159_sv2v_reg ;
  assign \piso.data_r [158] = \piso.data_r_158_sv2v_reg ;
  assign \piso.data_r [157] = \piso.data_r_157_sv2v_reg ;
  assign \piso.data_r [156] = \piso.data_r_156_sv2v_reg ;
  assign \piso.data_r [155] = \piso.data_r_155_sv2v_reg ;
  assign \piso.data_r [154] = \piso.data_r_154_sv2v_reg ;
  assign \piso.data_r [153] = \piso.data_r_153_sv2v_reg ;
  assign \piso.data_r [152] = \piso.data_r_152_sv2v_reg ;
  assign \piso.data_r [151] = \piso.data_r_151_sv2v_reg ;
  assign \piso.data_r [150] = \piso.data_r_150_sv2v_reg ;
  assign \piso.data_r [149] = \piso.data_r_149_sv2v_reg ;
  assign \piso.data_r [148] = \piso.data_r_148_sv2v_reg ;
  assign \piso.data_r [147] = \piso.data_r_147_sv2v_reg ;
  assign \piso.data_r [146] = \piso.data_r_146_sv2v_reg ;
  assign \piso.data_r [145] = \piso.data_r_145_sv2v_reg ;
  assign \piso.data_r [144] = \piso.data_r_144_sv2v_reg ;
  assign \piso.data_r [143] = \piso.data_r_143_sv2v_reg ;
  assign \piso.data_r [142] = \piso.data_r_142_sv2v_reg ;
  assign \piso.data_r [141] = \piso.data_r_141_sv2v_reg ;
  assign \piso.data_r [140] = \piso.data_r_140_sv2v_reg ;
  assign \piso.data_r [139] = \piso.data_r_139_sv2v_reg ;
  assign \piso.data_r [138] = \piso.data_r_138_sv2v_reg ;
  assign \piso.data_r [137] = \piso.data_r_137_sv2v_reg ;
  assign \piso.data_r [136] = \piso.data_r_136_sv2v_reg ;
  assign \piso.data_r [135] = \piso.data_r_135_sv2v_reg ;
  assign \piso.data_r [134] = \piso.data_r_134_sv2v_reg ;
  assign \piso.data_r [133] = \piso.data_r_133_sv2v_reg ;
  assign \piso.data_r [132] = \piso.data_r_132_sv2v_reg ;
  assign \piso.data_r [131] = \piso.data_r_131_sv2v_reg ;
  assign \piso.data_r [130] = \piso.data_r_130_sv2v_reg ;
  assign \piso.data_r [129] = \piso.data_r_129_sv2v_reg ;
  assign \piso.data_r [128] = \piso.data_r_128_sv2v_reg ;
  assign \piso.data_r [127] = \piso.data_r_127_sv2v_reg ;
  assign \piso.data_r [126] = \piso.data_r_126_sv2v_reg ;
  assign \piso.data_r [125] = \piso.data_r_125_sv2v_reg ;
  assign \piso.data_r [124] = \piso.data_r_124_sv2v_reg ;
  assign \piso.data_r [123] = \piso.data_r_123_sv2v_reg ;
  assign \piso.data_r [122] = \piso.data_r_122_sv2v_reg ;
  assign \piso.data_r [121] = \piso.data_r_121_sv2v_reg ;
  assign \piso.data_r [120] = \piso.data_r_120_sv2v_reg ;
  assign \piso.data_r [119] = \piso.data_r_119_sv2v_reg ;
  assign \piso.data_r [118] = \piso.data_r_118_sv2v_reg ;
  assign \piso.data_r [117] = \piso.data_r_117_sv2v_reg ;
  assign \piso.data_r [116] = \piso.data_r_116_sv2v_reg ;
  assign \piso.data_r [115] = \piso.data_r_115_sv2v_reg ;
  assign \piso.data_r [114] = \piso.data_r_114_sv2v_reg ;
  assign \piso.data_r [113] = \piso.data_r_113_sv2v_reg ;
  assign \piso.data_r [112] = \piso.data_r_112_sv2v_reg ;
  assign \piso.data_r [111] = \piso.data_r_111_sv2v_reg ;
  assign \piso.data_r [110] = \piso.data_r_110_sv2v_reg ;
  assign \piso.data_r [109] = \piso.data_r_109_sv2v_reg ;
  assign \piso.data_r [108] = \piso.data_r_108_sv2v_reg ;
  assign \piso.data_r [107] = \piso.data_r_107_sv2v_reg ;
  assign \piso.data_r [106] = \piso.data_r_106_sv2v_reg ;
  assign \piso.data_r [105] = \piso.data_r_105_sv2v_reg ;
  assign \piso.data_r [104] = \piso.data_r_104_sv2v_reg ;
  assign \piso.data_r [103] = \piso.data_r_103_sv2v_reg ;
  assign \piso.data_r [102] = \piso.data_r_102_sv2v_reg ;
  assign \piso.data_r [101] = \piso.data_r_101_sv2v_reg ;
  assign \piso.data_r [100] = \piso.data_r_100_sv2v_reg ;
  assign \piso.data_r [99] = \piso.data_r_99_sv2v_reg ;
  assign \piso.data_r [98] = \piso.data_r_98_sv2v_reg ;
  assign \piso.data_r [97] = \piso.data_r_97_sv2v_reg ;
  assign \piso.data_r [96] = \piso.data_r_96_sv2v_reg ;
  assign \piso.data_r [95] = \piso.data_r_95_sv2v_reg ;
  assign \piso.data_r [94] = \piso.data_r_94_sv2v_reg ;
  assign \piso.data_r [93] = \piso.data_r_93_sv2v_reg ;
  assign \piso.data_r [92] = \piso.data_r_92_sv2v_reg ;
  assign \piso.data_r [91] = \piso.data_r_91_sv2v_reg ;
  assign \piso.data_r [90] = \piso.data_r_90_sv2v_reg ;
  assign \piso.data_r [89] = \piso.data_r_89_sv2v_reg ;
  assign \piso.data_r [88] = \piso.data_r_88_sv2v_reg ;
  assign \piso.data_r [87] = \piso.data_r_87_sv2v_reg ;
  assign \piso.data_r [86] = \piso.data_r_86_sv2v_reg ;
  assign \piso.data_r [85] = \piso.data_r_85_sv2v_reg ;
  assign \piso.data_r [84] = \piso.data_r_84_sv2v_reg ;
  assign \piso.data_r [83] = \piso.data_r_83_sv2v_reg ;
  assign \piso.data_r [82] = \piso.data_r_82_sv2v_reg ;
  assign \piso.data_r [81] = \piso.data_r_81_sv2v_reg ;
  assign \piso.data_r [80] = \piso.data_r_80_sv2v_reg ;
  assign \piso.data_r [79] = \piso.data_r_79_sv2v_reg ;
  assign \piso.data_r [78] = \piso.data_r_78_sv2v_reg ;
  assign \piso.data_r [77] = \piso.data_r_77_sv2v_reg ;
  assign \piso.data_r [76] = \piso.data_r_76_sv2v_reg ;
  assign \piso.data_r [75] = \piso.data_r_75_sv2v_reg ;
  assign \piso.data_r [74] = \piso.data_r_74_sv2v_reg ;
  assign \piso.data_r [73] = \piso.data_r_73_sv2v_reg ;
  assign \piso.data_r [72] = \piso.data_r_72_sv2v_reg ;
  assign \piso.data_r [71] = \piso.data_r_71_sv2v_reg ;
  assign \piso.data_r [70] = \piso.data_r_70_sv2v_reg ;
  assign \piso.data_r [69] = \piso.data_r_69_sv2v_reg ;
  assign \piso.data_r [68] = \piso.data_r_68_sv2v_reg ;
  assign \piso.data_r [67] = \piso.data_r_67_sv2v_reg ;
  assign \piso.data_r [66] = \piso.data_r_66_sv2v_reg ;
  assign \piso.data_r [65] = \piso.data_r_65_sv2v_reg ;
  assign \piso.data_r [64] = \piso.data_r_64_sv2v_reg ;
  assign \piso.data_r [63] = \piso.data_r_63_sv2v_reg ;
  assign \piso.data_r [62] = \piso.data_r_62_sv2v_reg ;
  assign \piso.data_r [61] = \piso.data_r_61_sv2v_reg ;
  assign \piso.data_r [60] = \piso.data_r_60_sv2v_reg ;
  assign \piso.data_r [59] = \piso.data_r_59_sv2v_reg ;
  assign \piso.data_r [58] = \piso.data_r_58_sv2v_reg ;
  assign \piso.data_r [57] = \piso.data_r_57_sv2v_reg ;
  assign \piso.data_r [56] = \piso.data_r_56_sv2v_reg ;
  assign \piso.data_r [55] = \piso.data_r_55_sv2v_reg ;
  assign \piso.data_r [54] = \piso.data_r_54_sv2v_reg ;
  assign \piso.data_r [53] = \piso.data_r_53_sv2v_reg ;
  assign \piso.data_r [52] = \piso.data_r_52_sv2v_reg ;
  assign \piso.data_r [51] = \piso.data_r_51_sv2v_reg ;
  assign \piso.data_r [50] = \piso.data_r_50_sv2v_reg ;
  assign \piso.data_r [49] = \piso.data_r_49_sv2v_reg ;
  assign \piso.data_r [48] = \piso.data_r_48_sv2v_reg ;
  assign \piso.data_r [47] = \piso.data_r_47_sv2v_reg ;
  assign \piso.data_r [46] = \piso.data_r_46_sv2v_reg ;
  assign \piso.data_r [45] = \piso.data_r_45_sv2v_reg ;
  assign \piso.data_r [44] = \piso.data_r_44_sv2v_reg ;
  assign \piso.data_r [43] = \piso.data_r_43_sv2v_reg ;
  assign \piso.data_r [42] = \piso.data_r_42_sv2v_reg ;
  assign \piso.data_r [41] = \piso.data_r_41_sv2v_reg ;
  assign \piso.data_r [40] = \piso.data_r_40_sv2v_reg ;
  assign \piso.data_r [39] = \piso.data_r_39_sv2v_reg ;
  assign \piso.data_r [38] = \piso.data_r_38_sv2v_reg ;
  assign \piso.data_r [37] = \piso.data_r_37_sv2v_reg ;
  assign \piso.data_r [36] = \piso.data_r_36_sv2v_reg ;
  assign \piso.data_r [35] = \piso.data_r_35_sv2v_reg ;
  assign \piso.data_r [34] = \piso.data_r_34_sv2v_reg ;
  assign \piso.data_r [33] = \piso.data_r_33_sv2v_reg ;
  assign \piso.data_r [32] = \piso.data_r_32_sv2v_reg ;
  assign \piso.data_r [31] = \piso.data_r_31_sv2v_reg ;
  assign \piso.data_r [30] = \piso.data_r_30_sv2v_reg ;
  assign \piso.data_r [29] = \piso.data_r_29_sv2v_reg ;
  assign \piso.data_r [28] = \piso.data_r_28_sv2v_reg ;
  assign \piso.data_r [27] = \piso.data_r_27_sv2v_reg ;
  assign \piso.data_r [26] = \piso.data_r_26_sv2v_reg ;
  assign \piso.data_r [25] = \piso.data_r_25_sv2v_reg ;
  assign \piso.data_r [24] = \piso.data_r_24_sv2v_reg ;
  assign \piso.data_r [23] = \piso.data_r_23_sv2v_reg ;
  assign \piso.data_r [22] = \piso.data_r_22_sv2v_reg ;
  assign \piso.data_r [21] = \piso.data_r_21_sv2v_reg ;
  assign \piso.data_r [20] = \piso.data_r_20_sv2v_reg ;
  assign \piso.data_r [19] = \piso.data_r_19_sv2v_reg ;
  assign \piso.data_r [18] = \piso.data_r_18_sv2v_reg ;
  assign \piso.data_r [17] = \piso.data_r_17_sv2v_reg ;
  assign \piso.data_r [16] = \piso.data_r_16_sv2v_reg ;
  assign \piso.data_r [15] = \piso.data_r_15_sv2v_reg ;
  assign \piso.data_r [14] = \piso.data_r_14_sv2v_reg ;
  assign \piso.data_r [13] = \piso.data_r_13_sv2v_reg ;
  assign \piso.data_r [12] = \piso.data_r_12_sv2v_reg ;
  assign \piso.data_r [11] = \piso.data_r_11_sv2v_reg ;
  assign \piso.data_r [10] = \piso.data_r_10_sv2v_reg ;
  assign \piso.data_r [9] = \piso.data_r_9_sv2v_reg ;
  assign \piso.data_r [8] = \piso.data_r_8_sv2v_reg ;
  assign \piso.data_r [7] = \piso.data_r_7_sv2v_reg ;
  assign \piso.data_r [6] = \piso.data_r_6_sv2v_reg ;
  assign \piso.data_r [5] = \piso.data_r_5_sv2v_reg ;
  assign \piso.data_r [4] = \piso.data_r_4_sv2v_reg ;
  assign \piso.data_r [3] = \piso.data_r_3_sv2v_reg ;
  assign \piso.data_r [2] = \piso.data_r_2_sv2v_reg ;
  assign \piso.data_r [1] = \piso.data_r_1_sv2v_reg ;
  assign \piso.data_r [0] = \piso.data_r_0_sv2v_reg ;
  assign \piso.shift_ctr_r [6] = \piso.shift_ctr_r_6_sv2v_reg ;
  assign \piso.shift_ctr_r [5] = \piso.shift_ctr_r_5_sv2v_reg ;
  assign \piso.shift_ctr_r [4] = \piso.shift_ctr_r_4_sv2v_reg ;
  assign \piso.shift_ctr_r [3] = \piso.shift_ctr_r_3_sv2v_reg ;
  assign \piso.shift_ctr_r [2] = \piso.shift_ctr_r_2_sv2v_reg ;
  assign \piso.shift_ctr_r [1] = \piso.shift_ctr_r_1_sv2v_reg ;
  assign \piso.shift_ctr_r [0] = \piso.shift_ctr_r_0_sv2v_reg ;

  bsg_array_reverse_width_p32_els_p128
  \piso.hi2lo.bar 
  (
    .i(data_i),
    .o(\piso.data_li )
  );

  assign data_o[31] = (N156)? \piso.data_r [31] : 
                      (N158)? \piso.data_r [63] : 
                      (N160)? \piso.data_r [95] : 
                      (N162)? \piso.data_r [127] : 
                      (N164)? \piso.data_r [159] : 
                      (N166)? \piso.data_r [191] : 
                      (N168)? \piso.data_r [223] : 
                      (N170)? \piso.data_r [255] : 
                      (N172)? \piso.data_r [287] : 
                      (N174)? \piso.data_r [319] : 
                      (N176)? \piso.data_r [351] : 
                      (N178)? \piso.data_r [383] : 
                      (N180)? \piso.data_r [415] : 
                      (N182)? \piso.data_r [447] : 
                      (N184)? \piso.data_r [479] : 
                      (N186)? \piso.data_r [511] : 
                      (N188)? \piso.data_r [543] : 
                      (N190)? \piso.data_r [575] : 
                      (N192)? \piso.data_r [607] : 
                      (N194)? \piso.data_r [639] : 
                      (N196)? \piso.data_r [671] : 
                      (N198)? \piso.data_r [703] : 
                      (N200)? \piso.data_r [735] : 
                      (N202)? \piso.data_r [767] : 
                      (N204)? \piso.data_r [799] : 
                      (N206)? \piso.data_r [831] : 
                      (N208)? \piso.data_r [863] : 
                      (N210)? \piso.data_r [895] : 
                      (N212)? \piso.data_r [927] : 
                      (N214)? \piso.data_r [959] : 
                      (N216)? \piso.data_r [991] : 
                      (N218)? \piso.data_r [1023] : 
                      (N220)? \piso.data_r [1055] : 
                      (N222)? \piso.data_r [1087] : 
                      (N224)? \piso.data_r [1119] : 
                      (N226)? \piso.data_r [1151] : 
                      (N228)? \piso.data_r [1183] : 
                      (N230)? \piso.data_r [1215] : 
                      (N232)? \piso.data_r [1247] : 
                      (N234)? \piso.data_r [1279] : 
                      (N236)? \piso.data_r [1311] : 
                      (N238)? \piso.data_r [1343] : 
                      (N240)? \piso.data_r [1375] : 
                      (N242)? \piso.data_r [1407] : 
                      (N244)? \piso.data_r [1439] : 
                      (N246)? \piso.data_r [1471] : 
                      (N248)? \piso.data_r [1503] : 
                      (N250)? \piso.data_r [1535] : 
                      (N252)? \piso.data_r [1567] : 
                      (N254)? \piso.data_r [1599] : 
                      (N256)? \piso.data_r [1631] : 
                      (N258)? \piso.data_r [1663] : 
                      (N260)? \piso.data_r [1695] : 
                      (N262)? \piso.data_r [1727] : 
                      (N264)? \piso.data_r [1759] : 
                      (N266)? \piso.data_r [1791] : 
                      (N268)? \piso.data_r [1823] : 
                      (N270)? \piso.data_r [1855] : 
                      (N272)? \piso.data_r [1887] : 
                      (N274)? \piso.data_r [1919] : 
                      (N276)? \piso.data_r [1951] : 
                      (N278)? \piso.data_r [1983] : 
                      (N280)? \piso.data_r [2015] : 
                      (N282)? \piso.data_r [2047] : 
                      (N157)? \piso.data_r [2079] : 
                      (N159)? \piso.data_r [2111] : 
                      (N161)? \piso.data_r [2143] : 
                      (N163)? \piso.data_r [2175] : 
                      (N165)? \piso.data_r [2207] : 
                      (N167)? \piso.data_r [2239] : 
                      (N169)? \piso.data_r [2271] : 
                      (N171)? \piso.data_r [2303] : 
                      (N173)? \piso.data_r [2335] : 
                      (N175)? \piso.data_r [2367] : 
                      (N177)? \piso.data_r [2399] : 
                      (N179)? \piso.data_r [2431] : 
                      (N181)? \piso.data_r [2463] : 
                      (N183)? \piso.data_r [2495] : 
                      (N185)? \piso.data_r [2527] : 
                      (N187)? \piso.data_r [2559] : 
                      (N189)? \piso.data_r [2591] : 
                      (N191)? \piso.data_r [2623] : 
                      (N193)? \piso.data_r [2655] : 
                      (N195)? \piso.data_r [2687] : 
                      (N197)? \piso.data_r [2719] : 
                      (N199)? \piso.data_r [2751] : 
                      (N201)? \piso.data_r [2783] : 
                      (N203)? \piso.data_r [2815] : 
                      (N205)? \piso.data_r [2847] : 
                      (N207)? \piso.data_r [2879] : 
                      (N209)? \piso.data_r [2911] : 
                      (N211)? \piso.data_r [2943] : 
                      (N213)? \piso.data_r [2975] : 
                      (N215)? \piso.data_r [3007] : 
                      (N217)? \piso.data_r [3039] : 
                      (N219)? \piso.data_r [3071] : 
                      (N221)? \piso.data_r [3103] : 
                      (N223)? \piso.data_r [3135] : 
                      (N225)? \piso.data_r [3167] : 
                      (N227)? \piso.data_r [3199] : 
                      (N229)? \piso.data_r [3231] : 
                      (N231)? \piso.data_r [3263] : 
                      (N233)? \piso.data_r [3295] : 
                      (N235)? \piso.data_r [3327] : 
                      (N237)? \piso.data_r [3359] : 
                      (N239)? \piso.data_r [3391] : 
                      (N241)? \piso.data_r [3423] : 
                      (N243)? \piso.data_r [3455] : 
                      (N245)? \piso.data_r [3487] : 
                      (N247)? \piso.data_r [3519] : 
                      (N249)? \piso.data_r [3551] : 
                      (N251)? \piso.data_r [3583] : 
                      (N253)? \piso.data_r [3615] : 
                      (N255)? \piso.data_r [3647] : 
                      (N257)? \piso.data_r [3679] : 
                      (N259)? \piso.data_r [3711] : 
                      (N261)? \piso.data_r [3743] : 
                      (N263)? \piso.data_r [3775] : 
                      (N265)? \piso.data_r [3807] : 
                      (N267)? \piso.data_r [3839] : 
                      (N269)? \piso.data_r [3871] : 
                      (N271)? \piso.data_r [3903] : 
                      (N273)? \piso.data_r [3935] : 
                      (N275)? \piso.data_r [3967] : 
                      (N277)? \piso.data_r [3999] : 
                      (N279)? \piso.data_r [4031] : 
                      (N281)? \piso.data_r [4063] : 
                      (N283)? \piso.data_r [4095] : 1'b0;
  assign data_o[30] = (N156)? \piso.data_r [30] : 
                      (N158)? \piso.data_r [62] : 
                      (N160)? \piso.data_r [94] : 
                      (N162)? \piso.data_r [126] : 
                      (N164)? \piso.data_r [158] : 
                      (N166)? \piso.data_r [190] : 
                      (N168)? \piso.data_r [222] : 
                      (N170)? \piso.data_r [254] : 
                      (N172)? \piso.data_r [286] : 
                      (N174)? \piso.data_r [318] : 
                      (N176)? \piso.data_r [350] : 
                      (N178)? \piso.data_r [382] : 
                      (N180)? \piso.data_r [414] : 
                      (N182)? \piso.data_r [446] : 
                      (N184)? \piso.data_r [478] : 
                      (N186)? \piso.data_r [510] : 
                      (N188)? \piso.data_r [542] : 
                      (N190)? \piso.data_r [574] : 
                      (N192)? \piso.data_r [606] : 
                      (N194)? \piso.data_r [638] : 
                      (N196)? \piso.data_r [670] : 
                      (N198)? \piso.data_r [702] : 
                      (N200)? \piso.data_r [734] : 
                      (N202)? \piso.data_r [766] : 
                      (N204)? \piso.data_r [798] : 
                      (N206)? \piso.data_r [830] : 
                      (N208)? \piso.data_r [862] : 
                      (N210)? \piso.data_r [894] : 
                      (N212)? \piso.data_r [926] : 
                      (N214)? \piso.data_r [958] : 
                      (N216)? \piso.data_r [990] : 
                      (N218)? \piso.data_r [1022] : 
                      (N220)? \piso.data_r [1054] : 
                      (N222)? \piso.data_r [1086] : 
                      (N224)? \piso.data_r [1118] : 
                      (N226)? \piso.data_r [1150] : 
                      (N228)? \piso.data_r [1182] : 
                      (N230)? \piso.data_r [1214] : 
                      (N232)? \piso.data_r [1246] : 
                      (N234)? \piso.data_r [1278] : 
                      (N236)? \piso.data_r [1310] : 
                      (N238)? \piso.data_r [1342] : 
                      (N240)? \piso.data_r [1374] : 
                      (N242)? \piso.data_r [1406] : 
                      (N244)? \piso.data_r [1438] : 
                      (N246)? \piso.data_r [1470] : 
                      (N248)? \piso.data_r [1502] : 
                      (N250)? \piso.data_r [1534] : 
                      (N252)? \piso.data_r [1566] : 
                      (N254)? \piso.data_r [1598] : 
                      (N256)? \piso.data_r [1630] : 
                      (N258)? \piso.data_r [1662] : 
                      (N260)? \piso.data_r [1694] : 
                      (N262)? \piso.data_r [1726] : 
                      (N264)? \piso.data_r [1758] : 
                      (N266)? \piso.data_r [1790] : 
                      (N268)? \piso.data_r [1822] : 
                      (N270)? \piso.data_r [1854] : 
                      (N272)? \piso.data_r [1886] : 
                      (N274)? \piso.data_r [1918] : 
                      (N276)? \piso.data_r [1950] : 
                      (N278)? \piso.data_r [1982] : 
                      (N280)? \piso.data_r [2014] : 
                      (N282)? \piso.data_r [2046] : 
                      (N157)? \piso.data_r [2078] : 
                      (N159)? \piso.data_r [2110] : 
                      (N161)? \piso.data_r [2142] : 
                      (N163)? \piso.data_r [2174] : 
                      (N165)? \piso.data_r [2206] : 
                      (N167)? \piso.data_r [2238] : 
                      (N169)? \piso.data_r [2270] : 
                      (N171)? \piso.data_r [2302] : 
                      (N173)? \piso.data_r [2334] : 
                      (N175)? \piso.data_r [2366] : 
                      (N177)? \piso.data_r [2398] : 
                      (N179)? \piso.data_r [2430] : 
                      (N181)? \piso.data_r [2462] : 
                      (N183)? \piso.data_r [2494] : 
                      (N185)? \piso.data_r [2526] : 
                      (N187)? \piso.data_r [2558] : 
                      (N189)? \piso.data_r [2590] : 
                      (N191)? \piso.data_r [2622] : 
                      (N193)? \piso.data_r [2654] : 
                      (N195)? \piso.data_r [2686] : 
                      (N197)? \piso.data_r [2718] : 
                      (N199)? \piso.data_r [2750] : 
                      (N201)? \piso.data_r [2782] : 
                      (N203)? \piso.data_r [2814] : 
                      (N205)? \piso.data_r [2846] : 
                      (N207)? \piso.data_r [2878] : 
                      (N209)? \piso.data_r [2910] : 
                      (N211)? \piso.data_r [2942] : 
                      (N213)? \piso.data_r [2974] : 
                      (N215)? \piso.data_r [3006] : 
                      (N217)? \piso.data_r [3038] : 
                      (N219)? \piso.data_r [3070] : 
                      (N221)? \piso.data_r [3102] : 
                      (N223)? \piso.data_r [3134] : 
                      (N225)? \piso.data_r [3166] : 
                      (N227)? \piso.data_r [3198] : 
                      (N229)? \piso.data_r [3230] : 
                      (N231)? \piso.data_r [3262] : 
                      (N233)? \piso.data_r [3294] : 
                      (N235)? \piso.data_r [3326] : 
                      (N237)? \piso.data_r [3358] : 
                      (N239)? \piso.data_r [3390] : 
                      (N241)? \piso.data_r [3422] : 
                      (N243)? \piso.data_r [3454] : 
                      (N245)? \piso.data_r [3486] : 
                      (N247)? \piso.data_r [3518] : 
                      (N249)? \piso.data_r [3550] : 
                      (N251)? \piso.data_r [3582] : 
                      (N253)? \piso.data_r [3614] : 
                      (N255)? \piso.data_r [3646] : 
                      (N257)? \piso.data_r [3678] : 
                      (N259)? \piso.data_r [3710] : 
                      (N261)? \piso.data_r [3742] : 
                      (N263)? \piso.data_r [3774] : 
                      (N265)? \piso.data_r [3806] : 
                      (N267)? \piso.data_r [3838] : 
                      (N269)? \piso.data_r [3870] : 
                      (N271)? \piso.data_r [3902] : 
                      (N273)? \piso.data_r [3934] : 
                      (N275)? \piso.data_r [3966] : 
                      (N277)? \piso.data_r [3998] : 
                      (N279)? \piso.data_r [4030] : 
                      (N281)? \piso.data_r [4062] : 
                      (N283)? \piso.data_r [4094] : 1'b0;
  assign data_o[29] = (N156)? \piso.data_r [29] : 
                      (N158)? \piso.data_r [61] : 
                      (N160)? \piso.data_r [93] : 
                      (N162)? \piso.data_r [125] : 
                      (N164)? \piso.data_r [157] : 
                      (N166)? \piso.data_r [189] : 
                      (N168)? \piso.data_r [221] : 
                      (N170)? \piso.data_r [253] : 
                      (N172)? \piso.data_r [285] : 
                      (N174)? \piso.data_r [317] : 
                      (N176)? \piso.data_r [349] : 
                      (N178)? \piso.data_r [381] : 
                      (N180)? \piso.data_r [413] : 
                      (N182)? \piso.data_r [445] : 
                      (N184)? \piso.data_r [477] : 
                      (N186)? \piso.data_r [509] : 
                      (N188)? \piso.data_r [541] : 
                      (N190)? \piso.data_r [573] : 
                      (N192)? \piso.data_r [605] : 
                      (N194)? \piso.data_r [637] : 
                      (N196)? \piso.data_r [669] : 
                      (N198)? \piso.data_r [701] : 
                      (N200)? \piso.data_r [733] : 
                      (N202)? \piso.data_r [765] : 
                      (N204)? \piso.data_r [797] : 
                      (N206)? \piso.data_r [829] : 
                      (N208)? \piso.data_r [861] : 
                      (N210)? \piso.data_r [893] : 
                      (N212)? \piso.data_r [925] : 
                      (N214)? \piso.data_r [957] : 
                      (N216)? \piso.data_r [989] : 
                      (N218)? \piso.data_r [1021] : 
                      (N220)? \piso.data_r [1053] : 
                      (N222)? \piso.data_r [1085] : 
                      (N224)? \piso.data_r [1117] : 
                      (N226)? \piso.data_r [1149] : 
                      (N228)? \piso.data_r [1181] : 
                      (N230)? \piso.data_r [1213] : 
                      (N232)? \piso.data_r [1245] : 
                      (N234)? \piso.data_r [1277] : 
                      (N236)? \piso.data_r [1309] : 
                      (N238)? \piso.data_r [1341] : 
                      (N240)? \piso.data_r [1373] : 
                      (N242)? \piso.data_r [1405] : 
                      (N244)? \piso.data_r [1437] : 
                      (N246)? \piso.data_r [1469] : 
                      (N248)? \piso.data_r [1501] : 
                      (N250)? \piso.data_r [1533] : 
                      (N252)? \piso.data_r [1565] : 
                      (N254)? \piso.data_r [1597] : 
                      (N256)? \piso.data_r [1629] : 
                      (N258)? \piso.data_r [1661] : 
                      (N260)? \piso.data_r [1693] : 
                      (N262)? \piso.data_r [1725] : 
                      (N264)? \piso.data_r [1757] : 
                      (N266)? \piso.data_r [1789] : 
                      (N268)? \piso.data_r [1821] : 
                      (N270)? \piso.data_r [1853] : 
                      (N272)? \piso.data_r [1885] : 
                      (N274)? \piso.data_r [1917] : 
                      (N276)? \piso.data_r [1949] : 
                      (N278)? \piso.data_r [1981] : 
                      (N280)? \piso.data_r [2013] : 
                      (N282)? \piso.data_r [2045] : 
                      (N157)? \piso.data_r [2077] : 
                      (N159)? \piso.data_r [2109] : 
                      (N161)? \piso.data_r [2141] : 
                      (N163)? \piso.data_r [2173] : 
                      (N165)? \piso.data_r [2205] : 
                      (N167)? \piso.data_r [2237] : 
                      (N169)? \piso.data_r [2269] : 
                      (N171)? \piso.data_r [2301] : 
                      (N173)? \piso.data_r [2333] : 
                      (N175)? \piso.data_r [2365] : 
                      (N177)? \piso.data_r [2397] : 
                      (N179)? \piso.data_r [2429] : 
                      (N181)? \piso.data_r [2461] : 
                      (N183)? \piso.data_r [2493] : 
                      (N185)? \piso.data_r [2525] : 
                      (N187)? \piso.data_r [2557] : 
                      (N189)? \piso.data_r [2589] : 
                      (N191)? \piso.data_r [2621] : 
                      (N193)? \piso.data_r [2653] : 
                      (N195)? \piso.data_r [2685] : 
                      (N197)? \piso.data_r [2717] : 
                      (N199)? \piso.data_r [2749] : 
                      (N201)? \piso.data_r [2781] : 
                      (N203)? \piso.data_r [2813] : 
                      (N205)? \piso.data_r [2845] : 
                      (N207)? \piso.data_r [2877] : 
                      (N209)? \piso.data_r [2909] : 
                      (N211)? \piso.data_r [2941] : 
                      (N213)? \piso.data_r [2973] : 
                      (N215)? \piso.data_r [3005] : 
                      (N217)? \piso.data_r [3037] : 
                      (N219)? \piso.data_r [3069] : 
                      (N221)? \piso.data_r [3101] : 
                      (N223)? \piso.data_r [3133] : 
                      (N225)? \piso.data_r [3165] : 
                      (N227)? \piso.data_r [3197] : 
                      (N229)? \piso.data_r [3229] : 
                      (N231)? \piso.data_r [3261] : 
                      (N233)? \piso.data_r [3293] : 
                      (N235)? \piso.data_r [3325] : 
                      (N237)? \piso.data_r [3357] : 
                      (N239)? \piso.data_r [3389] : 
                      (N241)? \piso.data_r [3421] : 
                      (N243)? \piso.data_r [3453] : 
                      (N245)? \piso.data_r [3485] : 
                      (N247)? \piso.data_r [3517] : 
                      (N249)? \piso.data_r [3549] : 
                      (N251)? \piso.data_r [3581] : 
                      (N253)? \piso.data_r [3613] : 
                      (N255)? \piso.data_r [3645] : 
                      (N257)? \piso.data_r [3677] : 
                      (N259)? \piso.data_r [3709] : 
                      (N261)? \piso.data_r [3741] : 
                      (N263)? \piso.data_r [3773] : 
                      (N265)? \piso.data_r [3805] : 
                      (N267)? \piso.data_r [3837] : 
                      (N269)? \piso.data_r [3869] : 
                      (N271)? \piso.data_r [3901] : 
                      (N273)? \piso.data_r [3933] : 
                      (N275)? \piso.data_r [3965] : 
                      (N277)? \piso.data_r [3997] : 
                      (N279)? \piso.data_r [4029] : 
                      (N281)? \piso.data_r [4061] : 
                      (N283)? \piso.data_r [4093] : 1'b0;
  assign data_o[28] = (N156)? \piso.data_r [28] : 
                      (N158)? \piso.data_r [60] : 
                      (N160)? \piso.data_r [92] : 
                      (N162)? \piso.data_r [124] : 
                      (N164)? \piso.data_r [156] : 
                      (N166)? \piso.data_r [188] : 
                      (N168)? \piso.data_r [220] : 
                      (N170)? \piso.data_r [252] : 
                      (N172)? \piso.data_r [284] : 
                      (N174)? \piso.data_r [316] : 
                      (N176)? \piso.data_r [348] : 
                      (N178)? \piso.data_r [380] : 
                      (N180)? \piso.data_r [412] : 
                      (N182)? \piso.data_r [444] : 
                      (N184)? \piso.data_r [476] : 
                      (N186)? \piso.data_r [508] : 
                      (N188)? \piso.data_r [540] : 
                      (N190)? \piso.data_r [572] : 
                      (N192)? \piso.data_r [604] : 
                      (N194)? \piso.data_r [636] : 
                      (N196)? \piso.data_r [668] : 
                      (N198)? \piso.data_r [700] : 
                      (N200)? \piso.data_r [732] : 
                      (N202)? \piso.data_r [764] : 
                      (N204)? \piso.data_r [796] : 
                      (N206)? \piso.data_r [828] : 
                      (N208)? \piso.data_r [860] : 
                      (N210)? \piso.data_r [892] : 
                      (N212)? \piso.data_r [924] : 
                      (N214)? \piso.data_r [956] : 
                      (N216)? \piso.data_r [988] : 
                      (N218)? \piso.data_r [1020] : 
                      (N220)? \piso.data_r [1052] : 
                      (N222)? \piso.data_r [1084] : 
                      (N224)? \piso.data_r [1116] : 
                      (N226)? \piso.data_r [1148] : 
                      (N228)? \piso.data_r [1180] : 
                      (N230)? \piso.data_r [1212] : 
                      (N232)? \piso.data_r [1244] : 
                      (N234)? \piso.data_r [1276] : 
                      (N236)? \piso.data_r [1308] : 
                      (N238)? \piso.data_r [1340] : 
                      (N240)? \piso.data_r [1372] : 
                      (N242)? \piso.data_r [1404] : 
                      (N244)? \piso.data_r [1436] : 
                      (N246)? \piso.data_r [1468] : 
                      (N248)? \piso.data_r [1500] : 
                      (N250)? \piso.data_r [1532] : 
                      (N252)? \piso.data_r [1564] : 
                      (N254)? \piso.data_r [1596] : 
                      (N256)? \piso.data_r [1628] : 
                      (N258)? \piso.data_r [1660] : 
                      (N260)? \piso.data_r [1692] : 
                      (N262)? \piso.data_r [1724] : 
                      (N264)? \piso.data_r [1756] : 
                      (N266)? \piso.data_r [1788] : 
                      (N268)? \piso.data_r [1820] : 
                      (N270)? \piso.data_r [1852] : 
                      (N272)? \piso.data_r [1884] : 
                      (N274)? \piso.data_r [1916] : 
                      (N276)? \piso.data_r [1948] : 
                      (N278)? \piso.data_r [1980] : 
                      (N280)? \piso.data_r [2012] : 
                      (N282)? \piso.data_r [2044] : 
                      (N157)? \piso.data_r [2076] : 
                      (N159)? \piso.data_r [2108] : 
                      (N161)? \piso.data_r [2140] : 
                      (N163)? \piso.data_r [2172] : 
                      (N165)? \piso.data_r [2204] : 
                      (N167)? \piso.data_r [2236] : 
                      (N169)? \piso.data_r [2268] : 
                      (N171)? \piso.data_r [2300] : 
                      (N173)? \piso.data_r [2332] : 
                      (N175)? \piso.data_r [2364] : 
                      (N177)? \piso.data_r [2396] : 
                      (N179)? \piso.data_r [2428] : 
                      (N181)? \piso.data_r [2460] : 
                      (N183)? \piso.data_r [2492] : 
                      (N185)? \piso.data_r [2524] : 
                      (N187)? \piso.data_r [2556] : 
                      (N189)? \piso.data_r [2588] : 
                      (N191)? \piso.data_r [2620] : 
                      (N193)? \piso.data_r [2652] : 
                      (N195)? \piso.data_r [2684] : 
                      (N197)? \piso.data_r [2716] : 
                      (N199)? \piso.data_r [2748] : 
                      (N201)? \piso.data_r [2780] : 
                      (N203)? \piso.data_r [2812] : 
                      (N205)? \piso.data_r [2844] : 
                      (N207)? \piso.data_r [2876] : 
                      (N209)? \piso.data_r [2908] : 
                      (N211)? \piso.data_r [2940] : 
                      (N213)? \piso.data_r [2972] : 
                      (N215)? \piso.data_r [3004] : 
                      (N217)? \piso.data_r [3036] : 
                      (N219)? \piso.data_r [3068] : 
                      (N221)? \piso.data_r [3100] : 
                      (N223)? \piso.data_r [3132] : 
                      (N225)? \piso.data_r [3164] : 
                      (N227)? \piso.data_r [3196] : 
                      (N229)? \piso.data_r [3228] : 
                      (N231)? \piso.data_r [3260] : 
                      (N233)? \piso.data_r [3292] : 
                      (N235)? \piso.data_r [3324] : 
                      (N237)? \piso.data_r [3356] : 
                      (N239)? \piso.data_r [3388] : 
                      (N241)? \piso.data_r [3420] : 
                      (N243)? \piso.data_r [3452] : 
                      (N245)? \piso.data_r [3484] : 
                      (N247)? \piso.data_r [3516] : 
                      (N249)? \piso.data_r [3548] : 
                      (N251)? \piso.data_r [3580] : 
                      (N253)? \piso.data_r [3612] : 
                      (N255)? \piso.data_r [3644] : 
                      (N257)? \piso.data_r [3676] : 
                      (N259)? \piso.data_r [3708] : 
                      (N261)? \piso.data_r [3740] : 
                      (N263)? \piso.data_r [3772] : 
                      (N265)? \piso.data_r [3804] : 
                      (N267)? \piso.data_r [3836] : 
                      (N269)? \piso.data_r [3868] : 
                      (N271)? \piso.data_r [3900] : 
                      (N273)? \piso.data_r [3932] : 
                      (N275)? \piso.data_r [3964] : 
                      (N277)? \piso.data_r [3996] : 
                      (N279)? \piso.data_r [4028] : 
                      (N281)? \piso.data_r [4060] : 
                      (N283)? \piso.data_r [4092] : 1'b0;
  assign data_o[27] = (N156)? \piso.data_r [27] : 
                      (N158)? \piso.data_r [59] : 
                      (N160)? \piso.data_r [91] : 
                      (N162)? \piso.data_r [123] : 
                      (N164)? \piso.data_r [155] : 
                      (N166)? \piso.data_r [187] : 
                      (N168)? \piso.data_r [219] : 
                      (N170)? \piso.data_r [251] : 
                      (N172)? \piso.data_r [283] : 
                      (N174)? \piso.data_r [315] : 
                      (N176)? \piso.data_r [347] : 
                      (N178)? \piso.data_r [379] : 
                      (N180)? \piso.data_r [411] : 
                      (N182)? \piso.data_r [443] : 
                      (N184)? \piso.data_r [475] : 
                      (N186)? \piso.data_r [507] : 
                      (N188)? \piso.data_r [539] : 
                      (N190)? \piso.data_r [571] : 
                      (N192)? \piso.data_r [603] : 
                      (N194)? \piso.data_r [635] : 
                      (N196)? \piso.data_r [667] : 
                      (N198)? \piso.data_r [699] : 
                      (N200)? \piso.data_r [731] : 
                      (N202)? \piso.data_r [763] : 
                      (N204)? \piso.data_r [795] : 
                      (N206)? \piso.data_r [827] : 
                      (N208)? \piso.data_r [859] : 
                      (N210)? \piso.data_r [891] : 
                      (N212)? \piso.data_r [923] : 
                      (N214)? \piso.data_r [955] : 
                      (N216)? \piso.data_r [987] : 
                      (N218)? \piso.data_r [1019] : 
                      (N220)? \piso.data_r [1051] : 
                      (N222)? \piso.data_r [1083] : 
                      (N224)? \piso.data_r [1115] : 
                      (N226)? \piso.data_r [1147] : 
                      (N228)? \piso.data_r [1179] : 
                      (N230)? \piso.data_r [1211] : 
                      (N232)? \piso.data_r [1243] : 
                      (N234)? \piso.data_r [1275] : 
                      (N236)? \piso.data_r [1307] : 
                      (N238)? \piso.data_r [1339] : 
                      (N240)? \piso.data_r [1371] : 
                      (N242)? \piso.data_r [1403] : 
                      (N244)? \piso.data_r [1435] : 
                      (N246)? \piso.data_r [1467] : 
                      (N248)? \piso.data_r [1499] : 
                      (N250)? \piso.data_r [1531] : 
                      (N252)? \piso.data_r [1563] : 
                      (N254)? \piso.data_r [1595] : 
                      (N256)? \piso.data_r [1627] : 
                      (N258)? \piso.data_r [1659] : 
                      (N260)? \piso.data_r [1691] : 
                      (N262)? \piso.data_r [1723] : 
                      (N264)? \piso.data_r [1755] : 
                      (N266)? \piso.data_r [1787] : 
                      (N268)? \piso.data_r [1819] : 
                      (N270)? \piso.data_r [1851] : 
                      (N272)? \piso.data_r [1883] : 
                      (N274)? \piso.data_r [1915] : 
                      (N276)? \piso.data_r [1947] : 
                      (N278)? \piso.data_r [1979] : 
                      (N280)? \piso.data_r [2011] : 
                      (N282)? \piso.data_r [2043] : 
                      (N157)? \piso.data_r [2075] : 
                      (N159)? \piso.data_r [2107] : 
                      (N161)? \piso.data_r [2139] : 
                      (N163)? \piso.data_r [2171] : 
                      (N165)? \piso.data_r [2203] : 
                      (N167)? \piso.data_r [2235] : 
                      (N169)? \piso.data_r [2267] : 
                      (N171)? \piso.data_r [2299] : 
                      (N173)? \piso.data_r [2331] : 
                      (N175)? \piso.data_r [2363] : 
                      (N177)? \piso.data_r [2395] : 
                      (N179)? \piso.data_r [2427] : 
                      (N181)? \piso.data_r [2459] : 
                      (N183)? \piso.data_r [2491] : 
                      (N185)? \piso.data_r [2523] : 
                      (N187)? \piso.data_r [2555] : 
                      (N189)? \piso.data_r [2587] : 
                      (N191)? \piso.data_r [2619] : 
                      (N193)? \piso.data_r [2651] : 
                      (N195)? \piso.data_r [2683] : 
                      (N197)? \piso.data_r [2715] : 
                      (N199)? \piso.data_r [2747] : 
                      (N201)? \piso.data_r [2779] : 
                      (N203)? \piso.data_r [2811] : 
                      (N205)? \piso.data_r [2843] : 
                      (N207)? \piso.data_r [2875] : 
                      (N209)? \piso.data_r [2907] : 
                      (N211)? \piso.data_r [2939] : 
                      (N213)? \piso.data_r [2971] : 
                      (N215)? \piso.data_r [3003] : 
                      (N217)? \piso.data_r [3035] : 
                      (N219)? \piso.data_r [3067] : 
                      (N221)? \piso.data_r [3099] : 
                      (N223)? \piso.data_r [3131] : 
                      (N225)? \piso.data_r [3163] : 
                      (N227)? \piso.data_r [3195] : 
                      (N229)? \piso.data_r [3227] : 
                      (N231)? \piso.data_r [3259] : 
                      (N233)? \piso.data_r [3291] : 
                      (N235)? \piso.data_r [3323] : 
                      (N237)? \piso.data_r [3355] : 
                      (N239)? \piso.data_r [3387] : 
                      (N241)? \piso.data_r [3419] : 
                      (N243)? \piso.data_r [3451] : 
                      (N245)? \piso.data_r [3483] : 
                      (N247)? \piso.data_r [3515] : 
                      (N249)? \piso.data_r [3547] : 
                      (N251)? \piso.data_r [3579] : 
                      (N253)? \piso.data_r [3611] : 
                      (N255)? \piso.data_r [3643] : 
                      (N257)? \piso.data_r [3675] : 
                      (N259)? \piso.data_r [3707] : 
                      (N261)? \piso.data_r [3739] : 
                      (N263)? \piso.data_r [3771] : 
                      (N265)? \piso.data_r [3803] : 
                      (N267)? \piso.data_r [3835] : 
                      (N269)? \piso.data_r [3867] : 
                      (N271)? \piso.data_r [3899] : 
                      (N273)? \piso.data_r [3931] : 
                      (N275)? \piso.data_r [3963] : 
                      (N277)? \piso.data_r [3995] : 
                      (N279)? \piso.data_r [4027] : 
                      (N281)? \piso.data_r [4059] : 
                      (N283)? \piso.data_r [4091] : 1'b0;
  assign data_o[26] = (N156)? \piso.data_r [26] : 
                      (N158)? \piso.data_r [58] : 
                      (N160)? \piso.data_r [90] : 
                      (N162)? \piso.data_r [122] : 
                      (N164)? \piso.data_r [154] : 
                      (N166)? \piso.data_r [186] : 
                      (N168)? \piso.data_r [218] : 
                      (N170)? \piso.data_r [250] : 
                      (N172)? \piso.data_r [282] : 
                      (N174)? \piso.data_r [314] : 
                      (N176)? \piso.data_r [346] : 
                      (N178)? \piso.data_r [378] : 
                      (N180)? \piso.data_r [410] : 
                      (N182)? \piso.data_r [442] : 
                      (N184)? \piso.data_r [474] : 
                      (N186)? \piso.data_r [506] : 
                      (N188)? \piso.data_r [538] : 
                      (N190)? \piso.data_r [570] : 
                      (N192)? \piso.data_r [602] : 
                      (N194)? \piso.data_r [634] : 
                      (N196)? \piso.data_r [666] : 
                      (N198)? \piso.data_r [698] : 
                      (N200)? \piso.data_r [730] : 
                      (N202)? \piso.data_r [762] : 
                      (N204)? \piso.data_r [794] : 
                      (N206)? \piso.data_r [826] : 
                      (N208)? \piso.data_r [858] : 
                      (N210)? \piso.data_r [890] : 
                      (N212)? \piso.data_r [922] : 
                      (N214)? \piso.data_r [954] : 
                      (N216)? \piso.data_r [986] : 
                      (N218)? \piso.data_r [1018] : 
                      (N220)? \piso.data_r [1050] : 
                      (N222)? \piso.data_r [1082] : 
                      (N224)? \piso.data_r [1114] : 
                      (N226)? \piso.data_r [1146] : 
                      (N228)? \piso.data_r [1178] : 
                      (N230)? \piso.data_r [1210] : 
                      (N232)? \piso.data_r [1242] : 
                      (N234)? \piso.data_r [1274] : 
                      (N236)? \piso.data_r [1306] : 
                      (N238)? \piso.data_r [1338] : 
                      (N240)? \piso.data_r [1370] : 
                      (N242)? \piso.data_r [1402] : 
                      (N244)? \piso.data_r [1434] : 
                      (N246)? \piso.data_r [1466] : 
                      (N248)? \piso.data_r [1498] : 
                      (N250)? \piso.data_r [1530] : 
                      (N252)? \piso.data_r [1562] : 
                      (N254)? \piso.data_r [1594] : 
                      (N256)? \piso.data_r [1626] : 
                      (N258)? \piso.data_r [1658] : 
                      (N260)? \piso.data_r [1690] : 
                      (N262)? \piso.data_r [1722] : 
                      (N264)? \piso.data_r [1754] : 
                      (N266)? \piso.data_r [1786] : 
                      (N268)? \piso.data_r [1818] : 
                      (N270)? \piso.data_r [1850] : 
                      (N272)? \piso.data_r [1882] : 
                      (N274)? \piso.data_r [1914] : 
                      (N276)? \piso.data_r [1946] : 
                      (N278)? \piso.data_r [1978] : 
                      (N280)? \piso.data_r [2010] : 
                      (N282)? \piso.data_r [2042] : 
                      (N157)? \piso.data_r [2074] : 
                      (N159)? \piso.data_r [2106] : 
                      (N161)? \piso.data_r [2138] : 
                      (N163)? \piso.data_r [2170] : 
                      (N165)? \piso.data_r [2202] : 
                      (N167)? \piso.data_r [2234] : 
                      (N169)? \piso.data_r [2266] : 
                      (N171)? \piso.data_r [2298] : 
                      (N173)? \piso.data_r [2330] : 
                      (N175)? \piso.data_r [2362] : 
                      (N177)? \piso.data_r [2394] : 
                      (N179)? \piso.data_r [2426] : 
                      (N181)? \piso.data_r [2458] : 
                      (N183)? \piso.data_r [2490] : 
                      (N185)? \piso.data_r [2522] : 
                      (N187)? \piso.data_r [2554] : 
                      (N189)? \piso.data_r [2586] : 
                      (N191)? \piso.data_r [2618] : 
                      (N193)? \piso.data_r [2650] : 
                      (N195)? \piso.data_r [2682] : 
                      (N197)? \piso.data_r [2714] : 
                      (N199)? \piso.data_r [2746] : 
                      (N201)? \piso.data_r [2778] : 
                      (N203)? \piso.data_r [2810] : 
                      (N205)? \piso.data_r [2842] : 
                      (N207)? \piso.data_r [2874] : 
                      (N209)? \piso.data_r [2906] : 
                      (N211)? \piso.data_r [2938] : 
                      (N213)? \piso.data_r [2970] : 
                      (N215)? \piso.data_r [3002] : 
                      (N217)? \piso.data_r [3034] : 
                      (N219)? \piso.data_r [3066] : 
                      (N221)? \piso.data_r [3098] : 
                      (N223)? \piso.data_r [3130] : 
                      (N225)? \piso.data_r [3162] : 
                      (N227)? \piso.data_r [3194] : 
                      (N229)? \piso.data_r [3226] : 
                      (N231)? \piso.data_r [3258] : 
                      (N233)? \piso.data_r [3290] : 
                      (N235)? \piso.data_r [3322] : 
                      (N237)? \piso.data_r [3354] : 
                      (N239)? \piso.data_r [3386] : 
                      (N241)? \piso.data_r [3418] : 
                      (N243)? \piso.data_r [3450] : 
                      (N245)? \piso.data_r [3482] : 
                      (N247)? \piso.data_r [3514] : 
                      (N249)? \piso.data_r [3546] : 
                      (N251)? \piso.data_r [3578] : 
                      (N253)? \piso.data_r [3610] : 
                      (N255)? \piso.data_r [3642] : 
                      (N257)? \piso.data_r [3674] : 
                      (N259)? \piso.data_r [3706] : 
                      (N261)? \piso.data_r [3738] : 
                      (N263)? \piso.data_r [3770] : 
                      (N265)? \piso.data_r [3802] : 
                      (N267)? \piso.data_r [3834] : 
                      (N269)? \piso.data_r [3866] : 
                      (N271)? \piso.data_r [3898] : 
                      (N273)? \piso.data_r [3930] : 
                      (N275)? \piso.data_r [3962] : 
                      (N277)? \piso.data_r [3994] : 
                      (N279)? \piso.data_r [4026] : 
                      (N281)? \piso.data_r [4058] : 
                      (N283)? \piso.data_r [4090] : 1'b0;
  assign data_o[25] = (N156)? \piso.data_r [25] : 
                      (N158)? \piso.data_r [57] : 
                      (N160)? \piso.data_r [89] : 
                      (N162)? \piso.data_r [121] : 
                      (N164)? \piso.data_r [153] : 
                      (N166)? \piso.data_r [185] : 
                      (N168)? \piso.data_r [217] : 
                      (N170)? \piso.data_r [249] : 
                      (N172)? \piso.data_r [281] : 
                      (N174)? \piso.data_r [313] : 
                      (N176)? \piso.data_r [345] : 
                      (N178)? \piso.data_r [377] : 
                      (N180)? \piso.data_r [409] : 
                      (N182)? \piso.data_r [441] : 
                      (N184)? \piso.data_r [473] : 
                      (N186)? \piso.data_r [505] : 
                      (N188)? \piso.data_r [537] : 
                      (N190)? \piso.data_r [569] : 
                      (N192)? \piso.data_r [601] : 
                      (N194)? \piso.data_r [633] : 
                      (N196)? \piso.data_r [665] : 
                      (N198)? \piso.data_r [697] : 
                      (N200)? \piso.data_r [729] : 
                      (N202)? \piso.data_r [761] : 
                      (N204)? \piso.data_r [793] : 
                      (N206)? \piso.data_r [825] : 
                      (N208)? \piso.data_r [857] : 
                      (N210)? \piso.data_r [889] : 
                      (N212)? \piso.data_r [921] : 
                      (N214)? \piso.data_r [953] : 
                      (N216)? \piso.data_r [985] : 
                      (N218)? \piso.data_r [1017] : 
                      (N220)? \piso.data_r [1049] : 
                      (N222)? \piso.data_r [1081] : 
                      (N224)? \piso.data_r [1113] : 
                      (N226)? \piso.data_r [1145] : 
                      (N228)? \piso.data_r [1177] : 
                      (N230)? \piso.data_r [1209] : 
                      (N232)? \piso.data_r [1241] : 
                      (N234)? \piso.data_r [1273] : 
                      (N236)? \piso.data_r [1305] : 
                      (N238)? \piso.data_r [1337] : 
                      (N240)? \piso.data_r [1369] : 
                      (N242)? \piso.data_r [1401] : 
                      (N244)? \piso.data_r [1433] : 
                      (N246)? \piso.data_r [1465] : 
                      (N248)? \piso.data_r [1497] : 
                      (N250)? \piso.data_r [1529] : 
                      (N252)? \piso.data_r [1561] : 
                      (N254)? \piso.data_r [1593] : 
                      (N256)? \piso.data_r [1625] : 
                      (N258)? \piso.data_r [1657] : 
                      (N260)? \piso.data_r [1689] : 
                      (N262)? \piso.data_r [1721] : 
                      (N264)? \piso.data_r [1753] : 
                      (N266)? \piso.data_r [1785] : 
                      (N268)? \piso.data_r [1817] : 
                      (N270)? \piso.data_r [1849] : 
                      (N272)? \piso.data_r [1881] : 
                      (N274)? \piso.data_r [1913] : 
                      (N276)? \piso.data_r [1945] : 
                      (N278)? \piso.data_r [1977] : 
                      (N280)? \piso.data_r [2009] : 
                      (N282)? \piso.data_r [2041] : 
                      (N157)? \piso.data_r [2073] : 
                      (N159)? \piso.data_r [2105] : 
                      (N161)? \piso.data_r [2137] : 
                      (N163)? \piso.data_r [2169] : 
                      (N165)? \piso.data_r [2201] : 
                      (N167)? \piso.data_r [2233] : 
                      (N169)? \piso.data_r [2265] : 
                      (N171)? \piso.data_r [2297] : 
                      (N173)? \piso.data_r [2329] : 
                      (N175)? \piso.data_r [2361] : 
                      (N177)? \piso.data_r [2393] : 
                      (N179)? \piso.data_r [2425] : 
                      (N181)? \piso.data_r [2457] : 
                      (N183)? \piso.data_r [2489] : 
                      (N185)? \piso.data_r [2521] : 
                      (N187)? \piso.data_r [2553] : 
                      (N189)? \piso.data_r [2585] : 
                      (N191)? \piso.data_r [2617] : 
                      (N193)? \piso.data_r [2649] : 
                      (N195)? \piso.data_r [2681] : 
                      (N197)? \piso.data_r [2713] : 
                      (N199)? \piso.data_r [2745] : 
                      (N201)? \piso.data_r [2777] : 
                      (N203)? \piso.data_r [2809] : 
                      (N205)? \piso.data_r [2841] : 
                      (N207)? \piso.data_r [2873] : 
                      (N209)? \piso.data_r [2905] : 
                      (N211)? \piso.data_r [2937] : 
                      (N213)? \piso.data_r [2969] : 
                      (N215)? \piso.data_r [3001] : 
                      (N217)? \piso.data_r [3033] : 
                      (N219)? \piso.data_r [3065] : 
                      (N221)? \piso.data_r [3097] : 
                      (N223)? \piso.data_r [3129] : 
                      (N225)? \piso.data_r [3161] : 
                      (N227)? \piso.data_r [3193] : 
                      (N229)? \piso.data_r [3225] : 
                      (N231)? \piso.data_r [3257] : 
                      (N233)? \piso.data_r [3289] : 
                      (N235)? \piso.data_r [3321] : 
                      (N237)? \piso.data_r [3353] : 
                      (N239)? \piso.data_r [3385] : 
                      (N241)? \piso.data_r [3417] : 
                      (N243)? \piso.data_r [3449] : 
                      (N245)? \piso.data_r [3481] : 
                      (N247)? \piso.data_r [3513] : 
                      (N249)? \piso.data_r [3545] : 
                      (N251)? \piso.data_r [3577] : 
                      (N253)? \piso.data_r [3609] : 
                      (N255)? \piso.data_r [3641] : 
                      (N257)? \piso.data_r [3673] : 
                      (N259)? \piso.data_r [3705] : 
                      (N261)? \piso.data_r [3737] : 
                      (N263)? \piso.data_r [3769] : 
                      (N265)? \piso.data_r [3801] : 
                      (N267)? \piso.data_r [3833] : 
                      (N269)? \piso.data_r [3865] : 
                      (N271)? \piso.data_r [3897] : 
                      (N273)? \piso.data_r [3929] : 
                      (N275)? \piso.data_r [3961] : 
                      (N277)? \piso.data_r [3993] : 
                      (N279)? \piso.data_r [4025] : 
                      (N281)? \piso.data_r [4057] : 
                      (N283)? \piso.data_r [4089] : 1'b0;
  assign data_o[24] = (N156)? \piso.data_r [24] : 
                      (N158)? \piso.data_r [56] : 
                      (N160)? \piso.data_r [88] : 
                      (N162)? \piso.data_r [120] : 
                      (N164)? \piso.data_r [152] : 
                      (N166)? \piso.data_r [184] : 
                      (N168)? \piso.data_r [216] : 
                      (N170)? \piso.data_r [248] : 
                      (N172)? \piso.data_r [280] : 
                      (N174)? \piso.data_r [312] : 
                      (N176)? \piso.data_r [344] : 
                      (N178)? \piso.data_r [376] : 
                      (N180)? \piso.data_r [408] : 
                      (N182)? \piso.data_r [440] : 
                      (N184)? \piso.data_r [472] : 
                      (N186)? \piso.data_r [504] : 
                      (N188)? \piso.data_r [536] : 
                      (N190)? \piso.data_r [568] : 
                      (N192)? \piso.data_r [600] : 
                      (N194)? \piso.data_r [632] : 
                      (N196)? \piso.data_r [664] : 
                      (N198)? \piso.data_r [696] : 
                      (N200)? \piso.data_r [728] : 
                      (N202)? \piso.data_r [760] : 
                      (N204)? \piso.data_r [792] : 
                      (N206)? \piso.data_r [824] : 
                      (N208)? \piso.data_r [856] : 
                      (N210)? \piso.data_r [888] : 
                      (N212)? \piso.data_r [920] : 
                      (N214)? \piso.data_r [952] : 
                      (N216)? \piso.data_r [984] : 
                      (N218)? \piso.data_r [1016] : 
                      (N220)? \piso.data_r [1048] : 
                      (N222)? \piso.data_r [1080] : 
                      (N224)? \piso.data_r [1112] : 
                      (N226)? \piso.data_r [1144] : 
                      (N228)? \piso.data_r [1176] : 
                      (N230)? \piso.data_r [1208] : 
                      (N232)? \piso.data_r [1240] : 
                      (N234)? \piso.data_r [1272] : 
                      (N236)? \piso.data_r [1304] : 
                      (N238)? \piso.data_r [1336] : 
                      (N240)? \piso.data_r [1368] : 
                      (N242)? \piso.data_r [1400] : 
                      (N244)? \piso.data_r [1432] : 
                      (N246)? \piso.data_r [1464] : 
                      (N248)? \piso.data_r [1496] : 
                      (N250)? \piso.data_r [1528] : 
                      (N252)? \piso.data_r [1560] : 
                      (N254)? \piso.data_r [1592] : 
                      (N256)? \piso.data_r [1624] : 
                      (N258)? \piso.data_r [1656] : 
                      (N260)? \piso.data_r [1688] : 
                      (N262)? \piso.data_r [1720] : 
                      (N264)? \piso.data_r [1752] : 
                      (N266)? \piso.data_r [1784] : 
                      (N268)? \piso.data_r [1816] : 
                      (N270)? \piso.data_r [1848] : 
                      (N272)? \piso.data_r [1880] : 
                      (N274)? \piso.data_r [1912] : 
                      (N276)? \piso.data_r [1944] : 
                      (N278)? \piso.data_r [1976] : 
                      (N280)? \piso.data_r [2008] : 
                      (N282)? \piso.data_r [2040] : 
                      (N157)? \piso.data_r [2072] : 
                      (N159)? \piso.data_r [2104] : 
                      (N161)? \piso.data_r [2136] : 
                      (N163)? \piso.data_r [2168] : 
                      (N165)? \piso.data_r [2200] : 
                      (N167)? \piso.data_r [2232] : 
                      (N169)? \piso.data_r [2264] : 
                      (N171)? \piso.data_r [2296] : 
                      (N173)? \piso.data_r [2328] : 
                      (N175)? \piso.data_r [2360] : 
                      (N177)? \piso.data_r [2392] : 
                      (N179)? \piso.data_r [2424] : 
                      (N181)? \piso.data_r [2456] : 
                      (N183)? \piso.data_r [2488] : 
                      (N185)? \piso.data_r [2520] : 
                      (N187)? \piso.data_r [2552] : 
                      (N189)? \piso.data_r [2584] : 
                      (N191)? \piso.data_r [2616] : 
                      (N193)? \piso.data_r [2648] : 
                      (N195)? \piso.data_r [2680] : 
                      (N197)? \piso.data_r [2712] : 
                      (N199)? \piso.data_r [2744] : 
                      (N201)? \piso.data_r [2776] : 
                      (N203)? \piso.data_r [2808] : 
                      (N205)? \piso.data_r [2840] : 
                      (N207)? \piso.data_r [2872] : 
                      (N209)? \piso.data_r [2904] : 
                      (N211)? \piso.data_r [2936] : 
                      (N213)? \piso.data_r [2968] : 
                      (N215)? \piso.data_r [3000] : 
                      (N217)? \piso.data_r [3032] : 
                      (N219)? \piso.data_r [3064] : 
                      (N221)? \piso.data_r [3096] : 
                      (N223)? \piso.data_r [3128] : 
                      (N225)? \piso.data_r [3160] : 
                      (N227)? \piso.data_r [3192] : 
                      (N229)? \piso.data_r [3224] : 
                      (N231)? \piso.data_r [3256] : 
                      (N233)? \piso.data_r [3288] : 
                      (N235)? \piso.data_r [3320] : 
                      (N237)? \piso.data_r [3352] : 
                      (N239)? \piso.data_r [3384] : 
                      (N241)? \piso.data_r [3416] : 
                      (N243)? \piso.data_r [3448] : 
                      (N245)? \piso.data_r [3480] : 
                      (N247)? \piso.data_r [3512] : 
                      (N249)? \piso.data_r [3544] : 
                      (N251)? \piso.data_r [3576] : 
                      (N253)? \piso.data_r [3608] : 
                      (N255)? \piso.data_r [3640] : 
                      (N257)? \piso.data_r [3672] : 
                      (N259)? \piso.data_r [3704] : 
                      (N261)? \piso.data_r [3736] : 
                      (N263)? \piso.data_r [3768] : 
                      (N265)? \piso.data_r [3800] : 
                      (N267)? \piso.data_r [3832] : 
                      (N269)? \piso.data_r [3864] : 
                      (N271)? \piso.data_r [3896] : 
                      (N273)? \piso.data_r [3928] : 
                      (N275)? \piso.data_r [3960] : 
                      (N277)? \piso.data_r [3992] : 
                      (N279)? \piso.data_r [4024] : 
                      (N281)? \piso.data_r [4056] : 
                      (N283)? \piso.data_r [4088] : 1'b0;
  assign data_o[23] = (N156)? \piso.data_r [23] : 
                      (N158)? \piso.data_r [55] : 
                      (N160)? \piso.data_r [87] : 
                      (N162)? \piso.data_r [119] : 
                      (N164)? \piso.data_r [151] : 
                      (N166)? \piso.data_r [183] : 
                      (N168)? \piso.data_r [215] : 
                      (N170)? \piso.data_r [247] : 
                      (N172)? \piso.data_r [279] : 
                      (N174)? \piso.data_r [311] : 
                      (N176)? \piso.data_r [343] : 
                      (N178)? \piso.data_r [375] : 
                      (N180)? \piso.data_r [407] : 
                      (N182)? \piso.data_r [439] : 
                      (N184)? \piso.data_r [471] : 
                      (N186)? \piso.data_r [503] : 
                      (N188)? \piso.data_r [535] : 
                      (N190)? \piso.data_r [567] : 
                      (N192)? \piso.data_r [599] : 
                      (N194)? \piso.data_r [631] : 
                      (N196)? \piso.data_r [663] : 
                      (N198)? \piso.data_r [695] : 
                      (N200)? \piso.data_r [727] : 
                      (N202)? \piso.data_r [759] : 
                      (N204)? \piso.data_r [791] : 
                      (N206)? \piso.data_r [823] : 
                      (N208)? \piso.data_r [855] : 
                      (N210)? \piso.data_r [887] : 
                      (N212)? \piso.data_r [919] : 
                      (N214)? \piso.data_r [951] : 
                      (N216)? \piso.data_r [983] : 
                      (N218)? \piso.data_r [1015] : 
                      (N220)? \piso.data_r [1047] : 
                      (N222)? \piso.data_r [1079] : 
                      (N224)? \piso.data_r [1111] : 
                      (N226)? \piso.data_r [1143] : 
                      (N228)? \piso.data_r [1175] : 
                      (N230)? \piso.data_r [1207] : 
                      (N232)? \piso.data_r [1239] : 
                      (N234)? \piso.data_r [1271] : 
                      (N236)? \piso.data_r [1303] : 
                      (N238)? \piso.data_r [1335] : 
                      (N240)? \piso.data_r [1367] : 
                      (N242)? \piso.data_r [1399] : 
                      (N244)? \piso.data_r [1431] : 
                      (N246)? \piso.data_r [1463] : 
                      (N248)? \piso.data_r [1495] : 
                      (N250)? \piso.data_r [1527] : 
                      (N252)? \piso.data_r [1559] : 
                      (N254)? \piso.data_r [1591] : 
                      (N256)? \piso.data_r [1623] : 
                      (N258)? \piso.data_r [1655] : 
                      (N260)? \piso.data_r [1687] : 
                      (N262)? \piso.data_r [1719] : 
                      (N264)? \piso.data_r [1751] : 
                      (N266)? \piso.data_r [1783] : 
                      (N268)? \piso.data_r [1815] : 
                      (N270)? \piso.data_r [1847] : 
                      (N272)? \piso.data_r [1879] : 
                      (N274)? \piso.data_r [1911] : 
                      (N276)? \piso.data_r [1943] : 
                      (N278)? \piso.data_r [1975] : 
                      (N280)? \piso.data_r [2007] : 
                      (N282)? \piso.data_r [2039] : 
                      (N157)? \piso.data_r [2071] : 
                      (N159)? \piso.data_r [2103] : 
                      (N161)? \piso.data_r [2135] : 
                      (N163)? \piso.data_r [2167] : 
                      (N165)? \piso.data_r [2199] : 
                      (N167)? \piso.data_r [2231] : 
                      (N169)? \piso.data_r [2263] : 
                      (N171)? \piso.data_r [2295] : 
                      (N173)? \piso.data_r [2327] : 
                      (N175)? \piso.data_r [2359] : 
                      (N177)? \piso.data_r [2391] : 
                      (N179)? \piso.data_r [2423] : 
                      (N181)? \piso.data_r [2455] : 
                      (N183)? \piso.data_r [2487] : 
                      (N185)? \piso.data_r [2519] : 
                      (N187)? \piso.data_r [2551] : 
                      (N189)? \piso.data_r [2583] : 
                      (N191)? \piso.data_r [2615] : 
                      (N193)? \piso.data_r [2647] : 
                      (N195)? \piso.data_r [2679] : 
                      (N197)? \piso.data_r [2711] : 
                      (N199)? \piso.data_r [2743] : 
                      (N201)? \piso.data_r [2775] : 
                      (N203)? \piso.data_r [2807] : 
                      (N205)? \piso.data_r [2839] : 
                      (N207)? \piso.data_r [2871] : 
                      (N209)? \piso.data_r [2903] : 
                      (N211)? \piso.data_r [2935] : 
                      (N213)? \piso.data_r [2967] : 
                      (N215)? \piso.data_r [2999] : 
                      (N217)? \piso.data_r [3031] : 
                      (N219)? \piso.data_r [3063] : 
                      (N221)? \piso.data_r [3095] : 
                      (N223)? \piso.data_r [3127] : 
                      (N225)? \piso.data_r [3159] : 
                      (N227)? \piso.data_r [3191] : 
                      (N229)? \piso.data_r [3223] : 
                      (N231)? \piso.data_r [3255] : 
                      (N233)? \piso.data_r [3287] : 
                      (N235)? \piso.data_r [3319] : 
                      (N237)? \piso.data_r [3351] : 
                      (N239)? \piso.data_r [3383] : 
                      (N241)? \piso.data_r [3415] : 
                      (N243)? \piso.data_r [3447] : 
                      (N245)? \piso.data_r [3479] : 
                      (N247)? \piso.data_r [3511] : 
                      (N249)? \piso.data_r [3543] : 
                      (N251)? \piso.data_r [3575] : 
                      (N253)? \piso.data_r [3607] : 
                      (N255)? \piso.data_r [3639] : 
                      (N257)? \piso.data_r [3671] : 
                      (N259)? \piso.data_r [3703] : 
                      (N261)? \piso.data_r [3735] : 
                      (N263)? \piso.data_r [3767] : 
                      (N265)? \piso.data_r [3799] : 
                      (N267)? \piso.data_r [3831] : 
                      (N269)? \piso.data_r [3863] : 
                      (N271)? \piso.data_r [3895] : 
                      (N273)? \piso.data_r [3927] : 
                      (N275)? \piso.data_r [3959] : 
                      (N277)? \piso.data_r [3991] : 
                      (N279)? \piso.data_r [4023] : 
                      (N281)? \piso.data_r [4055] : 
                      (N283)? \piso.data_r [4087] : 1'b0;
  assign data_o[22] = (N156)? \piso.data_r [22] : 
                      (N158)? \piso.data_r [54] : 
                      (N160)? \piso.data_r [86] : 
                      (N162)? \piso.data_r [118] : 
                      (N164)? \piso.data_r [150] : 
                      (N166)? \piso.data_r [182] : 
                      (N168)? \piso.data_r [214] : 
                      (N170)? \piso.data_r [246] : 
                      (N172)? \piso.data_r [278] : 
                      (N174)? \piso.data_r [310] : 
                      (N176)? \piso.data_r [342] : 
                      (N178)? \piso.data_r [374] : 
                      (N180)? \piso.data_r [406] : 
                      (N182)? \piso.data_r [438] : 
                      (N184)? \piso.data_r [470] : 
                      (N186)? \piso.data_r [502] : 
                      (N188)? \piso.data_r [534] : 
                      (N190)? \piso.data_r [566] : 
                      (N192)? \piso.data_r [598] : 
                      (N194)? \piso.data_r [630] : 
                      (N196)? \piso.data_r [662] : 
                      (N198)? \piso.data_r [694] : 
                      (N200)? \piso.data_r [726] : 
                      (N202)? \piso.data_r [758] : 
                      (N204)? \piso.data_r [790] : 
                      (N206)? \piso.data_r [822] : 
                      (N208)? \piso.data_r [854] : 
                      (N210)? \piso.data_r [886] : 
                      (N212)? \piso.data_r [918] : 
                      (N214)? \piso.data_r [950] : 
                      (N216)? \piso.data_r [982] : 
                      (N218)? \piso.data_r [1014] : 
                      (N220)? \piso.data_r [1046] : 
                      (N222)? \piso.data_r [1078] : 
                      (N224)? \piso.data_r [1110] : 
                      (N226)? \piso.data_r [1142] : 
                      (N228)? \piso.data_r [1174] : 
                      (N230)? \piso.data_r [1206] : 
                      (N232)? \piso.data_r [1238] : 
                      (N234)? \piso.data_r [1270] : 
                      (N236)? \piso.data_r [1302] : 
                      (N238)? \piso.data_r [1334] : 
                      (N240)? \piso.data_r [1366] : 
                      (N242)? \piso.data_r [1398] : 
                      (N244)? \piso.data_r [1430] : 
                      (N246)? \piso.data_r [1462] : 
                      (N248)? \piso.data_r [1494] : 
                      (N250)? \piso.data_r [1526] : 
                      (N252)? \piso.data_r [1558] : 
                      (N254)? \piso.data_r [1590] : 
                      (N256)? \piso.data_r [1622] : 
                      (N258)? \piso.data_r [1654] : 
                      (N260)? \piso.data_r [1686] : 
                      (N262)? \piso.data_r [1718] : 
                      (N264)? \piso.data_r [1750] : 
                      (N266)? \piso.data_r [1782] : 
                      (N268)? \piso.data_r [1814] : 
                      (N270)? \piso.data_r [1846] : 
                      (N272)? \piso.data_r [1878] : 
                      (N274)? \piso.data_r [1910] : 
                      (N276)? \piso.data_r [1942] : 
                      (N278)? \piso.data_r [1974] : 
                      (N280)? \piso.data_r [2006] : 
                      (N282)? \piso.data_r [2038] : 
                      (N157)? \piso.data_r [2070] : 
                      (N159)? \piso.data_r [2102] : 
                      (N161)? \piso.data_r [2134] : 
                      (N163)? \piso.data_r [2166] : 
                      (N165)? \piso.data_r [2198] : 
                      (N167)? \piso.data_r [2230] : 
                      (N169)? \piso.data_r [2262] : 
                      (N171)? \piso.data_r [2294] : 
                      (N173)? \piso.data_r [2326] : 
                      (N175)? \piso.data_r [2358] : 
                      (N177)? \piso.data_r [2390] : 
                      (N179)? \piso.data_r [2422] : 
                      (N181)? \piso.data_r [2454] : 
                      (N183)? \piso.data_r [2486] : 
                      (N185)? \piso.data_r [2518] : 
                      (N187)? \piso.data_r [2550] : 
                      (N189)? \piso.data_r [2582] : 
                      (N191)? \piso.data_r [2614] : 
                      (N193)? \piso.data_r [2646] : 
                      (N195)? \piso.data_r [2678] : 
                      (N197)? \piso.data_r [2710] : 
                      (N199)? \piso.data_r [2742] : 
                      (N201)? \piso.data_r [2774] : 
                      (N203)? \piso.data_r [2806] : 
                      (N205)? \piso.data_r [2838] : 
                      (N207)? \piso.data_r [2870] : 
                      (N209)? \piso.data_r [2902] : 
                      (N211)? \piso.data_r [2934] : 
                      (N213)? \piso.data_r [2966] : 
                      (N215)? \piso.data_r [2998] : 
                      (N217)? \piso.data_r [3030] : 
                      (N219)? \piso.data_r [3062] : 
                      (N221)? \piso.data_r [3094] : 
                      (N223)? \piso.data_r [3126] : 
                      (N225)? \piso.data_r [3158] : 
                      (N227)? \piso.data_r [3190] : 
                      (N229)? \piso.data_r [3222] : 
                      (N231)? \piso.data_r [3254] : 
                      (N233)? \piso.data_r [3286] : 
                      (N235)? \piso.data_r [3318] : 
                      (N237)? \piso.data_r [3350] : 
                      (N239)? \piso.data_r [3382] : 
                      (N241)? \piso.data_r [3414] : 
                      (N243)? \piso.data_r [3446] : 
                      (N245)? \piso.data_r [3478] : 
                      (N247)? \piso.data_r [3510] : 
                      (N249)? \piso.data_r [3542] : 
                      (N251)? \piso.data_r [3574] : 
                      (N253)? \piso.data_r [3606] : 
                      (N255)? \piso.data_r [3638] : 
                      (N257)? \piso.data_r [3670] : 
                      (N259)? \piso.data_r [3702] : 
                      (N261)? \piso.data_r [3734] : 
                      (N263)? \piso.data_r [3766] : 
                      (N265)? \piso.data_r [3798] : 
                      (N267)? \piso.data_r [3830] : 
                      (N269)? \piso.data_r [3862] : 
                      (N271)? \piso.data_r [3894] : 
                      (N273)? \piso.data_r [3926] : 
                      (N275)? \piso.data_r [3958] : 
                      (N277)? \piso.data_r [3990] : 
                      (N279)? \piso.data_r [4022] : 
                      (N281)? \piso.data_r [4054] : 
                      (N283)? \piso.data_r [4086] : 1'b0;
  assign data_o[21] = (N156)? \piso.data_r [21] : 
                      (N158)? \piso.data_r [53] : 
                      (N160)? \piso.data_r [85] : 
                      (N162)? \piso.data_r [117] : 
                      (N164)? \piso.data_r [149] : 
                      (N166)? \piso.data_r [181] : 
                      (N168)? \piso.data_r [213] : 
                      (N170)? \piso.data_r [245] : 
                      (N172)? \piso.data_r [277] : 
                      (N174)? \piso.data_r [309] : 
                      (N176)? \piso.data_r [341] : 
                      (N178)? \piso.data_r [373] : 
                      (N180)? \piso.data_r [405] : 
                      (N182)? \piso.data_r [437] : 
                      (N184)? \piso.data_r [469] : 
                      (N186)? \piso.data_r [501] : 
                      (N188)? \piso.data_r [533] : 
                      (N190)? \piso.data_r [565] : 
                      (N192)? \piso.data_r [597] : 
                      (N194)? \piso.data_r [629] : 
                      (N196)? \piso.data_r [661] : 
                      (N198)? \piso.data_r [693] : 
                      (N200)? \piso.data_r [725] : 
                      (N202)? \piso.data_r [757] : 
                      (N204)? \piso.data_r [789] : 
                      (N206)? \piso.data_r [821] : 
                      (N208)? \piso.data_r [853] : 
                      (N210)? \piso.data_r [885] : 
                      (N212)? \piso.data_r [917] : 
                      (N214)? \piso.data_r [949] : 
                      (N216)? \piso.data_r [981] : 
                      (N218)? \piso.data_r [1013] : 
                      (N220)? \piso.data_r [1045] : 
                      (N222)? \piso.data_r [1077] : 
                      (N224)? \piso.data_r [1109] : 
                      (N226)? \piso.data_r [1141] : 
                      (N228)? \piso.data_r [1173] : 
                      (N230)? \piso.data_r [1205] : 
                      (N232)? \piso.data_r [1237] : 
                      (N234)? \piso.data_r [1269] : 
                      (N236)? \piso.data_r [1301] : 
                      (N238)? \piso.data_r [1333] : 
                      (N240)? \piso.data_r [1365] : 
                      (N242)? \piso.data_r [1397] : 
                      (N244)? \piso.data_r [1429] : 
                      (N246)? \piso.data_r [1461] : 
                      (N248)? \piso.data_r [1493] : 
                      (N250)? \piso.data_r [1525] : 
                      (N252)? \piso.data_r [1557] : 
                      (N254)? \piso.data_r [1589] : 
                      (N256)? \piso.data_r [1621] : 
                      (N258)? \piso.data_r [1653] : 
                      (N260)? \piso.data_r [1685] : 
                      (N262)? \piso.data_r [1717] : 
                      (N264)? \piso.data_r [1749] : 
                      (N266)? \piso.data_r [1781] : 
                      (N268)? \piso.data_r [1813] : 
                      (N270)? \piso.data_r [1845] : 
                      (N272)? \piso.data_r [1877] : 
                      (N274)? \piso.data_r [1909] : 
                      (N276)? \piso.data_r [1941] : 
                      (N278)? \piso.data_r [1973] : 
                      (N280)? \piso.data_r [2005] : 
                      (N282)? \piso.data_r [2037] : 
                      (N157)? \piso.data_r [2069] : 
                      (N159)? \piso.data_r [2101] : 
                      (N161)? \piso.data_r [2133] : 
                      (N163)? \piso.data_r [2165] : 
                      (N165)? \piso.data_r [2197] : 
                      (N167)? \piso.data_r [2229] : 
                      (N169)? \piso.data_r [2261] : 
                      (N171)? \piso.data_r [2293] : 
                      (N173)? \piso.data_r [2325] : 
                      (N175)? \piso.data_r [2357] : 
                      (N177)? \piso.data_r [2389] : 
                      (N179)? \piso.data_r [2421] : 
                      (N181)? \piso.data_r [2453] : 
                      (N183)? \piso.data_r [2485] : 
                      (N185)? \piso.data_r [2517] : 
                      (N187)? \piso.data_r [2549] : 
                      (N189)? \piso.data_r [2581] : 
                      (N191)? \piso.data_r [2613] : 
                      (N193)? \piso.data_r [2645] : 
                      (N195)? \piso.data_r [2677] : 
                      (N197)? \piso.data_r [2709] : 
                      (N199)? \piso.data_r [2741] : 
                      (N201)? \piso.data_r [2773] : 
                      (N203)? \piso.data_r [2805] : 
                      (N205)? \piso.data_r [2837] : 
                      (N207)? \piso.data_r [2869] : 
                      (N209)? \piso.data_r [2901] : 
                      (N211)? \piso.data_r [2933] : 
                      (N213)? \piso.data_r [2965] : 
                      (N215)? \piso.data_r [2997] : 
                      (N217)? \piso.data_r [3029] : 
                      (N219)? \piso.data_r [3061] : 
                      (N221)? \piso.data_r [3093] : 
                      (N223)? \piso.data_r [3125] : 
                      (N225)? \piso.data_r [3157] : 
                      (N227)? \piso.data_r [3189] : 
                      (N229)? \piso.data_r [3221] : 
                      (N231)? \piso.data_r [3253] : 
                      (N233)? \piso.data_r [3285] : 
                      (N235)? \piso.data_r [3317] : 
                      (N237)? \piso.data_r [3349] : 
                      (N239)? \piso.data_r [3381] : 
                      (N241)? \piso.data_r [3413] : 
                      (N243)? \piso.data_r [3445] : 
                      (N245)? \piso.data_r [3477] : 
                      (N247)? \piso.data_r [3509] : 
                      (N249)? \piso.data_r [3541] : 
                      (N251)? \piso.data_r [3573] : 
                      (N253)? \piso.data_r [3605] : 
                      (N255)? \piso.data_r [3637] : 
                      (N257)? \piso.data_r [3669] : 
                      (N259)? \piso.data_r [3701] : 
                      (N261)? \piso.data_r [3733] : 
                      (N263)? \piso.data_r [3765] : 
                      (N265)? \piso.data_r [3797] : 
                      (N267)? \piso.data_r [3829] : 
                      (N269)? \piso.data_r [3861] : 
                      (N271)? \piso.data_r [3893] : 
                      (N273)? \piso.data_r [3925] : 
                      (N275)? \piso.data_r [3957] : 
                      (N277)? \piso.data_r [3989] : 
                      (N279)? \piso.data_r [4021] : 
                      (N281)? \piso.data_r [4053] : 
                      (N283)? \piso.data_r [4085] : 1'b0;
  assign data_o[20] = (N156)? \piso.data_r [20] : 
                      (N158)? \piso.data_r [52] : 
                      (N160)? \piso.data_r [84] : 
                      (N162)? \piso.data_r [116] : 
                      (N164)? \piso.data_r [148] : 
                      (N166)? \piso.data_r [180] : 
                      (N168)? \piso.data_r [212] : 
                      (N170)? \piso.data_r [244] : 
                      (N172)? \piso.data_r [276] : 
                      (N174)? \piso.data_r [308] : 
                      (N176)? \piso.data_r [340] : 
                      (N178)? \piso.data_r [372] : 
                      (N180)? \piso.data_r [404] : 
                      (N182)? \piso.data_r [436] : 
                      (N184)? \piso.data_r [468] : 
                      (N186)? \piso.data_r [500] : 
                      (N188)? \piso.data_r [532] : 
                      (N190)? \piso.data_r [564] : 
                      (N192)? \piso.data_r [596] : 
                      (N194)? \piso.data_r [628] : 
                      (N196)? \piso.data_r [660] : 
                      (N198)? \piso.data_r [692] : 
                      (N200)? \piso.data_r [724] : 
                      (N202)? \piso.data_r [756] : 
                      (N204)? \piso.data_r [788] : 
                      (N206)? \piso.data_r [820] : 
                      (N208)? \piso.data_r [852] : 
                      (N210)? \piso.data_r [884] : 
                      (N212)? \piso.data_r [916] : 
                      (N214)? \piso.data_r [948] : 
                      (N216)? \piso.data_r [980] : 
                      (N218)? \piso.data_r [1012] : 
                      (N220)? \piso.data_r [1044] : 
                      (N222)? \piso.data_r [1076] : 
                      (N224)? \piso.data_r [1108] : 
                      (N226)? \piso.data_r [1140] : 
                      (N228)? \piso.data_r [1172] : 
                      (N230)? \piso.data_r [1204] : 
                      (N232)? \piso.data_r [1236] : 
                      (N234)? \piso.data_r [1268] : 
                      (N236)? \piso.data_r [1300] : 
                      (N238)? \piso.data_r [1332] : 
                      (N240)? \piso.data_r [1364] : 
                      (N242)? \piso.data_r [1396] : 
                      (N244)? \piso.data_r [1428] : 
                      (N246)? \piso.data_r [1460] : 
                      (N248)? \piso.data_r [1492] : 
                      (N250)? \piso.data_r [1524] : 
                      (N252)? \piso.data_r [1556] : 
                      (N254)? \piso.data_r [1588] : 
                      (N256)? \piso.data_r [1620] : 
                      (N258)? \piso.data_r [1652] : 
                      (N260)? \piso.data_r [1684] : 
                      (N262)? \piso.data_r [1716] : 
                      (N264)? \piso.data_r [1748] : 
                      (N266)? \piso.data_r [1780] : 
                      (N268)? \piso.data_r [1812] : 
                      (N270)? \piso.data_r [1844] : 
                      (N272)? \piso.data_r [1876] : 
                      (N274)? \piso.data_r [1908] : 
                      (N276)? \piso.data_r [1940] : 
                      (N278)? \piso.data_r [1972] : 
                      (N280)? \piso.data_r [2004] : 
                      (N282)? \piso.data_r [2036] : 
                      (N157)? \piso.data_r [2068] : 
                      (N159)? \piso.data_r [2100] : 
                      (N161)? \piso.data_r [2132] : 
                      (N163)? \piso.data_r [2164] : 
                      (N165)? \piso.data_r [2196] : 
                      (N167)? \piso.data_r [2228] : 
                      (N169)? \piso.data_r [2260] : 
                      (N171)? \piso.data_r [2292] : 
                      (N173)? \piso.data_r [2324] : 
                      (N175)? \piso.data_r [2356] : 
                      (N177)? \piso.data_r [2388] : 
                      (N179)? \piso.data_r [2420] : 
                      (N181)? \piso.data_r [2452] : 
                      (N183)? \piso.data_r [2484] : 
                      (N185)? \piso.data_r [2516] : 
                      (N187)? \piso.data_r [2548] : 
                      (N189)? \piso.data_r [2580] : 
                      (N191)? \piso.data_r [2612] : 
                      (N193)? \piso.data_r [2644] : 
                      (N195)? \piso.data_r [2676] : 
                      (N197)? \piso.data_r [2708] : 
                      (N199)? \piso.data_r [2740] : 
                      (N201)? \piso.data_r [2772] : 
                      (N203)? \piso.data_r [2804] : 
                      (N205)? \piso.data_r [2836] : 
                      (N207)? \piso.data_r [2868] : 
                      (N209)? \piso.data_r [2900] : 
                      (N211)? \piso.data_r [2932] : 
                      (N213)? \piso.data_r [2964] : 
                      (N215)? \piso.data_r [2996] : 
                      (N217)? \piso.data_r [3028] : 
                      (N219)? \piso.data_r [3060] : 
                      (N221)? \piso.data_r [3092] : 
                      (N223)? \piso.data_r [3124] : 
                      (N225)? \piso.data_r [3156] : 
                      (N227)? \piso.data_r [3188] : 
                      (N229)? \piso.data_r [3220] : 
                      (N231)? \piso.data_r [3252] : 
                      (N233)? \piso.data_r [3284] : 
                      (N235)? \piso.data_r [3316] : 
                      (N237)? \piso.data_r [3348] : 
                      (N239)? \piso.data_r [3380] : 
                      (N241)? \piso.data_r [3412] : 
                      (N243)? \piso.data_r [3444] : 
                      (N245)? \piso.data_r [3476] : 
                      (N247)? \piso.data_r [3508] : 
                      (N249)? \piso.data_r [3540] : 
                      (N251)? \piso.data_r [3572] : 
                      (N253)? \piso.data_r [3604] : 
                      (N255)? \piso.data_r [3636] : 
                      (N257)? \piso.data_r [3668] : 
                      (N259)? \piso.data_r [3700] : 
                      (N261)? \piso.data_r [3732] : 
                      (N263)? \piso.data_r [3764] : 
                      (N265)? \piso.data_r [3796] : 
                      (N267)? \piso.data_r [3828] : 
                      (N269)? \piso.data_r [3860] : 
                      (N271)? \piso.data_r [3892] : 
                      (N273)? \piso.data_r [3924] : 
                      (N275)? \piso.data_r [3956] : 
                      (N277)? \piso.data_r [3988] : 
                      (N279)? \piso.data_r [4020] : 
                      (N281)? \piso.data_r [4052] : 
                      (N283)? \piso.data_r [4084] : 1'b0;
  assign data_o[19] = (N156)? \piso.data_r [19] : 
                      (N158)? \piso.data_r [51] : 
                      (N160)? \piso.data_r [83] : 
                      (N162)? \piso.data_r [115] : 
                      (N164)? \piso.data_r [147] : 
                      (N166)? \piso.data_r [179] : 
                      (N168)? \piso.data_r [211] : 
                      (N170)? \piso.data_r [243] : 
                      (N172)? \piso.data_r [275] : 
                      (N174)? \piso.data_r [307] : 
                      (N176)? \piso.data_r [339] : 
                      (N178)? \piso.data_r [371] : 
                      (N180)? \piso.data_r [403] : 
                      (N182)? \piso.data_r [435] : 
                      (N184)? \piso.data_r [467] : 
                      (N186)? \piso.data_r [499] : 
                      (N188)? \piso.data_r [531] : 
                      (N190)? \piso.data_r [563] : 
                      (N192)? \piso.data_r [595] : 
                      (N194)? \piso.data_r [627] : 
                      (N196)? \piso.data_r [659] : 
                      (N198)? \piso.data_r [691] : 
                      (N200)? \piso.data_r [723] : 
                      (N202)? \piso.data_r [755] : 
                      (N204)? \piso.data_r [787] : 
                      (N206)? \piso.data_r [819] : 
                      (N208)? \piso.data_r [851] : 
                      (N210)? \piso.data_r [883] : 
                      (N212)? \piso.data_r [915] : 
                      (N214)? \piso.data_r [947] : 
                      (N216)? \piso.data_r [979] : 
                      (N218)? \piso.data_r [1011] : 
                      (N220)? \piso.data_r [1043] : 
                      (N222)? \piso.data_r [1075] : 
                      (N224)? \piso.data_r [1107] : 
                      (N226)? \piso.data_r [1139] : 
                      (N228)? \piso.data_r [1171] : 
                      (N230)? \piso.data_r [1203] : 
                      (N232)? \piso.data_r [1235] : 
                      (N234)? \piso.data_r [1267] : 
                      (N236)? \piso.data_r [1299] : 
                      (N238)? \piso.data_r [1331] : 
                      (N240)? \piso.data_r [1363] : 
                      (N242)? \piso.data_r [1395] : 
                      (N244)? \piso.data_r [1427] : 
                      (N246)? \piso.data_r [1459] : 
                      (N248)? \piso.data_r [1491] : 
                      (N250)? \piso.data_r [1523] : 
                      (N252)? \piso.data_r [1555] : 
                      (N254)? \piso.data_r [1587] : 
                      (N256)? \piso.data_r [1619] : 
                      (N258)? \piso.data_r [1651] : 
                      (N260)? \piso.data_r [1683] : 
                      (N262)? \piso.data_r [1715] : 
                      (N264)? \piso.data_r [1747] : 
                      (N266)? \piso.data_r [1779] : 
                      (N268)? \piso.data_r [1811] : 
                      (N270)? \piso.data_r [1843] : 
                      (N272)? \piso.data_r [1875] : 
                      (N274)? \piso.data_r [1907] : 
                      (N276)? \piso.data_r [1939] : 
                      (N278)? \piso.data_r [1971] : 
                      (N280)? \piso.data_r [2003] : 
                      (N282)? \piso.data_r [2035] : 
                      (N157)? \piso.data_r [2067] : 
                      (N159)? \piso.data_r [2099] : 
                      (N161)? \piso.data_r [2131] : 
                      (N163)? \piso.data_r [2163] : 
                      (N165)? \piso.data_r [2195] : 
                      (N167)? \piso.data_r [2227] : 
                      (N169)? \piso.data_r [2259] : 
                      (N171)? \piso.data_r [2291] : 
                      (N173)? \piso.data_r [2323] : 
                      (N175)? \piso.data_r [2355] : 
                      (N177)? \piso.data_r [2387] : 
                      (N179)? \piso.data_r [2419] : 
                      (N181)? \piso.data_r [2451] : 
                      (N183)? \piso.data_r [2483] : 
                      (N185)? \piso.data_r [2515] : 
                      (N187)? \piso.data_r [2547] : 
                      (N189)? \piso.data_r [2579] : 
                      (N191)? \piso.data_r [2611] : 
                      (N193)? \piso.data_r [2643] : 
                      (N195)? \piso.data_r [2675] : 
                      (N197)? \piso.data_r [2707] : 
                      (N199)? \piso.data_r [2739] : 
                      (N201)? \piso.data_r [2771] : 
                      (N203)? \piso.data_r [2803] : 
                      (N205)? \piso.data_r [2835] : 
                      (N207)? \piso.data_r [2867] : 
                      (N209)? \piso.data_r [2899] : 
                      (N211)? \piso.data_r [2931] : 
                      (N213)? \piso.data_r [2963] : 
                      (N215)? \piso.data_r [2995] : 
                      (N217)? \piso.data_r [3027] : 
                      (N219)? \piso.data_r [3059] : 
                      (N221)? \piso.data_r [3091] : 
                      (N223)? \piso.data_r [3123] : 
                      (N225)? \piso.data_r [3155] : 
                      (N227)? \piso.data_r [3187] : 
                      (N229)? \piso.data_r [3219] : 
                      (N231)? \piso.data_r [3251] : 
                      (N233)? \piso.data_r [3283] : 
                      (N235)? \piso.data_r [3315] : 
                      (N237)? \piso.data_r [3347] : 
                      (N239)? \piso.data_r [3379] : 
                      (N241)? \piso.data_r [3411] : 
                      (N243)? \piso.data_r [3443] : 
                      (N245)? \piso.data_r [3475] : 
                      (N247)? \piso.data_r [3507] : 
                      (N249)? \piso.data_r [3539] : 
                      (N251)? \piso.data_r [3571] : 
                      (N253)? \piso.data_r [3603] : 
                      (N255)? \piso.data_r [3635] : 
                      (N257)? \piso.data_r [3667] : 
                      (N259)? \piso.data_r [3699] : 
                      (N261)? \piso.data_r [3731] : 
                      (N263)? \piso.data_r [3763] : 
                      (N265)? \piso.data_r [3795] : 
                      (N267)? \piso.data_r [3827] : 
                      (N269)? \piso.data_r [3859] : 
                      (N271)? \piso.data_r [3891] : 
                      (N273)? \piso.data_r [3923] : 
                      (N275)? \piso.data_r [3955] : 
                      (N277)? \piso.data_r [3987] : 
                      (N279)? \piso.data_r [4019] : 
                      (N281)? \piso.data_r [4051] : 
                      (N283)? \piso.data_r [4083] : 1'b0;
  assign data_o[18] = (N156)? \piso.data_r [18] : 
                      (N158)? \piso.data_r [50] : 
                      (N160)? \piso.data_r [82] : 
                      (N162)? \piso.data_r [114] : 
                      (N164)? \piso.data_r [146] : 
                      (N166)? \piso.data_r [178] : 
                      (N168)? \piso.data_r [210] : 
                      (N170)? \piso.data_r [242] : 
                      (N172)? \piso.data_r [274] : 
                      (N174)? \piso.data_r [306] : 
                      (N176)? \piso.data_r [338] : 
                      (N178)? \piso.data_r [370] : 
                      (N180)? \piso.data_r [402] : 
                      (N182)? \piso.data_r [434] : 
                      (N184)? \piso.data_r [466] : 
                      (N186)? \piso.data_r [498] : 
                      (N188)? \piso.data_r [530] : 
                      (N190)? \piso.data_r [562] : 
                      (N192)? \piso.data_r [594] : 
                      (N194)? \piso.data_r [626] : 
                      (N196)? \piso.data_r [658] : 
                      (N198)? \piso.data_r [690] : 
                      (N200)? \piso.data_r [722] : 
                      (N202)? \piso.data_r [754] : 
                      (N204)? \piso.data_r [786] : 
                      (N206)? \piso.data_r [818] : 
                      (N208)? \piso.data_r [850] : 
                      (N210)? \piso.data_r [882] : 
                      (N212)? \piso.data_r [914] : 
                      (N214)? \piso.data_r [946] : 
                      (N216)? \piso.data_r [978] : 
                      (N218)? \piso.data_r [1010] : 
                      (N220)? \piso.data_r [1042] : 
                      (N222)? \piso.data_r [1074] : 
                      (N224)? \piso.data_r [1106] : 
                      (N226)? \piso.data_r [1138] : 
                      (N228)? \piso.data_r [1170] : 
                      (N230)? \piso.data_r [1202] : 
                      (N232)? \piso.data_r [1234] : 
                      (N234)? \piso.data_r [1266] : 
                      (N236)? \piso.data_r [1298] : 
                      (N238)? \piso.data_r [1330] : 
                      (N240)? \piso.data_r [1362] : 
                      (N242)? \piso.data_r [1394] : 
                      (N244)? \piso.data_r [1426] : 
                      (N246)? \piso.data_r [1458] : 
                      (N248)? \piso.data_r [1490] : 
                      (N250)? \piso.data_r [1522] : 
                      (N252)? \piso.data_r [1554] : 
                      (N254)? \piso.data_r [1586] : 
                      (N256)? \piso.data_r [1618] : 
                      (N258)? \piso.data_r [1650] : 
                      (N260)? \piso.data_r [1682] : 
                      (N262)? \piso.data_r [1714] : 
                      (N264)? \piso.data_r [1746] : 
                      (N266)? \piso.data_r [1778] : 
                      (N268)? \piso.data_r [1810] : 
                      (N270)? \piso.data_r [1842] : 
                      (N272)? \piso.data_r [1874] : 
                      (N274)? \piso.data_r [1906] : 
                      (N276)? \piso.data_r [1938] : 
                      (N278)? \piso.data_r [1970] : 
                      (N280)? \piso.data_r [2002] : 
                      (N282)? \piso.data_r [2034] : 
                      (N157)? \piso.data_r [2066] : 
                      (N159)? \piso.data_r [2098] : 
                      (N161)? \piso.data_r [2130] : 
                      (N163)? \piso.data_r [2162] : 
                      (N165)? \piso.data_r [2194] : 
                      (N167)? \piso.data_r [2226] : 
                      (N169)? \piso.data_r [2258] : 
                      (N171)? \piso.data_r [2290] : 
                      (N173)? \piso.data_r [2322] : 
                      (N175)? \piso.data_r [2354] : 
                      (N177)? \piso.data_r [2386] : 
                      (N179)? \piso.data_r [2418] : 
                      (N181)? \piso.data_r [2450] : 
                      (N183)? \piso.data_r [2482] : 
                      (N185)? \piso.data_r [2514] : 
                      (N187)? \piso.data_r [2546] : 
                      (N189)? \piso.data_r [2578] : 
                      (N191)? \piso.data_r [2610] : 
                      (N193)? \piso.data_r [2642] : 
                      (N195)? \piso.data_r [2674] : 
                      (N197)? \piso.data_r [2706] : 
                      (N199)? \piso.data_r [2738] : 
                      (N201)? \piso.data_r [2770] : 
                      (N203)? \piso.data_r [2802] : 
                      (N205)? \piso.data_r [2834] : 
                      (N207)? \piso.data_r [2866] : 
                      (N209)? \piso.data_r [2898] : 
                      (N211)? \piso.data_r [2930] : 
                      (N213)? \piso.data_r [2962] : 
                      (N215)? \piso.data_r [2994] : 
                      (N217)? \piso.data_r [3026] : 
                      (N219)? \piso.data_r [3058] : 
                      (N221)? \piso.data_r [3090] : 
                      (N223)? \piso.data_r [3122] : 
                      (N225)? \piso.data_r [3154] : 
                      (N227)? \piso.data_r [3186] : 
                      (N229)? \piso.data_r [3218] : 
                      (N231)? \piso.data_r [3250] : 
                      (N233)? \piso.data_r [3282] : 
                      (N235)? \piso.data_r [3314] : 
                      (N237)? \piso.data_r [3346] : 
                      (N239)? \piso.data_r [3378] : 
                      (N241)? \piso.data_r [3410] : 
                      (N243)? \piso.data_r [3442] : 
                      (N245)? \piso.data_r [3474] : 
                      (N247)? \piso.data_r [3506] : 
                      (N249)? \piso.data_r [3538] : 
                      (N251)? \piso.data_r [3570] : 
                      (N253)? \piso.data_r [3602] : 
                      (N255)? \piso.data_r [3634] : 
                      (N257)? \piso.data_r [3666] : 
                      (N259)? \piso.data_r [3698] : 
                      (N261)? \piso.data_r [3730] : 
                      (N263)? \piso.data_r [3762] : 
                      (N265)? \piso.data_r [3794] : 
                      (N267)? \piso.data_r [3826] : 
                      (N269)? \piso.data_r [3858] : 
                      (N271)? \piso.data_r [3890] : 
                      (N273)? \piso.data_r [3922] : 
                      (N275)? \piso.data_r [3954] : 
                      (N277)? \piso.data_r [3986] : 
                      (N279)? \piso.data_r [4018] : 
                      (N281)? \piso.data_r [4050] : 
                      (N283)? \piso.data_r [4082] : 1'b0;
  assign data_o[17] = (N156)? \piso.data_r [17] : 
                      (N158)? \piso.data_r [49] : 
                      (N160)? \piso.data_r [81] : 
                      (N162)? \piso.data_r [113] : 
                      (N164)? \piso.data_r [145] : 
                      (N166)? \piso.data_r [177] : 
                      (N168)? \piso.data_r [209] : 
                      (N170)? \piso.data_r [241] : 
                      (N172)? \piso.data_r [273] : 
                      (N174)? \piso.data_r [305] : 
                      (N176)? \piso.data_r [337] : 
                      (N178)? \piso.data_r [369] : 
                      (N180)? \piso.data_r [401] : 
                      (N182)? \piso.data_r [433] : 
                      (N184)? \piso.data_r [465] : 
                      (N186)? \piso.data_r [497] : 
                      (N188)? \piso.data_r [529] : 
                      (N190)? \piso.data_r [561] : 
                      (N192)? \piso.data_r [593] : 
                      (N194)? \piso.data_r [625] : 
                      (N196)? \piso.data_r [657] : 
                      (N198)? \piso.data_r [689] : 
                      (N200)? \piso.data_r [721] : 
                      (N202)? \piso.data_r [753] : 
                      (N204)? \piso.data_r [785] : 
                      (N206)? \piso.data_r [817] : 
                      (N208)? \piso.data_r [849] : 
                      (N210)? \piso.data_r [881] : 
                      (N212)? \piso.data_r [913] : 
                      (N214)? \piso.data_r [945] : 
                      (N216)? \piso.data_r [977] : 
                      (N218)? \piso.data_r [1009] : 
                      (N220)? \piso.data_r [1041] : 
                      (N222)? \piso.data_r [1073] : 
                      (N224)? \piso.data_r [1105] : 
                      (N226)? \piso.data_r [1137] : 
                      (N228)? \piso.data_r [1169] : 
                      (N230)? \piso.data_r [1201] : 
                      (N232)? \piso.data_r [1233] : 
                      (N234)? \piso.data_r [1265] : 
                      (N236)? \piso.data_r [1297] : 
                      (N238)? \piso.data_r [1329] : 
                      (N240)? \piso.data_r [1361] : 
                      (N242)? \piso.data_r [1393] : 
                      (N244)? \piso.data_r [1425] : 
                      (N246)? \piso.data_r [1457] : 
                      (N248)? \piso.data_r [1489] : 
                      (N250)? \piso.data_r [1521] : 
                      (N252)? \piso.data_r [1553] : 
                      (N254)? \piso.data_r [1585] : 
                      (N256)? \piso.data_r [1617] : 
                      (N258)? \piso.data_r [1649] : 
                      (N260)? \piso.data_r [1681] : 
                      (N262)? \piso.data_r [1713] : 
                      (N264)? \piso.data_r [1745] : 
                      (N266)? \piso.data_r [1777] : 
                      (N268)? \piso.data_r [1809] : 
                      (N270)? \piso.data_r [1841] : 
                      (N272)? \piso.data_r [1873] : 
                      (N274)? \piso.data_r [1905] : 
                      (N276)? \piso.data_r [1937] : 
                      (N278)? \piso.data_r [1969] : 
                      (N280)? \piso.data_r [2001] : 
                      (N282)? \piso.data_r [2033] : 
                      (N157)? \piso.data_r [2065] : 
                      (N159)? \piso.data_r [2097] : 
                      (N161)? \piso.data_r [2129] : 
                      (N163)? \piso.data_r [2161] : 
                      (N165)? \piso.data_r [2193] : 
                      (N167)? \piso.data_r [2225] : 
                      (N169)? \piso.data_r [2257] : 
                      (N171)? \piso.data_r [2289] : 
                      (N173)? \piso.data_r [2321] : 
                      (N175)? \piso.data_r [2353] : 
                      (N177)? \piso.data_r [2385] : 
                      (N179)? \piso.data_r [2417] : 
                      (N181)? \piso.data_r [2449] : 
                      (N183)? \piso.data_r [2481] : 
                      (N185)? \piso.data_r [2513] : 
                      (N187)? \piso.data_r [2545] : 
                      (N189)? \piso.data_r [2577] : 
                      (N191)? \piso.data_r [2609] : 
                      (N193)? \piso.data_r [2641] : 
                      (N195)? \piso.data_r [2673] : 
                      (N197)? \piso.data_r [2705] : 
                      (N199)? \piso.data_r [2737] : 
                      (N201)? \piso.data_r [2769] : 
                      (N203)? \piso.data_r [2801] : 
                      (N205)? \piso.data_r [2833] : 
                      (N207)? \piso.data_r [2865] : 
                      (N209)? \piso.data_r [2897] : 
                      (N211)? \piso.data_r [2929] : 
                      (N213)? \piso.data_r [2961] : 
                      (N215)? \piso.data_r [2993] : 
                      (N217)? \piso.data_r [3025] : 
                      (N219)? \piso.data_r [3057] : 
                      (N221)? \piso.data_r [3089] : 
                      (N223)? \piso.data_r [3121] : 
                      (N225)? \piso.data_r [3153] : 
                      (N227)? \piso.data_r [3185] : 
                      (N229)? \piso.data_r [3217] : 
                      (N231)? \piso.data_r [3249] : 
                      (N233)? \piso.data_r [3281] : 
                      (N235)? \piso.data_r [3313] : 
                      (N237)? \piso.data_r [3345] : 
                      (N239)? \piso.data_r [3377] : 
                      (N241)? \piso.data_r [3409] : 
                      (N243)? \piso.data_r [3441] : 
                      (N245)? \piso.data_r [3473] : 
                      (N247)? \piso.data_r [3505] : 
                      (N249)? \piso.data_r [3537] : 
                      (N251)? \piso.data_r [3569] : 
                      (N253)? \piso.data_r [3601] : 
                      (N255)? \piso.data_r [3633] : 
                      (N257)? \piso.data_r [3665] : 
                      (N259)? \piso.data_r [3697] : 
                      (N261)? \piso.data_r [3729] : 
                      (N263)? \piso.data_r [3761] : 
                      (N265)? \piso.data_r [3793] : 
                      (N267)? \piso.data_r [3825] : 
                      (N269)? \piso.data_r [3857] : 
                      (N271)? \piso.data_r [3889] : 
                      (N273)? \piso.data_r [3921] : 
                      (N275)? \piso.data_r [3953] : 
                      (N277)? \piso.data_r [3985] : 
                      (N279)? \piso.data_r [4017] : 
                      (N281)? \piso.data_r [4049] : 
                      (N283)? \piso.data_r [4081] : 1'b0;
  assign data_o[16] = (N156)? \piso.data_r [16] : 
                      (N158)? \piso.data_r [48] : 
                      (N160)? \piso.data_r [80] : 
                      (N162)? \piso.data_r [112] : 
                      (N164)? \piso.data_r [144] : 
                      (N166)? \piso.data_r [176] : 
                      (N168)? \piso.data_r [208] : 
                      (N170)? \piso.data_r [240] : 
                      (N172)? \piso.data_r [272] : 
                      (N174)? \piso.data_r [304] : 
                      (N176)? \piso.data_r [336] : 
                      (N178)? \piso.data_r [368] : 
                      (N180)? \piso.data_r [400] : 
                      (N182)? \piso.data_r [432] : 
                      (N184)? \piso.data_r [464] : 
                      (N186)? \piso.data_r [496] : 
                      (N188)? \piso.data_r [528] : 
                      (N190)? \piso.data_r [560] : 
                      (N192)? \piso.data_r [592] : 
                      (N194)? \piso.data_r [624] : 
                      (N196)? \piso.data_r [656] : 
                      (N198)? \piso.data_r [688] : 
                      (N200)? \piso.data_r [720] : 
                      (N202)? \piso.data_r [752] : 
                      (N204)? \piso.data_r [784] : 
                      (N206)? \piso.data_r [816] : 
                      (N208)? \piso.data_r [848] : 
                      (N210)? \piso.data_r [880] : 
                      (N212)? \piso.data_r [912] : 
                      (N214)? \piso.data_r [944] : 
                      (N216)? \piso.data_r [976] : 
                      (N218)? \piso.data_r [1008] : 
                      (N220)? \piso.data_r [1040] : 
                      (N222)? \piso.data_r [1072] : 
                      (N224)? \piso.data_r [1104] : 
                      (N226)? \piso.data_r [1136] : 
                      (N228)? \piso.data_r [1168] : 
                      (N230)? \piso.data_r [1200] : 
                      (N232)? \piso.data_r [1232] : 
                      (N234)? \piso.data_r [1264] : 
                      (N236)? \piso.data_r [1296] : 
                      (N238)? \piso.data_r [1328] : 
                      (N240)? \piso.data_r [1360] : 
                      (N242)? \piso.data_r [1392] : 
                      (N244)? \piso.data_r [1424] : 
                      (N246)? \piso.data_r [1456] : 
                      (N248)? \piso.data_r [1488] : 
                      (N250)? \piso.data_r [1520] : 
                      (N252)? \piso.data_r [1552] : 
                      (N254)? \piso.data_r [1584] : 
                      (N256)? \piso.data_r [1616] : 
                      (N258)? \piso.data_r [1648] : 
                      (N260)? \piso.data_r [1680] : 
                      (N262)? \piso.data_r [1712] : 
                      (N264)? \piso.data_r [1744] : 
                      (N266)? \piso.data_r [1776] : 
                      (N268)? \piso.data_r [1808] : 
                      (N270)? \piso.data_r [1840] : 
                      (N272)? \piso.data_r [1872] : 
                      (N274)? \piso.data_r [1904] : 
                      (N276)? \piso.data_r [1936] : 
                      (N278)? \piso.data_r [1968] : 
                      (N280)? \piso.data_r [2000] : 
                      (N282)? \piso.data_r [2032] : 
                      (N157)? \piso.data_r [2064] : 
                      (N159)? \piso.data_r [2096] : 
                      (N161)? \piso.data_r [2128] : 
                      (N163)? \piso.data_r [2160] : 
                      (N165)? \piso.data_r [2192] : 
                      (N167)? \piso.data_r [2224] : 
                      (N169)? \piso.data_r [2256] : 
                      (N171)? \piso.data_r [2288] : 
                      (N173)? \piso.data_r [2320] : 
                      (N175)? \piso.data_r [2352] : 
                      (N177)? \piso.data_r [2384] : 
                      (N179)? \piso.data_r [2416] : 
                      (N181)? \piso.data_r [2448] : 
                      (N183)? \piso.data_r [2480] : 
                      (N185)? \piso.data_r [2512] : 
                      (N187)? \piso.data_r [2544] : 
                      (N189)? \piso.data_r [2576] : 
                      (N191)? \piso.data_r [2608] : 
                      (N193)? \piso.data_r [2640] : 
                      (N195)? \piso.data_r [2672] : 
                      (N197)? \piso.data_r [2704] : 
                      (N199)? \piso.data_r [2736] : 
                      (N201)? \piso.data_r [2768] : 
                      (N203)? \piso.data_r [2800] : 
                      (N205)? \piso.data_r [2832] : 
                      (N207)? \piso.data_r [2864] : 
                      (N209)? \piso.data_r [2896] : 
                      (N211)? \piso.data_r [2928] : 
                      (N213)? \piso.data_r [2960] : 
                      (N215)? \piso.data_r [2992] : 
                      (N217)? \piso.data_r [3024] : 
                      (N219)? \piso.data_r [3056] : 
                      (N221)? \piso.data_r [3088] : 
                      (N223)? \piso.data_r [3120] : 
                      (N225)? \piso.data_r [3152] : 
                      (N227)? \piso.data_r [3184] : 
                      (N229)? \piso.data_r [3216] : 
                      (N231)? \piso.data_r [3248] : 
                      (N233)? \piso.data_r [3280] : 
                      (N235)? \piso.data_r [3312] : 
                      (N237)? \piso.data_r [3344] : 
                      (N239)? \piso.data_r [3376] : 
                      (N241)? \piso.data_r [3408] : 
                      (N243)? \piso.data_r [3440] : 
                      (N245)? \piso.data_r [3472] : 
                      (N247)? \piso.data_r [3504] : 
                      (N249)? \piso.data_r [3536] : 
                      (N251)? \piso.data_r [3568] : 
                      (N253)? \piso.data_r [3600] : 
                      (N255)? \piso.data_r [3632] : 
                      (N257)? \piso.data_r [3664] : 
                      (N259)? \piso.data_r [3696] : 
                      (N261)? \piso.data_r [3728] : 
                      (N263)? \piso.data_r [3760] : 
                      (N265)? \piso.data_r [3792] : 
                      (N267)? \piso.data_r [3824] : 
                      (N269)? \piso.data_r [3856] : 
                      (N271)? \piso.data_r [3888] : 
                      (N273)? \piso.data_r [3920] : 
                      (N275)? \piso.data_r [3952] : 
                      (N277)? \piso.data_r [3984] : 
                      (N279)? \piso.data_r [4016] : 
                      (N281)? \piso.data_r [4048] : 
                      (N283)? \piso.data_r [4080] : 1'b0;
  assign data_o[15] = (N156)? \piso.data_r [15] : 
                      (N158)? \piso.data_r [47] : 
                      (N160)? \piso.data_r [79] : 
                      (N162)? \piso.data_r [111] : 
                      (N164)? \piso.data_r [143] : 
                      (N166)? \piso.data_r [175] : 
                      (N168)? \piso.data_r [207] : 
                      (N170)? \piso.data_r [239] : 
                      (N172)? \piso.data_r [271] : 
                      (N174)? \piso.data_r [303] : 
                      (N176)? \piso.data_r [335] : 
                      (N178)? \piso.data_r [367] : 
                      (N180)? \piso.data_r [399] : 
                      (N182)? \piso.data_r [431] : 
                      (N184)? \piso.data_r [463] : 
                      (N186)? \piso.data_r [495] : 
                      (N188)? \piso.data_r [527] : 
                      (N190)? \piso.data_r [559] : 
                      (N192)? \piso.data_r [591] : 
                      (N194)? \piso.data_r [623] : 
                      (N196)? \piso.data_r [655] : 
                      (N198)? \piso.data_r [687] : 
                      (N200)? \piso.data_r [719] : 
                      (N202)? \piso.data_r [751] : 
                      (N204)? \piso.data_r [783] : 
                      (N206)? \piso.data_r [815] : 
                      (N208)? \piso.data_r [847] : 
                      (N210)? \piso.data_r [879] : 
                      (N212)? \piso.data_r [911] : 
                      (N214)? \piso.data_r [943] : 
                      (N216)? \piso.data_r [975] : 
                      (N218)? \piso.data_r [1007] : 
                      (N220)? \piso.data_r [1039] : 
                      (N222)? \piso.data_r [1071] : 
                      (N224)? \piso.data_r [1103] : 
                      (N226)? \piso.data_r [1135] : 
                      (N228)? \piso.data_r [1167] : 
                      (N230)? \piso.data_r [1199] : 
                      (N232)? \piso.data_r [1231] : 
                      (N234)? \piso.data_r [1263] : 
                      (N236)? \piso.data_r [1295] : 
                      (N238)? \piso.data_r [1327] : 
                      (N240)? \piso.data_r [1359] : 
                      (N242)? \piso.data_r [1391] : 
                      (N244)? \piso.data_r [1423] : 
                      (N246)? \piso.data_r [1455] : 
                      (N248)? \piso.data_r [1487] : 
                      (N250)? \piso.data_r [1519] : 
                      (N252)? \piso.data_r [1551] : 
                      (N254)? \piso.data_r [1583] : 
                      (N256)? \piso.data_r [1615] : 
                      (N258)? \piso.data_r [1647] : 
                      (N260)? \piso.data_r [1679] : 
                      (N262)? \piso.data_r [1711] : 
                      (N264)? \piso.data_r [1743] : 
                      (N266)? \piso.data_r [1775] : 
                      (N268)? \piso.data_r [1807] : 
                      (N270)? \piso.data_r [1839] : 
                      (N272)? \piso.data_r [1871] : 
                      (N274)? \piso.data_r [1903] : 
                      (N276)? \piso.data_r [1935] : 
                      (N278)? \piso.data_r [1967] : 
                      (N280)? \piso.data_r [1999] : 
                      (N282)? \piso.data_r [2031] : 
                      (N157)? \piso.data_r [2063] : 
                      (N159)? \piso.data_r [2095] : 
                      (N161)? \piso.data_r [2127] : 
                      (N163)? \piso.data_r [2159] : 
                      (N165)? \piso.data_r [2191] : 
                      (N167)? \piso.data_r [2223] : 
                      (N169)? \piso.data_r [2255] : 
                      (N171)? \piso.data_r [2287] : 
                      (N173)? \piso.data_r [2319] : 
                      (N175)? \piso.data_r [2351] : 
                      (N177)? \piso.data_r [2383] : 
                      (N179)? \piso.data_r [2415] : 
                      (N181)? \piso.data_r [2447] : 
                      (N183)? \piso.data_r [2479] : 
                      (N185)? \piso.data_r [2511] : 
                      (N187)? \piso.data_r [2543] : 
                      (N189)? \piso.data_r [2575] : 
                      (N191)? \piso.data_r [2607] : 
                      (N193)? \piso.data_r [2639] : 
                      (N195)? \piso.data_r [2671] : 
                      (N197)? \piso.data_r [2703] : 
                      (N199)? \piso.data_r [2735] : 
                      (N201)? \piso.data_r [2767] : 
                      (N203)? \piso.data_r [2799] : 
                      (N205)? \piso.data_r [2831] : 
                      (N207)? \piso.data_r [2863] : 
                      (N209)? \piso.data_r [2895] : 
                      (N211)? \piso.data_r [2927] : 
                      (N213)? \piso.data_r [2959] : 
                      (N215)? \piso.data_r [2991] : 
                      (N217)? \piso.data_r [3023] : 
                      (N219)? \piso.data_r [3055] : 
                      (N221)? \piso.data_r [3087] : 
                      (N223)? \piso.data_r [3119] : 
                      (N225)? \piso.data_r [3151] : 
                      (N227)? \piso.data_r [3183] : 
                      (N229)? \piso.data_r [3215] : 
                      (N231)? \piso.data_r [3247] : 
                      (N233)? \piso.data_r [3279] : 
                      (N235)? \piso.data_r [3311] : 
                      (N237)? \piso.data_r [3343] : 
                      (N239)? \piso.data_r [3375] : 
                      (N241)? \piso.data_r [3407] : 
                      (N243)? \piso.data_r [3439] : 
                      (N245)? \piso.data_r [3471] : 
                      (N247)? \piso.data_r [3503] : 
                      (N249)? \piso.data_r [3535] : 
                      (N251)? \piso.data_r [3567] : 
                      (N253)? \piso.data_r [3599] : 
                      (N255)? \piso.data_r [3631] : 
                      (N257)? \piso.data_r [3663] : 
                      (N259)? \piso.data_r [3695] : 
                      (N261)? \piso.data_r [3727] : 
                      (N263)? \piso.data_r [3759] : 
                      (N265)? \piso.data_r [3791] : 
                      (N267)? \piso.data_r [3823] : 
                      (N269)? \piso.data_r [3855] : 
                      (N271)? \piso.data_r [3887] : 
                      (N273)? \piso.data_r [3919] : 
                      (N275)? \piso.data_r [3951] : 
                      (N277)? \piso.data_r [3983] : 
                      (N279)? \piso.data_r [4015] : 
                      (N281)? \piso.data_r [4047] : 
                      (N283)? \piso.data_r [4079] : 1'b0;
  assign data_o[14] = (N156)? \piso.data_r [14] : 
                      (N158)? \piso.data_r [46] : 
                      (N160)? \piso.data_r [78] : 
                      (N162)? \piso.data_r [110] : 
                      (N164)? \piso.data_r [142] : 
                      (N166)? \piso.data_r [174] : 
                      (N168)? \piso.data_r [206] : 
                      (N170)? \piso.data_r [238] : 
                      (N172)? \piso.data_r [270] : 
                      (N174)? \piso.data_r [302] : 
                      (N176)? \piso.data_r [334] : 
                      (N178)? \piso.data_r [366] : 
                      (N180)? \piso.data_r [398] : 
                      (N182)? \piso.data_r [430] : 
                      (N184)? \piso.data_r [462] : 
                      (N186)? \piso.data_r [494] : 
                      (N188)? \piso.data_r [526] : 
                      (N190)? \piso.data_r [558] : 
                      (N192)? \piso.data_r [590] : 
                      (N194)? \piso.data_r [622] : 
                      (N196)? \piso.data_r [654] : 
                      (N198)? \piso.data_r [686] : 
                      (N200)? \piso.data_r [718] : 
                      (N202)? \piso.data_r [750] : 
                      (N204)? \piso.data_r [782] : 
                      (N206)? \piso.data_r [814] : 
                      (N208)? \piso.data_r [846] : 
                      (N210)? \piso.data_r [878] : 
                      (N212)? \piso.data_r [910] : 
                      (N214)? \piso.data_r [942] : 
                      (N216)? \piso.data_r [974] : 
                      (N218)? \piso.data_r [1006] : 
                      (N220)? \piso.data_r [1038] : 
                      (N222)? \piso.data_r [1070] : 
                      (N224)? \piso.data_r [1102] : 
                      (N226)? \piso.data_r [1134] : 
                      (N228)? \piso.data_r [1166] : 
                      (N230)? \piso.data_r [1198] : 
                      (N232)? \piso.data_r [1230] : 
                      (N234)? \piso.data_r [1262] : 
                      (N236)? \piso.data_r [1294] : 
                      (N238)? \piso.data_r [1326] : 
                      (N240)? \piso.data_r [1358] : 
                      (N242)? \piso.data_r [1390] : 
                      (N244)? \piso.data_r [1422] : 
                      (N246)? \piso.data_r [1454] : 
                      (N248)? \piso.data_r [1486] : 
                      (N250)? \piso.data_r [1518] : 
                      (N252)? \piso.data_r [1550] : 
                      (N254)? \piso.data_r [1582] : 
                      (N256)? \piso.data_r [1614] : 
                      (N258)? \piso.data_r [1646] : 
                      (N260)? \piso.data_r [1678] : 
                      (N262)? \piso.data_r [1710] : 
                      (N264)? \piso.data_r [1742] : 
                      (N266)? \piso.data_r [1774] : 
                      (N268)? \piso.data_r [1806] : 
                      (N270)? \piso.data_r [1838] : 
                      (N272)? \piso.data_r [1870] : 
                      (N274)? \piso.data_r [1902] : 
                      (N276)? \piso.data_r [1934] : 
                      (N278)? \piso.data_r [1966] : 
                      (N280)? \piso.data_r [1998] : 
                      (N282)? \piso.data_r [2030] : 
                      (N157)? \piso.data_r [2062] : 
                      (N159)? \piso.data_r [2094] : 
                      (N161)? \piso.data_r [2126] : 
                      (N163)? \piso.data_r [2158] : 
                      (N165)? \piso.data_r [2190] : 
                      (N167)? \piso.data_r [2222] : 
                      (N169)? \piso.data_r [2254] : 
                      (N171)? \piso.data_r [2286] : 
                      (N173)? \piso.data_r [2318] : 
                      (N175)? \piso.data_r [2350] : 
                      (N177)? \piso.data_r [2382] : 
                      (N179)? \piso.data_r [2414] : 
                      (N181)? \piso.data_r [2446] : 
                      (N183)? \piso.data_r [2478] : 
                      (N185)? \piso.data_r [2510] : 
                      (N187)? \piso.data_r [2542] : 
                      (N189)? \piso.data_r [2574] : 
                      (N191)? \piso.data_r [2606] : 
                      (N193)? \piso.data_r [2638] : 
                      (N195)? \piso.data_r [2670] : 
                      (N197)? \piso.data_r [2702] : 
                      (N199)? \piso.data_r [2734] : 
                      (N201)? \piso.data_r [2766] : 
                      (N203)? \piso.data_r [2798] : 
                      (N205)? \piso.data_r [2830] : 
                      (N207)? \piso.data_r [2862] : 
                      (N209)? \piso.data_r [2894] : 
                      (N211)? \piso.data_r [2926] : 
                      (N213)? \piso.data_r [2958] : 
                      (N215)? \piso.data_r [2990] : 
                      (N217)? \piso.data_r [3022] : 
                      (N219)? \piso.data_r [3054] : 
                      (N221)? \piso.data_r [3086] : 
                      (N223)? \piso.data_r [3118] : 
                      (N225)? \piso.data_r [3150] : 
                      (N227)? \piso.data_r [3182] : 
                      (N229)? \piso.data_r [3214] : 
                      (N231)? \piso.data_r [3246] : 
                      (N233)? \piso.data_r [3278] : 
                      (N235)? \piso.data_r [3310] : 
                      (N237)? \piso.data_r [3342] : 
                      (N239)? \piso.data_r [3374] : 
                      (N241)? \piso.data_r [3406] : 
                      (N243)? \piso.data_r [3438] : 
                      (N245)? \piso.data_r [3470] : 
                      (N247)? \piso.data_r [3502] : 
                      (N249)? \piso.data_r [3534] : 
                      (N251)? \piso.data_r [3566] : 
                      (N253)? \piso.data_r [3598] : 
                      (N255)? \piso.data_r [3630] : 
                      (N257)? \piso.data_r [3662] : 
                      (N259)? \piso.data_r [3694] : 
                      (N261)? \piso.data_r [3726] : 
                      (N263)? \piso.data_r [3758] : 
                      (N265)? \piso.data_r [3790] : 
                      (N267)? \piso.data_r [3822] : 
                      (N269)? \piso.data_r [3854] : 
                      (N271)? \piso.data_r [3886] : 
                      (N273)? \piso.data_r [3918] : 
                      (N275)? \piso.data_r [3950] : 
                      (N277)? \piso.data_r [3982] : 
                      (N279)? \piso.data_r [4014] : 
                      (N281)? \piso.data_r [4046] : 
                      (N283)? \piso.data_r [4078] : 1'b0;
  assign data_o[13] = (N156)? \piso.data_r [13] : 
                      (N158)? \piso.data_r [45] : 
                      (N160)? \piso.data_r [77] : 
                      (N162)? \piso.data_r [109] : 
                      (N164)? \piso.data_r [141] : 
                      (N166)? \piso.data_r [173] : 
                      (N168)? \piso.data_r [205] : 
                      (N170)? \piso.data_r [237] : 
                      (N172)? \piso.data_r [269] : 
                      (N174)? \piso.data_r [301] : 
                      (N176)? \piso.data_r [333] : 
                      (N178)? \piso.data_r [365] : 
                      (N180)? \piso.data_r [397] : 
                      (N182)? \piso.data_r [429] : 
                      (N184)? \piso.data_r [461] : 
                      (N186)? \piso.data_r [493] : 
                      (N188)? \piso.data_r [525] : 
                      (N190)? \piso.data_r [557] : 
                      (N192)? \piso.data_r [589] : 
                      (N194)? \piso.data_r [621] : 
                      (N196)? \piso.data_r [653] : 
                      (N198)? \piso.data_r [685] : 
                      (N200)? \piso.data_r [717] : 
                      (N202)? \piso.data_r [749] : 
                      (N204)? \piso.data_r [781] : 
                      (N206)? \piso.data_r [813] : 
                      (N208)? \piso.data_r [845] : 
                      (N210)? \piso.data_r [877] : 
                      (N212)? \piso.data_r [909] : 
                      (N214)? \piso.data_r [941] : 
                      (N216)? \piso.data_r [973] : 
                      (N218)? \piso.data_r [1005] : 
                      (N220)? \piso.data_r [1037] : 
                      (N222)? \piso.data_r [1069] : 
                      (N224)? \piso.data_r [1101] : 
                      (N226)? \piso.data_r [1133] : 
                      (N228)? \piso.data_r [1165] : 
                      (N230)? \piso.data_r [1197] : 
                      (N232)? \piso.data_r [1229] : 
                      (N234)? \piso.data_r [1261] : 
                      (N236)? \piso.data_r [1293] : 
                      (N238)? \piso.data_r [1325] : 
                      (N240)? \piso.data_r [1357] : 
                      (N242)? \piso.data_r [1389] : 
                      (N244)? \piso.data_r [1421] : 
                      (N246)? \piso.data_r [1453] : 
                      (N248)? \piso.data_r [1485] : 
                      (N250)? \piso.data_r [1517] : 
                      (N252)? \piso.data_r [1549] : 
                      (N254)? \piso.data_r [1581] : 
                      (N256)? \piso.data_r [1613] : 
                      (N258)? \piso.data_r [1645] : 
                      (N260)? \piso.data_r [1677] : 
                      (N262)? \piso.data_r [1709] : 
                      (N264)? \piso.data_r [1741] : 
                      (N266)? \piso.data_r [1773] : 
                      (N268)? \piso.data_r [1805] : 
                      (N270)? \piso.data_r [1837] : 
                      (N272)? \piso.data_r [1869] : 
                      (N274)? \piso.data_r [1901] : 
                      (N276)? \piso.data_r [1933] : 
                      (N278)? \piso.data_r [1965] : 
                      (N280)? \piso.data_r [1997] : 
                      (N282)? \piso.data_r [2029] : 
                      (N157)? \piso.data_r [2061] : 
                      (N159)? \piso.data_r [2093] : 
                      (N161)? \piso.data_r [2125] : 
                      (N163)? \piso.data_r [2157] : 
                      (N165)? \piso.data_r [2189] : 
                      (N167)? \piso.data_r [2221] : 
                      (N169)? \piso.data_r [2253] : 
                      (N171)? \piso.data_r [2285] : 
                      (N173)? \piso.data_r [2317] : 
                      (N175)? \piso.data_r [2349] : 
                      (N177)? \piso.data_r [2381] : 
                      (N179)? \piso.data_r [2413] : 
                      (N181)? \piso.data_r [2445] : 
                      (N183)? \piso.data_r [2477] : 
                      (N185)? \piso.data_r [2509] : 
                      (N187)? \piso.data_r [2541] : 
                      (N189)? \piso.data_r [2573] : 
                      (N191)? \piso.data_r [2605] : 
                      (N193)? \piso.data_r [2637] : 
                      (N195)? \piso.data_r [2669] : 
                      (N197)? \piso.data_r [2701] : 
                      (N199)? \piso.data_r [2733] : 
                      (N201)? \piso.data_r [2765] : 
                      (N203)? \piso.data_r [2797] : 
                      (N205)? \piso.data_r [2829] : 
                      (N207)? \piso.data_r [2861] : 
                      (N209)? \piso.data_r [2893] : 
                      (N211)? \piso.data_r [2925] : 
                      (N213)? \piso.data_r [2957] : 
                      (N215)? \piso.data_r [2989] : 
                      (N217)? \piso.data_r [3021] : 
                      (N219)? \piso.data_r [3053] : 
                      (N221)? \piso.data_r [3085] : 
                      (N223)? \piso.data_r [3117] : 
                      (N225)? \piso.data_r [3149] : 
                      (N227)? \piso.data_r [3181] : 
                      (N229)? \piso.data_r [3213] : 
                      (N231)? \piso.data_r [3245] : 
                      (N233)? \piso.data_r [3277] : 
                      (N235)? \piso.data_r [3309] : 
                      (N237)? \piso.data_r [3341] : 
                      (N239)? \piso.data_r [3373] : 
                      (N241)? \piso.data_r [3405] : 
                      (N243)? \piso.data_r [3437] : 
                      (N245)? \piso.data_r [3469] : 
                      (N247)? \piso.data_r [3501] : 
                      (N249)? \piso.data_r [3533] : 
                      (N251)? \piso.data_r [3565] : 
                      (N253)? \piso.data_r [3597] : 
                      (N255)? \piso.data_r [3629] : 
                      (N257)? \piso.data_r [3661] : 
                      (N259)? \piso.data_r [3693] : 
                      (N261)? \piso.data_r [3725] : 
                      (N263)? \piso.data_r [3757] : 
                      (N265)? \piso.data_r [3789] : 
                      (N267)? \piso.data_r [3821] : 
                      (N269)? \piso.data_r [3853] : 
                      (N271)? \piso.data_r [3885] : 
                      (N273)? \piso.data_r [3917] : 
                      (N275)? \piso.data_r [3949] : 
                      (N277)? \piso.data_r [3981] : 
                      (N279)? \piso.data_r [4013] : 
                      (N281)? \piso.data_r [4045] : 
                      (N283)? \piso.data_r [4077] : 1'b0;
  assign data_o[12] = (N156)? \piso.data_r [12] : 
                      (N158)? \piso.data_r [44] : 
                      (N160)? \piso.data_r [76] : 
                      (N162)? \piso.data_r [108] : 
                      (N164)? \piso.data_r [140] : 
                      (N166)? \piso.data_r [172] : 
                      (N168)? \piso.data_r [204] : 
                      (N170)? \piso.data_r [236] : 
                      (N172)? \piso.data_r [268] : 
                      (N174)? \piso.data_r [300] : 
                      (N176)? \piso.data_r [332] : 
                      (N178)? \piso.data_r [364] : 
                      (N180)? \piso.data_r [396] : 
                      (N182)? \piso.data_r [428] : 
                      (N184)? \piso.data_r [460] : 
                      (N186)? \piso.data_r [492] : 
                      (N188)? \piso.data_r [524] : 
                      (N190)? \piso.data_r [556] : 
                      (N192)? \piso.data_r [588] : 
                      (N194)? \piso.data_r [620] : 
                      (N196)? \piso.data_r [652] : 
                      (N198)? \piso.data_r [684] : 
                      (N200)? \piso.data_r [716] : 
                      (N202)? \piso.data_r [748] : 
                      (N204)? \piso.data_r [780] : 
                      (N206)? \piso.data_r [812] : 
                      (N208)? \piso.data_r [844] : 
                      (N210)? \piso.data_r [876] : 
                      (N212)? \piso.data_r [908] : 
                      (N214)? \piso.data_r [940] : 
                      (N216)? \piso.data_r [972] : 
                      (N218)? \piso.data_r [1004] : 
                      (N220)? \piso.data_r [1036] : 
                      (N222)? \piso.data_r [1068] : 
                      (N224)? \piso.data_r [1100] : 
                      (N226)? \piso.data_r [1132] : 
                      (N228)? \piso.data_r [1164] : 
                      (N230)? \piso.data_r [1196] : 
                      (N232)? \piso.data_r [1228] : 
                      (N234)? \piso.data_r [1260] : 
                      (N236)? \piso.data_r [1292] : 
                      (N238)? \piso.data_r [1324] : 
                      (N240)? \piso.data_r [1356] : 
                      (N242)? \piso.data_r [1388] : 
                      (N244)? \piso.data_r [1420] : 
                      (N246)? \piso.data_r [1452] : 
                      (N248)? \piso.data_r [1484] : 
                      (N250)? \piso.data_r [1516] : 
                      (N252)? \piso.data_r [1548] : 
                      (N254)? \piso.data_r [1580] : 
                      (N256)? \piso.data_r [1612] : 
                      (N258)? \piso.data_r [1644] : 
                      (N260)? \piso.data_r [1676] : 
                      (N262)? \piso.data_r [1708] : 
                      (N264)? \piso.data_r [1740] : 
                      (N266)? \piso.data_r [1772] : 
                      (N268)? \piso.data_r [1804] : 
                      (N270)? \piso.data_r [1836] : 
                      (N272)? \piso.data_r [1868] : 
                      (N274)? \piso.data_r [1900] : 
                      (N276)? \piso.data_r [1932] : 
                      (N278)? \piso.data_r [1964] : 
                      (N280)? \piso.data_r [1996] : 
                      (N282)? \piso.data_r [2028] : 
                      (N157)? \piso.data_r [2060] : 
                      (N159)? \piso.data_r [2092] : 
                      (N161)? \piso.data_r [2124] : 
                      (N163)? \piso.data_r [2156] : 
                      (N165)? \piso.data_r [2188] : 
                      (N167)? \piso.data_r [2220] : 
                      (N169)? \piso.data_r [2252] : 
                      (N171)? \piso.data_r [2284] : 
                      (N173)? \piso.data_r [2316] : 
                      (N175)? \piso.data_r [2348] : 
                      (N177)? \piso.data_r [2380] : 
                      (N179)? \piso.data_r [2412] : 
                      (N181)? \piso.data_r [2444] : 
                      (N183)? \piso.data_r [2476] : 
                      (N185)? \piso.data_r [2508] : 
                      (N187)? \piso.data_r [2540] : 
                      (N189)? \piso.data_r [2572] : 
                      (N191)? \piso.data_r [2604] : 
                      (N193)? \piso.data_r [2636] : 
                      (N195)? \piso.data_r [2668] : 
                      (N197)? \piso.data_r [2700] : 
                      (N199)? \piso.data_r [2732] : 
                      (N201)? \piso.data_r [2764] : 
                      (N203)? \piso.data_r [2796] : 
                      (N205)? \piso.data_r [2828] : 
                      (N207)? \piso.data_r [2860] : 
                      (N209)? \piso.data_r [2892] : 
                      (N211)? \piso.data_r [2924] : 
                      (N213)? \piso.data_r [2956] : 
                      (N215)? \piso.data_r [2988] : 
                      (N217)? \piso.data_r [3020] : 
                      (N219)? \piso.data_r [3052] : 
                      (N221)? \piso.data_r [3084] : 
                      (N223)? \piso.data_r [3116] : 
                      (N225)? \piso.data_r [3148] : 
                      (N227)? \piso.data_r [3180] : 
                      (N229)? \piso.data_r [3212] : 
                      (N231)? \piso.data_r [3244] : 
                      (N233)? \piso.data_r [3276] : 
                      (N235)? \piso.data_r [3308] : 
                      (N237)? \piso.data_r [3340] : 
                      (N239)? \piso.data_r [3372] : 
                      (N241)? \piso.data_r [3404] : 
                      (N243)? \piso.data_r [3436] : 
                      (N245)? \piso.data_r [3468] : 
                      (N247)? \piso.data_r [3500] : 
                      (N249)? \piso.data_r [3532] : 
                      (N251)? \piso.data_r [3564] : 
                      (N253)? \piso.data_r [3596] : 
                      (N255)? \piso.data_r [3628] : 
                      (N257)? \piso.data_r [3660] : 
                      (N259)? \piso.data_r [3692] : 
                      (N261)? \piso.data_r [3724] : 
                      (N263)? \piso.data_r [3756] : 
                      (N265)? \piso.data_r [3788] : 
                      (N267)? \piso.data_r [3820] : 
                      (N269)? \piso.data_r [3852] : 
                      (N271)? \piso.data_r [3884] : 
                      (N273)? \piso.data_r [3916] : 
                      (N275)? \piso.data_r [3948] : 
                      (N277)? \piso.data_r [3980] : 
                      (N279)? \piso.data_r [4012] : 
                      (N281)? \piso.data_r [4044] : 
                      (N283)? \piso.data_r [4076] : 1'b0;
  assign data_o[11] = (N156)? \piso.data_r [11] : 
                      (N158)? \piso.data_r [43] : 
                      (N160)? \piso.data_r [75] : 
                      (N162)? \piso.data_r [107] : 
                      (N164)? \piso.data_r [139] : 
                      (N166)? \piso.data_r [171] : 
                      (N168)? \piso.data_r [203] : 
                      (N170)? \piso.data_r [235] : 
                      (N172)? \piso.data_r [267] : 
                      (N174)? \piso.data_r [299] : 
                      (N176)? \piso.data_r [331] : 
                      (N178)? \piso.data_r [363] : 
                      (N180)? \piso.data_r [395] : 
                      (N182)? \piso.data_r [427] : 
                      (N184)? \piso.data_r [459] : 
                      (N186)? \piso.data_r [491] : 
                      (N188)? \piso.data_r [523] : 
                      (N190)? \piso.data_r [555] : 
                      (N192)? \piso.data_r [587] : 
                      (N194)? \piso.data_r [619] : 
                      (N196)? \piso.data_r [651] : 
                      (N198)? \piso.data_r [683] : 
                      (N200)? \piso.data_r [715] : 
                      (N202)? \piso.data_r [747] : 
                      (N204)? \piso.data_r [779] : 
                      (N206)? \piso.data_r [811] : 
                      (N208)? \piso.data_r [843] : 
                      (N210)? \piso.data_r [875] : 
                      (N212)? \piso.data_r [907] : 
                      (N214)? \piso.data_r [939] : 
                      (N216)? \piso.data_r [971] : 
                      (N218)? \piso.data_r [1003] : 
                      (N220)? \piso.data_r [1035] : 
                      (N222)? \piso.data_r [1067] : 
                      (N224)? \piso.data_r [1099] : 
                      (N226)? \piso.data_r [1131] : 
                      (N228)? \piso.data_r [1163] : 
                      (N230)? \piso.data_r [1195] : 
                      (N232)? \piso.data_r [1227] : 
                      (N234)? \piso.data_r [1259] : 
                      (N236)? \piso.data_r [1291] : 
                      (N238)? \piso.data_r [1323] : 
                      (N240)? \piso.data_r [1355] : 
                      (N242)? \piso.data_r [1387] : 
                      (N244)? \piso.data_r [1419] : 
                      (N246)? \piso.data_r [1451] : 
                      (N248)? \piso.data_r [1483] : 
                      (N250)? \piso.data_r [1515] : 
                      (N252)? \piso.data_r [1547] : 
                      (N254)? \piso.data_r [1579] : 
                      (N256)? \piso.data_r [1611] : 
                      (N258)? \piso.data_r [1643] : 
                      (N260)? \piso.data_r [1675] : 
                      (N262)? \piso.data_r [1707] : 
                      (N264)? \piso.data_r [1739] : 
                      (N266)? \piso.data_r [1771] : 
                      (N268)? \piso.data_r [1803] : 
                      (N270)? \piso.data_r [1835] : 
                      (N272)? \piso.data_r [1867] : 
                      (N274)? \piso.data_r [1899] : 
                      (N276)? \piso.data_r [1931] : 
                      (N278)? \piso.data_r [1963] : 
                      (N280)? \piso.data_r [1995] : 
                      (N282)? \piso.data_r [2027] : 
                      (N157)? \piso.data_r [2059] : 
                      (N159)? \piso.data_r [2091] : 
                      (N161)? \piso.data_r [2123] : 
                      (N163)? \piso.data_r [2155] : 
                      (N165)? \piso.data_r [2187] : 
                      (N167)? \piso.data_r [2219] : 
                      (N169)? \piso.data_r [2251] : 
                      (N171)? \piso.data_r [2283] : 
                      (N173)? \piso.data_r [2315] : 
                      (N175)? \piso.data_r [2347] : 
                      (N177)? \piso.data_r [2379] : 
                      (N179)? \piso.data_r [2411] : 
                      (N181)? \piso.data_r [2443] : 
                      (N183)? \piso.data_r [2475] : 
                      (N185)? \piso.data_r [2507] : 
                      (N187)? \piso.data_r [2539] : 
                      (N189)? \piso.data_r [2571] : 
                      (N191)? \piso.data_r [2603] : 
                      (N193)? \piso.data_r [2635] : 
                      (N195)? \piso.data_r [2667] : 
                      (N197)? \piso.data_r [2699] : 
                      (N199)? \piso.data_r [2731] : 
                      (N201)? \piso.data_r [2763] : 
                      (N203)? \piso.data_r [2795] : 
                      (N205)? \piso.data_r [2827] : 
                      (N207)? \piso.data_r [2859] : 
                      (N209)? \piso.data_r [2891] : 
                      (N211)? \piso.data_r [2923] : 
                      (N213)? \piso.data_r [2955] : 
                      (N215)? \piso.data_r [2987] : 
                      (N217)? \piso.data_r [3019] : 
                      (N219)? \piso.data_r [3051] : 
                      (N221)? \piso.data_r [3083] : 
                      (N223)? \piso.data_r [3115] : 
                      (N225)? \piso.data_r [3147] : 
                      (N227)? \piso.data_r [3179] : 
                      (N229)? \piso.data_r [3211] : 
                      (N231)? \piso.data_r [3243] : 
                      (N233)? \piso.data_r [3275] : 
                      (N235)? \piso.data_r [3307] : 
                      (N237)? \piso.data_r [3339] : 
                      (N239)? \piso.data_r [3371] : 
                      (N241)? \piso.data_r [3403] : 
                      (N243)? \piso.data_r [3435] : 
                      (N245)? \piso.data_r [3467] : 
                      (N247)? \piso.data_r [3499] : 
                      (N249)? \piso.data_r [3531] : 
                      (N251)? \piso.data_r [3563] : 
                      (N253)? \piso.data_r [3595] : 
                      (N255)? \piso.data_r [3627] : 
                      (N257)? \piso.data_r [3659] : 
                      (N259)? \piso.data_r [3691] : 
                      (N261)? \piso.data_r [3723] : 
                      (N263)? \piso.data_r [3755] : 
                      (N265)? \piso.data_r [3787] : 
                      (N267)? \piso.data_r [3819] : 
                      (N269)? \piso.data_r [3851] : 
                      (N271)? \piso.data_r [3883] : 
                      (N273)? \piso.data_r [3915] : 
                      (N275)? \piso.data_r [3947] : 
                      (N277)? \piso.data_r [3979] : 
                      (N279)? \piso.data_r [4011] : 
                      (N281)? \piso.data_r [4043] : 
                      (N283)? \piso.data_r [4075] : 1'b0;
  assign data_o[10] = (N156)? \piso.data_r [10] : 
                      (N158)? \piso.data_r [42] : 
                      (N160)? \piso.data_r [74] : 
                      (N162)? \piso.data_r [106] : 
                      (N164)? \piso.data_r [138] : 
                      (N166)? \piso.data_r [170] : 
                      (N168)? \piso.data_r [202] : 
                      (N170)? \piso.data_r [234] : 
                      (N172)? \piso.data_r [266] : 
                      (N174)? \piso.data_r [298] : 
                      (N176)? \piso.data_r [330] : 
                      (N178)? \piso.data_r [362] : 
                      (N180)? \piso.data_r [394] : 
                      (N182)? \piso.data_r [426] : 
                      (N184)? \piso.data_r [458] : 
                      (N186)? \piso.data_r [490] : 
                      (N188)? \piso.data_r [522] : 
                      (N190)? \piso.data_r [554] : 
                      (N192)? \piso.data_r [586] : 
                      (N194)? \piso.data_r [618] : 
                      (N196)? \piso.data_r [650] : 
                      (N198)? \piso.data_r [682] : 
                      (N200)? \piso.data_r [714] : 
                      (N202)? \piso.data_r [746] : 
                      (N204)? \piso.data_r [778] : 
                      (N206)? \piso.data_r [810] : 
                      (N208)? \piso.data_r [842] : 
                      (N210)? \piso.data_r [874] : 
                      (N212)? \piso.data_r [906] : 
                      (N214)? \piso.data_r [938] : 
                      (N216)? \piso.data_r [970] : 
                      (N218)? \piso.data_r [1002] : 
                      (N220)? \piso.data_r [1034] : 
                      (N222)? \piso.data_r [1066] : 
                      (N224)? \piso.data_r [1098] : 
                      (N226)? \piso.data_r [1130] : 
                      (N228)? \piso.data_r [1162] : 
                      (N230)? \piso.data_r [1194] : 
                      (N232)? \piso.data_r [1226] : 
                      (N234)? \piso.data_r [1258] : 
                      (N236)? \piso.data_r [1290] : 
                      (N238)? \piso.data_r [1322] : 
                      (N240)? \piso.data_r [1354] : 
                      (N242)? \piso.data_r [1386] : 
                      (N244)? \piso.data_r [1418] : 
                      (N246)? \piso.data_r [1450] : 
                      (N248)? \piso.data_r [1482] : 
                      (N250)? \piso.data_r [1514] : 
                      (N252)? \piso.data_r [1546] : 
                      (N254)? \piso.data_r [1578] : 
                      (N256)? \piso.data_r [1610] : 
                      (N258)? \piso.data_r [1642] : 
                      (N260)? \piso.data_r [1674] : 
                      (N262)? \piso.data_r [1706] : 
                      (N264)? \piso.data_r [1738] : 
                      (N266)? \piso.data_r [1770] : 
                      (N268)? \piso.data_r [1802] : 
                      (N270)? \piso.data_r [1834] : 
                      (N272)? \piso.data_r [1866] : 
                      (N274)? \piso.data_r [1898] : 
                      (N276)? \piso.data_r [1930] : 
                      (N278)? \piso.data_r [1962] : 
                      (N280)? \piso.data_r [1994] : 
                      (N282)? \piso.data_r [2026] : 
                      (N157)? \piso.data_r [2058] : 
                      (N159)? \piso.data_r [2090] : 
                      (N161)? \piso.data_r [2122] : 
                      (N163)? \piso.data_r [2154] : 
                      (N165)? \piso.data_r [2186] : 
                      (N167)? \piso.data_r [2218] : 
                      (N169)? \piso.data_r [2250] : 
                      (N171)? \piso.data_r [2282] : 
                      (N173)? \piso.data_r [2314] : 
                      (N175)? \piso.data_r [2346] : 
                      (N177)? \piso.data_r [2378] : 
                      (N179)? \piso.data_r [2410] : 
                      (N181)? \piso.data_r [2442] : 
                      (N183)? \piso.data_r [2474] : 
                      (N185)? \piso.data_r [2506] : 
                      (N187)? \piso.data_r [2538] : 
                      (N189)? \piso.data_r [2570] : 
                      (N191)? \piso.data_r [2602] : 
                      (N193)? \piso.data_r [2634] : 
                      (N195)? \piso.data_r [2666] : 
                      (N197)? \piso.data_r [2698] : 
                      (N199)? \piso.data_r [2730] : 
                      (N201)? \piso.data_r [2762] : 
                      (N203)? \piso.data_r [2794] : 
                      (N205)? \piso.data_r [2826] : 
                      (N207)? \piso.data_r [2858] : 
                      (N209)? \piso.data_r [2890] : 
                      (N211)? \piso.data_r [2922] : 
                      (N213)? \piso.data_r [2954] : 
                      (N215)? \piso.data_r [2986] : 
                      (N217)? \piso.data_r [3018] : 
                      (N219)? \piso.data_r [3050] : 
                      (N221)? \piso.data_r [3082] : 
                      (N223)? \piso.data_r [3114] : 
                      (N225)? \piso.data_r [3146] : 
                      (N227)? \piso.data_r [3178] : 
                      (N229)? \piso.data_r [3210] : 
                      (N231)? \piso.data_r [3242] : 
                      (N233)? \piso.data_r [3274] : 
                      (N235)? \piso.data_r [3306] : 
                      (N237)? \piso.data_r [3338] : 
                      (N239)? \piso.data_r [3370] : 
                      (N241)? \piso.data_r [3402] : 
                      (N243)? \piso.data_r [3434] : 
                      (N245)? \piso.data_r [3466] : 
                      (N247)? \piso.data_r [3498] : 
                      (N249)? \piso.data_r [3530] : 
                      (N251)? \piso.data_r [3562] : 
                      (N253)? \piso.data_r [3594] : 
                      (N255)? \piso.data_r [3626] : 
                      (N257)? \piso.data_r [3658] : 
                      (N259)? \piso.data_r [3690] : 
                      (N261)? \piso.data_r [3722] : 
                      (N263)? \piso.data_r [3754] : 
                      (N265)? \piso.data_r [3786] : 
                      (N267)? \piso.data_r [3818] : 
                      (N269)? \piso.data_r [3850] : 
                      (N271)? \piso.data_r [3882] : 
                      (N273)? \piso.data_r [3914] : 
                      (N275)? \piso.data_r [3946] : 
                      (N277)? \piso.data_r [3978] : 
                      (N279)? \piso.data_r [4010] : 
                      (N281)? \piso.data_r [4042] : 
                      (N283)? \piso.data_r [4074] : 1'b0;
  assign data_o[9] = (N156)? \piso.data_r [9] : 
                     (N158)? \piso.data_r [41] : 
                     (N160)? \piso.data_r [73] : 
                     (N162)? \piso.data_r [105] : 
                     (N164)? \piso.data_r [137] : 
                     (N166)? \piso.data_r [169] : 
                     (N168)? \piso.data_r [201] : 
                     (N170)? \piso.data_r [233] : 
                     (N172)? \piso.data_r [265] : 
                     (N174)? \piso.data_r [297] : 
                     (N176)? \piso.data_r [329] : 
                     (N178)? \piso.data_r [361] : 
                     (N180)? \piso.data_r [393] : 
                     (N182)? \piso.data_r [425] : 
                     (N184)? \piso.data_r [457] : 
                     (N186)? \piso.data_r [489] : 
                     (N188)? \piso.data_r [521] : 
                     (N190)? \piso.data_r [553] : 
                     (N192)? \piso.data_r [585] : 
                     (N194)? \piso.data_r [617] : 
                     (N196)? \piso.data_r [649] : 
                     (N198)? \piso.data_r [681] : 
                     (N200)? \piso.data_r [713] : 
                     (N202)? \piso.data_r [745] : 
                     (N204)? \piso.data_r [777] : 
                     (N206)? \piso.data_r [809] : 
                     (N208)? \piso.data_r [841] : 
                     (N210)? \piso.data_r [873] : 
                     (N212)? \piso.data_r [905] : 
                     (N214)? \piso.data_r [937] : 
                     (N216)? \piso.data_r [969] : 
                     (N218)? \piso.data_r [1001] : 
                     (N220)? \piso.data_r [1033] : 
                     (N222)? \piso.data_r [1065] : 
                     (N224)? \piso.data_r [1097] : 
                     (N226)? \piso.data_r [1129] : 
                     (N228)? \piso.data_r [1161] : 
                     (N230)? \piso.data_r [1193] : 
                     (N232)? \piso.data_r [1225] : 
                     (N234)? \piso.data_r [1257] : 
                     (N236)? \piso.data_r [1289] : 
                     (N238)? \piso.data_r [1321] : 
                     (N240)? \piso.data_r [1353] : 
                     (N242)? \piso.data_r [1385] : 
                     (N244)? \piso.data_r [1417] : 
                     (N246)? \piso.data_r [1449] : 
                     (N248)? \piso.data_r [1481] : 
                     (N250)? \piso.data_r [1513] : 
                     (N252)? \piso.data_r [1545] : 
                     (N254)? \piso.data_r [1577] : 
                     (N256)? \piso.data_r [1609] : 
                     (N258)? \piso.data_r [1641] : 
                     (N260)? \piso.data_r [1673] : 
                     (N262)? \piso.data_r [1705] : 
                     (N264)? \piso.data_r [1737] : 
                     (N266)? \piso.data_r [1769] : 
                     (N268)? \piso.data_r [1801] : 
                     (N270)? \piso.data_r [1833] : 
                     (N272)? \piso.data_r [1865] : 
                     (N274)? \piso.data_r [1897] : 
                     (N276)? \piso.data_r [1929] : 
                     (N278)? \piso.data_r [1961] : 
                     (N280)? \piso.data_r [1993] : 
                     (N282)? \piso.data_r [2025] : 
                     (N157)? \piso.data_r [2057] : 
                     (N159)? \piso.data_r [2089] : 
                     (N161)? \piso.data_r [2121] : 
                     (N163)? \piso.data_r [2153] : 
                     (N165)? \piso.data_r [2185] : 
                     (N167)? \piso.data_r [2217] : 
                     (N169)? \piso.data_r [2249] : 
                     (N171)? \piso.data_r [2281] : 
                     (N173)? \piso.data_r [2313] : 
                     (N175)? \piso.data_r [2345] : 
                     (N177)? \piso.data_r [2377] : 
                     (N179)? \piso.data_r [2409] : 
                     (N181)? \piso.data_r [2441] : 
                     (N183)? \piso.data_r [2473] : 
                     (N185)? \piso.data_r [2505] : 
                     (N187)? \piso.data_r [2537] : 
                     (N189)? \piso.data_r [2569] : 
                     (N191)? \piso.data_r [2601] : 
                     (N193)? \piso.data_r [2633] : 
                     (N195)? \piso.data_r [2665] : 
                     (N197)? \piso.data_r [2697] : 
                     (N199)? \piso.data_r [2729] : 
                     (N201)? \piso.data_r [2761] : 
                     (N203)? \piso.data_r [2793] : 
                     (N205)? \piso.data_r [2825] : 
                     (N207)? \piso.data_r [2857] : 
                     (N209)? \piso.data_r [2889] : 
                     (N211)? \piso.data_r [2921] : 
                     (N213)? \piso.data_r [2953] : 
                     (N215)? \piso.data_r [2985] : 
                     (N217)? \piso.data_r [3017] : 
                     (N219)? \piso.data_r [3049] : 
                     (N221)? \piso.data_r [3081] : 
                     (N223)? \piso.data_r [3113] : 
                     (N225)? \piso.data_r [3145] : 
                     (N227)? \piso.data_r [3177] : 
                     (N229)? \piso.data_r [3209] : 
                     (N231)? \piso.data_r [3241] : 
                     (N233)? \piso.data_r [3273] : 
                     (N235)? \piso.data_r [3305] : 
                     (N237)? \piso.data_r [3337] : 
                     (N239)? \piso.data_r [3369] : 
                     (N241)? \piso.data_r [3401] : 
                     (N243)? \piso.data_r [3433] : 
                     (N245)? \piso.data_r [3465] : 
                     (N247)? \piso.data_r [3497] : 
                     (N249)? \piso.data_r [3529] : 
                     (N251)? \piso.data_r [3561] : 
                     (N253)? \piso.data_r [3593] : 
                     (N255)? \piso.data_r [3625] : 
                     (N257)? \piso.data_r [3657] : 
                     (N259)? \piso.data_r [3689] : 
                     (N261)? \piso.data_r [3721] : 
                     (N263)? \piso.data_r [3753] : 
                     (N265)? \piso.data_r [3785] : 
                     (N267)? \piso.data_r [3817] : 
                     (N269)? \piso.data_r [3849] : 
                     (N271)? \piso.data_r [3881] : 
                     (N273)? \piso.data_r [3913] : 
                     (N275)? \piso.data_r [3945] : 
                     (N277)? \piso.data_r [3977] : 
                     (N279)? \piso.data_r [4009] : 
                     (N281)? \piso.data_r [4041] : 
                     (N283)? \piso.data_r [4073] : 1'b0;
  assign data_o[8] = (N156)? \piso.data_r [8] : 
                     (N158)? \piso.data_r [40] : 
                     (N160)? \piso.data_r [72] : 
                     (N162)? \piso.data_r [104] : 
                     (N164)? \piso.data_r [136] : 
                     (N166)? \piso.data_r [168] : 
                     (N168)? \piso.data_r [200] : 
                     (N170)? \piso.data_r [232] : 
                     (N172)? \piso.data_r [264] : 
                     (N174)? \piso.data_r [296] : 
                     (N176)? \piso.data_r [328] : 
                     (N178)? \piso.data_r [360] : 
                     (N180)? \piso.data_r [392] : 
                     (N182)? \piso.data_r [424] : 
                     (N184)? \piso.data_r [456] : 
                     (N186)? \piso.data_r [488] : 
                     (N188)? \piso.data_r [520] : 
                     (N190)? \piso.data_r [552] : 
                     (N192)? \piso.data_r [584] : 
                     (N194)? \piso.data_r [616] : 
                     (N196)? \piso.data_r [648] : 
                     (N198)? \piso.data_r [680] : 
                     (N200)? \piso.data_r [712] : 
                     (N202)? \piso.data_r [744] : 
                     (N204)? \piso.data_r [776] : 
                     (N206)? \piso.data_r [808] : 
                     (N208)? \piso.data_r [840] : 
                     (N210)? \piso.data_r [872] : 
                     (N212)? \piso.data_r [904] : 
                     (N214)? \piso.data_r [936] : 
                     (N216)? \piso.data_r [968] : 
                     (N218)? \piso.data_r [1000] : 
                     (N220)? \piso.data_r [1032] : 
                     (N222)? \piso.data_r [1064] : 
                     (N224)? \piso.data_r [1096] : 
                     (N226)? \piso.data_r [1128] : 
                     (N228)? \piso.data_r [1160] : 
                     (N230)? \piso.data_r [1192] : 
                     (N232)? \piso.data_r [1224] : 
                     (N234)? \piso.data_r [1256] : 
                     (N236)? \piso.data_r [1288] : 
                     (N238)? \piso.data_r [1320] : 
                     (N240)? \piso.data_r [1352] : 
                     (N242)? \piso.data_r [1384] : 
                     (N244)? \piso.data_r [1416] : 
                     (N246)? \piso.data_r [1448] : 
                     (N248)? \piso.data_r [1480] : 
                     (N250)? \piso.data_r [1512] : 
                     (N252)? \piso.data_r [1544] : 
                     (N254)? \piso.data_r [1576] : 
                     (N256)? \piso.data_r [1608] : 
                     (N258)? \piso.data_r [1640] : 
                     (N260)? \piso.data_r [1672] : 
                     (N262)? \piso.data_r [1704] : 
                     (N264)? \piso.data_r [1736] : 
                     (N266)? \piso.data_r [1768] : 
                     (N268)? \piso.data_r [1800] : 
                     (N270)? \piso.data_r [1832] : 
                     (N272)? \piso.data_r [1864] : 
                     (N274)? \piso.data_r [1896] : 
                     (N276)? \piso.data_r [1928] : 
                     (N278)? \piso.data_r [1960] : 
                     (N280)? \piso.data_r [1992] : 
                     (N282)? \piso.data_r [2024] : 
                     (N157)? \piso.data_r [2056] : 
                     (N159)? \piso.data_r [2088] : 
                     (N161)? \piso.data_r [2120] : 
                     (N163)? \piso.data_r [2152] : 
                     (N165)? \piso.data_r [2184] : 
                     (N167)? \piso.data_r [2216] : 
                     (N169)? \piso.data_r [2248] : 
                     (N171)? \piso.data_r [2280] : 
                     (N173)? \piso.data_r [2312] : 
                     (N175)? \piso.data_r [2344] : 
                     (N177)? \piso.data_r [2376] : 
                     (N179)? \piso.data_r [2408] : 
                     (N181)? \piso.data_r [2440] : 
                     (N183)? \piso.data_r [2472] : 
                     (N185)? \piso.data_r [2504] : 
                     (N187)? \piso.data_r [2536] : 
                     (N189)? \piso.data_r [2568] : 
                     (N191)? \piso.data_r [2600] : 
                     (N193)? \piso.data_r [2632] : 
                     (N195)? \piso.data_r [2664] : 
                     (N197)? \piso.data_r [2696] : 
                     (N199)? \piso.data_r [2728] : 
                     (N201)? \piso.data_r [2760] : 
                     (N203)? \piso.data_r [2792] : 
                     (N205)? \piso.data_r [2824] : 
                     (N207)? \piso.data_r [2856] : 
                     (N209)? \piso.data_r [2888] : 
                     (N211)? \piso.data_r [2920] : 
                     (N213)? \piso.data_r [2952] : 
                     (N215)? \piso.data_r [2984] : 
                     (N217)? \piso.data_r [3016] : 
                     (N219)? \piso.data_r [3048] : 
                     (N221)? \piso.data_r [3080] : 
                     (N223)? \piso.data_r [3112] : 
                     (N225)? \piso.data_r [3144] : 
                     (N227)? \piso.data_r [3176] : 
                     (N229)? \piso.data_r [3208] : 
                     (N231)? \piso.data_r [3240] : 
                     (N233)? \piso.data_r [3272] : 
                     (N235)? \piso.data_r [3304] : 
                     (N237)? \piso.data_r [3336] : 
                     (N239)? \piso.data_r [3368] : 
                     (N241)? \piso.data_r [3400] : 
                     (N243)? \piso.data_r [3432] : 
                     (N245)? \piso.data_r [3464] : 
                     (N247)? \piso.data_r [3496] : 
                     (N249)? \piso.data_r [3528] : 
                     (N251)? \piso.data_r [3560] : 
                     (N253)? \piso.data_r [3592] : 
                     (N255)? \piso.data_r [3624] : 
                     (N257)? \piso.data_r [3656] : 
                     (N259)? \piso.data_r [3688] : 
                     (N261)? \piso.data_r [3720] : 
                     (N263)? \piso.data_r [3752] : 
                     (N265)? \piso.data_r [3784] : 
                     (N267)? \piso.data_r [3816] : 
                     (N269)? \piso.data_r [3848] : 
                     (N271)? \piso.data_r [3880] : 
                     (N273)? \piso.data_r [3912] : 
                     (N275)? \piso.data_r [3944] : 
                     (N277)? \piso.data_r [3976] : 
                     (N279)? \piso.data_r [4008] : 
                     (N281)? \piso.data_r [4040] : 
                     (N283)? \piso.data_r [4072] : 1'b0;
  assign data_o[7] = (N156)? \piso.data_r [7] : 
                     (N158)? \piso.data_r [39] : 
                     (N160)? \piso.data_r [71] : 
                     (N162)? \piso.data_r [103] : 
                     (N164)? \piso.data_r [135] : 
                     (N166)? \piso.data_r [167] : 
                     (N168)? \piso.data_r [199] : 
                     (N170)? \piso.data_r [231] : 
                     (N172)? \piso.data_r [263] : 
                     (N174)? \piso.data_r [295] : 
                     (N176)? \piso.data_r [327] : 
                     (N178)? \piso.data_r [359] : 
                     (N180)? \piso.data_r [391] : 
                     (N182)? \piso.data_r [423] : 
                     (N184)? \piso.data_r [455] : 
                     (N186)? \piso.data_r [487] : 
                     (N188)? \piso.data_r [519] : 
                     (N190)? \piso.data_r [551] : 
                     (N192)? \piso.data_r [583] : 
                     (N194)? \piso.data_r [615] : 
                     (N196)? \piso.data_r [647] : 
                     (N198)? \piso.data_r [679] : 
                     (N200)? \piso.data_r [711] : 
                     (N202)? \piso.data_r [743] : 
                     (N204)? \piso.data_r [775] : 
                     (N206)? \piso.data_r [807] : 
                     (N208)? \piso.data_r [839] : 
                     (N210)? \piso.data_r [871] : 
                     (N212)? \piso.data_r [903] : 
                     (N214)? \piso.data_r [935] : 
                     (N216)? \piso.data_r [967] : 
                     (N218)? \piso.data_r [999] : 
                     (N220)? \piso.data_r [1031] : 
                     (N222)? \piso.data_r [1063] : 
                     (N224)? \piso.data_r [1095] : 
                     (N226)? \piso.data_r [1127] : 
                     (N228)? \piso.data_r [1159] : 
                     (N230)? \piso.data_r [1191] : 
                     (N232)? \piso.data_r [1223] : 
                     (N234)? \piso.data_r [1255] : 
                     (N236)? \piso.data_r [1287] : 
                     (N238)? \piso.data_r [1319] : 
                     (N240)? \piso.data_r [1351] : 
                     (N242)? \piso.data_r [1383] : 
                     (N244)? \piso.data_r [1415] : 
                     (N246)? \piso.data_r [1447] : 
                     (N248)? \piso.data_r [1479] : 
                     (N250)? \piso.data_r [1511] : 
                     (N252)? \piso.data_r [1543] : 
                     (N254)? \piso.data_r [1575] : 
                     (N256)? \piso.data_r [1607] : 
                     (N258)? \piso.data_r [1639] : 
                     (N260)? \piso.data_r [1671] : 
                     (N262)? \piso.data_r [1703] : 
                     (N264)? \piso.data_r [1735] : 
                     (N266)? \piso.data_r [1767] : 
                     (N268)? \piso.data_r [1799] : 
                     (N270)? \piso.data_r [1831] : 
                     (N272)? \piso.data_r [1863] : 
                     (N274)? \piso.data_r [1895] : 
                     (N276)? \piso.data_r [1927] : 
                     (N278)? \piso.data_r [1959] : 
                     (N280)? \piso.data_r [1991] : 
                     (N282)? \piso.data_r [2023] : 
                     (N157)? \piso.data_r [2055] : 
                     (N159)? \piso.data_r [2087] : 
                     (N161)? \piso.data_r [2119] : 
                     (N163)? \piso.data_r [2151] : 
                     (N165)? \piso.data_r [2183] : 
                     (N167)? \piso.data_r [2215] : 
                     (N169)? \piso.data_r [2247] : 
                     (N171)? \piso.data_r [2279] : 
                     (N173)? \piso.data_r [2311] : 
                     (N175)? \piso.data_r [2343] : 
                     (N177)? \piso.data_r [2375] : 
                     (N179)? \piso.data_r [2407] : 
                     (N181)? \piso.data_r [2439] : 
                     (N183)? \piso.data_r [2471] : 
                     (N185)? \piso.data_r [2503] : 
                     (N187)? \piso.data_r [2535] : 
                     (N189)? \piso.data_r [2567] : 
                     (N191)? \piso.data_r [2599] : 
                     (N193)? \piso.data_r [2631] : 
                     (N195)? \piso.data_r [2663] : 
                     (N197)? \piso.data_r [2695] : 
                     (N199)? \piso.data_r [2727] : 
                     (N201)? \piso.data_r [2759] : 
                     (N203)? \piso.data_r [2791] : 
                     (N205)? \piso.data_r [2823] : 
                     (N207)? \piso.data_r [2855] : 
                     (N209)? \piso.data_r [2887] : 
                     (N211)? \piso.data_r [2919] : 
                     (N213)? \piso.data_r [2951] : 
                     (N215)? \piso.data_r [2983] : 
                     (N217)? \piso.data_r [3015] : 
                     (N219)? \piso.data_r [3047] : 
                     (N221)? \piso.data_r [3079] : 
                     (N223)? \piso.data_r [3111] : 
                     (N225)? \piso.data_r [3143] : 
                     (N227)? \piso.data_r [3175] : 
                     (N229)? \piso.data_r [3207] : 
                     (N231)? \piso.data_r [3239] : 
                     (N233)? \piso.data_r [3271] : 
                     (N235)? \piso.data_r [3303] : 
                     (N237)? \piso.data_r [3335] : 
                     (N239)? \piso.data_r [3367] : 
                     (N241)? \piso.data_r [3399] : 
                     (N243)? \piso.data_r [3431] : 
                     (N245)? \piso.data_r [3463] : 
                     (N247)? \piso.data_r [3495] : 
                     (N249)? \piso.data_r [3527] : 
                     (N251)? \piso.data_r [3559] : 
                     (N253)? \piso.data_r [3591] : 
                     (N255)? \piso.data_r [3623] : 
                     (N257)? \piso.data_r [3655] : 
                     (N259)? \piso.data_r [3687] : 
                     (N261)? \piso.data_r [3719] : 
                     (N263)? \piso.data_r [3751] : 
                     (N265)? \piso.data_r [3783] : 
                     (N267)? \piso.data_r [3815] : 
                     (N269)? \piso.data_r [3847] : 
                     (N271)? \piso.data_r [3879] : 
                     (N273)? \piso.data_r [3911] : 
                     (N275)? \piso.data_r [3943] : 
                     (N277)? \piso.data_r [3975] : 
                     (N279)? \piso.data_r [4007] : 
                     (N281)? \piso.data_r [4039] : 
                     (N283)? \piso.data_r [4071] : 1'b0;
  assign data_o[6] = (N156)? \piso.data_r [6] : 
                     (N158)? \piso.data_r [38] : 
                     (N160)? \piso.data_r [70] : 
                     (N162)? \piso.data_r [102] : 
                     (N164)? \piso.data_r [134] : 
                     (N166)? \piso.data_r [166] : 
                     (N168)? \piso.data_r [198] : 
                     (N170)? \piso.data_r [230] : 
                     (N172)? \piso.data_r [262] : 
                     (N174)? \piso.data_r [294] : 
                     (N176)? \piso.data_r [326] : 
                     (N178)? \piso.data_r [358] : 
                     (N180)? \piso.data_r [390] : 
                     (N182)? \piso.data_r [422] : 
                     (N184)? \piso.data_r [454] : 
                     (N186)? \piso.data_r [486] : 
                     (N188)? \piso.data_r [518] : 
                     (N190)? \piso.data_r [550] : 
                     (N192)? \piso.data_r [582] : 
                     (N194)? \piso.data_r [614] : 
                     (N196)? \piso.data_r [646] : 
                     (N198)? \piso.data_r [678] : 
                     (N200)? \piso.data_r [710] : 
                     (N202)? \piso.data_r [742] : 
                     (N204)? \piso.data_r [774] : 
                     (N206)? \piso.data_r [806] : 
                     (N208)? \piso.data_r [838] : 
                     (N210)? \piso.data_r [870] : 
                     (N212)? \piso.data_r [902] : 
                     (N214)? \piso.data_r [934] : 
                     (N216)? \piso.data_r [966] : 
                     (N218)? \piso.data_r [998] : 
                     (N220)? \piso.data_r [1030] : 
                     (N222)? \piso.data_r [1062] : 
                     (N224)? \piso.data_r [1094] : 
                     (N226)? \piso.data_r [1126] : 
                     (N228)? \piso.data_r [1158] : 
                     (N230)? \piso.data_r [1190] : 
                     (N232)? \piso.data_r [1222] : 
                     (N234)? \piso.data_r [1254] : 
                     (N236)? \piso.data_r [1286] : 
                     (N238)? \piso.data_r [1318] : 
                     (N240)? \piso.data_r [1350] : 
                     (N242)? \piso.data_r [1382] : 
                     (N244)? \piso.data_r [1414] : 
                     (N246)? \piso.data_r [1446] : 
                     (N248)? \piso.data_r [1478] : 
                     (N250)? \piso.data_r [1510] : 
                     (N252)? \piso.data_r [1542] : 
                     (N254)? \piso.data_r [1574] : 
                     (N256)? \piso.data_r [1606] : 
                     (N258)? \piso.data_r [1638] : 
                     (N260)? \piso.data_r [1670] : 
                     (N262)? \piso.data_r [1702] : 
                     (N264)? \piso.data_r [1734] : 
                     (N266)? \piso.data_r [1766] : 
                     (N268)? \piso.data_r [1798] : 
                     (N270)? \piso.data_r [1830] : 
                     (N272)? \piso.data_r [1862] : 
                     (N274)? \piso.data_r [1894] : 
                     (N276)? \piso.data_r [1926] : 
                     (N278)? \piso.data_r [1958] : 
                     (N280)? \piso.data_r [1990] : 
                     (N282)? \piso.data_r [2022] : 
                     (N157)? \piso.data_r [2054] : 
                     (N159)? \piso.data_r [2086] : 
                     (N161)? \piso.data_r [2118] : 
                     (N163)? \piso.data_r [2150] : 
                     (N165)? \piso.data_r [2182] : 
                     (N167)? \piso.data_r [2214] : 
                     (N169)? \piso.data_r [2246] : 
                     (N171)? \piso.data_r [2278] : 
                     (N173)? \piso.data_r [2310] : 
                     (N175)? \piso.data_r [2342] : 
                     (N177)? \piso.data_r [2374] : 
                     (N179)? \piso.data_r [2406] : 
                     (N181)? \piso.data_r [2438] : 
                     (N183)? \piso.data_r [2470] : 
                     (N185)? \piso.data_r [2502] : 
                     (N187)? \piso.data_r [2534] : 
                     (N189)? \piso.data_r [2566] : 
                     (N191)? \piso.data_r [2598] : 
                     (N193)? \piso.data_r [2630] : 
                     (N195)? \piso.data_r [2662] : 
                     (N197)? \piso.data_r [2694] : 
                     (N199)? \piso.data_r [2726] : 
                     (N201)? \piso.data_r [2758] : 
                     (N203)? \piso.data_r [2790] : 
                     (N205)? \piso.data_r [2822] : 
                     (N207)? \piso.data_r [2854] : 
                     (N209)? \piso.data_r [2886] : 
                     (N211)? \piso.data_r [2918] : 
                     (N213)? \piso.data_r [2950] : 
                     (N215)? \piso.data_r [2982] : 
                     (N217)? \piso.data_r [3014] : 
                     (N219)? \piso.data_r [3046] : 
                     (N221)? \piso.data_r [3078] : 
                     (N223)? \piso.data_r [3110] : 
                     (N225)? \piso.data_r [3142] : 
                     (N227)? \piso.data_r [3174] : 
                     (N229)? \piso.data_r [3206] : 
                     (N231)? \piso.data_r [3238] : 
                     (N233)? \piso.data_r [3270] : 
                     (N235)? \piso.data_r [3302] : 
                     (N237)? \piso.data_r [3334] : 
                     (N239)? \piso.data_r [3366] : 
                     (N241)? \piso.data_r [3398] : 
                     (N243)? \piso.data_r [3430] : 
                     (N245)? \piso.data_r [3462] : 
                     (N247)? \piso.data_r [3494] : 
                     (N249)? \piso.data_r [3526] : 
                     (N251)? \piso.data_r [3558] : 
                     (N253)? \piso.data_r [3590] : 
                     (N255)? \piso.data_r [3622] : 
                     (N257)? \piso.data_r [3654] : 
                     (N259)? \piso.data_r [3686] : 
                     (N261)? \piso.data_r [3718] : 
                     (N263)? \piso.data_r [3750] : 
                     (N265)? \piso.data_r [3782] : 
                     (N267)? \piso.data_r [3814] : 
                     (N269)? \piso.data_r [3846] : 
                     (N271)? \piso.data_r [3878] : 
                     (N273)? \piso.data_r [3910] : 
                     (N275)? \piso.data_r [3942] : 
                     (N277)? \piso.data_r [3974] : 
                     (N279)? \piso.data_r [4006] : 
                     (N281)? \piso.data_r [4038] : 
                     (N283)? \piso.data_r [4070] : 1'b0;
  assign data_o[5] = (N156)? \piso.data_r [5] : 
                     (N158)? \piso.data_r [37] : 
                     (N160)? \piso.data_r [69] : 
                     (N162)? \piso.data_r [101] : 
                     (N164)? \piso.data_r [133] : 
                     (N166)? \piso.data_r [165] : 
                     (N168)? \piso.data_r [197] : 
                     (N170)? \piso.data_r [229] : 
                     (N172)? \piso.data_r [261] : 
                     (N174)? \piso.data_r [293] : 
                     (N176)? \piso.data_r [325] : 
                     (N178)? \piso.data_r [357] : 
                     (N180)? \piso.data_r [389] : 
                     (N182)? \piso.data_r [421] : 
                     (N184)? \piso.data_r [453] : 
                     (N186)? \piso.data_r [485] : 
                     (N188)? \piso.data_r [517] : 
                     (N190)? \piso.data_r [549] : 
                     (N192)? \piso.data_r [581] : 
                     (N194)? \piso.data_r [613] : 
                     (N196)? \piso.data_r [645] : 
                     (N198)? \piso.data_r [677] : 
                     (N200)? \piso.data_r [709] : 
                     (N202)? \piso.data_r [741] : 
                     (N204)? \piso.data_r [773] : 
                     (N206)? \piso.data_r [805] : 
                     (N208)? \piso.data_r [837] : 
                     (N210)? \piso.data_r [869] : 
                     (N212)? \piso.data_r [901] : 
                     (N214)? \piso.data_r [933] : 
                     (N216)? \piso.data_r [965] : 
                     (N218)? \piso.data_r [997] : 
                     (N220)? \piso.data_r [1029] : 
                     (N222)? \piso.data_r [1061] : 
                     (N224)? \piso.data_r [1093] : 
                     (N226)? \piso.data_r [1125] : 
                     (N228)? \piso.data_r [1157] : 
                     (N230)? \piso.data_r [1189] : 
                     (N232)? \piso.data_r [1221] : 
                     (N234)? \piso.data_r [1253] : 
                     (N236)? \piso.data_r [1285] : 
                     (N238)? \piso.data_r [1317] : 
                     (N240)? \piso.data_r [1349] : 
                     (N242)? \piso.data_r [1381] : 
                     (N244)? \piso.data_r [1413] : 
                     (N246)? \piso.data_r [1445] : 
                     (N248)? \piso.data_r [1477] : 
                     (N250)? \piso.data_r [1509] : 
                     (N252)? \piso.data_r [1541] : 
                     (N254)? \piso.data_r [1573] : 
                     (N256)? \piso.data_r [1605] : 
                     (N258)? \piso.data_r [1637] : 
                     (N260)? \piso.data_r [1669] : 
                     (N262)? \piso.data_r [1701] : 
                     (N264)? \piso.data_r [1733] : 
                     (N266)? \piso.data_r [1765] : 
                     (N268)? \piso.data_r [1797] : 
                     (N270)? \piso.data_r [1829] : 
                     (N272)? \piso.data_r [1861] : 
                     (N274)? \piso.data_r [1893] : 
                     (N276)? \piso.data_r [1925] : 
                     (N278)? \piso.data_r [1957] : 
                     (N280)? \piso.data_r [1989] : 
                     (N282)? \piso.data_r [2021] : 
                     (N157)? \piso.data_r [2053] : 
                     (N159)? \piso.data_r [2085] : 
                     (N161)? \piso.data_r [2117] : 
                     (N163)? \piso.data_r [2149] : 
                     (N165)? \piso.data_r [2181] : 
                     (N167)? \piso.data_r [2213] : 
                     (N169)? \piso.data_r [2245] : 
                     (N171)? \piso.data_r [2277] : 
                     (N173)? \piso.data_r [2309] : 
                     (N175)? \piso.data_r [2341] : 
                     (N177)? \piso.data_r [2373] : 
                     (N179)? \piso.data_r [2405] : 
                     (N181)? \piso.data_r [2437] : 
                     (N183)? \piso.data_r [2469] : 
                     (N185)? \piso.data_r [2501] : 
                     (N187)? \piso.data_r [2533] : 
                     (N189)? \piso.data_r [2565] : 
                     (N191)? \piso.data_r [2597] : 
                     (N193)? \piso.data_r [2629] : 
                     (N195)? \piso.data_r [2661] : 
                     (N197)? \piso.data_r [2693] : 
                     (N199)? \piso.data_r [2725] : 
                     (N201)? \piso.data_r [2757] : 
                     (N203)? \piso.data_r [2789] : 
                     (N205)? \piso.data_r [2821] : 
                     (N207)? \piso.data_r [2853] : 
                     (N209)? \piso.data_r [2885] : 
                     (N211)? \piso.data_r [2917] : 
                     (N213)? \piso.data_r [2949] : 
                     (N215)? \piso.data_r [2981] : 
                     (N217)? \piso.data_r [3013] : 
                     (N219)? \piso.data_r [3045] : 
                     (N221)? \piso.data_r [3077] : 
                     (N223)? \piso.data_r [3109] : 
                     (N225)? \piso.data_r [3141] : 
                     (N227)? \piso.data_r [3173] : 
                     (N229)? \piso.data_r [3205] : 
                     (N231)? \piso.data_r [3237] : 
                     (N233)? \piso.data_r [3269] : 
                     (N235)? \piso.data_r [3301] : 
                     (N237)? \piso.data_r [3333] : 
                     (N239)? \piso.data_r [3365] : 
                     (N241)? \piso.data_r [3397] : 
                     (N243)? \piso.data_r [3429] : 
                     (N245)? \piso.data_r [3461] : 
                     (N247)? \piso.data_r [3493] : 
                     (N249)? \piso.data_r [3525] : 
                     (N251)? \piso.data_r [3557] : 
                     (N253)? \piso.data_r [3589] : 
                     (N255)? \piso.data_r [3621] : 
                     (N257)? \piso.data_r [3653] : 
                     (N259)? \piso.data_r [3685] : 
                     (N261)? \piso.data_r [3717] : 
                     (N263)? \piso.data_r [3749] : 
                     (N265)? \piso.data_r [3781] : 
                     (N267)? \piso.data_r [3813] : 
                     (N269)? \piso.data_r [3845] : 
                     (N271)? \piso.data_r [3877] : 
                     (N273)? \piso.data_r [3909] : 
                     (N275)? \piso.data_r [3941] : 
                     (N277)? \piso.data_r [3973] : 
                     (N279)? \piso.data_r [4005] : 
                     (N281)? \piso.data_r [4037] : 
                     (N283)? \piso.data_r [4069] : 1'b0;
  assign data_o[4] = (N156)? \piso.data_r [4] : 
                     (N158)? \piso.data_r [36] : 
                     (N160)? \piso.data_r [68] : 
                     (N162)? \piso.data_r [100] : 
                     (N164)? \piso.data_r [132] : 
                     (N166)? \piso.data_r [164] : 
                     (N168)? \piso.data_r [196] : 
                     (N170)? \piso.data_r [228] : 
                     (N172)? \piso.data_r [260] : 
                     (N174)? \piso.data_r [292] : 
                     (N176)? \piso.data_r [324] : 
                     (N178)? \piso.data_r [356] : 
                     (N180)? \piso.data_r [388] : 
                     (N182)? \piso.data_r [420] : 
                     (N184)? \piso.data_r [452] : 
                     (N186)? \piso.data_r [484] : 
                     (N188)? \piso.data_r [516] : 
                     (N190)? \piso.data_r [548] : 
                     (N192)? \piso.data_r [580] : 
                     (N194)? \piso.data_r [612] : 
                     (N196)? \piso.data_r [644] : 
                     (N198)? \piso.data_r [676] : 
                     (N200)? \piso.data_r [708] : 
                     (N202)? \piso.data_r [740] : 
                     (N204)? \piso.data_r [772] : 
                     (N206)? \piso.data_r [804] : 
                     (N208)? \piso.data_r [836] : 
                     (N210)? \piso.data_r [868] : 
                     (N212)? \piso.data_r [900] : 
                     (N214)? \piso.data_r [932] : 
                     (N216)? \piso.data_r [964] : 
                     (N218)? \piso.data_r [996] : 
                     (N220)? \piso.data_r [1028] : 
                     (N222)? \piso.data_r [1060] : 
                     (N224)? \piso.data_r [1092] : 
                     (N226)? \piso.data_r [1124] : 
                     (N228)? \piso.data_r [1156] : 
                     (N230)? \piso.data_r [1188] : 
                     (N232)? \piso.data_r [1220] : 
                     (N234)? \piso.data_r [1252] : 
                     (N236)? \piso.data_r [1284] : 
                     (N238)? \piso.data_r [1316] : 
                     (N240)? \piso.data_r [1348] : 
                     (N242)? \piso.data_r [1380] : 
                     (N244)? \piso.data_r [1412] : 
                     (N246)? \piso.data_r [1444] : 
                     (N248)? \piso.data_r [1476] : 
                     (N250)? \piso.data_r [1508] : 
                     (N252)? \piso.data_r [1540] : 
                     (N254)? \piso.data_r [1572] : 
                     (N256)? \piso.data_r [1604] : 
                     (N258)? \piso.data_r [1636] : 
                     (N260)? \piso.data_r [1668] : 
                     (N262)? \piso.data_r [1700] : 
                     (N264)? \piso.data_r [1732] : 
                     (N266)? \piso.data_r [1764] : 
                     (N268)? \piso.data_r [1796] : 
                     (N270)? \piso.data_r [1828] : 
                     (N272)? \piso.data_r [1860] : 
                     (N274)? \piso.data_r [1892] : 
                     (N276)? \piso.data_r [1924] : 
                     (N278)? \piso.data_r [1956] : 
                     (N280)? \piso.data_r [1988] : 
                     (N282)? \piso.data_r [2020] : 
                     (N157)? \piso.data_r [2052] : 
                     (N159)? \piso.data_r [2084] : 
                     (N161)? \piso.data_r [2116] : 
                     (N163)? \piso.data_r [2148] : 
                     (N165)? \piso.data_r [2180] : 
                     (N167)? \piso.data_r [2212] : 
                     (N169)? \piso.data_r [2244] : 
                     (N171)? \piso.data_r [2276] : 
                     (N173)? \piso.data_r [2308] : 
                     (N175)? \piso.data_r [2340] : 
                     (N177)? \piso.data_r [2372] : 
                     (N179)? \piso.data_r [2404] : 
                     (N181)? \piso.data_r [2436] : 
                     (N183)? \piso.data_r [2468] : 
                     (N185)? \piso.data_r [2500] : 
                     (N187)? \piso.data_r [2532] : 
                     (N189)? \piso.data_r [2564] : 
                     (N191)? \piso.data_r [2596] : 
                     (N193)? \piso.data_r [2628] : 
                     (N195)? \piso.data_r [2660] : 
                     (N197)? \piso.data_r [2692] : 
                     (N199)? \piso.data_r [2724] : 
                     (N201)? \piso.data_r [2756] : 
                     (N203)? \piso.data_r [2788] : 
                     (N205)? \piso.data_r [2820] : 
                     (N207)? \piso.data_r [2852] : 
                     (N209)? \piso.data_r [2884] : 
                     (N211)? \piso.data_r [2916] : 
                     (N213)? \piso.data_r [2948] : 
                     (N215)? \piso.data_r [2980] : 
                     (N217)? \piso.data_r [3012] : 
                     (N219)? \piso.data_r [3044] : 
                     (N221)? \piso.data_r [3076] : 
                     (N223)? \piso.data_r [3108] : 
                     (N225)? \piso.data_r [3140] : 
                     (N227)? \piso.data_r [3172] : 
                     (N229)? \piso.data_r [3204] : 
                     (N231)? \piso.data_r [3236] : 
                     (N233)? \piso.data_r [3268] : 
                     (N235)? \piso.data_r [3300] : 
                     (N237)? \piso.data_r [3332] : 
                     (N239)? \piso.data_r [3364] : 
                     (N241)? \piso.data_r [3396] : 
                     (N243)? \piso.data_r [3428] : 
                     (N245)? \piso.data_r [3460] : 
                     (N247)? \piso.data_r [3492] : 
                     (N249)? \piso.data_r [3524] : 
                     (N251)? \piso.data_r [3556] : 
                     (N253)? \piso.data_r [3588] : 
                     (N255)? \piso.data_r [3620] : 
                     (N257)? \piso.data_r [3652] : 
                     (N259)? \piso.data_r [3684] : 
                     (N261)? \piso.data_r [3716] : 
                     (N263)? \piso.data_r [3748] : 
                     (N265)? \piso.data_r [3780] : 
                     (N267)? \piso.data_r [3812] : 
                     (N269)? \piso.data_r [3844] : 
                     (N271)? \piso.data_r [3876] : 
                     (N273)? \piso.data_r [3908] : 
                     (N275)? \piso.data_r [3940] : 
                     (N277)? \piso.data_r [3972] : 
                     (N279)? \piso.data_r [4004] : 
                     (N281)? \piso.data_r [4036] : 
                     (N283)? \piso.data_r [4068] : 1'b0;
  assign data_o[3] = (N156)? \piso.data_r [3] : 
                     (N158)? \piso.data_r [35] : 
                     (N160)? \piso.data_r [67] : 
                     (N162)? \piso.data_r [99] : 
                     (N164)? \piso.data_r [131] : 
                     (N166)? \piso.data_r [163] : 
                     (N168)? \piso.data_r [195] : 
                     (N170)? \piso.data_r [227] : 
                     (N172)? \piso.data_r [259] : 
                     (N174)? \piso.data_r [291] : 
                     (N176)? \piso.data_r [323] : 
                     (N178)? \piso.data_r [355] : 
                     (N180)? \piso.data_r [387] : 
                     (N182)? \piso.data_r [419] : 
                     (N184)? \piso.data_r [451] : 
                     (N186)? \piso.data_r [483] : 
                     (N188)? \piso.data_r [515] : 
                     (N190)? \piso.data_r [547] : 
                     (N192)? \piso.data_r [579] : 
                     (N194)? \piso.data_r [611] : 
                     (N196)? \piso.data_r [643] : 
                     (N198)? \piso.data_r [675] : 
                     (N200)? \piso.data_r [707] : 
                     (N202)? \piso.data_r [739] : 
                     (N204)? \piso.data_r [771] : 
                     (N206)? \piso.data_r [803] : 
                     (N208)? \piso.data_r [835] : 
                     (N210)? \piso.data_r [867] : 
                     (N212)? \piso.data_r [899] : 
                     (N214)? \piso.data_r [931] : 
                     (N216)? \piso.data_r [963] : 
                     (N218)? \piso.data_r [995] : 
                     (N220)? \piso.data_r [1027] : 
                     (N222)? \piso.data_r [1059] : 
                     (N224)? \piso.data_r [1091] : 
                     (N226)? \piso.data_r [1123] : 
                     (N228)? \piso.data_r [1155] : 
                     (N230)? \piso.data_r [1187] : 
                     (N232)? \piso.data_r [1219] : 
                     (N234)? \piso.data_r [1251] : 
                     (N236)? \piso.data_r [1283] : 
                     (N238)? \piso.data_r [1315] : 
                     (N240)? \piso.data_r [1347] : 
                     (N242)? \piso.data_r [1379] : 
                     (N244)? \piso.data_r [1411] : 
                     (N246)? \piso.data_r [1443] : 
                     (N248)? \piso.data_r [1475] : 
                     (N250)? \piso.data_r [1507] : 
                     (N252)? \piso.data_r [1539] : 
                     (N254)? \piso.data_r [1571] : 
                     (N256)? \piso.data_r [1603] : 
                     (N258)? \piso.data_r [1635] : 
                     (N260)? \piso.data_r [1667] : 
                     (N262)? \piso.data_r [1699] : 
                     (N264)? \piso.data_r [1731] : 
                     (N266)? \piso.data_r [1763] : 
                     (N268)? \piso.data_r [1795] : 
                     (N270)? \piso.data_r [1827] : 
                     (N272)? \piso.data_r [1859] : 
                     (N274)? \piso.data_r [1891] : 
                     (N276)? \piso.data_r [1923] : 
                     (N278)? \piso.data_r [1955] : 
                     (N280)? \piso.data_r [1987] : 
                     (N282)? \piso.data_r [2019] : 
                     (N157)? \piso.data_r [2051] : 
                     (N159)? \piso.data_r [2083] : 
                     (N161)? \piso.data_r [2115] : 
                     (N163)? \piso.data_r [2147] : 
                     (N165)? \piso.data_r [2179] : 
                     (N167)? \piso.data_r [2211] : 
                     (N169)? \piso.data_r [2243] : 
                     (N171)? \piso.data_r [2275] : 
                     (N173)? \piso.data_r [2307] : 
                     (N175)? \piso.data_r [2339] : 
                     (N177)? \piso.data_r [2371] : 
                     (N179)? \piso.data_r [2403] : 
                     (N181)? \piso.data_r [2435] : 
                     (N183)? \piso.data_r [2467] : 
                     (N185)? \piso.data_r [2499] : 
                     (N187)? \piso.data_r [2531] : 
                     (N189)? \piso.data_r [2563] : 
                     (N191)? \piso.data_r [2595] : 
                     (N193)? \piso.data_r [2627] : 
                     (N195)? \piso.data_r [2659] : 
                     (N197)? \piso.data_r [2691] : 
                     (N199)? \piso.data_r [2723] : 
                     (N201)? \piso.data_r [2755] : 
                     (N203)? \piso.data_r [2787] : 
                     (N205)? \piso.data_r [2819] : 
                     (N207)? \piso.data_r [2851] : 
                     (N209)? \piso.data_r [2883] : 
                     (N211)? \piso.data_r [2915] : 
                     (N213)? \piso.data_r [2947] : 
                     (N215)? \piso.data_r [2979] : 
                     (N217)? \piso.data_r [3011] : 
                     (N219)? \piso.data_r [3043] : 
                     (N221)? \piso.data_r [3075] : 
                     (N223)? \piso.data_r [3107] : 
                     (N225)? \piso.data_r [3139] : 
                     (N227)? \piso.data_r [3171] : 
                     (N229)? \piso.data_r [3203] : 
                     (N231)? \piso.data_r [3235] : 
                     (N233)? \piso.data_r [3267] : 
                     (N235)? \piso.data_r [3299] : 
                     (N237)? \piso.data_r [3331] : 
                     (N239)? \piso.data_r [3363] : 
                     (N241)? \piso.data_r [3395] : 
                     (N243)? \piso.data_r [3427] : 
                     (N245)? \piso.data_r [3459] : 
                     (N247)? \piso.data_r [3491] : 
                     (N249)? \piso.data_r [3523] : 
                     (N251)? \piso.data_r [3555] : 
                     (N253)? \piso.data_r [3587] : 
                     (N255)? \piso.data_r [3619] : 
                     (N257)? \piso.data_r [3651] : 
                     (N259)? \piso.data_r [3683] : 
                     (N261)? \piso.data_r [3715] : 
                     (N263)? \piso.data_r [3747] : 
                     (N265)? \piso.data_r [3779] : 
                     (N267)? \piso.data_r [3811] : 
                     (N269)? \piso.data_r [3843] : 
                     (N271)? \piso.data_r [3875] : 
                     (N273)? \piso.data_r [3907] : 
                     (N275)? \piso.data_r [3939] : 
                     (N277)? \piso.data_r [3971] : 
                     (N279)? \piso.data_r [4003] : 
                     (N281)? \piso.data_r [4035] : 
                     (N283)? \piso.data_r [4067] : 1'b0;
  assign data_o[2] = (N156)? \piso.data_r [2] : 
                     (N158)? \piso.data_r [34] : 
                     (N160)? \piso.data_r [66] : 
                     (N162)? \piso.data_r [98] : 
                     (N164)? \piso.data_r [130] : 
                     (N166)? \piso.data_r [162] : 
                     (N168)? \piso.data_r [194] : 
                     (N170)? \piso.data_r [226] : 
                     (N172)? \piso.data_r [258] : 
                     (N174)? \piso.data_r [290] : 
                     (N176)? \piso.data_r [322] : 
                     (N178)? \piso.data_r [354] : 
                     (N180)? \piso.data_r [386] : 
                     (N182)? \piso.data_r [418] : 
                     (N184)? \piso.data_r [450] : 
                     (N186)? \piso.data_r [482] : 
                     (N188)? \piso.data_r [514] : 
                     (N190)? \piso.data_r [546] : 
                     (N192)? \piso.data_r [578] : 
                     (N194)? \piso.data_r [610] : 
                     (N196)? \piso.data_r [642] : 
                     (N198)? \piso.data_r [674] : 
                     (N200)? \piso.data_r [706] : 
                     (N202)? \piso.data_r [738] : 
                     (N204)? \piso.data_r [770] : 
                     (N206)? \piso.data_r [802] : 
                     (N208)? \piso.data_r [834] : 
                     (N210)? \piso.data_r [866] : 
                     (N212)? \piso.data_r [898] : 
                     (N214)? \piso.data_r [930] : 
                     (N216)? \piso.data_r [962] : 
                     (N218)? \piso.data_r [994] : 
                     (N220)? \piso.data_r [1026] : 
                     (N222)? \piso.data_r [1058] : 
                     (N224)? \piso.data_r [1090] : 
                     (N226)? \piso.data_r [1122] : 
                     (N228)? \piso.data_r [1154] : 
                     (N230)? \piso.data_r [1186] : 
                     (N232)? \piso.data_r [1218] : 
                     (N234)? \piso.data_r [1250] : 
                     (N236)? \piso.data_r [1282] : 
                     (N238)? \piso.data_r [1314] : 
                     (N240)? \piso.data_r [1346] : 
                     (N242)? \piso.data_r [1378] : 
                     (N244)? \piso.data_r [1410] : 
                     (N246)? \piso.data_r [1442] : 
                     (N248)? \piso.data_r [1474] : 
                     (N250)? \piso.data_r [1506] : 
                     (N252)? \piso.data_r [1538] : 
                     (N254)? \piso.data_r [1570] : 
                     (N256)? \piso.data_r [1602] : 
                     (N258)? \piso.data_r [1634] : 
                     (N260)? \piso.data_r [1666] : 
                     (N262)? \piso.data_r [1698] : 
                     (N264)? \piso.data_r [1730] : 
                     (N266)? \piso.data_r [1762] : 
                     (N268)? \piso.data_r [1794] : 
                     (N270)? \piso.data_r [1826] : 
                     (N272)? \piso.data_r [1858] : 
                     (N274)? \piso.data_r [1890] : 
                     (N276)? \piso.data_r [1922] : 
                     (N278)? \piso.data_r [1954] : 
                     (N280)? \piso.data_r [1986] : 
                     (N282)? \piso.data_r [2018] : 
                     (N157)? \piso.data_r [2050] : 
                     (N159)? \piso.data_r [2082] : 
                     (N161)? \piso.data_r [2114] : 
                     (N163)? \piso.data_r [2146] : 
                     (N165)? \piso.data_r [2178] : 
                     (N167)? \piso.data_r [2210] : 
                     (N169)? \piso.data_r [2242] : 
                     (N171)? \piso.data_r [2274] : 
                     (N173)? \piso.data_r [2306] : 
                     (N175)? \piso.data_r [2338] : 
                     (N177)? \piso.data_r [2370] : 
                     (N179)? \piso.data_r [2402] : 
                     (N181)? \piso.data_r [2434] : 
                     (N183)? \piso.data_r [2466] : 
                     (N185)? \piso.data_r [2498] : 
                     (N187)? \piso.data_r [2530] : 
                     (N189)? \piso.data_r [2562] : 
                     (N191)? \piso.data_r [2594] : 
                     (N193)? \piso.data_r [2626] : 
                     (N195)? \piso.data_r [2658] : 
                     (N197)? \piso.data_r [2690] : 
                     (N199)? \piso.data_r [2722] : 
                     (N201)? \piso.data_r [2754] : 
                     (N203)? \piso.data_r [2786] : 
                     (N205)? \piso.data_r [2818] : 
                     (N207)? \piso.data_r [2850] : 
                     (N209)? \piso.data_r [2882] : 
                     (N211)? \piso.data_r [2914] : 
                     (N213)? \piso.data_r [2946] : 
                     (N215)? \piso.data_r [2978] : 
                     (N217)? \piso.data_r [3010] : 
                     (N219)? \piso.data_r [3042] : 
                     (N221)? \piso.data_r [3074] : 
                     (N223)? \piso.data_r [3106] : 
                     (N225)? \piso.data_r [3138] : 
                     (N227)? \piso.data_r [3170] : 
                     (N229)? \piso.data_r [3202] : 
                     (N231)? \piso.data_r [3234] : 
                     (N233)? \piso.data_r [3266] : 
                     (N235)? \piso.data_r [3298] : 
                     (N237)? \piso.data_r [3330] : 
                     (N239)? \piso.data_r [3362] : 
                     (N241)? \piso.data_r [3394] : 
                     (N243)? \piso.data_r [3426] : 
                     (N245)? \piso.data_r [3458] : 
                     (N247)? \piso.data_r [3490] : 
                     (N249)? \piso.data_r [3522] : 
                     (N251)? \piso.data_r [3554] : 
                     (N253)? \piso.data_r [3586] : 
                     (N255)? \piso.data_r [3618] : 
                     (N257)? \piso.data_r [3650] : 
                     (N259)? \piso.data_r [3682] : 
                     (N261)? \piso.data_r [3714] : 
                     (N263)? \piso.data_r [3746] : 
                     (N265)? \piso.data_r [3778] : 
                     (N267)? \piso.data_r [3810] : 
                     (N269)? \piso.data_r [3842] : 
                     (N271)? \piso.data_r [3874] : 
                     (N273)? \piso.data_r [3906] : 
                     (N275)? \piso.data_r [3938] : 
                     (N277)? \piso.data_r [3970] : 
                     (N279)? \piso.data_r [4002] : 
                     (N281)? \piso.data_r [4034] : 
                     (N283)? \piso.data_r [4066] : 1'b0;
  assign data_o[1] = (N156)? \piso.data_r [1] : 
                     (N158)? \piso.data_r [33] : 
                     (N160)? \piso.data_r [65] : 
                     (N162)? \piso.data_r [97] : 
                     (N164)? \piso.data_r [129] : 
                     (N166)? \piso.data_r [161] : 
                     (N168)? \piso.data_r [193] : 
                     (N170)? \piso.data_r [225] : 
                     (N172)? \piso.data_r [257] : 
                     (N174)? \piso.data_r [289] : 
                     (N176)? \piso.data_r [321] : 
                     (N178)? \piso.data_r [353] : 
                     (N180)? \piso.data_r [385] : 
                     (N182)? \piso.data_r [417] : 
                     (N184)? \piso.data_r [449] : 
                     (N186)? \piso.data_r [481] : 
                     (N188)? \piso.data_r [513] : 
                     (N190)? \piso.data_r [545] : 
                     (N192)? \piso.data_r [577] : 
                     (N194)? \piso.data_r [609] : 
                     (N196)? \piso.data_r [641] : 
                     (N198)? \piso.data_r [673] : 
                     (N200)? \piso.data_r [705] : 
                     (N202)? \piso.data_r [737] : 
                     (N204)? \piso.data_r [769] : 
                     (N206)? \piso.data_r [801] : 
                     (N208)? \piso.data_r [833] : 
                     (N210)? \piso.data_r [865] : 
                     (N212)? \piso.data_r [897] : 
                     (N214)? \piso.data_r [929] : 
                     (N216)? \piso.data_r [961] : 
                     (N218)? \piso.data_r [993] : 
                     (N220)? \piso.data_r [1025] : 
                     (N222)? \piso.data_r [1057] : 
                     (N224)? \piso.data_r [1089] : 
                     (N226)? \piso.data_r [1121] : 
                     (N228)? \piso.data_r [1153] : 
                     (N230)? \piso.data_r [1185] : 
                     (N232)? \piso.data_r [1217] : 
                     (N234)? \piso.data_r [1249] : 
                     (N236)? \piso.data_r [1281] : 
                     (N238)? \piso.data_r [1313] : 
                     (N240)? \piso.data_r [1345] : 
                     (N242)? \piso.data_r [1377] : 
                     (N244)? \piso.data_r [1409] : 
                     (N246)? \piso.data_r [1441] : 
                     (N248)? \piso.data_r [1473] : 
                     (N250)? \piso.data_r [1505] : 
                     (N252)? \piso.data_r [1537] : 
                     (N254)? \piso.data_r [1569] : 
                     (N256)? \piso.data_r [1601] : 
                     (N258)? \piso.data_r [1633] : 
                     (N260)? \piso.data_r [1665] : 
                     (N262)? \piso.data_r [1697] : 
                     (N264)? \piso.data_r [1729] : 
                     (N266)? \piso.data_r [1761] : 
                     (N268)? \piso.data_r [1793] : 
                     (N270)? \piso.data_r [1825] : 
                     (N272)? \piso.data_r [1857] : 
                     (N274)? \piso.data_r [1889] : 
                     (N276)? \piso.data_r [1921] : 
                     (N278)? \piso.data_r [1953] : 
                     (N280)? \piso.data_r [1985] : 
                     (N282)? \piso.data_r [2017] : 
                     (N157)? \piso.data_r [2049] : 
                     (N159)? \piso.data_r [2081] : 
                     (N161)? \piso.data_r [2113] : 
                     (N163)? \piso.data_r [2145] : 
                     (N165)? \piso.data_r [2177] : 
                     (N167)? \piso.data_r [2209] : 
                     (N169)? \piso.data_r [2241] : 
                     (N171)? \piso.data_r [2273] : 
                     (N173)? \piso.data_r [2305] : 
                     (N175)? \piso.data_r [2337] : 
                     (N177)? \piso.data_r [2369] : 
                     (N179)? \piso.data_r [2401] : 
                     (N181)? \piso.data_r [2433] : 
                     (N183)? \piso.data_r [2465] : 
                     (N185)? \piso.data_r [2497] : 
                     (N187)? \piso.data_r [2529] : 
                     (N189)? \piso.data_r [2561] : 
                     (N191)? \piso.data_r [2593] : 
                     (N193)? \piso.data_r [2625] : 
                     (N195)? \piso.data_r [2657] : 
                     (N197)? \piso.data_r [2689] : 
                     (N199)? \piso.data_r [2721] : 
                     (N201)? \piso.data_r [2753] : 
                     (N203)? \piso.data_r [2785] : 
                     (N205)? \piso.data_r [2817] : 
                     (N207)? \piso.data_r [2849] : 
                     (N209)? \piso.data_r [2881] : 
                     (N211)? \piso.data_r [2913] : 
                     (N213)? \piso.data_r [2945] : 
                     (N215)? \piso.data_r [2977] : 
                     (N217)? \piso.data_r [3009] : 
                     (N219)? \piso.data_r [3041] : 
                     (N221)? \piso.data_r [3073] : 
                     (N223)? \piso.data_r [3105] : 
                     (N225)? \piso.data_r [3137] : 
                     (N227)? \piso.data_r [3169] : 
                     (N229)? \piso.data_r [3201] : 
                     (N231)? \piso.data_r [3233] : 
                     (N233)? \piso.data_r [3265] : 
                     (N235)? \piso.data_r [3297] : 
                     (N237)? \piso.data_r [3329] : 
                     (N239)? \piso.data_r [3361] : 
                     (N241)? \piso.data_r [3393] : 
                     (N243)? \piso.data_r [3425] : 
                     (N245)? \piso.data_r [3457] : 
                     (N247)? \piso.data_r [3489] : 
                     (N249)? \piso.data_r [3521] : 
                     (N251)? \piso.data_r [3553] : 
                     (N253)? \piso.data_r [3585] : 
                     (N255)? \piso.data_r [3617] : 
                     (N257)? \piso.data_r [3649] : 
                     (N259)? \piso.data_r [3681] : 
                     (N261)? \piso.data_r [3713] : 
                     (N263)? \piso.data_r [3745] : 
                     (N265)? \piso.data_r [3777] : 
                     (N267)? \piso.data_r [3809] : 
                     (N269)? \piso.data_r [3841] : 
                     (N271)? \piso.data_r [3873] : 
                     (N273)? \piso.data_r [3905] : 
                     (N275)? \piso.data_r [3937] : 
                     (N277)? \piso.data_r [3969] : 
                     (N279)? \piso.data_r [4001] : 
                     (N281)? \piso.data_r [4033] : 
                     (N283)? \piso.data_r [4065] : 1'b0;
  assign data_o[0] = (N156)? \piso.data_r [0] : 
                     (N158)? \piso.data_r [32] : 
                     (N160)? \piso.data_r [64] : 
                     (N162)? \piso.data_r [96] : 
                     (N164)? \piso.data_r [128] : 
                     (N166)? \piso.data_r [160] : 
                     (N168)? \piso.data_r [192] : 
                     (N170)? \piso.data_r [224] : 
                     (N172)? \piso.data_r [256] : 
                     (N174)? \piso.data_r [288] : 
                     (N176)? \piso.data_r [320] : 
                     (N178)? \piso.data_r [352] : 
                     (N180)? \piso.data_r [384] : 
                     (N182)? \piso.data_r [416] : 
                     (N184)? \piso.data_r [448] : 
                     (N186)? \piso.data_r [480] : 
                     (N188)? \piso.data_r [512] : 
                     (N190)? \piso.data_r [544] : 
                     (N192)? \piso.data_r [576] : 
                     (N194)? \piso.data_r [608] : 
                     (N196)? \piso.data_r [640] : 
                     (N198)? \piso.data_r [672] : 
                     (N200)? \piso.data_r [704] : 
                     (N202)? \piso.data_r [736] : 
                     (N204)? \piso.data_r [768] : 
                     (N206)? \piso.data_r [800] : 
                     (N208)? \piso.data_r [832] : 
                     (N210)? \piso.data_r [864] : 
                     (N212)? \piso.data_r [896] : 
                     (N214)? \piso.data_r [928] : 
                     (N216)? \piso.data_r [960] : 
                     (N218)? \piso.data_r [992] : 
                     (N220)? \piso.data_r [1024] : 
                     (N222)? \piso.data_r [1056] : 
                     (N224)? \piso.data_r [1088] : 
                     (N226)? \piso.data_r [1120] : 
                     (N228)? \piso.data_r [1152] : 
                     (N230)? \piso.data_r [1184] : 
                     (N232)? \piso.data_r [1216] : 
                     (N234)? \piso.data_r [1248] : 
                     (N236)? \piso.data_r [1280] : 
                     (N238)? \piso.data_r [1312] : 
                     (N240)? \piso.data_r [1344] : 
                     (N242)? \piso.data_r [1376] : 
                     (N244)? \piso.data_r [1408] : 
                     (N246)? \piso.data_r [1440] : 
                     (N248)? \piso.data_r [1472] : 
                     (N250)? \piso.data_r [1504] : 
                     (N252)? \piso.data_r [1536] : 
                     (N254)? \piso.data_r [1568] : 
                     (N256)? \piso.data_r [1600] : 
                     (N258)? \piso.data_r [1632] : 
                     (N260)? \piso.data_r [1664] : 
                     (N262)? \piso.data_r [1696] : 
                     (N264)? \piso.data_r [1728] : 
                     (N266)? \piso.data_r [1760] : 
                     (N268)? \piso.data_r [1792] : 
                     (N270)? \piso.data_r [1824] : 
                     (N272)? \piso.data_r [1856] : 
                     (N274)? \piso.data_r [1888] : 
                     (N276)? \piso.data_r [1920] : 
                     (N278)? \piso.data_r [1952] : 
                     (N280)? \piso.data_r [1984] : 
                     (N282)? \piso.data_r [2016] : 
                     (N157)? \piso.data_r [2048] : 
                     (N159)? \piso.data_r [2080] : 
                     (N161)? \piso.data_r [2112] : 
                     (N163)? \piso.data_r [2144] : 
                     (N165)? \piso.data_r [2176] : 
                     (N167)? \piso.data_r [2208] : 
                     (N169)? \piso.data_r [2240] : 
                     (N171)? \piso.data_r [2272] : 
                     (N173)? \piso.data_r [2304] : 
                     (N175)? \piso.data_r [2336] : 
                     (N177)? \piso.data_r [2368] : 
                     (N179)? \piso.data_r [2400] : 
                     (N181)? \piso.data_r [2432] : 
                     (N183)? \piso.data_r [2464] : 
                     (N185)? \piso.data_r [2496] : 
                     (N187)? \piso.data_r [2528] : 
                     (N189)? \piso.data_r [2560] : 
                     (N191)? \piso.data_r [2592] : 
                     (N193)? \piso.data_r [2624] : 
                     (N195)? \piso.data_r [2656] : 
                     (N197)? \piso.data_r [2688] : 
                     (N199)? \piso.data_r [2720] : 
                     (N201)? \piso.data_r [2752] : 
                     (N203)? \piso.data_r [2784] : 
                     (N205)? \piso.data_r [2816] : 
                     (N207)? \piso.data_r [2848] : 
                     (N209)? \piso.data_r [2880] : 
                     (N211)? \piso.data_r [2912] : 
                     (N213)? \piso.data_r [2944] : 
                     (N215)? \piso.data_r [2976] : 
                     (N217)? \piso.data_r [3008] : 
                     (N219)? \piso.data_r [3040] : 
                     (N221)? \piso.data_r [3072] : 
                     (N223)? \piso.data_r [3104] : 
                     (N225)? \piso.data_r [3136] : 
                     (N227)? \piso.data_r [3168] : 
                     (N229)? \piso.data_r [3200] : 
                     (N231)? \piso.data_r [3232] : 
                     (N233)? \piso.data_r [3264] : 
                     (N235)? \piso.data_r [3296] : 
                     (N237)? \piso.data_r [3328] : 
                     (N239)? \piso.data_r [3360] : 
                     (N241)? \piso.data_r [3392] : 
                     (N243)? \piso.data_r [3424] : 
                     (N245)? \piso.data_r [3456] : 
                     (N247)? \piso.data_r [3488] : 
                     (N249)? \piso.data_r [3520] : 
                     (N251)? \piso.data_r [3552] : 
                     (N253)? \piso.data_r [3584] : 
                     (N255)? \piso.data_r [3616] : 
                     (N257)? \piso.data_r [3648] : 
                     (N259)? \piso.data_r [3680] : 
                     (N261)? \piso.data_r [3712] : 
                     (N263)? \piso.data_r [3744] : 
                     (N265)? \piso.data_r [3776] : 
                     (N267)? \piso.data_r [3808] : 
                     (N269)? \piso.data_r [3840] : 
                     (N271)? \piso.data_r [3872] : 
                     (N273)? \piso.data_r [3904] : 
                     (N275)? \piso.data_r [3936] : 
                     (N277)? \piso.data_r [3968] : 
                     (N279)? \piso.data_r [4000] : 
                     (N281)? \piso.data_r [4032] : 
                     (N283)? \piso.data_r [4064] : 1'b0;
  assign N286 = ~valid_o;
  assign N287 = \piso.shift_ctr_r [5] & \piso.shift_ctr_r [6];
  assign N288 = \piso.shift_ctr_r [4] & N287;
  assign N289 = \piso.shift_ctr_r [3] & N288;
  assign N290 = \piso.shift_ctr_r [2] & N289;
  assign N291 = \piso.shift_ctr_r [1] & N290;
  assign N292 = \piso.shift_ctr_r [0] & N291;
  assign { N24, N23, N22, N21, N20, N19, N18 } = \piso.shift_ctr_r  + 1'b1;
  assign \piso.state_n [0] = (N0)? 1'b1 : 
                             (N5)? 1'b0 : 1'b0;
  assign N0 = N2;
  assign { N15, N14, N13, N12, N11, N10, N9 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N8)? { N24, N23, N22, N21, N20, N19, N18 } : 1'b0;
  assign N1 = N7;
  assign \piso.done_tx_n  = N293 & yumi_i;
  assign N293 = valid_o & N292;
  assign ready_o = N286 | \piso.done_tx_n ;
  assign N2 = ready_o & valid_i;
  assign N3 = \piso.done_tx_n  | N2;
  assign N4 = ~N2;
  assign N5 = \piso.done_tx_n  & N4;
  assign N6 = ready_o & valid_i;
  assign N7 = ready_o & valid_i;
  assign N8 = ~N7;
  assign N16 = N294 & N295;
  assign N294 = valid_o & yumi_i;
  assign N295 = ~\piso.done_tx_n ;
  assign N17 = ~N16;
  assign N25 = ~\piso.shift_ctr_r [0];
  assign N26 = ~\piso.shift_ctr_r [1];
  assign N27 = N25 & N26;
  assign N28 = N25 & \piso.shift_ctr_r [1];
  assign N29 = \piso.shift_ctr_r [0] & N26;
  assign N30 = \piso.shift_ctr_r [0] & \piso.shift_ctr_r [1];
  assign N31 = ~\piso.shift_ctr_r [2];
  assign N32 = N27 & N31;
  assign N33 = N27 & \piso.shift_ctr_r [2];
  assign N34 = N29 & N31;
  assign N35 = N29 & \piso.shift_ctr_r [2];
  assign N36 = N28 & N31;
  assign N37 = N28 & \piso.shift_ctr_r [2];
  assign N38 = N30 & N31;
  assign N39 = N30 & \piso.shift_ctr_r [2];
  assign N40 = ~\piso.shift_ctr_r [3];
  assign N41 = N32 & N40;
  assign N42 = N32 & \piso.shift_ctr_r [3];
  assign N43 = N34 & N40;
  assign N44 = N34 & \piso.shift_ctr_r [3];
  assign N45 = N36 & N40;
  assign N46 = N36 & \piso.shift_ctr_r [3];
  assign N47 = N38 & N40;
  assign N48 = N38 & \piso.shift_ctr_r [3];
  assign N49 = N33 & N40;
  assign N50 = N33 & \piso.shift_ctr_r [3];
  assign N51 = N35 & N40;
  assign N52 = N35 & \piso.shift_ctr_r [3];
  assign N53 = N37 & N40;
  assign N54 = N37 & \piso.shift_ctr_r [3];
  assign N55 = N39 & N40;
  assign N56 = N39 & \piso.shift_ctr_r [3];
  assign N57 = ~\piso.shift_ctr_r [4];
  assign N58 = N41 & N57;
  assign N59 = N41 & \piso.shift_ctr_r [4];
  assign N60 = N43 & N57;
  assign N61 = N43 & \piso.shift_ctr_r [4];
  assign N62 = N45 & N57;
  assign N63 = N45 & \piso.shift_ctr_r [4];
  assign N64 = N47 & N57;
  assign N65 = N47 & \piso.shift_ctr_r [4];
  assign N66 = N49 & N57;
  assign N67 = N49 & \piso.shift_ctr_r [4];
  assign N68 = N51 & N57;
  assign N69 = N51 & \piso.shift_ctr_r [4];
  assign N70 = N53 & N57;
  assign N71 = N53 & \piso.shift_ctr_r [4];
  assign N72 = N55 & N57;
  assign N73 = N55 & \piso.shift_ctr_r [4];
  assign N74 = N42 & N57;
  assign N75 = N42 & \piso.shift_ctr_r [4];
  assign N76 = N44 & N57;
  assign N77 = N44 & \piso.shift_ctr_r [4];
  assign N78 = N46 & N57;
  assign N79 = N46 & \piso.shift_ctr_r [4];
  assign N80 = N48 & N57;
  assign N81 = N48 & \piso.shift_ctr_r [4];
  assign N82 = N50 & N57;
  assign N83 = N50 & \piso.shift_ctr_r [4];
  assign N84 = N52 & N57;
  assign N85 = N52 & \piso.shift_ctr_r [4];
  assign N86 = N54 & N57;
  assign N87 = N54 & \piso.shift_ctr_r [4];
  assign N88 = N56 & N57;
  assign N89 = N56 & \piso.shift_ctr_r [4];
  assign N90 = ~\piso.shift_ctr_r [5];
  assign N91 = N58 & N90;
  assign N92 = N58 & \piso.shift_ctr_r [5];
  assign N93 = N60 & N90;
  assign N94 = N60 & \piso.shift_ctr_r [5];
  assign N95 = N62 & N90;
  assign N96 = N62 & \piso.shift_ctr_r [5];
  assign N97 = N64 & N90;
  assign N98 = N64 & \piso.shift_ctr_r [5];
  assign N99 = N66 & N90;
  assign N100 = N66 & \piso.shift_ctr_r [5];
  assign N101 = N68 & N90;
  assign N102 = N68 & \piso.shift_ctr_r [5];
  assign N103 = N70 & N90;
  assign N104 = N70 & \piso.shift_ctr_r [5];
  assign N105 = N72 & N90;
  assign N106 = N72 & \piso.shift_ctr_r [5];
  assign N107 = N74 & N90;
  assign N108 = N74 & \piso.shift_ctr_r [5];
  assign N109 = N76 & N90;
  assign N110 = N76 & \piso.shift_ctr_r [5];
  assign N111 = N78 & N90;
  assign N112 = N78 & \piso.shift_ctr_r [5];
  assign N113 = N80 & N90;
  assign N114 = N80 & \piso.shift_ctr_r [5];
  assign N115 = N82 & N90;
  assign N116 = N82 & \piso.shift_ctr_r [5];
  assign N117 = N84 & N90;
  assign N118 = N84 & \piso.shift_ctr_r [5];
  assign N119 = N86 & N90;
  assign N120 = N86 & \piso.shift_ctr_r [5];
  assign N121 = N88 & N90;
  assign N122 = N88 & \piso.shift_ctr_r [5];
  assign N123 = N59 & N90;
  assign N124 = N59 & \piso.shift_ctr_r [5];
  assign N125 = N61 & N90;
  assign N126 = N61 & \piso.shift_ctr_r [5];
  assign N127 = N63 & N90;
  assign N128 = N63 & \piso.shift_ctr_r [5];
  assign N129 = N65 & N90;
  assign N130 = N65 & \piso.shift_ctr_r [5];
  assign N131 = N67 & N90;
  assign N132 = N67 & \piso.shift_ctr_r [5];
  assign N133 = N69 & N90;
  assign N134 = N69 & \piso.shift_ctr_r [5];
  assign N135 = N71 & N90;
  assign N136 = N71 & \piso.shift_ctr_r [5];
  assign N137 = N73 & N90;
  assign N138 = N73 & \piso.shift_ctr_r [5];
  assign N139 = N75 & N90;
  assign N140 = N75 & \piso.shift_ctr_r [5];
  assign N141 = N77 & N90;
  assign N142 = N77 & \piso.shift_ctr_r [5];
  assign N143 = N79 & N90;
  assign N144 = N79 & \piso.shift_ctr_r [5];
  assign N145 = N81 & N90;
  assign N146 = N81 & \piso.shift_ctr_r [5];
  assign N147 = N83 & N90;
  assign N148 = N83 & \piso.shift_ctr_r [5];
  assign N149 = N85 & N90;
  assign N150 = N85 & \piso.shift_ctr_r [5];
  assign N151 = N87 & N90;
  assign N152 = N87 & \piso.shift_ctr_r [5];
  assign N153 = N89 & N90;
  assign N154 = N89 & \piso.shift_ctr_r [5];
  assign N155 = ~\piso.shift_ctr_r [6];
  assign N156 = N91 & N155;
  assign N157 = N91 & \piso.shift_ctr_r [6];
  assign N158 = N93 & N155;
  assign N159 = N93 & \piso.shift_ctr_r [6];
  assign N160 = N95 & N155;
  assign N161 = N95 & \piso.shift_ctr_r [6];
  assign N162 = N97 & N155;
  assign N163 = N97 & \piso.shift_ctr_r [6];
  assign N164 = N99 & N155;
  assign N165 = N99 & \piso.shift_ctr_r [6];
  assign N166 = N101 & N155;
  assign N167 = N101 & \piso.shift_ctr_r [6];
  assign N168 = N103 & N155;
  assign N169 = N103 & \piso.shift_ctr_r [6];
  assign N170 = N105 & N155;
  assign N171 = N105 & \piso.shift_ctr_r [6];
  assign N172 = N107 & N155;
  assign N173 = N107 & \piso.shift_ctr_r [6];
  assign N174 = N109 & N155;
  assign N175 = N109 & \piso.shift_ctr_r [6];
  assign N176 = N111 & N155;
  assign N177 = N111 & \piso.shift_ctr_r [6];
  assign N178 = N113 & N155;
  assign N179 = N113 & \piso.shift_ctr_r [6];
  assign N180 = N115 & N155;
  assign N181 = N115 & \piso.shift_ctr_r [6];
  assign N182 = N117 & N155;
  assign N183 = N117 & \piso.shift_ctr_r [6];
  assign N184 = N119 & N155;
  assign N185 = N119 & \piso.shift_ctr_r [6];
  assign N186 = N121 & N155;
  assign N187 = N121 & \piso.shift_ctr_r [6];
  assign N188 = N123 & N155;
  assign N189 = N123 & \piso.shift_ctr_r [6];
  assign N190 = N125 & N155;
  assign N191 = N125 & \piso.shift_ctr_r [6];
  assign N192 = N127 & N155;
  assign N193 = N127 & \piso.shift_ctr_r [6];
  assign N194 = N129 & N155;
  assign N195 = N129 & \piso.shift_ctr_r [6];
  assign N196 = N131 & N155;
  assign N197 = N131 & \piso.shift_ctr_r [6];
  assign N198 = N133 & N155;
  assign N199 = N133 & \piso.shift_ctr_r [6];
  assign N200 = N135 & N155;
  assign N201 = N135 & \piso.shift_ctr_r [6];
  assign N202 = N137 & N155;
  assign N203 = N137 & \piso.shift_ctr_r [6];
  assign N204 = N139 & N155;
  assign N205 = N139 & \piso.shift_ctr_r [6];
  assign N206 = N141 & N155;
  assign N207 = N141 & \piso.shift_ctr_r [6];
  assign N208 = N143 & N155;
  assign N209 = N143 & \piso.shift_ctr_r [6];
  assign N210 = N145 & N155;
  assign N211 = N145 & \piso.shift_ctr_r [6];
  assign N212 = N147 & N155;
  assign N213 = N147 & \piso.shift_ctr_r [6];
  assign N214 = N149 & N155;
  assign N215 = N149 & \piso.shift_ctr_r [6];
  assign N216 = N151 & N155;
  assign N217 = N151 & \piso.shift_ctr_r [6];
  assign N218 = N153 & N155;
  assign N219 = N153 & \piso.shift_ctr_r [6];
  assign N220 = N92 & N155;
  assign N221 = N92 & \piso.shift_ctr_r [6];
  assign N222 = N94 & N155;
  assign N223 = N94 & \piso.shift_ctr_r [6];
  assign N224 = N96 & N155;
  assign N225 = N96 & \piso.shift_ctr_r [6];
  assign N226 = N98 & N155;
  assign N227 = N98 & \piso.shift_ctr_r [6];
  assign N228 = N100 & N155;
  assign N229 = N100 & \piso.shift_ctr_r [6];
  assign N230 = N102 & N155;
  assign N231 = N102 & \piso.shift_ctr_r [6];
  assign N232 = N104 & N155;
  assign N233 = N104 & \piso.shift_ctr_r [6];
  assign N234 = N106 & N155;
  assign N235 = N106 & \piso.shift_ctr_r [6];
  assign N236 = N108 & N155;
  assign N237 = N108 & \piso.shift_ctr_r [6];
  assign N238 = N110 & N155;
  assign N239 = N110 & \piso.shift_ctr_r [6];
  assign N240 = N112 & N155;
  assign N241 = N112 & \piso.shift_ctr_r [6];
  assign N242 = N114 & N155;
  assign N243 = N114 & \piso.shift_ctr_r [6];
  assign N244 = N116 & N155;
  assign N245 = N116 & \piso.shift_ctr_r [6];
  assign N246 = N118 & N155;
  assign N247 = N118 & \piso.shift_ctr_r [6];
  assign N248 = N120 & N155;
  assign N249 = N120 & \piso.shift_ctr_r [6];
  assign N250 = N122 & N155;
  assign N251 = N122 & \piso.shift_ctr_r [6];
  assign N252 = N124 & N155;
  assign N253 = N124 & \piso.shift_ctr_r [6];
  assign N254 = N126 & N155;
  assign N255 = N126 & \piso.shift_ctr_r [6];
  assign N256 = N128 & N155;
  assign N257 = N128 & \piso.shift_ctr_r [6];
  assign N258 = N130 & N155;
  assign N259 = N130 & \piso.shift_ctr_r [6];
  assign N260 = N132 & N155;
  assign N261 = N132 & \piso.shift_ctr_r [6];
  assign N262 = N134 & N155;
  assign N263 = N134 & \piso.shift_ctr_r [6];
  assign N264 = N136 & N155;
  assign N265 = N136 & \piso.shift_ctr_r [6];
  assign N266 = N138 & N155;
  assign N267 = N138 & \piso.shift_ctr_r [6];
  assign N268 = N140 & N155;
  assign N269 = N140 & \piso.shift_ctr_r [6];
  assign N270 = N142 & N155;
  assign N271 = N142 & \piso.shift_ctr_r [6];
  assign N272 = N144 & N155;
  assign N273 = N144 & \piso.shift_ctr_r [6];
  assign N274 = N146 & N155;
  assign N275 = N146 & \piso.shift_ctr_r [6];
  assign N276 = N148 & N155;
  assign N277 = N148 & \piso.shift_ctr_r [6];
  assign N278 = N150 & N155;
  assign N279 = N150 & \piso.shift_ctr_r [6];
  assign N280 = N152 & N155;
  assign N281 = N152 & \piso.shift_ctr_r [6];
  assign N282 = N154 & N155;
  assign N283 = N154 & \piso.shift_ctr_r [6];
  assign N284 = N17 & N8;
  assign N285 = ~N284;

  always @(posedge clk_i) begin
    if(reset_i) begin
      valid_o_sv2v_reg <= 1'b0;
    end else if(N3) begin
      valid_o_sv2v_reg <= \piso.state_n [0];
    end 
    if(reset_i) begin
      \piso.data_r_4095_sv2v_reg  <= 1'b0;
      \piso.data_r_4094_sv2v_reg  <= 1'b0;
      \piso.data_r_4093_sv2v_reg  <= 1'b0;
      \piso.data_r_4092_sv2v_reg  <= 1'b0;
      \piso.data_r_4091_sv2v_reg  <= 1'b0;
      \piso.data_r_4090_sv2v_reg  <= 1'b0;
      \piso.data_r_4089_sv2v_reg  <= 1'b0;
      \piso.data_r_4088_sv2v_reg  <= 1'b0;
      \piso.data_r_4087_sv2v_reg  <= 1'b0;
      \piso.data_r_4086_sv2v_reg  <= 1'b0;
      \piso.data_r_4085_sv2v_reg  <= 1'b0;
      \piso.data_r_4084_sv2v_reg  <= 1'b0;
      \piso.data_r_4083_sv2v_reg  <= 1'b0;
      \piso.data_r_4082_sv2v_reg  <= 1'b0;
      \piso.data_r_4081_sv2v_reg  <= 1'b0;
      \piso.data_r_4080_sv2v_reg  <= 1'b0;
      \piso.data_r_4079_sv2v_reg  <= 1'b0;
      \piso.data_r_4078_sv2v_reg  <= 1'b0;
      \piso.data_r_4077_sv2v_reg  <= 1'b0;
      \piso.data_r_4076_sv2v_reg  <= 1'b0;
      \piso.data_r_4075_sv2v_reg  <= 1'b0;
      \piso.data_r_4074_sv2v_reg  <= 1'b0;
      \piso.data_r_4073_sv2v_reg  <= 1'b0;
      \piso.data_r_4072_sv2v_reg  <= 1'b0;
      \piso.data_r_4071_sv2v_reg  <= 1'b0;
      \piso.data_r_4070_sv2v_reg  <= 1'b0;
      \piso.data_r_4069_sv2v_reg  <= 1'b0;
      \piso.data_r_4068_sv2v_reg  <= 1'b0;
      \piso.data_r_4067_sv2v_reg  <= 1'b0;
      \piso.data_r_4066_sv2v_reg  <= 1'b0;
      \piso.data_r_4065_sv2v_reg  <= 1'b0;
      \piso.data_r_4064_sv2v_reg  <= 1'b0;
      \piso.data_r_4063_sv2v_reg  <= 1'b0;
      \piso.data_r_4062_sv2v_reg  <= 1'b0;
      \piso.data_r_4061_sv2v_reg  <= 1'b0;
      \piso.data_r_4060_sv2v_reg  <= 1'b0;
      \piso.data_r_4059_sv2v_reg  <= 1'b0;
      \piso.data_r_4058_sv2v_reg  <= 1'b0;
      \piso.data_r_4057_sv2v_reg  <= 1'b0;
      \piso.data_r_4056_sv2v_reg  <= 1'b0;
      \piso.data_r_4055_sv2v_reg  <= 1'b0;
      \piso.data_r_4054_sv2v_reg  <= 1'b0;
      \piso.data_r_4053_sv2v_reg  <= 1'b0;
      \piso.data_r_4052_sv2v_reg  <= 1'b0;
      \piso.data_r_4051_sv2v_reg  <= 1'b0;
      \piso.data_r_4050_sv2v_reg  <= 1'b0;
      \piso.data_r_4049_sv2v_reg  <= 1'b0;
      \piso.data_r_4048_sv2v_reg  <= 1'b0;
      \piso.data_r_4047_sv2v_reg  <= 1'b0;
      \piso.data_r_4046_sv2v_reg  <= 1'b0;
      \piso.data_r_4045_sv2v_reg  <= 1'b0;
      \piso.data_r_4044_sv2v_reg  <= 1'b0;
      \piso.data_r_4043_sv2v_reg  <= 1'b0;
      \piso.data_r_4042_sv2v_reg  <= 1'b0;
      \piso.data_r_4041_sv2v_reg  <= 1'b0;
      \piso.data_r_4040_sv2v_reg  <= 1'b0;
      \piso.data_r_4039_sv2v_reg  <= 1'b0;
      \piso.data_r_4038_sv2v_reg  <= 1'b0;
      \piso.data_r_4037_sv2v_reg  <= 1'b0;
      \piso.data_r_4036_sv2v_reg  <= 1'b0;
      \piso.data_r_4035_sv2v_reg  <= 1'b0;
      \piso.data_r_4034_sv2v_reg  <= 1'b0;
      \piso.data_r_4033_sv2v_reg  <= 1'b0;
      \piso.data_r_4032_sv2v_reg  <= 1'b0;
      \piso.data_r_4031_sv2v_reg  <= 1'b0;
      \piso.data_r_4030_sv2v_reg  <= 1'b0;
      \piso.data_r_4029_sv2v_reg  <= 1'b0;
      \piso.data_r_4028_sv2v_reg  <= 1'b0;
      \piso.data_r_4027_sv2v_reg  <= 1'b0;
      \piso.data_r_4026_sv2v_reg  <= 1'b0;
      \piso.data_r_4025_sv2v_reg  <= 1'b0;
      \piso.data_r_4024_sv2v_reg  <= 1'b0;
      \piso.data_r_4023_sv2v_reg  <= 1'b0;
      \piso.data_r_4022_sv2v_reg  <= 1'b0;
      \piso.data_r_4021_sv2v_reg  <= 1'b0;
      \piso.data_r_4020_sv2v_reg  <= 1'b0;
      \piso.data_r_4019_sv2v_reg  <= 1'b0;
      \piso.data_r_4018_sv2v_reg  <= 1'b0;
      \piso.data_r_4017_sv2v_reg  <= 1'b0;
      \piso.data_r_4016_sv2v_reg  <= 1'b0;
      \piso.data_r_4015_sv2v_reg  <= 1'b0;
      \piso.data_r_4014_sv2v_reg  <= 1'b0;
      \piso.data_r_4013_sv2v_reg  <= 1'b0;
      \piso.data_r_4012_sv2v_reg  <= 1'b0;
      \piso.data_r_4011_sv2v_reg  <= 1'b0;
      \piso.data_r_4010_sv2v_reg  <= 1'b0;
      \piso.data_r_4009_sv2v_reg  <= 1'b0;
      \piso.data_r_4008_sv2v_reg  <= 1'b0;
      \piso.data_r_4007_sv2v_reg  <= 1'b0;
      \piso.data_r_4006_sv2v_reg  <= 1'b0;
      \piso.data_r_4005_sv2v_reg  <= 1'b0;
      \piso.data_r_4004_sv2v_reg  <= 1'b0;
      \piso.data_r_4003_sv2v_reg  <= 1'b0;
      \piso.data_r_4002_sv2v_reg  <= 1'b0;
      \piso.data_r_4001_sv2v_reg  <= 1'b0;
      \piso.data_r_4000_sv2v_reg  <= 1'b0;
      \piso.data_r_3999_sv2v_reg  <= 1'b0;
      \piso.data_r_3998_sv2v_reg  <= 1'b0;
      \piso.data_r_3997_sv2v_reg  <= 1'b0;
      \piso.data_r_3996_sv2v_reg  <= 1'b0;
      \piso.data_r_3995_sv2v_reg  <= 1'b0;
      \piso.data_r_3994_sv2v_reg  <= 1'b0;
      \piso.data_r_3993_sv2v_reg  <= 1'b0;
      \piso.data_r_3992_sv2v_reg  <= 1'b0;
      \piso.data_r_3991_sv2v_reg  <= 1'b0;
      \piso.data_r_3990_sv2v_reg  <= 1'b0;
      \piso.data_r_3989_sv2v_reg  <= 1'b0;
      \piso.data_r_3988_sv2v_reg  <= 1'b0;
      \piso.data_r_3987_sv2v_reg  <= 1'b0;
      \piso.data_r_3986_sv2v_reg  <= 1'b0;
      \piso.data_r_3985_sv2v_reg  <= 1'b0;
      \piso.data_r_3984_sv2v_reg  <= 1'b0;
      \piso.data_r_3983_sv2v_reg  <= 1'b0;
      \piso.data_r_3982_sv2v_reg  <= 1'b0;
      \piso.data_r_3981_sv2v_reg  <= 1'b0;
      \piso.data_r_3980_sv2v_reg  <= 1'b0;
      \piso.data_r_3979_sv2v_reg  <= 1'b0;
      \piso.data_r_3978_sv2v_reg  <= 1'b0;
      \piso.data_r_3977_sv2v_reg  <= 1'b0;
      \piso.data_r_3976_sv2v_reg  <= 1'b0;
      \piso.data_r_3975_sv2v_reg  <= 1'b0;
      \piso.data_r_3974_sv2v_reg  <= 1'b0;
      \piso.data_r_3973_sv2v_reg  <= 1'b0;
      \piso.data_r_3972_sv2v_reg  <= 1'b0;
      \piso.data_r_3971_sv2v_reg  <= 1'b0;
      \piso.data_r_3970_sv2v_reg  <= 1'b0;
      \piso.data_r_3969_sv2v_reg  <= 1'b0;
      \piso.data_r_3968_sv2v_reg  <= 1'b0;
      \piso.data_r_3967_sv2v_reg  <= 1'b0;
      \piso.data_r_3966_sv2v_reg  <= 1'b0;
      \piso.data_r_3965_sv2v_reg  <= 1'b0;
      \piso.data_r_3964_sv2v_reg  <= 1'b0;
      \piso.data_r_3963_sv2v_reg  <= 1'b0;
      \piso.data_r_3962_sv2v_reg  <= 1'b0;
      \piso.data_r_3961_sv2v_reg  <= 1'b0;
      \piso.data_r_3960_sv2v_reg  <= 1'b0;
      \piso.data_r_3959_sv2v_reg  <= 1'b0;
      \piso.data_r_3958_sv2v_reg  <= 1'b0;
      \piso.data_r_3957_sv2v_reg  <= 1'b0;
      \piso.data_r_3956_sv2v_reg  <= 1'b0;
      \piso.data_r_3955_sv2v_reg  <= 1'b0;
      \piso.data_r_3954_sv2v_reg  <= 1'b0;
      \piso.data_r_3953_sv2v_reg  <= 1'b0;
      \piso.data_r_3952_sv2v_reg  <= 1'b0;
      \piso.data_r_3951_sv2v_reg  <= 1'b0;
      \piso.data_r_3950_sv2v_reg  <= 1'b0;
      \piso.data_r_3949_sv2v_reg  <= 1'b0;
      \piso.data_r_3948_sv2v_reg  <= 1'b0;
      \piso.data_r_3947_sv2v_reg  <= 1'b0;
      \piso.data_r_3946_sv2v_reg  <= 1'b0;
      \piso.data_r_3945_sv2v_reg  <= 1'b0;
      \piso.data_r_3944_sv2v_reg  <= 1'b0;
      \piso.data_r_3943_sv2v_reg  <= 1'b0;
      \piso.data_r_3942_sv2v_reg  <= 1'b0;
      \piso.data_r_3941_sv2v_reg  <= 1'b0;
      \piso.data_r_3940_sv2v_reg  <= 1'b0;
      \piso.data_r_3939_sv2v_reg  <= 1'b0;
      \piso.data_r_3938_sv2v_reg  <= 1'b0;
      \piso.data_r_3937_sv2v_reg  <= 1'b0;
      \piso.data_r_3936_sv2v_reg  <= 1'b0;
      \piso.data_r_3935_sv2v_reg  <= 1'b0;
      \piso.data_r_3934_sv2v_reg  <= 1'b0;
      \piso.data_r_3933_sv2v_reg  <= 1'b0;
      \piso.data_r_3932_sv2v_reg  <= 1'b0;
      \piso.data_r_3931_sv2v_reg  <= 1'b0;
      \piso.data_r_3930_sv2v_reg  <= 1'b0;
      \piso.data_r_3929_sv2v_reg  <= 1'b0;
      \piso.data_r_3928_sv2v_reg  <= 1'b0;
      \piso.data_r_3927_sv2v_reg  <= 1'b0;
      \piso.data_r_3926_sv2v_reg  <= 1'b0;
      \piso.data_r_3925_sv2v_reg  <= 1'b0;
      \piso.data_r_3924_sv2v_reg  <= 1'b0;
      \piso.data_r_3923_sv2v_reg  <= 1'b0;
      \piso.data_r_3922_sv2v_reg  <= 1'b0;
      \piso.data_r_3921_sv2v_reg  <= 1'b0;
      \piso.data_r_3920_sv2v_reg  <= 1'b0;
      \piso.data_r_3919_sv2v_reg  <= 1'b0;
      \piso.data_r_3918_sv2v_reg  <= 1'b0;
      \piso.data_r_3917_sv2v_reg  <= 1'b0;
      \piso.data_r_3916_sv2v_reg  <= 1'b0;
      \piso.data_r_3915_sv2v_reg  <= 1'b0;
      \piso.data_r_3914_sv2v_reg  <= 1'b0;
      \piso.data_r_3913_sv2v_reg  <= 1'b0;
      \piso.data_r_3912_sv2v_reg  <= 1'b0;
      \piso.data_r_3911_sv2v_reg  <= 1'b0;
      \piso.data_r_3910_sv2v_reg  <= 1'b0;
      \piso.data_r_3909_sv2v_reg  <= 1'b0;
      \piso.data_r_3908_sv2v_reg  <= 1'b0;
      \piso.data_r_3907_sv2v_reg  <= 1'b0;
      \piso.data_r_3906_sv2v_reg  <= 1'b0;
      \piso.data_r_3905_sv2v_reg  <= 1'b0;
      \piso.data_r_3904_sv2v_reg  <= 1'b0;
      \piso.data_r_3903_sv2v_reg  <= 1'b0;
      \piso.data_r_3902_sv2v_reg  <= 1'b0;
      \piso.data_r_3901_sv2v_reg  <= 1'b0;
      \piso.data_r_3900_sv2v_reg  <= 1'b0;
      \piso.data_r_3899_sv2v_reg  <= 1'b0;
      \piso.data_r_3898_sv2v_reg  <= 1'b0;
      \piso.data_r_3897_sv2v_reg  <= 1'b0;
      \piso.data_r_3896_sv2v_reg  <= 1'b0;
      \piso.data_r_3895_sv2v_reg  <= 1'b0;
      \piso.data_r_3894_sv2v_reg  <= 1'b0;
      \piso.data_r_3893_sv2v_reg  <= 1'b0;
      \piso.data_r_3892_sv2v_reg  <= 1'b0;
      \piso.data_r_3891_sv2v_reg  <= 1'b0;
      \piso.data_r_3890_sv2v_reg  <= 1'b0;
      \piso.data_r_3889_sv2v_reg  <= 1'b0;
      \piso.data_r_3888_sv2v_reg  <= 1'b0;
      \piso.data_r_3887_sv2v_reg  <= 1'b0;
      \piso.data_r_3886_sv2v_reg  <= 1'b0;
      \piso.data_r_3885_sv2v_reg  <= 1'b0;
      \piso.data_r_3884_sv2v_reg  <= 1'b0;
      \piso.data_r_3883_sv2v_reg  <= 1'b0;
      \piso.data_r_3882_sv2v_reg  <= 1'b0;
      \piso.data_r_3881_sv2v_reg  <= 1'b0;
      \piso.data_r_3880_sv2v_reg  <= 1'b0;
      \piso.data_r_3879_sv2v_reg  <= 1'b0;
      \piso.data_r_3878_sv2v_reg  <= 1'b0;
      \piso.data_r_3877_sv2v_reg  <= 1'b0;
      \piso.data_r_3876_sv2v_reg  <= 1'b0;
      \piso.data_r_3875_sv2v_reg  <= 1'b0;
      \piso.data_r_3874_sv2v_reg  <= 1'b0;
      \piso.data_r_3873_sv2v_reg  <= 1'b0;
      \piso.data_r_3872_sv2v_reg  <= 1'b0;
      \piso.data_r_3871_sv2v_reg  <= 1'b0;
      \piso.data_r_3870_sv2v_reg  <= 1'b0;
      \piso.data_r_3869_sv2v_reg  <= 1'b0;
      \piso.data_r_3868_sv2v_reg  <= 1'b0;
      \piso.data_r_3867_sv2v_reg  <= 1'b0;
      \piso.data_r_3866_sv2v_reg  <= 1'b0;
      \piso.data_r_3865_sv2v_reg  <= 1'b0;
      \piso.data_r_3864_sv2v_reg  <= 1'b0;
      \piso.data_r_3863_sv2v_reg  <= 1'b0;
      \piso.data_r_3862_sv2v_reg  <= 1'b0;
      \piso.data_r_3861_sv2v_reg  <= 1'b0;
      \piso.data_r_3860_sv2v_reg  <= 1'b0;
      \piso.data_r_3859_sv2v_reg  <= 1'b0;
      \piso.data_r_3858_sv2v_reg  <= 1'b0;
      \piso.data_r_3857_sv2v_reg  <= 1'b0;
      \piso.data_r_3856_sv2v_reg  <= 1'b0;
      \piso.data_r_3855_sv2v_reg  <= 1'b0;
      \piso.data_r_3854_sv2v_reg  <= 1'b0;
      \piso.data_r_3853_sv2v_reg  <= 1'b0;
      \piso.data_r_3852_sv2v_reg  <= 1'b0;
      \piso.data_r_3851_sv2v_reg  <= 1'b0;
      \piso.data_r_3850_sv2v_reg  <= 1'b0;
      \piso.data_r_3849_sv2v_reg  <= 1'b0;
      \piso.data_r_3848_sv2v_reg  <= 1'b0;
      \piso.data_r_3847_sv2v_reg  <= 1'b0;
      \piso.data_r_3846_sv2v_reg  <= 1'b0;
      \piso.data_r_3845_sv2v_reg  <= 1'b0;
      \piso.data_r_3844_sv2v_reg  <= 1'b0;
      \piso.data_r_3843_sv2v_reg  <= 1'b0;
      \piso.data_r_3842_sv2v_reg  <= 1'b0;
      \piso.data_r_3841_sv2v_reg  <= 1'b0;
      \piso.data_r_3840_sv2v_reg  <= 1'b0;
      \piso.data_r_3839_sv2v_reg  <= 1'b0;
      \piso.data_r_3838_sv2v_reg  <= 1'b0;
      \piso.data_r_3837_sv2v_reg  <= 1'b0;
      \piso.data_r_3836_sv2v_reg  <= 1'b0;
      \piso.data_r_3835_sv2v_reg  <= 1'b0;
      \piso.data_r_3834_sv2v_reg  <= 1'b0;
      \piso.data_r_3833_sv2v_reg  <= 1'b0;
      \piso.data_r_3832_sv2v_reg  <= 1'b0;
      \piso.data_r_3831_sv2v_reg  <= 1'b0;
      \piso.data_r_3830_sv2v_reg  <= 1'b0;
      \piso.data_r_3829_sv2v_reg  <= 1'b0;
      \piso.data_r_3828_sv2v_reg  <= 1'b0;
      \piso.data_r_3827_sv2v_reg  <= 1'b0;
      \piso.data_r_3826_sv2v_reg  <= 1'b0;
      \piso.data_r_3825_sv2v_reg  <= 1'b0;
      \piso.data_r_3824_sv2v_reg  <= 1'b0;
      \piso.data_r_3823_sv2v_reg  <= 1'b0;
      \piso.data_r_3822_sv2v_reg  <= 1'b0;
      \piso.data_r_3821_sv2v_reg  <= 1'b0;
      \piso.data_r_3820_sv2v_reg  <= 1'b0;
      \piso.data_r_3819_sv2v_reg  <= 1'b0;
      \piso.data_r_3818_sv2v_reg  <= 1'b0;
      \piso.data_r_3817_sv2v_reg  <= 1'b0;
      \piso.data_r_3816_sv2v_reg  <= 1'b0;
      \piso.data_r_3815_sv2v_reg  <= 1'b0;
      \piso.data_r_3814_sv2v_reg  <= 1'b0;
      \piso.data_r_3813_sv2v_reg  <= 1'b0;
      \piso.data_r_3812_sv2v_reg  <= 1'b0;
      \piso.data_r_3811_sv2v_reg  <= 1'b0;
      \piso.data_r_3810_sv2v_reg  <= 1'b0;
      \piso.data_r_3809_sv2v_reg  <= 1'b0;
      \piso.data_r_3808_sv2v_reg  <= 1'b0;
      \piso.data_r_3807_sv2v_reg  <= 1'b0;
      \piso.data_r_3806_sv2v_reg  <= 1'b0;
      \piso.data_r_3805_sv2v_reg  <= 1'b0;
      \piso.data_r_3804_sv2v_reg  <= 1'b0;
      \piso.data_r_3803_sv2v_reg  <= 1'b0;
      \piso.data_r_3802_sv2v_reg  <= 1'b0;
      \piso.data_r_3801_sv2v_reg  <= 1'b0;
      \piso.data_r_3800_sv2v_reg  <= 1'b0;
      \piso.data_r_3799_sv2v_reg  <= 1'b0;
      \piso.data_r_3798_sv2v_reg  <= 1'b0;
      \piso.data_r_3797_sv2v_reg  <= 1'b0;
      \piso.data_r_3796_sv2v_reg  <= 1'b0;
      \piso.data_r_3795_sv2v_reg  <= 1'b0;
      \piso.data_r_3794_sv2v_reg  <= 1'b0;
      \piso.data_r_3793_sv2v_reg  <= 1'b0;
      \piso.data_r_3792_sv2v_reg  <= 1'b0;
      \piso.data_r_3791_sv2v_reg  <= 1'b0;
      \piso.data_r_3790_sv2v_reg  <= 1'b0;
      \piso.data_r_3789_sv2v_reg  <= 1'b0;
      \piso.data_r_3788_sv2v_reg  <= 1'b0;
      \piso.data_r_3787_sv2v_reg  <= 1'b0;
      \piso.data_r_3786_sv2v_reg  <= 1'b0;
      \piso.data_r_3785_sv2v_reg  <= 1'b0;
      \piso.data_r_3784_sv2v_reg  <= 1'b0;
      \piso.data_r_3783_sv2v_reg  <= 1'b0;
      \piso.data_r_3782_sv2v_reg  <= 1'b0;
      \piso.data_r_3781_sv2v_reg  <= 1'b0;
      \piso.data_r_3780_sv2v_reg  <= 1'b0;
      \piso.data_r_3779_sv2v_reg  <= 1'b0;
      \piso.data_r_3778_sv2v_reg  <= 1'b0;
      \piso.data_r_3777_sv2v_reg  <= 1'b0;
      \piso.data_r_3776_sv2v_reg  <= 1'b0;
      \piso.data_r_3775_sv2v_reg  <= 1'b0;
      \piso.data_r_3774_sv2v_reg  <= 1'b0;
      \piso.data_r_3773_sv2v_reg  <= 1'b0;
      \piso.data_r_3772_sv2v_reg  <= 1'b0;
      \piso.data_r_3771_sv2v_reg  <= 1'b0;
      \piso.data_r_3770_sv2v_reg  <= 1'b0;
      \piso.data_r_3769_sv2v_reg  <= 1'b0;
      \piso.data_r_3768_sv2v_reg  <= 1'b0;
      \piso.data_r_3767_sv2v_reg  <= 1'b0;
      \piso.data_r_3766_sv2v_reg  <= 1'b0;
      \piso.data_r_3765_sv2v_reg  <= 1'b0;
      \piso.data_r_3764_sv2v_reg  <= 1'b0;
      \piso.data_r_3763_sv2v_reg  <= 1'b0;
      \piso.data_r_3762_sv2v_reg  <= 1'b0;
      \piso.data_r_3761_sv2v_reg  <= 1'b0;
      \piso.data_r_3760_sv2v_reg  <= 1'b0;
      \piso.data_r_3759_sv2v_reg  <= 1'b0;
      \piso.data_r_3758_sv2v_reg  <= 1'b0;
      \piso.data_r_3757_sv2v_reg  <= 1'b0;
      \piso.data_r_3756_sv2v_reg  <= 1'b0;
      \piso.data_r_3755_sv2v_reg  <= 1'b0;
      \piso.data_r_3754_sv2v_reg  <= 1'b0;
      \piso.data_r_3753_sv2v_reg  <= 1'b0;
      \piso.data_r_3752_sv2v_reg  <= 1'b0;
      \piso.data_r_3751_sv2v_reg  <= 1'b0;
      \piso.data_r_3750_sv2v_reg  <= 1'b0;
      \piso.data_r_3749_sv2v_reg  <= 1'b0;
      \piso.data_r_3748_sv2v_reg  <= 1'b0;
      \piso.data_r_3747_sv2v_reg  <= 1'b0;
      \piso.data_r_3746_sv2v_reg  <= 1'b0;
      \piso.data_r_3745_sv2v_reg  <= 1'b0;
      \piso.data_r_3744_sv2v_reg  <= 1'b0;
      \piso.data_r_3743_sv2v_reg  <= 1'b0;
      \piso.data_r_3742_sv2v_reg  <= 1'b0;
      \piso.data_r_3741_sv2v_reg  <= 1'b0;
      \piso.data_r_3740_sv2v_reg  <= 1'b0;
      \piso.data_r_3739_sv2v_reg  <= 1'b0;
      \piso.data_r_3738_sv2v_reg  <= 1'b0;
      \piso.data_r_3737_sv2v_reg  <= 1'b0;
      \piso.data_r_3736_sv2v_reg  <= 1'b0;
      \piso.data_r_3735_sv2v_reg  <= 1'b0;
      \piso.data_r_3734_sv2v_reg  <= 1'b0;
      \piso.data_r_3733_sv2v_reg  <= 1'b0;
      \piso.data_r_3732_sv2v_reg  <= 1'b0;
      \piso.data_r_3731_sv2v_reg  <= 1'b0;
      \piso.data_r_3730_sv2v_reg  <= 1'b0;
      \piso.data_r_3729_sv2v_reg  <= 1'b0;
      \piso.data_r_3728_sv2v_reg  <= 1'b0;
      \piso.data_r_3727_sv2v_reg  <= 1'b0;
      \piso.data_r_3726_sv2v_reg  <= 1'b0;
      \piso.data_r_3725_sv2v_reg  <= 1'b0;
      \piso.data_r_3724_sv2v_reg  <= 1'b0;
      \piso.data_r_3723_sv2v_reg  <= 1'b0;
      \piso.data_r_3722_sv2v_reg  <= 1'b0;
      \piso.data_r_3721_sv2v_reg  <= 1'b0;
      \piso.data_r_3720_sv2v_reg  <= 1'b0;
      \piso.data_r_3719_sv2v_reg  <= 1'b0;
      \piso.data_r_3718_sv2v_reg  <= 1'b0;
      \piso.data_r_3717_sv2v_reg  <= 1'b0;
      \piso.data_r_3716_sv2v_reg  <= 1'b0;
      \piso.data_r_3715_sv2v_reg  <= 1'b0;
      \piso.data_r_3714_sv2v_reg  <= 1'b0;
      \piso.data_r_3713_sv2v_reg  <= 1'b0;
      \piso.data_r_3712_sv2v_reg  <= 1'b0;
      \piso.data_r_3711_sv2v_reg  <= 1'b0;
      \piso.data_r_3710_sv2v_reg  <= 1'b0;
      \piso.data_r_3709_sv2v_reg  <= 1'b0;
      \piso.data_r_3708_sv2v_reg  <= 1'b0;
      \piso.data_r_3707_sv2v_reg  <= 1'b0;
      \piso.data_r_3706_sv2v_reg  <= 1'b0;
      \piso.data_r_3705_sv2v_reg  <= 1'b0;
      \piso.data_r_3704_sv2v_reg  <= 1'b0;
      \piso.data_r_3703_sv2v_reg  <= 1'b0;
      \piso.data_r_3702_sv2v_reg  <= 1'b0;
      \piso.data_r_3701_sv2v_reg  <= 1'b0;
      \piso.data_r_3700_sv2v_reg  <= 1'b0;
      \piso.data_r_3699_sv2v_reg  <= 1'b0;
      \piso.data_r_3698_sv2v_reg  <= 1'b0;
      \piso.data_r_3697_sv2v_reg  <= 1'b0;
      \piso.data_r_3696_sv2v_reg  <= 1'b0;
      \piso.data_r_3695_sv2v_reg  <= 1'b0;
      \piso.data_r_3694_sv2v_reg  <= 1'b0;
      \piso.data_r_3693_sv2v_reg  <= 1'b0;
      \piso.data_r_3692_sv2v_reg  <= 1'b0;
      \piso.data_r_3691_sv2v_reg  <= 1'b0;
      \piso.data_r_3690_sv2v_reg  <= 1'b0;
      \piso.data_r_3689_sv2v_reg  <= 1'b0;
      \piso.data_r_3688_sv2v_reg  <= 1'b0;
      \piso.data_r_3687_sv2v_reg  <= 1'b0;
      \piso.data_r_3686_sv2v_reg  <= 1'b0;
      \piso.data_r_3685_sv2v_reg  <= 1'b0;
      \piso.data_r_3684_sv2v_reg  <= 1'b0;
      \piso.data_r_3683_sv2v_reg  <= 1'b0;
      \piso.data_r_3682_sv2v_reg  <= 1'b0;
      \piso.data_r_3681_sv2v_reg  <= 1'b0;
      \piso.data_r_3680_sv2v_reg  <= 1'b0;
      \piso.data_r_3679_sv2v_reg  <= 1'b0;
      \piso.data_r_3678_sv2v_reg  <= 1'b0;
      \piso.data_r_3677_sv2v_reg  <= 1'b0;
      \piso.data_r_3676_sv2v_reg  <= 1'b0;
      \piso.data_r_3675_sv2v_reg  <= 1'b0;
      \piso.data_r_3674_sv2v_reg  <= 1'b0;
      \piso.data_r_3673_sv2v_reg  <= 1'b0;
      \piso.data_r_3672_sv2v_reg  <= 1'b0;
      \piso.data_r_3671_sv2v_reg  <= 1'b0;
      \piso.data_r_3670_sv2v_reg  <= 1'b0;
      \piso.data_r_3669_sv2v_reg  <= 1'b0;
      \piso.data_r_3668_sv2v_reg  <= 1'b0;
      \piso.data_r_3667_sv2v_reg  <= 1'b0;
      \piso.data_r_3666_sv2v_reg  <= 1'b0;
      \piso.data_r_3665_sv2v_reg  <= 1'b0;
      \piso.data_r_3664_sv2v_reg  <= 1'b0;
      \piso.data_r_3663_sv2v_reg  <= 1'b0;
      \piso.data_r_3662_sv2v_reg  <= 1'b0;
      \piso.data_r_3661_sv2v_reg  <= 1'b0;
      \piso.data_r_3660_sv2v_reg  <= 1'b0;
      \piso.data_r_3659_sv2v_reg  <= 1'b0;
      \piso.data_r_3658_sv2v_reg  <= 1'b0;
      \piso.data_r_3657_sv2v_reg  <= 1'b0;
      \piso.data_r_3656_sv2v_reg  <= 1'b0;
      \piso.data_r_3655_sv2v_reg  <= 1'b0;
      \piso.data_r_3654_sv2v_reg  <= 1'b0;
      \piso.data_r_3653_sv2v_reg  <= 1'b0;
      \piso.data_r_3652_sv2v_reg  <= 1'b0;
      \piso.data_r_3651_sv2v_reg  <= 1'b0;
      \piso.data_r_3650_sv2v_reg  <= 1'b0;
      \piso.data_r_3649_sv2v_reg  <= 1'b0;
      \piso.data_r_3648_sv2v_reg  <= 1'b0;
      \piso.data_r_3647_sv2v_reg  <= 1'b0;
      \piso.data_r_3646_sv2v_reg  <= 1'b0;
      \piso.data_r_3645_sv2v_reg  <= 1'b0;
      \piso.data_r_3644_sv2v_reg  <= 1'b0;
      \piso.data_r_3643_sv2v_reg  <= 1'b0;
      \piso.data_r_3642_sv2v_reg  <= 1'b0;
      \piso.data_r_3641_sv2v_reg  <= 1'b0;
      \piso.data_r_3640_sv2v_reg  <= 1'b0;
      \piso.data_r_3639_sv2v_reg  <= 1'b0;
      \piso.data_r_3638_sv2v_reg  <= 1'b0;
      \piso.data_r_3637_sv2v_reg  <= 1'b0;
      \piso.data_r_3636_sv2v_reg  <= 1'b0;
      \piso.data_r_3635_sv2v_reg  <= 1'b0;
      \piso.data_r_3634_sv2v_reg  <= 1'b0;
      \piso.data_r_3633_sv2v_reg  <= 1'b0;
      \piso.data_r_3632_sv2v_reg  <= 1'b0;
      \piso.data_r_3631_sv2v_reg  <= 1'b0;
      \piso.data_r_3630_sv2v_reg  <= 1'b0;
      \piso.data_r_3629_sv2v_reg  <= 1'b0;
      \piso.data_r_3628_sv2v_reg  <= 1'b0;
      \piso.data_r_3627_sv2v_reg  <= 1'b0;
      \piso.data_r_3626_sv2v_reg  <= 1'b0;
      \piso.data_r_3625_sv2v_reg  <= 1'b0;
      \piso.data_r_3624_sv2v_reg  <= 1'b0;
      \piso.data_r_3623_sv2v_reg  <= 1'b0;
      \piso.data_r_3622_sv2v_reg  <= 1'b0;
      \piso.data_r_3621_sv2v_reg  <= 1'b0;
      \piso.data_r_3620_sv2v_reg  <= 1'b0;
      \piso.data_r_3619_sv2v_reg  <= 1'b0;
      \piso.data_r_3618_sv2v_reg  <= 1'b0;
      \piso.data_r_3617_sv2v_reg  <= 1'b0;
      \piso.data_r_3616_sv2v_reg  <= 1'b0;
      \piso.data_r_3615_sv2v_reg  <= 1'b0;
      \piso.data_r_3614_sv2v_reg  <= 1'b0;
      \piso.data_r_3613_sv2v_reg  <= 1'b0;
      \piso.data_r_3612_sv2v_reg  <= 1'b0;
      \piso.data_r_3611_sv2v_reg  <= 1'b0;
      \piso.data_r_3610_sv2v_reg  <= 1'b0;
      \piso.data_r_3609_sv2v_reg  <= 1'b0;
      \piso.data_r_3608_sv2v_reg  <= 1'b0;
      \piso.data_r_3607_sv2v_reg  <= 1'b0;
      \piso.data_r_3606_sv2v_reg  <= 1'b0;
      \piso.data_r_3605_sv2v_reg  <= 1'b0;
      \piso.data_r_3604_sv2v_reg  <= 1'b0;
      \piso.data_r_3603_sv2v_reg  <= 1'b0;
      \piso.data_r_3602_sv2v_reg  <= 1'b0;
      \piso.data_r_3601_sv2v_reg  <= 1'b0;
      \piso.data_r_3600_sv2v_reg  <= 1'b0;
      \piso.data_r_3599_sv2v_reg  <= 1'b0;
      \piso.data_r_3598_sv2v_reg  <= 1'b0;
      \piso.data_r_3597_sv2v_reg  <= 1'b0;
      \piso.data_r_3596_sv2v_reg  <= 1'b0;
      \piso.data_r_3595_sv2v_reg  <= 1'b0;
      \piso.data_r_3594_sv2v_reg  <= 1'b0;
      \piso.data_r_3593_sv2v_reg  <= 1'b0;
      \piso.data_r_3592_sv2v_reg  <= 1'b0;
      \piso.data_r_3591_sv2v_reg  <= 1'b0;
      \piso.data_r_3590_sv2v_reg  <= 1'b0;
      \piso.data_r_3589_sv2v_reg  <= 1'b0;
      \piso.data_r_3588_sv2v_reg  <= 1'b0;
      \piso.data_r_3587_sv2v_reg  <= 1'b0;
      \piso.data_r_3586_sv2v_reg  <= 1'b0;
      \piso.data_r_3585_sv2v_reg  <= 1'b0;
      \piso.data_r_3584_sv2v_reg  <= 1'b0;
      \piso.data_r_3583_sv2v_reg  <= 1'b0;
      \piso.data_r_3582_sv2v_reg  <= 1'b0;
      \piso.data_r_3581_sv2v_reg  <= 1'b0;
      \piso.data_r_3580_sv2v_reg  <= 1'b0;
      \piso.data_r_3579_sv2v_reg  <= 1'b0;
      \piso.data_r_3578_sv2v_reg  <= 1'b0;
      \piso.data_r_3577_sv2v_reg  <= 1'b0;
      \piso.data_r_3576_sv2v_reg  <= 1'b0;
      \piso.data_r_3575_sv2v_reg  <= 1'b0;
      \piso.data_r_3574_sv2v_reg  <= 1'b0;
      \piso.data_r_3573_sv2v_reg  <= 1'b0;
      \piso.data_r_3572_sv2v_reg  <= 1'b0;
      \piso.data_r_3571_sv2v_reg  <= 1'b0;
      \piso.data_r_3570_sv2v_reg  <= 1'b0;
      \piso.data_r_3569_sv2v_reg  <= 1'b0;
      \piso.data_r_3568_sv2v_reg  <= 1'b0;
      \piso.data_r_3567_sv2v_reg  <= 1'b0;
      \piso.data_r_3566_sv2v_reg  <= 1'b0;
      \piso.data_r_3565_sv2v_reg  <= 1'b0;
      \piso.data_r_3564_sv2v_reg  <= 1'b0;
      \piso.data_r_3563_sv2v_reg  <= 1'b0;
      \piso.data_r_3562_sv2v_reg  <= 1'b0;
      \piso.data_r_3561_sv2v_reg  <= 1'b0;
      \piso.data_r_3560_sv2v_reg  <= 1'b0;
      \piso.data_r_3559_sv2v_reg  <= 1'b0;
      \piso.data_r_3558_sv2v_reg  <= 1'b0;
      \piso.data_r_3557_sv2v_reg  <= 1'b0;
      \piso.data_r_3556_sv2v_reg  <= 1'b0;
      \piso.data_r_3555_sv2v_reg  <= 1'b0;
      \piso.data_r_3554_sv2v_reg  <= 1'b0;
      \piso.data_r_3553_sv2v_reg  <= 1'b0;
      \piso.data_r_3552_sv2v_reg  <= 1'b0;
      \piso.data_r_3551_sv2v_reg  <= 1'b0;
      \piso.data_r_3550_sv2v_reg  <= 1'b0;
      \piso.data_r_3549_sv2v_reg  <= 1'b0;
      \piso.data_r_3548_sv2v_reg  <= 1'b0;
      \piso.data_r_3547_sv2v_reg  <= 1'b0;
      \piso.data_r_3546_sv2v_reg  <= 1'b0;
      \piso.data_r_3545_sv2v_reg  <= 1'b0;
      \piso.data_r_3544_sv2v_reg  <= 1'b0;
      \piso.data_r_3543_sv2v_reg  <= 1'b0;
      \piso.data_r_3542_sv2v_reg  <= 1'b0;
      \piso.data_r_3541_sv2v_reg  <= 1'b0;
      \piso.data_r_3540_sv2v_reg  <= 1'b0;
      \piso.data_r_3539_sv2v_reg  <= 1'b0;
      \piso.data_r_3538_sv2v_reg  <= 1'b0;
      \piso.data_r_3537_sv2v_reg  <= 1'b0;
      \piso.data_r_3536_sv2v_reg  <= 1'b0;
      \piso.data_r_3535_sv2v_reg  <= 1'b0;
      \piso.data_r_3534_sv2v_reg  <= 1'b0;
      \piso.data_r_3533_sv2v_reg  <= 1'b0;
      \piso.data_r_3532_sv2v_reg  <= 1'b0;
      \piso.data_r_3531_sv2v_reg  <= 1'b0;
      \piso.data_r_3530_sv2v_reg  <= 1'b0;
      \piso.data_r_3529_sv2v_reg  <= 1'b0;
      \piso.data_r_3528_sv2v_reg  <= 1'b0;
      \piso.data_r_3527_sv2v_reg  <= 1'b0;
      \piso.data_r_3526_sv2v_reg  <= 1'b0;
      \piso.data_r_3525_sv2v_reg  <= 1'b0;
      \piso.data_r_3524_sv2v_reg  <= 1'b0;
      \piso.data_r_3523_sv2v_reg  <= 1'b0;
      \piso.data_r_3522_sv2v_reg  <= 1'b0;
      \piso.data_r_3521_sv2v_reg  <= 1'b0;
      \piso.data_r_3520_sv2v_reg  <= 1'b0;
      \piso.data_r_3519_sv2v_reg  <= 1'b0;
      \piso.data_r_3518_sv2v_reg  <= 1'b0;
      \piso.data_r_3517_sv2v_reg  <= 1'b0;
      \piso.data_r_3516_sv2v_reg  <= 1'b0;
      \piso.data_r_3515_sv2v_reg  <= 1'b0;
      \piso.data_r_3514_sv2v_reg  <= 1'b0;
      \piso.data_r_3513_sv2v_reg  <= 1'b0;
      \piso.data_r_3512_sv2v_reg  <= 1'b0;
      \piso.data_r_3511_sv2v_reg  <= 1'b0;
      \piso.data_r_3510_sv2v_reg  <= 1'b0;
      \piso.data_r_3509_sv2v_reg  <= 1'b0;
      \piso.data_r_3508_sv2v_reg  <= 1'b0;
      \piso.data_r_3507_sv2v_reg  <= 1'b0;
      \piso.data_r_3506_sv2v_reg  <= 1'b0;
      \piso.data_r_3505_sv2v_reg  <= 1'b0;
      \piso.data_r_3504_sv2v_reg  <= 1'b0;
      \piso.data_r_3503_sv2v_reg  <= 1'b0;
      \piso.data_r_3502_sv2v_reg  <= 1'b0;
      \piso.data_r_3501_sv2v_reg  <= 1'b0;
      \piso.data_r_3500_sv2v_reg  <= 1'b0;
      \piso.data_r_3499_sv2v_reg  <= 1'b0;
      \piso.data_r_3498_sv2v_reg  <= 1'b0;
      \piso.data_r_3497_sv2v_reg  <= 1'b0;
      \piso.data_r_3496_sv2v_reg  <= 1'b0;
      \piso.data_r_3495_sv2v_reg  <= 1'b0;
      \piso.data_r_3494_sv2v_reg  <= 1'b0;
      \piso.data_r_3493_sv2v_reg  <= 1'b0;
      \piso.data_r_3492_sv2v_reg  <= 1'b0;
      \piso.data_r_3491_sv2v_reg  <= 1'b0;
      \piso.data_r_3490_sv2v_reg  <= 1'b0;
      \piso.data_r_3489_sv2v_reg  <= 1'b0;
      \piso.data_r_3488_sv2v_reg  <= 1'b0;
      \piso.data_r_3487_sv2v_reg  <= 1'b0;
      \piso.data_r_3486_sv2v_reg  <= 1'b0;
      \piso.data_r_3485_sv2v_reg  <= 1'b0;
      \piso.data_r_3484_sv2v_reg  <= 1'b0;
      \piso.data_r_3483_sv2v_reg  <= 1'b0;
      \piso.data_r_3482_sv2v_reg  <= 1'b0;
      \piso.data_r_3481_sv2v_reg  <= 1'b0;
      \piso.data_r_3480_sv2v_reg  <= 1'b0;
      \piso.data_r_3479_sv2v_reg  <= 1'b0;
      \piso.data_r_3478_sv2v_reg  <= 1'b0;
      \piso.data_r_3477_sv2v_reg  <= 1'b0;
      \piso.data_r_3476_sv2v_reg  <= 1'b0;
      \piso.data_r_3475_sv2v_reg  <= 1'b0;
      \piso.data_r_3474_sv2v_reg  <= 1'b0;
      \piso.data_r_3473_sv2v_reg  <= 1'b0;
      \piso.data_r_3472_sv2v_reg  <= 1'b0;
      \piso.data_r_3471_sv2v_reg  <= 1'b0;
      \piso.data_r_3470_sv2v_reg  <= 1'b0;
      \piso.data_r_3469_sv2v_reg  <= 1'b0;
      \piso.data_r_3468_sv2v_reg  <= 1'b0;
      \piso.data_r_3467_sv2v_reg  <= 1'b0;
      \piso.data_r_3466_sv2v_reg  <= 1'b0;
      \piso.data_r_3465_sv2v_reg  <= 1'b0;
      \piso.data_r_3464_sv2v_reg  <= 1'b0;
      \piso.data_r_3463_sv2v_reg  <= 1'b0;
      \piso.data_r_3462_sv2v_reg  <= 1'b0;
      \piso.data_r_3461_sv2v_reg  <= 1'b0;
      \piso.data_r_3460_sv2v_reg  <= 1'b0;
      \piso.data_r_3459_sv2v_reg  <= 1'b0;
      \piso.data_r_3458_sv2v_reg  <= 1'b0;
      \piso.data_r_3457_sv2v_reg  <= 1'b0;
      \piso.data_r_3456_sv2v_reg  <= 1'b0;
      \piso.data_r_3455_sv2v_reg  <= 1'b0;
      \piso.data_r_3454_sv2v_reg  <= 1'b0;
      \piso.data_r_3453_sv2v_reg  <= 1'b0;
      \piso.data_r_3452_sv2v_reg  <= 1'b0;
      \piso.data_r_3451_sv2v_reg  <= 1'b0;
      \piso.data_r_3450_sv2v_reg  <= 1'b0;
      \piso.data_r_3449_sv2v_reg  <= 1'b0;
      \piso.data_r_3448_sv2v_reg  <= 1'b0;
      \piso.data_r_3447_sv2v_reg  <= 1'b0;
      \piso.data_r_3446_sv2v_reg  <= 1'b0;
      \piso.data_r_3445_sv2v_reg  <= 1'b0;
      \piso.data_r_3444_sv2v_reg  <= 1'b0;
      \piso.data_r_3443_sv2v_reg  <= 1'b0;
      \piso.data_r_3442_sv2v_reg  <= 1'b0;
      \piso.data_r_3441_sv2v_reg  <= 1'b0;
      \piso.data_r_3440_sv2v_reg  <= 1'b0;
      \piso.data_r_3439_sv2v_reg  <= 1'b0;
      \piso.data_r_3438_sv2v_reg  <= 1'b0;
      \piso.data_r_3437_sv2v_reg  <= 1'b0;
      \piso.data_r_3436_sv2v_reg  <= 1'b0;
      \piso.data_r_3435_sv2v_reg  <= 1'b0;
      \piso.data_r_3434_sv2v_reg  <= 1'b0;
      \piso.data_r_3433_sv2v_reg  <= 1'b0;
      \piso.data_r_3432_sv2v_reg  <= 1'b0;
      \piso.data_r_3431_sv2v_reg  <= 1'b0;
      \piso.data_r_3430_sv2v_reg  <= 1'b0;
      \piso.data_r_3429_sv2v_reg  <= 1'b0;
      \piso.data_r_3428_sv2v_reg  <= 1'b0;
      \piso.data_r_3427_sv2v_reg  <= 1'b0;
      \piso.data_r_3426_sv2v_reg  <= 1'b0;
      \piso.data_r_3425_sv2v_reg  <= 1'b0;
      \piso.data_r_3424_sv2v_reg  <= 1'b0;
      \piso.data_r_3423_sv2v_reg  <= 1'b0;
      \piso.data_r_3422_sv2v_reg  <= 1'b0;
      \piso.data_r_3421_sv2v_reg  <= 1'b0;
      \piso.data_r_3420_sv2v_reg  <= 1'b0;
      \piso.data_r_3419_sv2v_reg  <= 1'b0;
      \piso.data_r_3418_sv2v_reg  <= 1'b0;
      \piso.data_r_3417_sv2v_reg  <= 1'b0;
      \piso.data_r_3416_sv2v_reg  <= 1'b0;
      \piso.data_r_3415_sv2v_reg  <= 1'b0;
      \piso.data_r_3414_sv2v_reg  <= 1'b0;
      \piso.data_r_3413_sv2v_reg  <= 1'b0;
      \piso.data_r_3412_sv2v_reg  <= 1'b0;
      \piso.data_r_3411_sv2v_reg  <= 1'b0;
      \piso.data_r_3410_sv2v_reg  <= 1'b0;
      \piso.data_r_3409_sv2v_reg  <= 1'b0;
      \piso.data_r_3408_sv2v_reg  <= 1'b0;
      \piso.data_r_3407_sv2v_reg  <= 1'b0;
      \piso.data_r_3406_sv2v_reg  <= 1'b0;
      \piso.data_r_3405_sv2v_reg  <= 1'b0;
      \piso.data_r_3404_sv2v_reg  <= 1'b0;
      \piso.data_r_3403_sv2v_reg  <= 1'b0;
      \piso.data_r_3402_sv2v_reg  <= 1'b0;
      \piso.data_r_3401_sv2v_reg  <= 1'b0;
      \piso.data_r_3400_sv2v_reg  <= 1'b0;
      \piso.data_r_3399_sv2v_reg  <= 1'b0;
      \piso.data_r_3398_sv2v_reg  <= 1'b0;
      \piso.data_r_3397_sv2v_reg  <= 1'b0;
      \piso.data_r_3396_sv2v_reg  <= 1'b0;
      \piso.data_r_3395_sv2v_reg  <= 1'b0;
      \piso.data_r_3394_sv2v_reg  <= 1'b0;
      \piso.data_r_3393_sv2v_reg  <= 1'b0;
      \piso.data_r_3392_sv2v_reg  <= 1'b0;
      \piso.data_r_3391_sv2v_reg  <= 1'b0;
      \piso.data_r_3390_sv2v_reg  <= 1'b0;
      \piso.data_r_3389_sv2v_reg  <= 1'b0;
      \piso.data_r_3388_sv2v_reg  <= 1'b0;
      \piso.data_r_3387_sv2v_reg  <= 1'b0;
      \piso.data_r_3386_sv2v_reg  <= 1'b0;
      \piso.data_r_3385_sv2v_reg  <= 1'b0;
      \piso.data_r_3384_sv2v_reg  <= 1'b0;
      \piso.data_r_3383_sv2v_reg  <= 1'b0;
      \piso.data_r_3382_sv2v_reg  <= 1'b0;
      \piso.data_r_3381_sv2v_reg  <= 1'b0;
      \piso.data_r_3380_sv2v_reg  <= 1'b0;
      \piso.data_r_3379_sv2v_reg  <= 1'b0;
      \piso.data_r_3378_sv2v_reg  <= 1'b0;
      \piso.data_r_3377_sv2v_reg  <= 1'b0;
      \piso.data_r_3376_sv2v_reg  <= 1'b0;
      \piso.data_r_3375_sv2v_reg  <= 1'b0;
      \piso.data_r_3374_sv2v_reg  <= 1'b0;
      \piso.data_r_3373_sv2v_reg  <= 1'b0;
      \piso.data_r_3372_sv2v_reg  <= 1'b0;
      \piso.data_r_3371_sv2v_reg  <= 1'b0;
      \piso.data_r_3370_sv2v_reg  <= 1'b0;
      \piso.data_r_3369_sv2v_reg  <= 1'b0;
      \piso.data_r_3368_sv2v_reg  <= 1'b0;
      \piso.data_r_3367_sv2v_reg  <= 1'b0;
      \piso.data_r_3366_sv2v_reg  <= 1'b0;
      \piso.data_r_3365_sv2v_reg  <= 1'b0;
      \piso.data_r_3364_sv2v_reg  <= 1'b0;
      \piso.data_r_3363_sv2v_reg  <= 1'b0;
      \piso.data_r_3362_sv2v_reg  <= 1'b0;
      \piso.data_r_3361_sv2v_reg  <= 1'b0;
      \piso.data_r_3360_sv2v_reg  <= 1'b0;
      \piso.data_r_3359_sv2v_reg  <= 1'b0;
      \piso.data_r_3358_sv2v_reg  <= 1'b0;
      \piso.data_r_3357_sv2v_reg  <= 1'b0;
      \piso.data_r_3356_sv2v_reg  <= 1'b0;
      \piso.data_r_3355_sv2v_reg  <= 1'b0;
      \piso.data_r_3354_sv2v_reg  <= 1'b0;
      \piso.data_r_3353_sv2v_reg  <= 1'b0;
      \piso.data_r_3352_sv2v_reg  <= 1'b0;
      \piso.data_r_3351_sv2v_reg  <= 1'b0;
      \piso.data_r_3350_sv2v_reg  <= 1'b0;
      \piso.data_r_3349_sv2v_reg  <= 1'b0;
      \piso.data_r_3348_sv2v_reg  <= 1'b0;
      \piso.data_r_3347_sv2v_reg  <= 1'b0;
      \piso.data_r_3346_sv2v_reg  <= 1'b0;
      \piso.data_r_3345_sv2v_reg  <= 1'b0;
      \piso.data_r_3344_sv2v_reg  <= 1'b0;
      \piso.data_r_3343_sv2v_reg  <= 1'b0;
      \piso.data_r_3342_sv2v_reg  <= 1'b0;
      \piso.data_r_3341_sv2v_reg  <= 1'b0;
      \piso.data_r_3340_sv2v_reg  <= 1'b0;
      \piso.data_r_3339_sv2v_reg  <= 1'b0;
      \piso.data_r_3338_sv2v_reg  <= 1'b0;
      \piso.data_r_3337_sv2v_reg  <= 1'b0;
      \piso.data_r_3336_sv2v_reg  <= 1'b0;
      \piso.data_r_3335_sv2v_reg  <= 1'b0;
      \piso.data_r_3334_sv2v_reg  <= 1'b0;
      \piso.data_r_3333_sv2v_reg  <= 1'b0;
      \piso.data_r_3332_sv2v_reg  <= 1'b0;
      \piso.data_r_3331_sv2v_reg  <= 1'b0;
      \piso.data_r_3330_sv2v_reg  <= 1'b0;
      \piso.data_r_3329_sv2v_reg  <= 1'b0;
      \piso.data_r_3328_sv2v_reg  <= 1'b0;
      \piso.data_r_3327_sv2v_reg  <= 1'b0;
      \piso.data_r_3326_sv2v_reg  <= 1'b0;
      \piso.data_r_3325_sv2v_reg  <= 1'b0;
      \piso.data_r_3324_sv2v_reg  <= 1'b0;
      \piso.data_r_3323_sv2v_reg  <= 1'b0;
      \piso.data_r_3322_sv2v_reg  <= 1'b0;
      \piso.data_r_3321_sv2v_reg  <= 1'b0;
      \piso.data_r_3320_sv2v_reg  <= 1'b0;
      \piso.data_r_3319_sv2v_reg  <= 1'b0;
      \piso.data_r_3318_sv2v_reg  <= 1'b0;
      \piso.data_r_3317_sv2v_reg  <= 1'b0;
      \piso.data_r_3316_sv2v_reg  <= 1'b0;
      \piso.data_r_3315_sv2v_reg  <= 1'b0;
      \piso.data_r_3314_sv2v_reg  <= 1'b0;
      \piso.data_r_3313_sv2v_reg  <= 1'b0;
      \piso.data_r_3312_sv2v_reg  <= 1'b0;
      \piso.data_r_3311_sv2v_reg  <= 1'b0;
      \piso.data_r_3310_sv2v_reg  <= 1'b0;
      \piso.data_r_3309_sv2v_reg  <= 1'b0;
      \piso.data_r_3308_sv2v_reg  <= 1'b0;
      \piso.data_r_3307_sv2v_reg  <= 1'b0;
      \piso.data_r_3306_sv2v_reg  <= 1'b0;
      \piso.data_r_3305_sv2v_reg  <= 1'b0;
      \piso.data_r_3304_sv2v_reg  <= 1'b0;
      \piso.data_r_3303_sv2v_reg  <= 1'b0;
      \piso.data_r_3302_sv2v_reg  <= 1'b0;
      \piso.data_r_3301_sv2v_reg  <= 1'b0;
      \piso.data_r_3300_sv2v_reg  <= 1'b0;
      \piso.data_r_3299_sv2v_reg  <= 1'b0;
      \piso.data_r_3298_sv2v_reg  <= 1'b0;
      \piso.data_r_3297_sv2v_reg  <= 1'b0;
      \piso.data_r_3296_sv2v_reg  <= 1'b0;
      \piso.data_r_3295_sv2v_reg  <= 1'b0;
      \piso.data_r_3294_sv2v_reg  <= 1'b0;
      \piso.data_r_3293_sv2v_reg  <= 1'b0;
      \piso.data_r_3292_sv2v_reg  <= 1'b0;
      \piso.data_r_3291_sv2v_reg  <= 1'b0;
      \piso.data_r_3290_sv2v_reg  <= 1'b0;
      \piso.data_r_3289_sv2v_reg  <= 1'b0;
      \piso.data_r_3288_sv2v_reg  <= 1'b0;
      \piso.data_r_3287_sv2v_reg  <= 1'b0;
      \piso.data_r_3286_sv2v_reg  <= 1'b0;
      \piso.data_r_3285_sv2v_reg  <= 1'b0;
      \piso.data_r_3284_sv2v_reg  <= 1'b0;
      \piso.data_r_3283_sv2v_reg  <= 1'b0;
      \piso.data_r_3282_sv2v_reg  <= 1'b0;
      \piso.data_r_3281_sv2v_reg  <= 1'b0;
      \piso.data_r_3280_sv2v_reg  <= 1'b0;
      \piso.data_r_3279_sv2v_reg  <= 1'b0;
      \piso.data_r_3278_sv2v_reg  <= 1'b0;
      \piso.data_r_3277_sv2v_reg  <= 1'b0;
      \piso.data_r_3276_sv2v_reg  <= 1'b0;
      \piso.data_r_3275_sv2v_reg  <= 1'b0;
      \piso.data_r_3274_sv2v_reg  <= 1'b0;
      \piso.data_r_3273_sv2v_reg  <= 1'b0;
      \piso.data_r_3272_sv2v_reg  <= 1'b0;
      \piso.data_r_3271_sv2v_reg  <= 1'b0;
      \piso.data_r_3270_sv2v_reg  <= 1'b0;
      \piso.data_r_3269_sv2v_reg  <= 1'b0;
      \piso.data_r_3268_sv2v_reg  <= 1'b0;
      \piso.data_r_3267_sv2v_reg  <= 1'b0;
      \piso.data_r_3266_sv2v_reg  <= 1'b0;
      \piso.data_r_3265_sv2v_reg  <= 1'b0;
      \piso.data_r_3264_sv2v_reg  <= 1'b0;
      \piso.data_r_3263_sv2v_reg  <= 1'b0;
      \piso.data_r_3262_sv2v_reg  <= 1'b0;
      \piso.data_r_3261_sv2v_reg  <= 1'b0;
      \piso.data_r_3260_sv2v_reg  <= 1'b0;
      \piso.data_r_3259_sv2v_reg  <= 1'b0;
      \piso.data_r_3258_sv2v_reg  <= 1'b0;
      \piso.data_r_3257_sv2v_reg  <= 1'b0;
      \piso.data_r_3256_sv2v_reg  <= 1'b0;
      \piso.data_r_3255_sv2v_reg  <= 1'b0;
      \piso.data_r_3254_sv2v_reg  <= 1'b0;
      \piso.data_r_3253_sv2v_reg  <= 1'b0;
      \piso.data_r_3252_sv2v_reg  <= 1'b0;
      \piso.data_r_3251_sv2v_reg  <= 1'b0;
      \piso.data_r_3250_sv2v_reg  <= 1'b0;
      \piso.data_r_3249_sv2v_reg  <= 1'b0;
      \piso.data_r_3248_sv2v_reg  <= 1'b0;
      \piso.data_r_3247_sv2v_reg  <= 1'b0;
      \piso.data_r_3246_sv2v_reg  <= 1'b0;
      \piso.data_r_3245_sv2v_reg  <= 1'b0;
      \piso.data_r_3244_sv2v_reg  <= 1'b0;
      \piso.data_r_3243_sv2v_reg  <= 1'b0;
      \piso.data_r_3242_sv2v_reg  <= 1'b0;
      \piso.data_r_3241_sv2v_reg  <= 1'b0;
      \piso.data_r_3240_sv2v_reg  <= 1'b0;
      \piso.data_r_3239_sv2v_reg  <= 1'b0;
      \piso.data_r_3238_sv2v_reg  <= 1'b0;
      \piso.data_r_3237_sv2v_reg  <= 1'b0;
      \piso.data_r_3236_sv2v_reg  <= 1'b0;
      \piso.data_r_3235_sv2v_reg  <= 1'b0;
      \piso.data_r_3234_sv2v_reg  <= 1'b0;
      \piso.data_r_3233_sv2v_reg  <= 1'b0;
      \piso.data_r_3232_sv2v_reg  <= 1'b0;
      \piso.data_r_3231_sv2v_reg  <= 1'b0;
      \piso.data_r_3230_sv2v_reg  <= 1'b0;
      \piso.data_r_3229_sv2v_reg  <= 1'b0;
      \piso.data_r_3228_sv2v_reg  <= 1'b0;
      \piso.data_r_3227_sv2v_reg  <= 1'b0;
      \piso.data_r_3226_sv2v_reg  <= 1'b0;
      \piso.data_r_3225_sv2v_reg  <= 1'b0;
      \piso.data_r_3224_sv2v_reg  <= 1'b0;
      \piso.data_r_3223_sv2v_reg  <= 1'b0;
      \piso.data_r_3222_sv2v_reg  <= 1'b0;
      \piso.data_r_3221_sv2v_reg  <= 1'b0;
      \piso.data_r_3220_sv2v_reg  <= 1'b0;
      \piso.data_r_3219_sv2v_reg  <= 1'b0;
      \piso.data_r_3218_sv2v_reg  <= 1'b0;
      \piso.data_r_3217_sv2v_reg  <= 1'b0;
      \piso.data_r_3216_sv2v_reg  <= 1'b0;
      \piso.data_r_3215_sv2v_reg  <= 1'b0;
      \piso.data_r_3214_sv2v_reg  <= 1'b0;
      \piso.data_r_3213_sv2v_reg  <= 1'b0;
      \piso.data_r_3212_sv2v_reg  <= 1'b0;
      \piso.data_r_3211_sv2v_reg  <= 1'b0;
      \piso.data_r_3210_sv2v_reg  <= 1'b0;
      \piso.data_r_3209_sv2v_reg  <= 1'b0;
      \piso.data_r_3208_sv2v_reg  <= 1'b0;
      \piso.data_r_3207_sv2v_reg  <= 1'b0;
      \piso.data_r_3206_sv2v_reg  <= 1'b0;
      \piso.data_r_3205_sv2v_reg  <= 1'b0;
      \piso.data_r_3204_sv2v_reg  <= 1'b0;
      \piso.data_r_3203_sv2v_reg  <= 1'b0;
      \piso.data_r_3202_sv2v_reg  <= 1'b0;
      \piso.data_r_3201_sv2v_reg  <= 1'b0;
      \piso.data_r_3200_sv2v_reg  <= 1'b0;
      \piso.data_r_3199_sv2v_reg  <= 1'b0;
      \piso.data_r_3198_sv2v_reg  <= 1'b0;
      \piso.data_r_3197_sv2v_reg  <= 1'b0;
      \piso.data_r_3196_sv2v_reg  <= 1'b0;
      \piso.data_r_3195_sv2v_reg  <= 1'b0;
      \piso.data_r_3194_sv2v_reg  <= 1'b0;
      \piso.data_r_3193_sv2v_reg  <= 1'b0;
      \piso.data_r_3192_sv2v_reg  <= 1'b0;
      \piso.data_r_3191_sv2v_reg  <= 1'b0;
      \piso.data_r_3190_sv2v_reg  <= 1'b0;
      \piso.data_r_3189_sv2v_reg  <= 1'b0;
      \piso.data_r_3188_sv2v_reg  <= 1'b0;
      \piso.data_r_3187_sv2v_reg  <= 1'b0;
      \piso.data_r_3186_sv2v_reg  <= 1'b0;
      \piso.data_r_3185_sv2v_reg  <= 1'b0;
      \piso.data_r_3184_sv2v_reg  <= 1'b0;
      \piso.data_r_3183_sv2v_reg  <= 1'b0;
      \piso.data_r_3182_sv2v_reg  <= 1'b0;
      \piso.data_r_3181_sv2v_reg  <= 1'b0;
      \piso.data_r_3180_sv2v_reg  <= 1'b0;
      \piso.data_r_3179_sv2v_reg  <= 1'b0;
      \piso.data_r_3178_sv2v_reg  <= 1'b0;
      \piso.data_r_3177_sv2v_reg  <= 1'b0;
      \piso.data_r_3176_sv2v_reg  <= 1'b0;
      \piso.data_r_3175_sv2v_reg  <= 1'b0;
      \piso.data_r_3174_sv2v_reg  <= 1'b0;
      \piso.data_r_3173_sv2v_reg  <= 1'b0;
      \piso.data_r_3172_sv2v_reg  <= 1'b0;
      \piso.data_r_3171_sv2v_reg  <= 1'b0;
      \piso.data_r_3170_sv2v_reg  <= 1'b0;
      \piso.data_r_3169_sv2v_reg  <= 1'b0;
      \piso.data_r_3168_sv2v_reg  <= 1'b0;
      \piso.data_r_3167_sv2v_reg  <= 1'b0;
      \piso.data_r_3166_sv2v_reg  <= 1'b0;
      \piso.data_r_3165_sv2v_reg  <= 1'b0;
      \piso.data_r_3164_sv2v_reg  <= 1'b0;
      \piso.data_r_3163_sv2v_reg  <= 1'b0;
      \piso.data_r_3162_sv2v_reg  <= 1'b0;
      \piso.data_r_3161_sv2v_reg  <= 1'b0;
      \piso.data_r_3160_sv2v_reg  <= 1'b0;
      \piso.data_r_3159_sv2v_reg  <= 1'b0;
      \piso.data_r_3158_sv2v_reg  <= 1'b0;
      \piso.data_r_3157_sv2v_reg  <= 1'b0;
      \piso.data_r_3156_sv2v_reg  <= 1'b0;
      \piso.data_r_3155_sv2v_reg  <= 1'b0;
      \piso.data_r_3154_sv2v_reg  <= 1'b0;
      \piso.data_r_3153_sv2v_reg  <= 1'b0;
      \piso.data_r_3152_sv2v_reg  <= 1'b0;
      \piso.data_r_3151_sv2v_reg  <= 1'b0;
      \piso.data_r_3150_sv2v_reg  <= 1'b0;
      \piso.data_r_3149_sv2v_reg  <= 1'b0;
      \piso.data_r_3148_sv2v_reg  <= 1'b0;
      \piso.data_r_3147_sv2v_reg  <= 1'b0;
      \piso.data_r_3146_sv2v_reg  <= 1'b0;
      \piso.data_r_3145_sv2v_reg  <= 1'b0;
      \piso.data_r_3144_sv2v_reg  <= 1'b0;
      \piso.data_r_3143_sv2v_reg  <= 1'b0;
      \piso.data_r_3142_sv2v_reg  <= 1'b0;
      \piso.data_r_3141_sv2v_reg  <= 1'b0;
      \piso.data_r_3140_sv2v_reg  <= 1'b0;
      \piso.data_r_3139_sv2v_reg  <= 1'b0;
      \piso.data_r_3138_sv2v_reg  <= 1'b0;
      \piso.data_r_3137_sv2v_reg  <= 1'b0;
      \piso.data_r_3136_sv2v_reg  <= 1'b0;
      \piso.data_r_3135_sv2v_reg  <= 1'b0;
      \piso.data_r_3134_sv2v_reg  <= 1'b0;
      \piso.data_r_3133_sv2v_reg  <= 1'b0;
      \piso.data_r_3132_sv2v_reg  <= 1'b0;
      \piso.data_r_3131_sv2v_reg  <= 1'b0;
      \piso.data_r_3130_sv2v_reg  <= 1'b0;
      \piso.data_r_3129_sv2v_reg  <= 1'b0;
      \piso.data_r_3128_sv2v_reg  <= 1'b0;
      \piso.data_r_3127_sv2v_reg  <= 1'b0;
      \piso.data_r_3126_sv2v_reg  <= 1'b0;
      \piso.data_r_3125_sv2v_reg  <= 1'b0;
      \piso.data_r_3124_sv2v_reg  <= 1'b0;
      \piso.data_r_3123_sv2v_reg  <= 1'b0;
      \piso.data_r_3122_sv2v_reg  <= 1'b0;
      \piso.data_r_3121_sv2v_reg  <= 1'b0;
      \piso.data_r_3120_sv2v_reg  <= 1'b0;
      \piso.data_r_3119_sv2v_reg  <= 1'b0;
      \piso.data_r_3118_sv2v_reg  <= 1'b0;
      \piso.data_r_3117_sv2v_reg  <= 1'b0;
      \piso.data_r_3116_sv2v_reg  <= 1'b0;
      \piso.data_r_3115_sv2v_reg  <= 1'b0;
      \piso.data_r_3114_sv2v_reg  <= 1'b0;
      \piso.data_r_3113_sv2v_reg  <= 1'b0;
      \piso.data_r_3112_sv2v_reg  <= 1'b0;
      \piso.data_r_3111_sv2v_reg  <= 1'b0;
      \piso.data_r_3110_sv2v_reg  <= 1'b0;
      \piso.data_r_3109_sv2v_reg  <= 1'b0;
      \piso.data_r_3108_sv2v_reg  <= 1'b0;
      \piso.data_r_3107_sv2v_reg  <= 1'b0;
      \piso.data_r_3106_sv2v_reg  <= 1'b0;
      \piso.data_r_3105_sv2v_reg  <= 1'b0;
      \piso.data_r_3104_sv2v_reg  <= 1'b0;
      \piso.data_r_3103_sv2v_reg  <= 1'b0;
      \piso.data_r_3102_sv2v_reg  <= 1'b0;
      \piso.data_r_3101_sv2v_reg  <= 1'b0;
      \piso.data_r_3100_sv2v_reg  <= 1'b0;
      \piso.data_r_3099_sv2v_reg  <= 1'b0;
      \piso.data_r_3098_sv2v_reg  <= 1'b0;
      \piso.data_r_3097_sv2v_reg  <= 1'b0;
      \piso.data_r_3096_sv2v_reg  <= 1'b0;
      \piso.data_r_3095_sv2v_reg  <= 1'b0;
      \piso.data_r_3094_sv2v_reg  <= 1'b0;
      \piso.data_r_3093_sv2v_reg  <= 1'b0;
      \piso.data_r_3092_sv2v_reg  <= 1'b0;
      \piso.data_r_3091_sv2v_reg  <= 1'b0;
      \piso.data_r_3090_sv2v_reg  <= 1'b0;
      \piso.data_r_3089_sv2v_reg  <= 1'b0;
      \piso.data_r_3088_sv2v_reg  <= 1'b0;
      \piso.data_r_3087_sv2v_reg  <= 1'b0;
      \piso.data_r_3086_sv2v_reg  <= 1'b0;
      \piso.data_r_3085_sv2v_reg  <= 1'b0;
      \piso.data_r_3084_sv2v_reg  <= 1'b0;
      \piso.data_r_3083_sv2v_reg  <= 1'b0;
      \piso.data_r_3082_sv2v_reg  <= 1'b0;
      \piso.data_r_3081_sv2v_reg  <= 1'b0;
      \piso.data_r_3080_sv2v_reg  <= 1'b0;
      \piso.data_r_3079_sv2v_reg  <= 1'b0;
      \piso.data_r_3078_sv2v_reg  <= 1'b0;
      \piso.data_r_3077_sv2v_reg  <= 1'b0;
      \piso.data_r_3076_sv2v_reg  <= 1'b0;
      \piso.data_r_3075_sv2v_reg  <= 1'b0;
      \piso.data_r_3074_sv2v_reg  <= 1'b0;
      \piso.data_r_3073_sv2v_reg  <= 1'b0;
      \piso.data_r_3072_sv2v_reg  <= 1'b0;
      \piso.data_r_3071_sv2v_reg  <= 1'b0;
      \piso.data_r_3070_sv2v_reg  <= 1'b0;
      \piso.data_r_3069_sv2v_reg  <= 1'b0;
      \piso.data_r_3068_sv2v_reg  <= 1'b0;
      \piso.data_r_3067_sv2v_reg  <= 1'b0;
      \piso.data_r_3066_sv2v_reg  <= 1'b0;
      \piso.data_r_3065_sv2v_reg  <= 1'b0;
      \piso.data_r_3064_sv2v_reg  <= 1'b0;
      \piso.data_r_3063_sv2v_reg  <= 1'b0;
      \piso.data_r_3062_sv2v_reg  <= 1'b0;
      \piso.data_r_3061_sv2v_reg  <= 1'b0;
      \piso.data_r_3060_sv2v_reg  <= 1'b0;
      \piso.data_r_3059_sv2v_reg  <= 1'b0;
      \piso.data_r_3058_sv2v_reg  <= 1'b0;
      \piso.data_r_3057_sv2v_reg  <= 1'b0;
      \piso.data_r_3056_sv2v_reg  <= 1'b0;
      \piso.data_r_3055_sv2v_reg  <= 1'b0;
      \piso.data_r_3054_sv2v_reg  <= 1'b0;
      \piso.data_r_3053_sv2v_reg  <= 1'b0;
      \piso.data_r_3052_sv2v_reg  <= 1'b0;
      \piso.data_r_3051_sv2v_reg  <= 1'b0;
      \piso.data_r_3050_sv2v_reg  <= 1'b0;
      \piso.data_r_3049_sv2v_reg  <= 1'b0;
      \piso.data_r_3048_sv2v_reg  <= 1'b0;
      \piso.data_r_3047_sv2v_reg  <= 1'b0;
      \piso.data_r_3046_sv2v_reg  <= 1'b0;
      \piso.data_r_3045_sv2v_reg  <= 1'b0;
      \piso.data_r_3044_sv2v_reg  <= 1'b0;
      \piso.data_r_3043_sv2v_reg  <= 1'b0;
      \piso.data_r_3042_sv2v_reg  <= 1'b0;
      \piso.data_r_3041_sv2v_reg  <= 1'b0;
      \piso.data_r_3040_sv2v_reg  <= 1'b0;
      \piso.data_r_3039_sv2v_reg  <= 1'b0;
      \piso.data_r_3038_sv2v_reg  <= 1'b0;
      \piso.data_r_3037_sv2v_reg  <= 1'b0;
      \piso.data_r_3036_sv2v_reg  <= 1'b0;
      \piso.data_r_3035_sv2v_reg  <= 1'b0;
      \piso.data_r_3034_sv2v_reg  <= 1'b0;
      \piso.data_r_3033_sv2v_reg  <= 1'b0;
      \piso.data_r_3032_sv2v_reg  <= 1'b0;
      \piso.data_r_3031_sv2v_reg  <= 1'b0;
      \piso.data_r_3030_sv2v_reg  <= 1'b0;
      \piso.data_r_3029_sv2v_reg  <= 1'b0;
      \piso.data_r_3028_sv2v_reg  <= 1'b0;
      \piso.data_r_3027_sv2v_reg  <= 1'b0;
      \piso.data_r_3026_sv2v_reg  <= 1'b0;
      \piso.data_r_3025_sv2v_reg  <= 1'b0;
      \piso.data_r_3024_sv2v_reg  <= 1'b0;
      \piso.data_r_3023_sv2v_reg  <= 1'b0;
      \piso.data_r_3022_sv2v_reg  <= 1'b0;
      \piso.data_r_3021_sv2v_reg  <= 1'b0;
      \piso.data_r_3020_sv2v_reg  <= 1'b0;
      \piso.data_r_3019_sv2v_reg  <= 1'b0;
      \piso.data_r_3018_sv2v_reg  <= 1'b0;
      \piso.data_r_3017_sv2v_reg  <= 1'b0;
      \piso.data_r_3016_sv2v_reg  <= 1'b0;
      \piso.data_r_3015_sv2v_reg  <= 1'b0;
      \piso.data_r_3014_sv2v_reg  <= 1'b0;
      \piso.data_r_3013_sv2v_reg  <= 1'b0;
      \piso.data_r_3012_sv2v_reg  <= 1'b0;
      \piso.data_r_3011_sv2v_reg  <= 1'b0;
      \piso.data_r_3010_sv2v_reg  <= 1'b0;
      \piso.data_r_3009_sv2v_reg  <= 1'b0;
      \piso.data_r_3008_sv2v_reg  <= 1'b0;
      \piso.data_r_3007_sv2v_reg  <= 1'b0;
      \piso.data_r_3006_sv2v_reg  <= 1'b0;
      \piso.data_r_3005_sv2v_reg  <= 1'b0;
      \piso.data_r_3004_sv2v_reg  <= 1'b0;
      \piso.data_r_3003_sv2v_reg  <= 1'b0;
      \piso.data_r_3002_sv2v_reg  <= 1'b0;
      \piso.data_r_3001_sv2v_reg  <= 1'b0;
      \piso.data_r_3000_sv2v_reg  <= 1'b0;
      \piso.data_r_2999_sv2v_reg  <= 1'b0;
      \piso.data_r_2998_sv2v_reg  <= 1'b0;
      \piso.data_r_2997_sv2v_reg  <= 1'b0;
      \piso.data_r_2996_sv2v_reg  <= 1'b0;
      \piso.data_r_2995_sv2v_reg  <= 1'b0;
      \piso.data_r_2994_sv2v_reg  <= 1'b0;
      \piso.data_r_2993_sv2v_reg  <= 1'b0;
      \piso.data_r_2992_sv2v_reg  <= 1'b0;
      \piso.data_r_2991_sv2v_reg  <= 1'b0;
      \piso.data_r_2990_sv2v_reg  <= 1'b0;
      \piso.data_r_2989_sv2v_reg  <= 1'b0;
      \piso.data_r_2988_sv2v_reg  <= 1'b0;
      \piso.data_r_2987_sv2v_reg  <= 1'b0;
      \piso.data_r_2986_sv2v_reg  <= 1'b0;
      \piso.data_r_2985_sv2v_reg  <= 1'b0;
      \piso.data_r_2984_sv2v_reg  <= 1'b0;
      \piso.data_r_2983_sv2v_reg  <= 1'b0;
      \piso.data_r_2982_sv2v_reg  <= 1'b0;
      \piso.data_r_2981_sv2v_reg  <= 1'b0;
      \piso.data_r_2980_sv2v_reg  <= 1'b0;
      \piso.data_r_2979_sv2v_reg  <= 1'b0;
      \piso.data_r_2978_sv2v_reg  <= 1'b0;
      \piso.data_r_2977_sv2v_reg  <= 1'b0;
      \piso.data_r_2976_sv2v_reg  <= 1'b0;
      \piso.data_r_2975_sv2v_reg  <= 1'b0;
      \piso.data_r_2974_sv2v_reg  <= 1'b0;
      \piso.data_r_2973_sv2v_reg  <= 1'b0;
      \piso.data_r_2972_sv2v_reg  <= 1'b0;
      \piso.data_r_2971_sv2v_reg  <= 1'b0;
      \piso.data_r_2970_sv2v_reg  <= 1'b0;
      \piso.data_r_2969_sv2v_reg  <= 1'b0;
      \piso.data_r_2968_sv2v_reg  <= 1'b0;
      \piso.data_r_2967_sv2v_reg  <= 1'b0;
      \piso.data_r_2966_sv2v_reg  <= 1'b0;
      \piso.data_r_2965_sv2v_reg  <= 1'b0;
      \piso.data_r_2964_sv2v_reg  <= 1'b0;
      \piso.data_r_2963_sv2v_reg  <= 1'b0;
      \piso.data_r_2962_sv2v_reg  <= 1'b0;
      \piso.data_r_2961_sv2v_reg  <= 1'b0;
      \piso.data_r_2960_sv2v_reg  <= 1'b0;
      \piso.data_r_2959_sv2v_reg  <= 1'b0;
      \piso.data_r_2958_sv2v_reg  <= 1'b0;
      \piso.data_r_2957_sv2v_reg  <= 1'b0;
      \piso.data_r_2956_sv2v_reg  <= 1'b0;
      \piso.data_r_2955_sv2v_reg  <= 1'b0;
      \piso.data_r_2954_sv2v_reg  <= 1'b0;
      \piso.data_r_2953_sv2v_reg  <= 1'b0;
      \piso.data_r_2952_sv2v_reg  <= 1'b0;
      \piso.data_r_2951_sv2v_reg  <= 1'b0;
      \piso.data_r_2950_sv2v_reg  <= 1'b0;
      \piso.data_r_2949_sv2v_reg  <= 1'b0;
      \piso.data_r_2948_sv2v_reg  <= 1'b0;
      \piso.data_r_2947_sv2v_reg  <= 1'b0;
      \piso.data_r_2946_sv2v_reg  <= 1'b0;
      \piso.data_r_2945_sv2v_reg  <= 1'b0;
      \piso.data_r_2944_sv2v_reg  <= 1'b0;
      \piso.data_r_2943_sv2v_reg  <= 1'b0;
      \piso.data_r_2942_sv2v_reg  <= 1'b0;
      \piso.data_r_2941_sv2v_reg  <= 1'b0;
      \piso.data_r_2940_sv2v_reg  <= 1'b0;
      \piso.data_r_2939_sv2v_reg  <= 1'b0;
      \piso.data_r_2938_sv2v_reg  <= 1'b0;
      \piso.data_r_2937_sv2v_reg  <= 1'b0;
      \piso.data_r_2936_sv2v_reg  <= 1'b0;
      \piso.data_r_2935_sv2v_reg  <= 1'b0;
      \piso.data_r_2934_sv2v_reg  <= 1'b0;
      \piso.data_r_2933_sv2v_reg  <= 1'b0;
      \piso.data_r_2932_sv2v_reg  <= 1'b0;
      \piso.data_r_2931_sv2v_reg  <= 1'b0;
      \piso.data_r_2930_sv2v_reg  <= 1'b0;
      \piso.data_r_2929_sv2v_reg  <= 1'b0;
      \piso.data_r_2928_sv2v_reg  <= 1'b0;
      \piso.data_r_2927_sv2v_reg  <= 1'b0;
      \piso.data_r_2926_sv2v_reg  <= 1'b0;
      \piso.data_r_2925_sv2v_reg  <= 1'b0;
      \piso.data_r_2924_sv2v_reg  <= 1'b0;
      \piso.data_r_2923_sv2v_reg  <= 1'b0;
      \piso.data_r_2922_sv2v_reg  <= 1'b0;
      \piso.data_r_2921_sv2v_reg  <= 1'b0;
      \piso.data_r_2920_sv2v_reg  <= 1'b0;
      \piso.data_r_2919_sv2v_reg  <= 1'b0;
      \piso.data_r_2918_sv2v_reg  <= 1'b0;
      \piso.data_r_2917_sv2v_reg  <= 1'b0;
      \piso.data_r_2916_sv2v_reg  <= 1'b0;
      \piso.data_r_2915_sv2v_reg  <= 1'b0;
      \piso.data_r_2914_sv2v_reg  <= 1'b0;
      \piso.data_r_2913_sv2v_reg  <= 1'b0;
      \piso.data_r_2912_sv2v_reg  <= 1'b0;
      \piso.data_r_2911_sv2v_reg  <= 1'b0;
      \piso.data_r_2910_sv2v_reg  <= 1'b0;
      \piso.data_r_2909_sv2v_reg  <= 1'b0;
      \piso.data_r_2908_sv2v_reg  <= 1'b0;
      \piso.data_r_2907_sv2v_reg  <= 1'b0;
      \piso.data_r_2906_sv2v_reg  <= 1'b0;
      \piso.data_r_2905_sv2v_reg  <= 1'b0;
      \piso.data_r_2904_sv2v_reg  <= 1'b0;
      \piso.data_r_2903_sv2v_reg  <= 1'b0;
      \piso.data_r_2902_sv2v_reg  <= 1'b0;
      \piso.data_r_2901_sv2v_reg  <= 1'b0;
      \piso.data_r_2900_sv2v_reg  <= 1'b0;
      \piso.data_r_2899_sv2v_reg  <= 1'b0;
      \piso.data_r_2898_sv2v_reg  <= 1'b0;
      \piso.data_r_2897_sv2v_reg  <= 1'b0;
      \piso.data_r_2896_sv2v_reg  <= 1'b0;
      \piso.data_r_2895_sv2v_reg  <= 1'b0;
      \piso.data_r_2894_sv2v_reg  <= 1'b0;
      \piso.data_r_2893_sv2v_reg  <= 1'b0;
      \piso.data_r_2892_sv2v_reg  <= 1'b0;
      \piso.data_r_2891_sv2v_reg  <= 1'b0;
      \piso.data_r_2890_sv2v_reg  <= 1'b0;
      \piso.data_r_2889_sv2v_reg  <= 1'b0;
      \piso.data_r_2888_sv2v_reg  <= 1'b0;
      \piso.data_r_2887_sv2v_reg  <= 1'b0;
      \piso.data_r_2886_sv2v_reg  <= 1'b0;
      \piso.data_r_2885_sv2v_reg  <= 1'b0;
      \piso.data_r_2884_sv2v_reg  <= 1'b0;
      \piso.data_r_2883_sv2v_reg  <= 1'b0;
      \piso.data_r_2882_sv2v_reg  <= 1'b0;
      \piso.data_r_2881_sv2v_reg  <= 1'b0;
      \piso.data_r_2880_sv2v_reg  <= 1'b0;
      \piso.data_r_2879_sv2v_reg  <= 1'b0;
      \piso.data_r_2878_sv2v_reg  <= 1'b0;
      \piso.data_r_2877_sv2v_reg  <= 1'b0;
      \piso.data_r_2876_sv2v_reg  <= 1'b0;
      \piso.data_r_2875_sv2v_reg  <= 1'b0;
      \piso.data_r_2874_sv2v_reg  <= 1'b0;
      \piso.data_r_2873_sv2v_reg  <= 1'b0;
      \piso.data_r_2872_sv2v_reg  <= 1'b0;
      \piso.data_r_2871_sv2v_reg  <= 1'b0;
      \piso.data_r_2870_sv2v_reg  <= 1'b0;
      \piso.data_r_2869_sv2v_reg  <= 1'b0;
      \piso.data_r_2868_sv2v_reg  <= 1'b0;
      \piso.data_r_2867_sv2v_reg  <= 1'b0;
      \piso.data_r_2866_sv2v_reg  <= 1'b0;
      \piso.data_r_2865_sv2v_reg  <= 1'b0;
      \piso.data_r_2864_sv2v_reg  <= 1'b0;
      \piso.data_r_2863_sv2v_reg  <= 1'b0;
      \piso.data_r_2862_sv2v_reg  <= 1'b0;
      \piso.data_r_2861_sv2v_reg  <= 1'b0;
      \piso.data_r_2860_sv2v_reg  <= 1'b0;
      \piso.data_r_2859_sv2v_reg  <= 1'b0;
      \piso.data_r_2858_sv2v_reg  <= 1'b0;
      \piso.data_r_2857_sv2v_reg  <= 1'b0;
      \piso.data_r_2856_sv2v_reg  <= 1'b0;
      \piso.data_r_2855_sv2v_reg  <= 1'b0;
      \piso.data_r_2854_sv2v_reg  <= 1'b0;
      \piso.data_r_2853_sv2v_reg  <= 1'b0;
      \piso.data_r_2852_sv2v_reg  <= 1'b0;
      \piso.data_r_2851_sv2v_reg  <= 1'b0;
      \piso.data_r_2850_sv2v_reg  <= 1'b0;
      \piso.data_r_2849_sv2v_reg  <= 1'b0;
      \piso.data_r_2848_sv2v_reg  <= 1'b0;
      \piso.data_r_2847_sv2v_reg  <= 1'b0;
      \piso.data_r_2846_sv2v_reg  <= 1'b0;
      \piso.data_r_2845_sv2v_reg  <= 1'b0;
      \piso.data_r_2844_sv2v_reg  <= 1'b0;
      \piso.data_r_2843_sv2v_reg  <= 1'b0;
      \piso.data_r_2842_sv2v_reg  <= 1'b0;
      \piso.data_r_2841_sv2v_reg  <= 1'b0;
      \piso.data_r_2840_sv2v_reg  <= 1'b0;
      \piso.data_r_2839_sv2v_reg  <= 1'b0;
      \piso.data_r_2838_sv2v_reg  <= 1'b0;
      \piso.data_r_2837_sv2v_reg  <= 1'b0;
      \piso.data_r_2836_sv2v_reg  <= 1'b0;
      \piso.data_r_2835_sv2v_reg  <= 1'b0;
      \piso.data_r_2834_sv2v_reg  <= 1'b0;
      \piso.data_r_2833_sv2v_reg  <= 1'b0;
      \piso.data_r_2832_sv2v_reg  <= 1'b0;
      \piso.data_r_2831_sv2v_reg  <= 1'b0;
      \piso.data_r_2830_sv2v_reg  <= 1'b0;
      \piso.data_r_2829_sv2v_reg  <= 1'b0;
      \piso.data_r_2828_sv2v_reg  <= 1'b0;
      \piso.data_r_2827_sv2v_reg  <= 1'b0;
      \piso.data_r_2826_sv2v_reg  <= 1'b0;
      \piso.data_r_2825_sv2v_reg  <= 1'b0;
      \piso.data_r_2824_sv2v_reg  <= 1'b0;
      \piso.data_r_2823_sv2v_reg  <= 1'b0;
      \piso.data_r_2822_sv2v_reg  <= 1'b0;
      \piso.data_r_2821_sv2v_reg  <= 1'b0;
      \piso.data_r_2820_sv2v_reg  <= 1'b0;
      \piso.data_r_2819_sv2v_reg  <= 1'b0;
      \piso.data_r_2818_sv2v_reg  <= 1'b0;
      \piso.data_r_2817_sv2v_reg  <= 1'b0;
      \piso.data_r_2816_sv2v_reg  <= 1'b0;
      \piso.data_r_2815_sv2v_reg  <= 1'b0;
      \piso.data_r_2814_sv2v_reg  <= 1'b0;
      \piso.data_r_2813_sv2v_reg  <= 1'b0;
      \piso.data_r_2812_sv2v_reg  <= 1'b0;
      \piso.data_r_2811_sv2v_reg  <= 1'b0;
      \piso.data_r_2810_sv2v_reg  <= 1'b0;
      \piso.data_r_2809_sv2v_reg  <= 1'b0;
      \piso.data_r_2808_sv2v_reg  <= 1'b0;
      \piso.data_r_2807_sv2v_reg  <= 1'b0;
      \piso.data_r_2806_sv2v_reg  <= 1'b0;
      \piso.data_r_2805_sv2v_reg  <= 1'b0;
      \piso.data_r_2804_sv2v_reg  <= 1'b0;
      \piso.data_r_2803_sv2v_reg  <= 1'b0;
      \piso.data_r_2802_sv2v_reg  <= 1'b0;
      \piso.data_r_2801_sv2v_reg  <= 1'b0;
      \piso.data_r_2800_sv2v_reg  <= 1'b0;
      \piso.data_r_2799_sv2v_reg  <= 1'b0;
      \piso.data_r_2798_sv2v_reg  <= 1'b0;
      \piso.data_r_2797_sv2v_reg  <= 1'b0;
      \piso.data_r_2796_sv2v_reg  <= 1'b0;
      \piso.data_r_2795_sv2v_reg  <= 1'b0;
      \piso.data_r_2794_sv2v_reg  <= 1'b0;
      \piso.data_r_2793_sv2v_reg  <= 1'b0;
      \piso.data_r_2792_sv2v_reg  <= 1'b0;
      \piso.data_r_2791_sv2v_reg  <= 1'b0;
      \piso.data_r_2790_sv2v_reg  <= 1'b0;
      \piso.data_r_2789_sv2v_reg  <= 1'b0;
      \piso.data_r_2788_sv2v_reg  <= 1'b0;
      \piso.data_r_2787_sv2v_reg  <= 1'b0;
      \piso.data_r_2786_sv2v_reg  <= 1'b0;
      \piso.data_r_2785_sv2v_reg  <= 1'b0;
      \piso.data_r_2784_sv2v_reg  <= 1'b0;
      \piso.data_r_2783_sv2v_reg  <= 1'b0;
      \piso.data_r_2782_sv2v_reg  <= 1'b0;
      \piso.data_r_2781_sv2v_reg  <= 1'b0;
      \piso.data_r_2780_sv2v_reg  <= 1'b0;
      \piso.data_r_2779_sv2v_reg  <= 1'b0;
      \piso.data_r_2778_sv2v_reg  <= 1'b0;
      \piso.data_r_2777_sv2v_reg  <= 1'b0;
      \piso.data_r_2776_sv2v_reg  <= 1'b0;
      \piso.data_r_2775_sv2v_reg  <= 1'b0;
      \piso.data_r_2774_sv2v_reg  <= 1'b0;
      \piso.data_r_2773_sv2v_reg  <= 1'b0;
      \piso.data_r_2772_sv2v_reg  <= 1'b0;
      \piso.data_r_2771_sv2v_reg  <= 1'b0;
      \piso.data_r_2770_sv2v_reg  <= 1'b0;
      \piso.data_r_2769_sv2v_reg  <= 1'b0;
      \piso.data_r_2768_sv2v_reg  <= 1'b0;
      \piso.data_r_2767_sv2v_reg  <= 1'b0;
      \piso.data_r_2766_sv2v_reg  <= 1'b0;
      \piso.data_r_2765_sv2v_reg  <= 1'b0;
      \piso.data_r_2764_sv2v_reg  <= 1'b0;
      \piso.data_r_2763_sv2v_reg  <= 1'b0;
      \piso.data_r_2762_sv2v_reg  <= 1'b0;
      \piso.data_r_2761_sv2v_reg  <= 1'b0;
      \piso.data_r_2760_sv2v_reg  <= 1'b0;
      \piso.data_r_2759_sv2v_reg  <= 1'b0;
      \piso.data_r_2758_sv2v_reg  <= 1'b0;
      \piso.data_r_2757_sv2v_reg  <= 1'b0;
      \piso.data_r_2756_sv2v_reg  <= 1'b0;
      \piso.data_r_2755_sv2v_reg  <= 1'b0;
      \piso.data_r_2754_sv2v_reg  <= 1'b0;
      \piso.data_r_2753_sv2v_reg  <= 1'b0;
      \piso.data_r_2752_sv2v_reg  <= 1'b0;
      \piso.data_r_2751_sv2v_reg  <= 1'b0;
      \piso.data_r_2750_sv2v_reg  <= 1'b0;
      \piso.data_r_2749_sv2v_reg  <= 1'b0;
      \piso.data_r_2748_sv2v_reg  <= 1'b0;
      \piso.data_r_2747_sv2v_reg  <= 1'b0;
      \piso.data_r_2746_sv2v_reg  <= 1'b0;
      \piso.data_r_2745_sv2v_reg  <= 1'b0;
      \piso.data_r_2744_sv2v_reg  <= 1'b0;
      \piso.data_r_2743_sv2v_reg  <= 1'b0;
      \piso.data_r_2742_sv2v_reg  <= 1'b0;
      \piso.data_r_2741_sv2v_reg  <= 1'b0;
      \piso.data_r_2740_sv2v_reg  <= 1'b0;
      \piso.data_r_2739_sv2v_reg  <= 1'b0;
      \piso.data_r_2738_sv2v_reg  <= 1'b0;
      \piso.data_r_2737_sv2v_reg  <= 1'b0;
      \piso.data_r_2736_sv2v_reg  <= 1'b0;
      \piso.data_r_2735_sv2v_reg  <= 1'b0;
      \piso.data_r_2734_sv2v_reg  <= 1'b0;
      \piso.data_r_2733_sv2v_reg  <= 1'b0;
      \piso.data_r_2732_sv2v_reg  <= 1'b0;
      \piso.data_r_2731_sv2v_reg  <= 1'b0;
      \piso.data_r_2730_sv2v_reg  <= 1'b0;
      \piso.data_r_2729_sv2v_reg  <= 1'b0;
      \piso.data_r_2728_sv2v_reg  <= 1'b0;
      \piso.data_r_2727_sv2v_reg  <= 1'b0;
      \piso.data_r_2726_sv2v_reg  <= 1'b0;
      \piso.data_r_2725_sv2v_reg  <= 1'b0;
      \piso.data_r_2724_sv2v_reg  <= 1'b0;
      \piso.data_r_2723_sv2v_reg  <= 1'b0;
      \piso.data_r_2722_sv2v_reg  <= 1'b0;
      \piso.data_r_2721_sv2v_reg  <= 1'b0;
      \piso.data_r_2720_sv2v_reg  <= 1'b0;
      \piso.data_r_2719_sv2v_reg  <= 1'b0;
      \piso.data_r_2718_sv2v_reg  <= 1'b0;
      \piso.data_r_2717_sv2v_reg  <= 1'b0;
      \piso.data_r_2716_sv2v_reg  <= 1'b0;
      \piso.data_r_2715_sv2v_reg  <= 1'b0;
      \piso.data_r_2714_sv2v_reg  <= 1'b0;
      \piso.data_r_2713_sv2v_reg  <= 1'b0;
      \piso.data_r_2712_sv2v_reg  <= 1'b0;
      \piso.data_r_2711_sv2v_reg  <= 1'b0;
      \piso.data_r_2710_sv2v_reg  <= 1'b0;
      \piso.data_r_2709_sv2v_reg  <= 1'b0;
      \piso.data_r_2708_sv2v_reg  <= 1'b0;
      \piso.data_r_2707_sv2v_reg  <= 1'b0;
      \piso.data_r_2706_sv2v_reg  <= 1'b0;
      \piso.data_r_2705_sv2v_reg  <= 1'b0;
      \piso.data_r_2704_sv2v_reg  <= 1'b0;
      \piso.data_r_2703_sv2v_reg  <= 1'b0;
      \piso.data_r_2702_sv2v_reg  <= 1'b0;
      \piso.data_r_2701_sv2v_reg  <= 1'b0;
      \piso.data_r_2700_sv2v_reg  <= 1'b0;
      \piso.data_r_2699_sv2v_reg  <= 1'b0;
      \piso.data_r_2698_sv2v_reg  <= 1'b0;
      \piso.data_r_2697_sv2v_reg  <= 1'b0;
      \piso.data_r_2696_sv2v_reg  <= 1'b0;
      \piso.data_r_2695_sv2v_reg  <= 1'b0;
      \piso.data_r_2694_sv2v_reg  <= 1'b0;
      \piso.data_r_2693_sv2v_reg  <= 1'b0;
      \piso.data_r_2692_sv2v_reg  <= 1'b0;
      \piso.data_r_2691_sv2v_reg  <= 1'b0;
      \piso.data_r_2690_sv2v_reg  <= 1'b0;
      \piso.data_r_2689_sv2v_reg  <= 1'b0;
      \piso.data_r_2688_sv2v_reg  <= 1'b0;
      \piso.data_r_2687_sv2v_reg  <= 1'b0;
      \piso.data_r_2686_sv2v_reg  <= 1'b0;
      \piso.data_r_2685_sv2v_reg  <= 1'b0;
      \piso.data_r_2684_sv2v_reg  <= 1'b0;
      \piso.data_r_2683_sv2v_reg  <= 1'b0;
      \piso.data_r_2682_sv2v_reg  <= 1'b0;
      \piso.data_r_2681_sv2v_reg  <= 1'b0;
      \piso.data_r_2680_sv2v_reg  <= 1'b0;
      \piso.data_r_2679_sv2v_reg  <= 1'b0;
      \piso.data_r_2678_sv2v_reg  <= 1'b0;
      \piso.data_r_2677_sv2v_reg  <= 1'b0;
      \piso.data_r_2676_sv2v_reg  <= 1'b0;
      \piso.data_r_2675_sv2v_reg  <= 1'b0;
      \piso.data_r_2674_sv2v_reg  <= 1'b0;
      \piso.data_r_2673_sv2v_reg  <= 1'b0;
      \piso.data_r_2672_sv2v_reg  <= 1'b0;
      \piso.data_r_2671_sv2v_reg  <= 1'b0;
      \piso.data_r_2670_sv2v_reg  <= 1'b0;
      \piso.data_r_2669_sv2v_reg  <= 1'b0;
      \piso.data_r_2668_sv2v_reg  <= 1'b0;
      \piso.data_r_2667_sv2v_reg  <= 1'b0;
      \piso.data_r_2666_sv2v_reg  <= 1'b0;
      \piso.data_r_2665_sv2v_reg  <= 1'b0;
      \piso.data_r_2664_sv2v_reg  <= 1'b0;
      \piso.data_r_2663_sv2v_reg  <= 1'b0;
      \piso.data_r_2662_sv2v_reg  <= 1'b0;
      \piso.data_r_2661_sv2v_reg  <= 1'b0;
      \piso.data_r_2660_sv2v_reg  <= 1'b0;
      \piso.data_r_2659_sv2v_reg  <= 1'b0;
      \piso.data_r_2658_sv2v_reg  <= 1'b0;
      \piso.data_r_2657_sv2v_reg  <= 1'b0;
      \piso.data_r_2656_sv2v_reg  <= 1'b0;
      \piso.data_r_2655_sv2v_reg  <= 1'b0;
      \piso.data_r_2654_sv2v_reg  <= 1'b0;
      \piso.data_r_2653_sv2v_reg  <= 1'b0;
      \piso.data_r_2652_sv2v_reg  <= 1'b0;
      \piso.data_r_2651_sv2v_reg  <= 1'b0;
      \piso.data_r_2650_sv2v_reg  <= 1'b0;
      \piso.data_r_2649_sv2v_reg  <= 1'b0;
      \piso.data_r_2648_sv2v_reg  <= 1'b0;
      \piso.data_r_2647_sv2v_reg  <= 1'b0;
      \piso.data_r_2646_sv2v_reg  <= 1'b0;
      \piso.data_r_2645_sv2v_reg  <= 1'b0;
      \piso.data_r_2644_sv2v_reg  <= 1'b0;
      \piso.data_r_2643_sv2v_reg  <= 1'b0;
      \piso.data_r_2642_sv2v_reg  <= 1'b0;
      \piso.data_r_2641_sv2v_reg  <= 1'b0;
      \piso.data_r_2640_sv2v_reg  <= 1'b0;
      \piso.data_r_2639_sv2v_reg  <= 1'b0;
      \piso.data_r_2638_sv2v_reg  <= 1'b0;
      \piso.data_r_2637_sv2v_reg  <= 1'b0;
      \piso.data_r_2636_sv2v_reg  <= 1'b0;
      \piso.data_r_2635_sv2v_reg  <= 1'b0;
      \piso.data_r_2634_sv2v_reg  <= 1'b0;
      \piso.data_r_2633_sv2v_reg  <= 1'b0;
      \piso.data_r_2632_sv2v_reg  <= 1'b0;
      \piso.data_r_2631_sv2v_reg  <= 1'b0;
      \piso.data_r_2630_sv2v_reg  <= 1'b0;
      \piso.data_r_2629_sv2v_reg  <= 1'b0;
      \piso.data_r_2628_sv2v_reg  <= 1'b0;
      \piso.data_r_2627_sv2v_reg  <= 1'b0;
      \piso.data_r_2626_sv2v_reg  <= 1'b0;
      \piso.data_r_2625_sv2v_reg  <= 1'b0;
      \piso.data_r_2624_sv2v_reg  <= 1'b0;
      \piso.data_r_2623_sv2v_reg  <= 1'b0;
      \piso.data_r_2622_sv2v_reg  <= 1'b0;
      \piso.data_r_2621_sv2v_reg  <= 1'b0;
      \piso.data_r_2620_sv2v_reg  <= 1'b0;
      \piso.data_r_2619_sv2v_reg  <= 1'b0;
      \piso.data_r_2618_sv2v_reg  <= 1'b0;
      \piso.data_r_2617_sv2v_reg  <= 1'b0;
      \piso.data_r_2616_sv2v_reg  <= 1'b0;
      \piso.data_r_2615_sv2v_reg  <= 1'b0;
      \piso.data_r_2614_sv2v_reg  <= 1'b0;
      \piso.data_r_2613_sv2v_reg  <= 1'b0;
      \piso.data_r_2612_sv2v_reg  <= 1'b0;
      \piso.data_r_2611_sv2v_reg  <= 1'b0;
      \piso.data_r_2610_sv2v_reg  <= 1'b0;
      \piso.data_r_2609_sv2v_reg  <= 1'b0;
      \piso.data_r_2608_sv2v_reg  <= 1'b0;
      \piso.data_r_2607_sv2v_reg  <= 1'b0;
      \piso.data_r_2606_sv2v_reg  <= 1'b0;
      \piso.data_r_2605_sv2v_reg  <= 1'b0;
      \piso.data_r_2604_sv2v_reg  <= 1'b0;
      \piso.data_r_2603_sv2v_reg  <= 1'b0;
      \piso.data_r_2602_sv2v_reg  <= 1'b0;
      \piso.data_r_2601_sv2v_reg  <= 1'b0;
      \piso.data_r_2600_sv2v_reg  <= 1'b0;
      \piso.data_r_2599_sv2v_reg  <= 1'b0;
      \piso.data_r_2598_sv2v_reg  <= 1'b0;
      \piso.data_r_2597_sv2v_reg  <= 1'b0;
      \piso.data_r_2596_sv2v_reg  <= 1'b0;
      \piso.data_r_2595_sv2v_reg  <= 1'b0;
      \piso.data_r_2594_sv2v_reg  <= 1'b0;
      \piso.data_r_2593_sv2v_reg  <= 1'b0;
      \piso.data_r_2592_sv2v_reg  <= 1'b0;
      \piso.data_r_2591_sv2v_reg  <= 1'b0;
      \piso.data_r_2590_sv2v_reg  <= 1'b0;
      \piso.data_r_2589_sv2v_reg  <= 1'b0;
      \piso.data_r_2588_sv2v_reg  <= 1'b0;
      \piso.data_r_2587_sv2v_reg  <= 1'b0;
      \piso.data_r_2586_sv2v_reg  <= 1'b0;
      \piso.data_r_2585_sv2v_reg  <= 1'b0;
      \piso.data_r_2584_sv2v_reg  <= 1'b0;
      \piso.data_r_2583_sv2v_reg  <= 1'b0;
      \piso.data_r_2582_sv2v_reg  <= 1'b0;
      \piso.data_r_2581_sv2v_reg  <= 1'b0;
      \piso.data_r_2580_sv2v_reg  <= 1'b0;
      \piso.data_r_2579_sv2v_reg  <= 1'b0;
      \piso.data_r_2578_sv2v_reg  <= 1'b0;
      \piso.data_r_2577_sv2v_reg  <= 1'b0;
      \piso.data_r_2576_sv2v_reg  <= 1'b0;
      \piso.data_r_2575_sv2v_reg  <= 1'b0;
      \piso.data_r_2574_sv2v_reg  <= 1'b0;
      \piso.data_r_2573_sv2v_reg  <= 1'b0;
      \piso.data_r_2572_sv2v_reg  <= 1'b0;
      \piso.data_r_2571_sv2v_reg  <= 1'b0;
      \piso.data_r_2570_sv2v_reg  <= 1'b0;
      \piso.data_r_2569_sv2v_reg  <= 1'b0;
      \piso.data_r_2568_sv2v_reg  <= 1'b0;
      \piso.data_r_2567_sv2v_reg  <= 1'b0;
      \piso.data_r_2566_sv2v_reg  <= 1'b0;
      \piso.data_r_2565_sv2v_reg  <= 1'b0;
      \piso.data_r_2564_sv2v_reg  <= 1'b0;
      \piso.data_r_2563_sv2v_reg  <= 1'b0;
      \piso.data_r_2562_sv2v_reg  <= 1'b0;
      \piso.data_r_2561_sv2v_reg  <= 1'b0;
      \piso.data_r_2560_sv2v_reg  <= 1'b0;
      \piso.data_r_2559_sv2v_reg  <= 1'b0;
      \piso.data_r_2558_sv2v_reg  <= 1'b0;
      \piso.data_r_2557_sv2v_reg  <= 1'b0;
      \piso.data_r_2556_sv2v_reg  <= 1'b0;
      \piso.data_r_2555_sv2v_reg  <= 1'b0;
      \piso.data_r_2554_sv2v_reg  <= 1'b0;
      \piso.data_r_2553_sv2v_reg  <= 1'b0;
      \piso.data_r_2552_sv2v_reg  <= 1'b0;
      \piso.data_r_2551_sv2v_reg  <= 1'b0;
      \piso.data_r_2550_sv2v_reg  <= 1'b0;
      \piso.data_r_2549_sv2v_reg  <= 1'b0;
      \piso.data_r_2548_sv2v_reg  <= 1'b0;
      \piso.data_r_2547_sv2v_reg  <= 1'b0;
      \piso.data_r_2546_sv2v_reg  <= 1'b0;
      \piso.data_r_2545_sv2v_reg  <= 1'b0;
      \piso.data_r_2544_sv2v_reg  <= 1'b0;
      \piso.data_r_2543_sv2v_reg  <= 1'b0;
      \piso.data_r_2542_sv2v_reg  <= 1'b0;
      \piso.data_r_2541_sv2v_reg  <= 1'b0;
      \piso.data_r_2540_sv2v_reg  <= 1'b0;
      \piso.data_r_2539_sv2v_reg  <= 1'b0;
      \piso.data_r_2538_sv2v_reg  <= 1'b0;
      \piso.data_r_2537_sv2v_reg  <= 1'b0;
      \piso.data_r_2536_sv2v_reg  <= 1'b0;
      \piso.data_r_2535_sv2v_reg  <= 1'b0;
      \piso.data_r_2534_sv2v_reg  <= 1'b0;
      \piso.data_r_2533_sv2v_reg  <= 1'b0;
      \piso.data_r_2532_sv2v_reg  <= 1'b0;
      \piso.data_r_2531_sv2v_reg  <= 1'b0;
      \piso.data_r_2530_sv2v_reg  <= 1'b0;
      \piso.data_r_2529_sv2v_reg  <= 1'b0;
      \piso.data_r_2528_sv2v_reg  <= 1'b0;
      \piso.data_r_2527_sv2v_reg  <= 1'b0;
      \piso.data_r_2526_sv2v_reg  <= 1'b0;
      \piso.data_r_2525_sv2v_reg  <= 1'b0;
      \piso.data_r_2524_sv2v_reg  <= 1'b0;
      \piso.data_r_2523_sv2v_reg  <= 1'b0;
      \piso.data_r_2522_sv2v_reg  <= 1'b0;
      \piso.data_r_2521_sv2v_reg  <= 1'b0;
      \piso.data_r_2520_sv2v_reg  <= 1'b0;
      \piso.data_r_2519_sv2v_reg  <= 1'b0;
      \piso.data_r_2518_sv2v_reg  <= 1'b0;
      \piso.data_r_2517_sv2v_reg  <= 1'b0;
      \piso.data_r_2516_sv2v_reg  <= 1'b0;
      \piso.data_r_2515_sv2v_reg  <= 1'b0;
      \piso.data_r_2514_sv2v_reg  <= 1'b0;
      \piso.data_r_2513_sv2v_reg  <= 1'b0;
      \piso.data_r_2512_sv2v_reg  <= 1'b0;
      \piso.data_r_2511_sv2v_reg  <= 1'b0;
      \piso.data_r_2510_sv2v_reg  <= 1'b0;
      \piso.data_r_2509_sv2v_reg  <= 1'b0;
      \piso.data_r_2508_sv2v_reg  <= 1'b0;
      \piso.data_r_2507_sv2v_reg  <= 1'b0;
      \piso.data_r_2506_sv2v_reg  <= 1'b0;
      \piso.data_r_2505_sv2v_reg  <= 1'b0;
      \piso.data_r_2504_sv2v_reg  <= 1'b0;
      \piso.data_r_2503_sv2v_reg  <= 1'b0;
      \piso.data_r_2502_sv2v_reg  <= 1'b0;
      \piso.data_r_2501_sv2v_reg  <= 1'b0;
      \piso.data_r_2500_sv2v_reg  <= 1'b0;
      \piso.data_r_2499_sv2v_reg  <= 1'b0;
      \piso.data_r_2498_sv2v_reg  <= 1'b0;
      \piso.data_r_2497_sv2v_reg  <= 1'b0;
      \piso.data_r_2496_sv2v_reg  <= 1'b0;
      \piso.data_r_2495_sv2v_reg  <= 1'b0;
      \piso.data_r_2494_sv2v_reg  <= 1'b0;
      \piso.data_r_2493_sv2v_reg  <= 1'b0;
      \piso.data_r_2492_sv2v_reg  <= 1'b0;
      \piso.data_r_2491_sv2v_reg  <= 1'b0;
      \piso.data_r_2490_sv2v_reg  <= 1'b0;
      \piso.data_r_2489_sv2v_reg  <= 1'b0;
      \piso.data_r_2488_sv2v_reg  <= 1'b0;
      \piso.data_r_2487_sv2v_reg  <= 1'b0;
      \piso.data_r_2486_sv2v_reg  <= 1'b0;
      \piso.data_r_2485_sv2v_reg  <= 1'b0;
      \piso.data_r_2484_sv2v_reg  <= 1'b0;
      \piso.data_r_2483_sv2v_reg  <= 1'b0;
      \piso.data_r_2482_sv2v_reg  <= 1'b0;
      \piso.data_r_2481_sv2v_reg  <= 1'b0;
      \piso.data_r_2480_sv2v_reg  <= 1'b0;
      \piso.data_r_2479_sv2v_reg  <= 1'b0;
      \piso.data_r_2478_sv2v_reg  <= 1'b0;
      \piso.data_r_2477_sv2v_reg  <= 1'b0;
      \piso.data_r_2476_sv2v_reg  <= 1'b0;
      \piso.data_r_2475_sv2v_reg  <= 1'b0;
      \piso.data_r_2474_sv2v_reg  <= 1'b0;
      \piso.data_r_2473_sv2v_reg  <= 1'b0;
      \piso.data_r_2472_sv2v_reg  <= 1'b0;
      \piso.data_r_2471_sv2v_reg  <= 1'b0;
      \piso.data_r_2470_sv2v_reg  <= 1'b0;
      \piso.data_r_2469_sv2v_reg  <= 1'b0;
      \piso.data_r_2468_sv2v_reg  <= 1'b0;
      \piso.data_r_2467_sv2v_reg  <= 1'b0;
      \piso.data_r_2466_sv2v_reg  <= 1'b0;
      \piso.data_r_2465_sv2v_reg  <= 1'b0;
      \piso.data_r_2464_sv2v_reg  <= 1'b0;
      \piso.data_r_2463_sv2v_reg  <= 1'b0;
      \piso.data_r_2462_sv2v_reg  <= 1'b0;
      \piso.data_r_2461_sv2v_reg  <= 1'b0;
      \piso.data_r_2460_sv2v_reg  <= 1'b0;
      \piso.data_r_2459_sv2v_reg  <= 1'b0;
      \piso.data_r_2458_sv2v_reg  <= 1'b0;
      \piso.data_r_2457_sv2v_reg  <= 1'b0;
      \piso.data_r_2456_sv2v_reg  <= 1'b0;
      \piso.data_r_2455_sv2v_reg  <= 1'b0;
      \piso.data_r_2454_sv2v_reg  <= 1'b0;
      \piso.data_r_2453_sv2v_reg  <= 1'b0;
      \piso.data_r_2452_sv2v_reg  <= 1'b0;
      \piso.data_r_2451_sv2v_reg  <= 1'b0;
      \piso.data_r_2450_sv2v_reg  <= 1'b0;
      \piso.data_r_2449_sv2v_reg  <= 1'b0;
      \piso.data_r_2448_sv2v_reg  <= 1'b0;
      \piso.data_r_2447_sv2v_reg  <= 1'b0;
      \piso.data_r_2446_sv2v_reg  <= 1'b0;
      \piso.data_r_2445_sv2v_reg  <= 1'b0;
      \piso.data_r_2444_sv2v_reg  <= 1'b0;
      \piso.data_r_2443_sv2v_reg  <= 1'b0;
      \piso.data_r_2442_sv2v_reg  <= 1'b0;
      \piso.data_r_2441_sv2v_reg  <= 1'b0;
      \piso.data_r_2440_sv2v_reg  <= 1'b0;
      \piso.data_r_2439_sv2v_reg  <= 1'b0;
      \piso.data_r_2438_sv2v_reg  <= 1'b0;
      \piso.data_r_2437_sv2v_reg  <= 1'b0;
      \piso.data_r_2436_sv2v_reg  <= 1'b0;
      \piso.data_r_2435_sv2v_reg  <= 1'b0;
      \piso.data_r_2434_sv2v_reg  <= 1'b0;
      \piso.data_r_2433_sv2v_reg  <= 1'b0;
      \piso.data_r_2432_sv2v_reg  <= 1'b0;
      \piso.data_r_2431_sv2v_reg  <= 1'b0;
      \piso.data_r_2430_sv2v_reg  <= 1'b0;
      \piso.data_r_2429_sv2v_reg  <= 1'b0;
      \piso.data_r_2428_sv2v_reg  <= 1'b0;
      \piso.data_r_2427_sv2v_reg  <= 1'b0;
      \piso.data_r_2426_sv2v_reg  <= 1'b0;
      \piso.data_r_2425_sv2v_reg  <= 1'b0;
      \piso.data_r_2424_sv2v_reg  <= 1'b0;
      \piso.data_r_2423_sv2v_reg  <= 1'b0;
      \piso.data_r_2422_sv2v_reg  <= 1'b0;
      \piso.data_r_2421_sv2v_reg  <= 1'b0;
      \piso.data_r_2420_sv2v_reg  <= 1'b0;
      \piso.data_r_2419_sv2v_reg  <= 1'b0;
      \piso.data_r_2418_sv2v_reg  <= 1'b0;
      \piso.data_r_2417_sv2v_reg  <= 1'b0;
      \piso.data_r_2416_sv2v_reg  <= 1'b0;
      \piso.data_r_2415_sv2v_reg  <= 1'b0;
      \piso.data_r_2414_sv2v_reg  <= 1'b0;
      \piso.data_r_2413_sv2v_reg  <= 1'b0;
      \piso.data_r_2412_sv2v_reg  <= 1'b0;
      \piso.data_r_2411_sv2v_reg  <= 1'b0;
      \piso.data_r_2410_sv2v_reg  <= 1'b0;
      \piso.data_r_2409_sv2v_reg  <= 1'b0;
      \piso.data_r_2408_sv2v_reg  <= 1'b0;
      \piso.data_r_2407_sv2v_reg  <= 1'b0;
      \piso.data_r_2406_sv2v_reg  <= 1'b0;
      \piso.data_r_2405_sv2v_reg  <= 1'b0;
      \piso.data_r_2404_sv2v_reg  <= 1'b0;
      \piso.data_r_2403_sv2v_reg  <= 1'b0;
      \piso.data_r_2402_sv2v_reg  <= 1'b0;
      \piso.data_r_2401_sv2v_reg  <= 1'b0;
      \piso.data_r_2400_sv2v_reg  <= 1'b0;
      \piso.data_r_2399_sv2v_reg  <= 1'b0;
      \piso.data_r_2398_sv2v_reg  <= 1'b0;
      \piso.data_r_2397_sv2v_reg  <= 1'b0;
      \piso.data_r_2396_sv2v_reg  <= 1'b0;
      \piso.data_r_2395_sv2v_reg  <= 1'b0;
      \piso.data_r_2394_sv2v_reg  <= 1'b0;
      \piso.data_r_2393_sv2v_reg  <= 1'b0;
      \piso.data_r_2392_sv2v_reg  <= 1'b0;
      \piso.data_r_2391_sv2v_reg  <= 1'b0;
      \piso.data_r_2390_sv2v_reg  <= 1'b0;
      \piso.data_r_2389_sv2v_reg  <= 1'b0;
      \piso.data_r_2388_sv2v_reg  <= 1'b0;
      \piso.data_r_2387_sv2v_reg  <= 1'b0;
      \piso.data_r_2386_sv2v_reg  <= 1'b0;
      \piso.data_r_2385_sv2v_reg  <= 1'b0;
      \piso.data_r_2384_sv2v_reg  <= 1'b0;
      \piso.data_r_2383_sv2v_reg  <= 1'b0;
      \piso.data_r_2382_sv2v_reg  <= 1'b0;
      \piso.data_r_2381_sv2v_reg  <= 1'b0;
      \piso.data_r_2380_sv2v_reg  <= 1'b0;
      \piso.data_r_2379_sv2v_reg  <= 1'b0;
      \piso.data_r_2378_sv2v_reg  <= 1'b0;
      \piso.data_r_2377_sv2v_reg  <= 1'b0;
      \piso.data_r_2376_sv2v_reg  <= 1'b0;
      \piso.data_r_2375_sv2v_reg  <= 1'b0;
      \piso.data_r_2374_sv2v_reg  <= 1'b0;
      \piso.data_r_2373_sv2v_reg  <= 1'b0;
      \piso.data_r_2372_sv2v_reg  <= 1'b0;
      \piso.data_r_2371_sv2v_reg  <= 1'b0;
      \piso.data_r_2370_sv2v_reg  <= 1'b0;
      \piso.data_r_2369_sv2v_reg  <= 1'b0;
      \piso.data_r_2368_sv2v_reg  <= 1'b0;
      \piso.data_r_2367_sv2v_reg  <= 1'b0;
      \piso.data_r_2366_sv2v_reg  <= 1'b0;
      \piso.data_r_2365_sv2v_reg  <= 1'b0;
      \piso.data_r_2364_sv2v_reg  <= 1'b0;
      \piso.data_r_2363_sv2v_reg  <= 1'b0;
      \piso.data_r_2362_sv2v_reg  <= 1'b0;
      \piso.data_r_2361_sv2v_reg  <= 1'b0;
      \piso.data_r_2360_sv2v_reg  <= 1'b0;
      \piso.data_r_2359_sv2v_reg  <= 1'b0;
      \piso.data_r_2358_sv2v_reg  <= 1'b0;
      \piso.data_r_2357_sv2v_reg  <= 1'b0;
      \piso.data_r_2356_sv2v_reg  <= 1'b0;
      \piso.data_r_2355_sv2v_reg  <= 1'b0;
      \piso.data_r_2354_sv2v_reg  <= 1'b0;
      \piso.data_r_2353_sv2v_reg  <= 1'b0;
      \piso.data_r_2352_sv2v_reg  <= 1'b0;
      \piso.data_r_2351_sv2v_reg  <= 1'b0;
      \piso.data_r_2350_sv2v_reg  <= 1'b0;
      \piso.data_r_2349_sv2v_reg  <= 1'b0;
      \piso.data_r_2348_sv2v_reg  <= 1'b0;
      \piso.data_r_2347_sv2v_reg  <= 1'b0;
      \piso.data_r_2346_sv2v_reg  <= 1'b0;
      \piso.data_r_2345_sv2v_reg  <= 1'b0;
      \piso.data_r_2344_sv2v_reg  <= 1'b0;
      \piso.data_r_2343_sv2v_reg  <= 1'b0;
      \piso.data_r_2342_sv2v_reg  <= 1'b0;
      \piso.data_r_2341_sv2v_reg  <= 1'b0;
      \piso.data_r_2340_sv2v_reg  <= 1'b0;
      \piso.data_r_2339_sv2v_reg  <= 1'b0;
      \piso.data_r_2338_sv2v_reg  <= 1'b0;
      \piso.data_r_2337_sv2v_reg  <= 1'b0;
      \piso.data_r_2336_sv2v_reg  <= 1'b0;
      \piso.data_r_2335_sv2v_reg  <= 1'b0;
      \piso.data_r_2334_sv2v_reg  <= 1'b0;
      \piso.data_r_2333_sv2v_reg  <= 1'b0;
      \piso.data_r_2332_sv2v_reg  <= 1'b0;
      \piso.data_r_2331_sv2v_reg  <= 1'b0;
      \piso.data_r_2330_sv2v_reg  <= 1'b0;
      \piso.data_r_2329_sv2v_reg  <= 1'b0;
      \piso.data_r_2328_sv2v_reg  <= 1'b0;
      \piso.data_r_2327_sv2v_reg  <= 1'b0;
      \piso.data_r_2326_sv2v_reg  <= 1'b0;
      \piso.data_r_2325_sv2v_reg  <= 1'b0;
      \piso.data_r_2324_sv2v_reg  <= 1'b0;
      \piso.data_r_2323_sv2v_reg  <= 1'b0;
      \piso.data_r_2322_sv2v_reg  <= 1'b0;
      \piso.data_r_2321_sv2v_reg  <= 1'b0;
      \piso.data_r_2320_sv2v_reg  <= 1'b0;
      \piso.data_r_2319_sv2v_reg  <= 1'b0;
      \piso.data_r_2318_sv2v_reg  <= 1'b0;
      \piso.data_r_2317_sv2v_reg  <= 1'b0;
      \piso.data_r_2316_sv2v_reg  <= 1'b0;
      \piso.data_r_2315_sv2v_reg  <= 1'b0;
      \piso.data_r_2314_sv2v_reg  <= 1'b0;
      \piso.data_r_2313_sv2v_reg  <= 1'b0;
      \piso.data_r_2312_sv2v_reg  <= 1'b0;
      \piso.data_r_2311_sv2v_reg  <= 1'b0;
      \piso.data_r_2310_sv2v_reg  <= 1'b0;
      \piso.data_r_2309_sv2v_reg  <= 1'b0;
      \piso.data_r_2308_sv2v_reg  <= 1'b0;
      \piso.data_r_2307_sv2v_reg  <= 1'b0;
      \piso.data_r_2306_sv2v_reg  <= 1'b0;
      \piso.data_r_2305_sv2v_reg  <= 1'b0;
      \piso.data_r_2304_sv2v_reg  <= 1'b0;
      \piso.data_r_2303_sv2v_reg  <= 1'b0;
      \piso.data_r_2302_sv2v_reg  <= 1'b0;
      \piso.data_r_2301_sv2v_reg  <= 1'b0;
      \piso.data_r_2300_sv2v_reg  <= 1'b0;
      \piso.data_r_2299_sv2v_reg  <= 1'b0;
      \piso.data_r_2298_sv2v_reg  <= 1'b0;
      \piso.data_r_2297_sv2v_reg  <= 1'b0;
      \piso.data_r_2296_sv2v_reg  <= 1'b0;
      \piso.data_r_2295_sv2v_reg  <= 1'b0;
      \piso.data_r_2294_sv2v_reg  <= 1'b0;
      \piso.data_r_2293_sv2v_reg  <= 1'b0;
      \piso.data_r_2292_sv2v_reg  <= 1'b0;
      \piso.data_r_2291_sv2v_reg  <= 1'b0;
      \piso.data_r_2290_sv2v_reg  <= 1'b0;
      \piso.data_r_2289_sv2v_reg  <= 1'b0;
      \piso.data_r_2288_sv2v_reg  <= 1'b0;
      \piso.data_r_2287_sv2v_reg  <= 1'b0;
      \piso.data_r_2286_sv2v_reg  <= 1'b0;
      \piso.data_r_2285_sv2v_reg  <= 1'b0;
      \piso.data_r_2284_sv2v_reg  <= 1'b0;
      \piso.data_r_2283_sv2v_reg  <= 1'b0;
      \piso.data_r_2282_sv2v_reg  <= 1'b0;
      \piso.data_r_2281_sv2v_reg  <= 1'b0;
      \piso.data_r_2280_sv2v_reg  <= 1'b0;
      \piso.data_r_2279_sv2v_reg  <= 1'b0;
      \piso.data_r_2278_sv2v_reg  <= 1'b0;
      \piso.data_r_2277_sv2v_reg  <= 1'b0;
      \piso.data_r_2276_sv2v_reg  <= 1'b0;
      \piso.data_r_2275_sv2v_reg  <= 1'b0;
      \piso.data_r_2274_sv2v_reg  <= 1'b0;
      \piso.data_r_2273_sv2v_reg  <= 1'b0;
      \piso.data_r_2272_sv2v_reg  <= 1'b0;
      \piso.data_r_2271_sv2v_reg  <= 1'b0;
      \piso.data_r_2270_sv2v_reg  <= 1'b0;
      \piso.data_r_2269_sv2v_reg  <= 1'b0;
      \piso.data_r_2268_sv2v_reg  <= 1'b0;
      \piso.data_r_2267_sv2v_reg  <= 1'b0;
      \piso.data_r_2266_sv2v_reg  <= 1'b0;
      \piso.data_r_2265_sv2v_reg  <= 1'b0;
      \piso.data_r_2264_sv2v_reg  <= 1'b0;
      \piso.data_r_2263_sv2v_reg  <= 1'b0;
      \piso.data_r_2262_sv2v_reg  <= 1'b0;
      \piso.data_r_2261_sv2v_reg  <= 1'b0;
      \piso.data_r_2260_sv2v_reg  <= 1'b0;
      \piso.data_r_2259_sv2v_reg  <= 1'b0;
      \piso.data_r_2258_sv2v_reg  <= 1'b0;
      \piso.data_r_2257_sv2v_reg  <= 1'b0;
      \piso.data_r_2256_sv2v_reg  <= 1'b0;
      \piso.data_r_2255_sv2v_reg  <= 1'b0;
      \piso.data_r_2254_sv2v_reg  <= 1'b0;
      \piso.data_r_2253_sv2v_reg  <= 1'b0;
      \piso.data_r_2252_sv2v_reg  <= 1'b0;
      \piso.data_r_2251_sv2v_reg  <= 1'b0;
      \piso.data_r_2250_sv2v_reg  <= 1'b0;
      \piso.data_r_2249_sv2v_reg  <= 1'b0;
      \piso.data_r_2248_sv2v_reg  <= 1'b0;
      \piso.data_r_2247_sv2v_reg  <= 1'b0;
      \piso.data_r_2246_sv2v_reg  <= 1'b0;
      \piso.data_r_2245_sv2v_reg  <= 1'b0;
      \piso.data_r_2244_sv2v_reg  <= 1'b0;
      \piso.data_r_2243_sv2v_reg  <= 1'b0;
      \piso.data_r_2242_sv2v_reg  <= 1'b0;
      \piso.data_r_2241_sv2v_reg  <= 1'b0;
      \piso.data_r_2240_sv2v_reg  <= 1'b0;
      \piso.data_r_2239_sv2v_reg  <= 1'b0;
      \piso.data_r_2238_sv2v_reg  <= 1'b0;
      \piso.data_r_2237_sv2v_reg  <= 1'b0;
      \piso.data_r_2236_sv2v_reg  <= 1'b0;
      \piso.data_r_2235_sv2v_reg  <= 1'b0;
      \piso.data_r_2234_sv2v_reg  <= 1'b0;
      \piso.data_r_2233_sv2v_reg  <= 1'b0;
      \piso.data_r_2232_sv2v_reg  <= 1'b0;
      \piso.data_r_2231_sv2v_reg  <= 1'b0;
      \piso.data_r_2230_sv2v_reg  <= 1'b0;
      \piso.data_r_2229_sv2v_reg  <= 1'b0;
      \piso.data_r_2228_sv2v_reg  <= 1'b0;
      \piso.data_r_2227_sv2v_reg  <= 1'b0;
      \piso.data_r_2226_sv2v_reg  <= 1'b0;
      \piso.data_r_2225_sv2v_reg  <= 1'b0;
      \piso.data_r_2224_sv2v_reg  <= 1'b0;
      \piso.data_r_2223_sv2v_reg  <= 1'b0;
      \piso.data_r_2222_sv2v_reg  <= 1'b0;
      \piso.data_r_2221_sv2v_reg  <= 1'b0;
      \piso.data_r_2220_sv2v_reg  <= 1'b0;
      \piso.data_r_2219_sv2v_reg  <= 1'b0;
      \piso.data_r_2218_sv2v_reg  <= 1'b0;
      \piso.data_r_2217_sv2v_reg  <= 1'b0;
      \piso.data_r_2216_sv2v_reg  <= 1'b0;
      \piso.data_r_2215_sv2v_reg  <= 1'b0;
      \piso.data_r_2214_sv2v_reg  <= 1'b0;
      \piso.data_r_2213_sv2v_reg  <= 1'b0;
      \piso.data_r_2212_sv2v_reg  <= 1'b0;
      \piso.data_r_2211_sv2v_reg  <= 1'b0;
      \piso.data_r_2210_sv2v_reg  <= 1'b0;
      \piso.data_r_2209_sv2v_reg  <= 1'b0;
      \piso.data_r_2208_sv2v_reg  <= 1'b0;
      \piso.data_r_2207_sv2v_reg  <= 1'b0;
      \piso.data_r_2206_sv2v_reg  <= 1'b0;
      \piso.data_r_2205_sv2v_reg  <= 1'b0;
      \piso.data_r_2204_sv2v_reg  <= 1'b0;
      \piso.data_r_2203_sv2v_reg  <= 1'b0;
      \piso.data_r_2202_sv2v_reg  <= 1'b0;
      \piso.data_r_2201_sv2v_reg  <= 1'b0;
      \piso.data_r_2200_sv2v_reg  <= 1'b0;
      \piso.data_r_2199_sv2v_reg  <= 1'b0;
      \piso.data_r_2198_sv2v_reg  <= 1'b0;
      \piso.data_r_2197_sv2v_reg  <= 1'b0;
      \piso.data_r_2196_sv2v_reg  <= 1'b0;
      \piso.data_r_2195_sv2v_reg  <= 1'b0;
      \piso.data_r_2194_sv2v_reg  <= 1'b0;
      \piso.data_r_2193_sv2v_reg  <= 1'b0;
      \piso.data_r_2192_sv2v_reg  <= 1'b0;
      \piso.data_r_2191_sv2v_reg  <= 1'b0;
      \piso.data_r_2190_sv2v_reg  <= 1'b0;
      \piso.data_r_2189_sv2v_reg  <= 1'b0;
      \piso.data_r_2188_sv2v_reg  <= 1'b0;
      \piso.data_r_2187_sv2v_reg  <= 1'b0;
      \piso.data_r_2186_sv2v_reg  <= 1'b0;
      \piso.data_r_2185_sv2v_reg  <= 1'b0;
      \piso.data_r_2184_sv2v_reg  <= 1'b0;
      \piso.data_r_2183_sv2v_reg  <= 1'b0;
      \piso.data_r_2182_sv2v_reg  <= 1'b0;
      \piso.data_r_2181_sv2v_reg  <= 1'b0;
      \piso.data_r_2180_sv2v_reg  <= 1'b0;
      \piso.data_r_2179_sv2v_reg  <= 1'b0;
      \piso.data_r_2178_sv2v_reg  <= 1'b0;
      \piso.data_r_2177_sv2v_reg  <= 1'b0;
      \piso.data_r_2176_sv2v_reg  <= 1'b0;
      \piso.data_r_2175_sv2v_reg  <= 1'b0;
      \piso.data_r_2174_sv2v_reg  <= 1'b0;
      \piso.data_r_2173_sv2v_reg  <= 1'b0;
      \piso.data_r_2172_sv2v_reg  <= 1'b0;
      \piso.data_r_2171_sv2v_reg  <= 1'b0;
      \piso.data_r_2170_sv2v_reg  <= 1'b0;
      \piso.data_r_2169_sv2v_reg  <= 1'b0;
      \piso.data_r_2168_sv2v_reg  <= 1'b0;
      \piso.data_r_2167_sv2v_reg  <= 1'b0;
      \piso.data_r_2166_sv2v_reg  <= 1'b0;
      \piso.data_r_2165_sv2v_reg  <= 1'b0;
      \piso.data_r_2164_sv2v_reg  <= 1'b0;
      \piso.data_r_2163_sv2v_reg  <= 1'b0;
      \piso.data_r_2162_sv2v_reg  <= 1'b0;
      \piso.data_r_2161_sv2v_reg  <= 1'b0;
      \piso.data_r_2160_sv2v_reg  <= 1'b0;
      \piso.data_r_2159_sv2v_reg  <= 1'b0;
      \piso.data_r_2158_sv2v_reg  <= 1'b0;
      \piso.data_r_2157_sv2v_reg  <= 1'b0;
      \piso.data_r_2156_sv2v_reg  <= 1'b0;
      \piso.data_r_2155_sv2v_reg  <= 1'b0;
      \piso.data_r_2154_sv2v_reg  <= 1'b0;
      \piso.data_r_2153_sv2v_reg  <= 1'b0;
      \piso.data_r_2152_sv2v_reg  <= 1'b0;
      \piso.data_r_2151_sv2v_reg  <= 1'b0;
      \piso.data_r_2150_sv2v_reg  <= 1'b0;
      \piso.data_r_2149_sv2v_reg  <= 1'b0;
      \piso.data_r_2148_sv2v_reg  <= 1'b0;
      \piso.data_r_2147_sv2v_reg  <= 1'b0;
      \piso.data_r_2146_sv2v_reg  <= 1'b0;
      \piso.data_r_2145_sv2v_reg  <= 1'b0;
      \piso.data_r_2144_sv2v_reg  <= 1'b0;
      \piso.data_r_2143_sv2v_reg  <= 1'b0;
      \piso.data_r_2142_sv2v_reg  <= 1'b0;
      \piso.data_r_2141_sv2v_reg  <= 1'b0;
      \piso.data_r_2140_sv2v_reg  <= 1'b0;
      \piso.data_r_2139_sv2v_reg  <= 1'b0;
      \piso.data_r_2138_sv2v_reg  <= 1'b0;
      \piso.data_r_2137_sv2v_reg  <= 1'b0;
      \piso.data_r_2136_sv2v_reg  <= 1'b0;
      \piso.data_r_2135_sv2v_reg  <= 1'b0;
      \piso.data_r_2134_sv2v_reg  <= 1'b0;
      \piso.data_r_2133_sv2v_reg  <= 1'b0;
      \piso.data_r_2132_sv2v_reg  <= 1'b0;
      \piso.data_r_2131_sv2v_reg  <= 1'b0;
      \piso.data_r_2130_sv2v_reg  <= 1'b0;
      \piso.data_r_2129_sv2v_reg  <= 1'b0;
      \piso.data_r_2128_sv2v_reg  <= 1'b0;
      \piso.data_r_2127_sv2v_reg  <= 1'b0;
      \piso.data_r_2126_sv2v_reg  <= 1'b0;
      \piso.data_r_2125_sv2v_reg  <= 1'b0;
      \piso.data_r_2124_sv2v_reg  <= 1'b0;
      \piso.data_r_2123_sv2v_reg  <= 1'b0;
      \piso.data_r_2122_sv2v_reg  <= 1'b0;
      \piso.data_r_2121_sv2v_reg  <= 1'b0;
      \piso.data_r_2120_sv2v_reg  <= 1'b0;
      \piso.data_r_2119_sv2v_reg  <= 1'b0;
      \piso.data_r_2118_sv2v_reg  <= 1'b0;
      \piso.data_r_2117_sv2v_reg  <= 1'b0;
      \piso.data_r_2116_sv2v_reg  <= 1'b0;
      \piso.data_r_2115_sv2v_reg  <= 1'b0;
      \piso.data_r_2114_sv2v_reg  <= 1'b0;
      \piso.data_r_2113_sv2v_reg  <= 1'b0;
      \piso.data_r_2112_sv2v_reg  <= 1'b0;
      \piso.data_r_2111_sv2v_reg  <= 1'b0;
      \piso.data_r_2110_sv2v_reg  <= 1'b0;
      \piso.data_r_2109_sv2v_reg  <= 1'b0;
      \piso.data_r_2108_sv2v_reg  <= 1'b0;
      \piso.data_r_2107_sv2v_reg  <= 1'b0;
      \piso.data_r_2106_sv2v_reg  <= 1'b0;
      \piso.data_r_2105_sv2v_reg  <= 1'b0;
      \piso.data_r_2104_sv2v_reg  <= 1'b0;
      \piso.data_r_2103_sv2v_reg  <= 1'b0;
      \piso.data_r_2102_sv2v_reg  <= 1'b0;
      \piso.data_r_2101_sv2v_reg  <= 1'b0;
      \piso.data_r_2100_sv2v_reg  <= 1'b0;
      \piso.data_r_2099_sv2v_reg  <= 1'b0;
      \piso.data_r_2098_sv2v_reg  <= 1'b0;
      \piso.data_r_2097_sv2v_reg  <= 1'b0;
      \piso.data_r_2096_sv2v_reg  <= 1'b0;
      \piso.data_r_2095_sv2v_reg  <= 1'b0;
      \piso.data_r_2094_sv2v_reg  <= 1'b0;
      \piso.data_r_2093_sv2v_reg  <= 1'b0;
      \piso.data_r_2092_sv2v_reg  <= 1'b0;
      \piso.data_r_2091_sv2v_reg  <= 1'b0;
      \piso.data_r_2090_sv2v_reg  <= 1'b0;
      \piso.data_r_2089_sv2v_reg  <= 1'b0;
      \piso.data_r_2088_sv2v_reg  <= 1'b0;
      \piso.data_r_2087_sv2v_reg  <= 1'b0;
      \piso.data_r_2086_sv2v_reg  <= 1'b0;
      \piso.data_r_2085_sv2v_reg  <= 1'b0;
      \piso.data_r_2084_sv2v_reg  <= 1'b0;
      \piso.data_r_2083_sv2v_reg  <= 1'b0;
      \piso.data_r_2082_sv2v_reg  <= 1'b0;
      \piso.data_r_2081_sv2v_reg  <= 1'b0;
      \piso.data_r_2080_sv2v_reg  <= 1'b0;
      \piso.data_r_2079_sv2v_reg  <= 1'b0;
      \piso.data_r_2078_sv2v_reg  <= 1'b0;
      \piso.data_r_2077_sv2v_reg  <= 1'b0;
      \piso.data_r_2076_sv2v_reg  <= 1'b0;
      \piso.data_r_2075_sv2v_reg  <= 1'b0;
      \piso.data_r_2074_sv2v_reg  <= 1'b0;
      \piso.data_r_2073_sv2v_reg  <= 1'b0;
      \piso.data_r_2072_sv2v_reg  <= 1'b0;
      \piso.data_r_2071_sv2v_reg  <= 1'b0;
      \piso.data_r_2070_sv2v_reg  <= 1'b0;
      \piso.data_r_2069_sv2v_reg  <= 1'b0;
      \piso.data_r_2068_sv2v_reg  <= 1'b0;
      \piso.data_r_2067_sv2v_reg  <= 1'b0;
      \piso.data_r_2066_sv2v_reg  <= 1'b0;
      \piso.data_r_2065_sv2v_reg  <= 1'b0;
      \piso.data_r_2064_sv2v_reg  <= 1'b0;
      \piso.data_r_2063_sv2v_reg  <= 1'b0;
      \piso.data_r_2062_sv2v_reg  <= 1'b0;
      \piso.data_r_2061_sv2v_reg  <= 1'b0;
      \piso.data_r_2060_sv2v_reg  <= 1'b0;
      \piso.data_r_2059_sv2v_reg  <= 1'b0;
      \piso.data_r_2058_sv2v_reg  <= 1'b0;
      \piso.data_r_2057_sv2v_reg  <= 1'b0;
      \piso.data_r_2056_sv2v_reg  <= 1'b0;
      \piso.data_r_2055_sv2v_reg  <= 1'b0;
      \piso.data_r_2054_sv2v_reg  <= 1'b0;
      \piso.data_r_2053_sv2v_reg  <= 1'b0;
      \piso.data_r_2052_sv2v_reg  <= 1'b0;
      \piso.data_r_2051_sv2v_reg  <= 1'b0;
      \piso.data_r_2050_sv2v_reg  <= 1'b0;
      \piso.data_r_2049_sv2v_reg  <= 1'b0;
      \piso.data_r_2048_sv2v_reg  <= 1'b0;
      \piso.data_r_2047_sv2v_reg  <= 1'b0;
      \piso.data_r_2046_sv2v_reg  <= 1'b0;
      \piso.data_r_2045_sv2v_reg  <= 1'b0;
      \piso.data_r_2044_sv2v_reg  <= 1'b0;
      \piso.data_r_2043_sv2v_reg  <= 1'b0;
      \piso.data_r_2042_sv2v_reg  <= 1'b0;
      \piso.data_r_2041_sv2v_reg  <= 1'b0;
      \piso.data_r_2040_sv2v_reg  <= 1'b0;
      \piso.data_r_2039_sv2v_reg  <= 1'b0;
      \piso.data_r_2038_sv2v_reg  <= 1'b0;
      \piso.data_r_2037_sv2v_reg  <= 1'b0;
      \piso.data_r_2036_sv2v_reg  <= 1'b0;
      \piso.data_r_2035_sv2v_reg  <= 1'b0;
      \piso.data_r_2034_sv2v_reg  <= 1'b0;
      \piso.data_r_2033_sv2v_reg  <= 1'b0;
      \piso.data_r_2032_sv2v_reg  <= 1'b0;
      \piso.data_r_2031_sv2v_reg  <= 1'b0;
      \piso.data_r_2030_sv2v_reg  <= 1'b0;
      \piso.data_r_2029_sv2v_reg  <= 1'b0;
      \piso.data_r_2028_sv2v_reg  <= 1'b0;
      \piso.data_r_2027_sv2v_reg  <= 1'b0;
      \piso.data_r_2026_sv2v_reg  <= 1'b0;
      \piso.data_r_2025_sv2v_reg  <= 1'b0;
      \piso.data_r_2024_sv2v_reg  <= 1'b0;
      \piso.data_r_2023_sv2v_reg  <= 1'b0;
      \piso.data_r_2022_sv2v_reg  <= 1'b0;
      \piso.data_r_2021_sv2v_reg  <= 1'b0;
      \piso.data_r_2020_sv2v_reg  <= 1'b0;
      \piso.data_r_2019_sv2v_reg  <= 1'b0;
      \piso.data_r_2018_sv2v_reg  <= 1'b0;
      \piso.data_r_2017_sv2v_reg  <= 1'b0;
      \piso.data_r_2016_sv2v_reg  <= 1'b0;
      \piso.data_r_2015_sv2v_reg  <= 1'b0;
      \piso.data_r_2014_sv2v_reg  <= 1'b0;
      \piso.data_r_2013_sv2v_reg  <= 1'b0;
      \piso.data_r_2012_sv2v_reg  <= 1'b0;
      \piso.data_r_2011_sv2v_reg  <= 1'b0;
      \piso.data_r_2010_sv2v_reg  <= 1'b0;
      \piso.data_r_2009_sv2v_reg  <= 1'b0;
      \piso.data_r_2008_sv2v_reg  <= 1'b0;
      \piso.data_r_2007_sv2v_reg  <= 1'b0;
      \piso.data_r_2006_sv2v_reg  <= 1'b0;
      \piso.data_r_2005_sv2v_reg  <= 1'b0;
      \piso.data_r_2004_sv2v_reg  <= 1'b0;
      \piso.data_r_2003_sv2v_reg  <= 1'b0;
      \piso.data_r_2002_sv2v_reg  <= 1'b0;
      \piso.data_r_2001_sv2v_reg  <= 1'b0;
      \piso.data_r_2000_sv2v_reg  <= 1'b0;
      \piso.data_r_1999_sv2v_reg  <= 1'b0;
      \piso.data_r_1998_sv2v_reg  <= 1'b0;
      \piso.data_r_1997_sv2v_reg  <= 1'b0;
      \piso.data_r_1996_sv2v_reg  <= 1'b0;
      \piso.data_r_1995_sv2v_reg  <= 1'b0;
      \piso.data_r_1994_sv2v_reg  <= 1'b0;
      \piso.data_r_1993_sv2v_reg  <= 1'b0;
      \piso.data_r_1992_sv2v_reg  <= 1'b0;
      \piso.data_r_1991_sv2v_reg  <= 1'b0;
      \piso.data_r_1990_sv2v_reg  <= 1'b0;
      \piso.data_r_1989_sv2v_reg  <= 1'b0;
      \piso.data_r_1988_sv2v_reg  <= 1'b0;
      \piso.data_r_1987_sv2v_reg  <= 1'b0;
      \piso.data_r_1986_sv2v_reg  <= 1'b0;
      \piso.data_r_1985_sv2v_reg  <= 1'b0;
      \piso.data_r_1984_sv2v_reg  <= 1'b0;
      \piso.data_r_1983_sv2v_reg  <= 1'b0;
      \piso.data_r_1982_sv2v_reg  <= 1'b0;
      \piso.data_r_1981_sv2v_reg  <= 1'b0;
      \piso.data_r_1980_sv2v_reg  <= 1'b0;
      \piso.data_r_1979_sv2v_reg  <= 1'b0;
      \piso.data_r_1978_sv2v_reg  <= 1'b0;
      \piso.data_r_1977_sv2v_reg  <= 1'b0;
      \piso.data_r_1976_sv2v_reg  <= 1'b0;
      \piso.data_r_1975_sv2v_reg  <= 1'b0;
      \piso.data_r_1974_sv2v_reg  <= 1'b0;
      \piso.data_r_1973_sv2v_reg  <= 1'b0;
      \piso.data_r_1972_sv2v_reg  <= 1'b0;
      \piso.data_r_1971_sv2v_reg  <= 1'b0;
      \piso.data_r_1970_sv2v_reg  <= 1'b0;
      \piso.data_r_1969_sv2v_reg  <= 1'b0;
      \piso.data_r_1968_sv2v_reg  <= 1'b0;
      \piso.data_r_1967_sv2v_reg  <= 1'b0;
      \piso.data_r_1966_sv2v_reg  <= 1'b0;
      \piso.data_r_1965_sv2v_reg  <= 1'b0;
      \piso.data_r_1964_sv2v_reg  <= 1'b0;
      \piso.data_r_1963_sv2v_reg  <= 1'b0;
      \piso.data_r_1962_sv2v_reg  <= 1'b0;
      \piso.data_r_1961_sv2v_reg  <= 1'b0;
      \piso.data_r_1960_sv2v_reg  <= 1'b0;
      \piso.data_r_1959_sv2v_reg  <= 1'b0;
      \piso.data_r_1958_sv2v_reg  <= 1'b0;
      \piso.data_r_1957_sv2v_reg  <= 1'b0;
      \piso.data_r_1956_sv2v_reg  <= 1'b0;
      \piso.data_r_1955_sv2v_reg  <= 1'b0;
      \piso.data_r_1954_sv2v_reg  <= 1'b0;
      \piso.data_r_1953_sv2v_reg  <= 1'b0;
      \piso.data_r_1952_sv2v_reg  <= 1'b0;
      \piso.data_r_1951_sv2v_reg  <= 1'b0;
      \piso.data_r_1950_sv2v_reg  <= 1'b0;
      \piso.data_r_1949_sv2v_reg  <= 1'b0;
      \piso.data_r_1948_sv2v_reg  <= 1'b0;
      \piso.data_r_1947_sv2v_reg  <= 1'b0;
      \piso.data_r_1946_sv2v_reg  <= 1'b0;
      \piso.data_r_1945_sv2v_reg  <= 1'b0;
      \piso.data_r_1944_sv2v_reg  <= 1'b0;
      \piso.data_r_1943_sv2v_reg  <= 1'b0;
      \piso.data_r_1942_sv2v_reg  <= 1'b0;
      \piso.data_r_1941_sv2v_reg  <= 1'b0;
      \piso.data_r_1940_sv2v_reg  <= 1'b0;
      \piso.data_r_1939_sv2v_reg  <= 1'b0;
      \piso.data_r_1938_sv2v_reg  <= 1'b0;
      \piso.data_r_1937_sv2v_reg  <= 1'b0;
      \piso.data_r_1936_sv2v_reg  <= 1'b0;
      \piso.data_r_1935_sv2v_reg  <= 1'b0;
      \piso.data_r_1934_sv2v_reg  <= 1'b0;
      \piso.data_r_1933_sv2v_reg  <= 1'b0;
      \piso.data_r_1932_sv2v_reg  <= 1'b0;
      \piso.data_r_1931_sv2v_reg  <= 1'b0;
      \piso.data_r_1930_sv2v_reg  <= 1'b0;
      \piso.data_r_1929_sv2v_reg  <= 1'b0;
      \piso.data_r_1928_sv2v_reg  <= 1'b0;
      \piso.data_r_1927_sv2v_reg  <= 1'b0;
      \piso.data_r_1926_sv2v_reg  <= 1'b0;
      \piso.data_r_1925_sv2v_reg  <= 1'b0;
      \piso.data_r_1924_sv2v_reg  <= 1'b0;
      \piso.data_r_1923_sv2v_reg  <= 1'b0;
      \piso.data_r_1922_sv2v_reg  <= 1'b0;
      \piso.data_r_1921_sv2v_reg  <= 1'b0;
      \piso.data_r_1920_sv2v_reg  <= 1'b0;
      \piso.data_r_1919_sv2v_reg  <= 1'b0;
      \piso.data_r_1918_sv2v_reg  <= 1'b0;
      \piso.data_r_1917_sv2v_reg  <= 1'b0;
      \piso.data_r_1916_sv2v_reg  <= 1'b0;
      \piso.data_r_1915_sv2v_reg  <= 1'b0;
      \piso.data_r_1914_sv2v_reg  <= 1'b0;
      \piso.data_r_1913_sv2v_reg  <= 1'b0;
      \piso.data_r_1912_sv2v_reg  <= 1'b0;
      \piso.data_r_1911_sv2v_reg  <= 1'b0;
      \piso.data_r_1910_sv2v_reg  <= 1'b0;
      \piso.data_r_1909_sv2v_reg  <= 1'b0;
      \piso.data_r_1908_sv2v_reg  <= 1'b0;
      \piso.data_r_1907_sv2v_reg  <= 1'b0;
      \piso.data_r_1906_sv2v_reg  <= 1'b0;
      \piso.data_r_1905_sv2v_reg  <= 1'b0;
      \piso.data_r_1904_sv2v_reg  <= 1'b0;
      \piso.data_r_1903_sv2v_reg  <= 1'b0;
      \piso.data_r_1902_sv2v_reg  <= 1'b0;
      \piso.data_r_1901_sv2v_reg  <= 1'b0;
      \piso.data_r_1900_sv2v_reg  <= 1'b0;
      \piso.data_r_1899_sv2v_reg  <= 1'b0;
      \piso.data_r_1898_sv2v_reg  <= 1'b0;
      \piso.data_r_1897_sv2v_reg  <= 1'b0;
      \piso.data_r_1896_sv2v_reg  <= 1'b0;
      \piso.data_r_1895_sv2v_reg  <= 1'b0;
      \piso.data_r_1894_sv2v_reg  <= 1'b0;
      \piso.data_r_1893_sv2v_reg  <= 1'b0;
      \piso.data_r_1892_sv2v_reg  <= 1'b0;
      \piso.data_r_1891_sv2v_reg  <= 1'b0;
      \piso.data_r_1890_sv2v_reg  <= 1'b0;
      \piso.data_r_1889_sv2v_reg  <= 1'b0;
      \piso.data_r_1888_sv2v_reg  <= 1'b0;
      \piso.data_r_1887_sv2v_reg  <= 1'b0;
      \piso.data_r_1886_sv2v_reg  <= 1'b0;
      \piso.data_r_1885_sv2v_reg  <= 1'b0;
      \piso.data_r_1884_sv2v_reg  <= 1'b0;
      \piso.data_r_1883_sv2v_reg  <= 1'b0;
      \piso.data_r_1882_sv2v_reg  <= 1'b0;
      \piso.data_r_1881_sv2v_reg  <= 1'b0;
      \piso.data_r_1880_sv2v_reg  <= 1'b0;
      \piso.data_r_1879_sv2v_reg  <= 1'b0;
      \piso.data_r_1878_sv2v_reg  <= 1'b0;
      \piso.data_r_1877_sv2v_reg  <= 1'b0;
      \piso.data_r_1876_sv2v_reg  <= 1'b0;
      \piso.data_r_1875_sv2v_reg  <= 1'b0;
      \piso.data_r_1874_sv2v_reg  <= 1'b0;
      \piso.data_r_1873_sv2v_reg  <= 1'b0;
      \piso.data_r_1872_sv2v_reg  <= 1'b0;
      \piso.data_r_1871_sv2v_reg  <= 1'b0;
      \piso.data_r_1870_sv2v_reg  <= 1'b0;
      \piso.data_r_1869_sv2v_reg  <= 1'b0;
      \piso.data_r_1868_sv2v_reg  <= 1'b0;
      \piso.data_r_1867_sv2v_reg  <= 1'b0;
      \piso.data_r_1866_sv2v_reg  <= 1'b0;
      \piso.data_r_1865_sv2v_reg  <= 1'b0;
      \piso.data_r_1864_sv2v_reg  <= 1'b0;
      \piso.data_r_1863_sv2v_reg  <= 1'b0;
      \piso.data_r_1862_sv2v_reg  <= 1'b0;
      \piso.data_r_1861_sv2v_reg  <= 1'b0;
      \piso.data_r_1860_sv2v_reg  <= 1'b0;
      \piso.data_r_1859_sv2v_reg  <= 1'b0;
      \piso.data_r_1858_sv2v_reg  <= 1'b0;
      \piso.data_r_1857_sv2v_reg  <= 1'b0;
      \piso.data_r_1856_sv2v_reg  <= 1'b0;
      \piso.data_r_1855_sv2v_reg  <= 1'b0;
      \piso.data_r_1854_sv2v_reg  <= 1'b0;
      \piso.data_r_1853_sv2v_reg  <= 1'b0;
      \piso.data_r_1852_sv2v_reg  <= 1'b0;
      \piso.data_r_1851_sv2v_reg  <= 1'b0;
      \piso.data_r_1850_sv2v_reg  <= 1'b0;
      \piso.data_r_1849_sv2v_reg  <= 1'b0;
      \piso.data_r_1848_sv2v_reg  <= 1'b0;
      \piso.data_r_1847_sv2v_reg  <= 1'b0;
      \piso.data_r_1846_sv2v_reg  <= 1'b0;
      \piso.data_r_1845_sv2v_reg  <= 1'b0;
      \piso.data_r_1844_sv2v_reg  <= 1'b0;
      \piso.data_r_1843_sv2v_reg  <= 1'b0;
      \piso.data_r_1842_sv2v_reg  <= 1'b0;
      \piso.data_r_1841_sv2v_reg  <= 1'b0;
      \piso.data_r_1840_sv2v_reg  <= 1'b0;
      \piso.data_r_1839_sv2v_reg  <= 1'b0;
      \piso.data_r_1838_sv2v_reg  <= 1'b0;
      \piso.data_r_1837_sv2v_reg  <= 1'b0;
      \piso.data_r_1836_sv2v_reg  <= 1'b0;
      \piso.data_r_1835_sv2v_reg  <= 1'b0;
      \piso.data_r_1834_sv2v_reg  <= 1'b0;
      \piso.data_r_1833_sv2v_reg  <= 1'b0;
      \piso.data_r_1832_sv2v_reg  <= 1'b0;
      \piso.data_r_1831_sv2v_reg  <= 1'b0;
      \piso.data_r_1830_sv2v_reg  <= 1'b0;
      \piso.data_r_1829_sv2v_reg  <= 1'b0;
      \piso.data_r_1828_sv2v_reg  <= 1'b0;
      \piso.data_r_1827_sv2v_reg  <= 1'b0;
      \piso.data_r_1826_sv2v_reg  <= 1'b0;
      \piso.data_r_1825_sv2v_reg  <= 1'b0;
      \piso.data_r_1824_sv2v_reg  <= 1'b0;
      \piso.data_r_1823_sv2v_reg  <= 1'b0;
      \piso.data_r_1822_sv2v_reg  <= 1'b0;
      \piso.data_r_1821_sv2v_reg  <= 1'b0;
      \piso.data_r_1820_sv2v_reg  <= 1'b0;
      \piso.data_r_1819_sv2v_reg  <= 1'b0;
      \piso.data_r_1818_sv2v_reg  <= 1'b0;
      \piso.data_r_1817_sv2v_reg  <= 1'b0;
      \piso.data_r_1816_sv2v_reg  <= 1'b0;
      \piso.data_r_1815_sv2v_reg  <= 1'b0;
      \piso.data_r_1814_sv2v_reg  <= 1'b0;
      \piso.data_r_1813_sv2v_reg  <= 1'b0;
      \piso.data_r_1812_sv2v_reg  <= 1'b0;
      \piso.data_r_1811_sv2v_reg  <= 1'b0;
      \piso.data_r_1810_sv2v_reg  <= 1'b0;
      \piso.data_r_1809_sv2v_reg  <= 1'b0;
      \piso.data_r_1808_sv2v_reg  <= 1'b0;
      \piso.data_r_1807_sv2v_reg  <= 1'b0;
      \piso.data_r_1806_sv2v_reg  <= 1'b0;
      \piso.data_r_1805_sv2v_reg  <= 1'b0;
      \piso.data_r_1804_sv2v_reg  <= 1'b0;
      \piso.data_r_1803_sv2v_reg  <= 1'b0;
      \piso.data_r_1802_sv2v_reg  <= 1'b0;
      \piso.data_r_1801_sv2v_reg  <= 1'b0;
      \piso.data_r_1800_sv2v_reg  <= 1'b0;
      \piso.data_r_1799_sv2v_reg  <= 1'b0;
      \piso.data_r_1798_sv2v_reg  <= 1'b0;
      \piso.data_r_1797_sv2v_reg  <= 1'b0;
      \piso.data_r_1796_sv2v_reg  <= 1'b0;
      \piso.data_r_1795_sv2v_reg  <= 1'b0;
      \piso.data_r_1794_sv2v_reg  <= 1'b0;
      \piso.data_r_1793_sv2v_reg  <= 1'b0;
      \piso.data_r_1792_sv2v_reg  <= 1'b0;
      \piso.data_r_1791_sv2v_reg  <= 1'b0;
      \piso.data_r_1790_sv2v_reg  <= 1'b0;
      \piso.data_r_1789_sv2v_reg  <= 1'b0;
      \piso.data_r_1788_sv2v_reg  <= 1'b0;
      \piso.data_r_1787_sv2v_reg  <= 1'b0;
      \piso.data_r_1786_sv2v_reg  <= 1'b0;
      \piso.data_r_1785_sv2v_reg  <= 1'b0;
      \piso.data_r_1784_sv2v_reg  <= 1'b0;
      \piso.data_r_1783_sv2v_reg  <= 1'b0;
      \piso.data_r_1782_sv2v_reg  <= 1'b0;
      \piso.data_r_1781_sv2v_reg  <= 1'b0;
      \piso.data_r_1780_sv2v_reg  <= 1'b0;
      \piso.data_r_1779_sv2v_reg  <= 1'b0;
      \piso.data_r_1778_sv2v_reg  <= 1'b0;
      \piso.data_r_1777_sv2v_reg  <= 1'b0;
      \piso.data_r_1776_sv2v_reg  <= 1'b0;
      \piso.data_r_1775_sv2v_reg  <= 1'b0;
      \piso.data_r_1774_sv2v_reg  <= 1'b0;
      \piso.data_r_1773_sv2v_reg  <= 1'b0;
      \piso.data_r_1772_sv2v_reg  <= 1'b0;
      \piso.data_r_1771_sv2v_reg  <= 1'b0;
      \piso.data_r_1770_sv2v_reg  <= 1'b0;
      \piso.data_r_1769_sv2v_reg  <= 1'b0;
      \piso.data_r_1768_sv2v_reg  <= 1'b0;
      \piso.data_r_1767_sv2v_reg  <= 1'b0;
      \piso.data_r_1766_sv2v_reg  <= 1'b0;
      \piso.data_r_1765_sv2v_reg  <= 1'b0;
      \piso.data_r_1764_sv2v_reg  <= 1'b0;
      \piso.data_r_1763_sv2v_reg  <= 1'b0;
      \piso.data_r_1762_sv2v_reg  <= 1'b0;
      \piso.data_r_1761_sv2v_reg  <= 1'b0;
      \piso.data_r_1760_sv2v_reg  <= 1'b0;
      \piso.data_r_1759_sv2v_reg  <= 1'b0;
      \piso.data_r_1758_sv2v_reg  <= 1'b0;
      \piso.data_r_1757_sv2v_reg  <= 1'b0;
      \piso.data_r_1756_sv2v_reg  <= 1'b0;
      \piso.data_r_1755_sv2v_reg  <= 1'b0;
      \piso.data_r_1754_sv2v_reg  <= 1'b0;
      \piso.data_r_1753_sv2v_reg  <= 1'b0;
      \piso.data_r_1752_sv2v_reg  <= 1'b0;
      \piso.data_r_1751_sv2v_reg  <= 1'b0;
      \piso.data_r_1750_sv2v_reg  <= 1'b0;
      \piso.data_r_1749_sv2v_reg  <= 1'b0;
      \piso.data_r_1748_sv2v_reg  <= 1'b0;
      \piso.data_r_1747_sv2v_reg  <= 1'b0;
      \piso.data_r_1746_sv2v_reg  <= 1'b0;
      \piso.data_r_1745_sv2v_reg  <= 1'b0;
      \piso.data_r_1744_sv2v_reg  <= 1'b0;
      \piso.data_r_1743_sv2v_reg  <= 1'b0;
      \piso.data_r_1742_sv2v_reg  <= 1'b0;
      \piso.data_r_1741_sv2v_reg  <= 1'b0;
      \piso.data_r_1740_sv2v_reg  <= 1'b0;
      \piso.data_r_1739_sv2v_reg  <= 1'b0;
      \piso.data_r_1738_sv2v_reg  <= 1'b0;
      \piso.data_r_1737_sv2v_reg  <= 1'b0;
      \piso.data_r_1736_sv2v_reg  <= 1'b0;
      \piso.data_r_1735_sv2v_reg  <= 1'b0;
      \piso.data_r_1734_sv2v_reg  <= 1'b0;
      \piso.data_r_1733_sv2v_reg  <= 1'b0;
      \piso.data_r_1732_sv2v_reg  <= 1'b0;
      \piso.data_r_1731_sv2v_reg  <= 1'b0;
      \piso.data_r_1730_sv2v_reg  <= 1'b0;
      \piso.data_r_1729_sv2v_reg  <= 1'b0;
      \piso.data_r_1728_sv2v_reg  <= 1'b0;
      \piso.data_r_1727_sv2v_reg  <= 1'b0;
      \piso.data_r_1726_sv2v_reg  <= 1'b0;
      \piso.data_r_1725_sv2v_reg  <= 1'b0;
      \piso.data_r_1724_sv2v_reg  <= 1'b0;
      \piso.data_r_1723_sv2v_reg  <= 1'b0;
      \piso.data_r_1722_sv2v_reg  <= 1'b0;
      \piso.data_r_1721_sv2v_reg  <= 1'b0;
      \piso.data_r_1720_sv2v_reg  <= 1'b0;
      \piso.data_r_1719_sv2v_reg  <= 1'b0;
      \piso.data_r_1718_sv2v_reg  <= 1'b0;
      \piso.data_r_1717_sv2v_reg  <= 1'b0;
      \piso.data_r_1716_sv2v_reg  <= 1'b0;
      \piso.data_r_1715_sv2v_reg  <= 1'b0;
      \piso.data_r_1714_sv2v_reg  <= 1'b0;
      \piso.data_r_1713_sv2v_reg  <= 1'b0;
      \piso.data_r_1712_sv2v_reg  <= 1'b0;
      \piso.data_r_1711_sv2v_reg  <= 1'b0;
      \piso.data_r_1710_sv2v_reg  <= 1'b0;
      \piso.data_r_1709_sv2v_reg  <= 1'b0;
      \piso.data_r_1708_sv2v_reg  <= 1'b0;
      \piso.data_r_1707_sv2v_reg  <= 1'b0;
      \piso.data_r_1706_sv2v_reg  <= 1'b0;
      \piso.data_r_1705_sv2v_reg  <= 1'b0;
      \piso.data_r_1704_sv2v_reg  <= 1'b0;
      \piso.data_r_1703_sv2v_reg  <= 1'b0;
      \piso.data_r_1702_sv2v_reg  <= 1'b0;
      \piso.data_r_1701_sv2v_reg  <= 1'b0;
      \piso.data_r_1700_sv2v_reg  <= 1'b0;
      \piso.data_r_1699_sv2v_reg  <= 1'b0;
      \piso.data_r_1698_sv2v_reg  <= 1'b0;
      \piso.data_r_1697_sv2v_reg  <= 1'b0;
      \piso.data_r_1696_sv2v_reg  <= 1'b0;
      \piso.data_r_1695_sv2v_reg  <= 1'b0;
      \piso.data_r_1694_sv2v_reg  <= 1'b0;
      \piso.data_r_1693_sv2v_reg  <= 1'b0;
      \piso.data_r_1692_sv2v_reg  <= 1'b0;
      \piso.data_r_1691_sv2v_reg  <= 1'b0;
      \piso.data_r_1690_sv2v_reg  <= 1'b0;
      \piso.data_r_1689_sv2v_reg  <= 1'b0;
      \piso.data_r_1688_sv2v_reg  <= 1'b0;
      \piso.data_r_1687_sv2v_reg  <= 1'b0;
      \piso.data_r_1686_sv2v_reg  <= 1'b0;
      \piso.data_r_1685_sv2v_reg  <= 1'b0;
      \piso.data_r_1684_sv2v_reg  <= 1'b0;
      \piso.data_r_1683_sv2v_reg  <= 1'b0;
      \piso.data_r_1682_sv2v_reg  <= 1'b0;
      \piso.data_r_1681_sv2v_reg  <= 1'b0;
      \piso.data_r_1680_sv2v_reg  <= 1'b0;
      \piso.data_r_1679_sv2v_reg  <= 1'b0;
      \piso.data_r_1678_sv2v_reg  <= 1'b0;
      \piso.data_r_1677_sv2v_reg  <= 1'b0;
      \piso.data_r_1676_sv2v_reg  <= 1'b0;
      \piso.data_r_1675_sv2v_reg  <= 1'b0;
      \piso.data_r_1674_sv2v_reg  <= 1'b0;
      \piso.data_r_1673_sv2v_reg  <= 1'b0;
      \piso.data_r_1672_sv2v_reg  <= 1'b0;
      \piso.data_r_1671_sv2v_reg  <= 1'b0;
      \piso.data_r_1670_sv2v_reg  <= 1'b0;
      \piso.data_r_1669_sv2v_reg  <= 1'b0;
      \piso.data_r_1668_sv2v_reg  <= 1'b0;
      \piso.data_r_1667_sv2v_reg  <= 1'b0;
      \piso.data_r_1666_sv2v_reg  <= 1'b0;
      \piso.data_r_1665_sv2v_reg  <= 1'b0;
      \piso.data_r_1664_sv2v_reg  <= 1'b0;
      \piso.data_r_1663_sv2v_reg  <= 1'b0;
      \piso.data_r_1662_sv2v_reg  <= 1'b0;
      \piso.data_r_1661_sv2v_reg  <= 1'b0;
      \piso.data_r_1660_sv2v_reg  <= 1'b0;
      \piso.data_r_1659_sv2v_reg  <= 1'b0;
      \piso.data_r_1658_sv2v_reg  <= 1'b0;
      \piso.data_r_1657_sv2v_reg  <= 1'b0;
      \piso.data_r_1656_sv2v_reg  <= 1'b0;
      \piso.data_r_1655_sv2v_reg  <= 1'b0;
      \piso.data_r_1654_sv2v_reg  <= 1'b0;
      \piso.data_r_1653_sv2v_reg  <= 1'b0;
      \piso.data_r_1652_sv2v_reg  <= 1'b0;
      \piso.data_r_1651_sv2v_reg  <= 1'b0;
      \piso.data_r_1650_sv2v_reg  <= 1'b0;
      \piso.data_r_1649_sv2v_reg  <= 1'b0;
      \piso.data_r_1648_sv2v_reg  <= 1'b0;
      \piso.data_r_1647_sv2v_reg  <= 1'b0;
      \piso.data_r_1646_sv2v_reg  <= 1'b0;
      \piso.data_r_1645_sv2v_reg  <= 1'b0;
      \piso.data_r_1644_sv2v_reg  <= 1'b0;
      \piso.data_r_1643_sv2v_reg  <= 1'b0;
      \piso.data_r_1642_sv2v_reg  <= 1'b0;
      \piso.data_r_1641_sv2v_reg  <= 1'b0;
      \piso.data_r_1640_sv2v_reg  <= 1'b0;
      \piso.data_r_1639_sv2v_reg  <= 1'b0;
      \piso.data_r_1638_sv2v_reg  <= 1'b0;
      \piso.data_r_1637_sv2v_reg  <= 1'b0;
      \piso.data_r_1636_sv2v_reg  <= 1'b0;
      \piso.data_r_1635_sv2v_reg  <= 1'b0;
      \piso.data_r_1634_sv2v_reg  <= 1'b0;
      \piso.data_r_1633_sv2v_reg  <= 1'b0;
      \piso.data_r_1632_sv2v_reg  <= 1'b0;
      \piso.data_r_1631_sv2v_reg  <= 1'b0;
      \piso.data_r_1630_sv2v_reg  <= 1'b0;
      \piso.data_r_1629_sv2v_reg  <= 1'b0;
      \piso.data_r_1628_sv2v_reg  <= 1'b0;
      \piso.data_r_1627_sv2v_reg  <= 1'b0;
      \piso.data_r_1626_sv2v_reg  <= 1'b0;
      \piso.data_r_1625_sv2v_reg  <= 1'b0;
      \piso.data_r_1624_sv2v_reg  <= 1'b0;
      \piso.data_r_1623_sv2v_reg  <= 1'b0;
      \piso.data_r_1622_sv2v_reg  <= 1'b0;
      \piso.data_r_1621_sv2v_reg  <= 1'b0;
      \piso.data_r_1620_sv2v_reg  <= 1'b0;
      \piso.data_r_1619_sv2v_reg  <= 1'b0;
      \piso.data_r_1618_sv2v_reg  <= 1'b0;
      \piso.data_r_1617_sv2v_reg  <= 1'b0;
      \piso.data_r_1616_sv2v_reg  <= 1'b0;
      \piso.data_r_1615_sv2v_reg  <= 1'b0;
      \piso.data_r_1614_sv2v_reg  <= 1'b0;
      \piso.data_r_1613_sv2v_reg  <= 1'b0;
      \piso.data_r_1612_sv2v_reg  <= 1'b0;
      \piso.data_r_1611_sv2v_reg  <= 1'b0;
      \piso.data_r_1610_sv2v_reg  <= 1'b0;
      \piso.data_r_1609_sv2v_reg  <= 1'b0;
      \piso.data_r_1608_sv2v_reg  <= 1'b0;
      \piso.data_r_1607_sv2v_reg  <= 1'b0;
      \piso.data_r_1606_sv2v_reg  <= 1'b0;
      \piso.data_r_1605_sv2v_reg  <= 1'b0;
      \piso.data_r_1604_sv2v_reg  <= 1'b0;
      \piso.data_r_1603_sv2v_reg  <= 1'b0;
      \piso.data_r_1602_sv2v_reg  <= 1'b0;
      \piso.data_r_1601_sv2v_reg  <= 1'b0;
      \piso.data_r_1600_sv2v_reg  <= 1'b0;
      \piso.data_r_1599_sv2v_reg  <= 1'b0;
      \piso.data_r_1598_sv2v_reg  <= 1'b0;
      \piso.data_r_1597_sv2v_reg  <= 1'b0;
      \piso.data_r_1596_sv2v_reg  <= 1'b0;
      \piso.data_r_1595_sv2v_reg  <= 1'b0;
      \piso.data_r_1594_sv2v_reg  <= 1'b0;
      \piso.data_r_1593_sv2v_reg  <= 1'b0;
      \piso.data_r_1592_sv2v_reg  <= 1'b0;
      \piso.data_r_1591_sv2v_reg  <= 1'b0;
      \piso.data_r_1590_sv2v_reg  <= 1'b0;
      \piso.data_r_1589_sv2v_reg  <= 1'b0;
      \piso.data_r_1588_sv2v_reg  <= 1'b0;
      \piso.data_r_1587_sv2v_reg  <= 1'b0;
      \piso.data_r_1586_sv2v_reg  <= 1'b0;
      \piso.data_r_1585_sv2v_reg  <= 1'b0;
      \piso.data_r_1584_sv2v_reg  <= 1'b0;
      \piso.data_r_1583_sv2v_reg  <= 1'b0;
      \piso.data_r_1582_sv2v_reg  <= 1'b0;
      \piso.data_r_1581_sv2v_reg  <= 1'b0;
      \piso.data_r_1580_sv2v_reg  <= 1'b0;
      \piso.data_r_1579_sv2v_reg  <= 1'b0;
      \piso.data_r_1578_sv2v_reg  <= 1'b0;
      \piso.data_r_1577_sv2v_reg  <= 1'b0;
      \piso.data_r_1576_sv2v_reg  <= 1'b0;
      \piso.data_r_1575_sv2v_reg  <= 1'b0;
      \piso.data_r_1574_sv2v_reg  <= 1'b0;
      \piso.data_r_1573_sv2v_reg  <= 1'b0;
      \piso.data_r_1572_sv2v_reg  <= 1'b0;
      \piso.data_r_1571_sv2v_reg  <= 1'b0;
      \piso.data_r_1570_sv2v_reg  <= 1'b0;
      \piso.data_r_1569_sv2v_reg  <= 1'b0;
      \piso.data_r_1568_sv2v_reg  <= 1'b0;
      \piso.data_r_1567_sv2v_reg  <= 1'b0;
      \piso.data_r_1566_sv2v_reg  <= 1'b0;
      \piso.data_r_1565_sv2v_reg  <= 1'b0;
      \piso.data_r_1564_sv2v_reg  <= 1'b0;
      \piso.data_r_1563_sv2v_reg  <= 1'b0;
      \piso.data_r_1562_sv2v_reg  <= 1'b0;
      \piso.data_r_1561_sv2v_reg  <= 1'b0;
      \piso.data_r_1560_sv2v_reg  <= 1'b0;
      \piso.data_r_1559_sv2v_reg  <= 1'b0;
      \piso.data_r_1558_sv2v_reg  <= 1'b0;
      \piso.data_r_1557_sv2v_reg  <= 1'b0;
      \piso.data_r_1556_sv2v_reg  <= 1'b0;
      \piso.data_r_1555_sv2v_reg  <= 1'b0;
      \piso.data_r_1554_sv2v_reg  <= 1'b0;
      \piso.data_r_1553_sv2v_reg  <= 1'b0;
      \piso.data_r_1552_sv2v_reg  <= 1'b0;
      \piso.data_r_1551_sv2v_reg  <= 1'b0;
      \piso.data_r_1550_sv2v_reg  <= 1'b0;
      \piso.data_r_1549_sv2v_reg  <= 1'b0;
      \piso.data_r_1548_sv2v_reg  <= 1'b0;
      \piso.data_r_1547_sv2v_reg  <= 1'b0;
      \piso.data_r_1546_sv2v_reg  <= 1'b0;
      \piso.data_r_1545_sv2v_reg  <= 1'b0;
      \piso.data_r_1544_sv2v_reg  <= 1'b0;
      \piso.data_r_1543_sv2v_reg  <= 1'b0;
      \piso.data_r_1542_sv2v_reg  <= 1'b0;
      \piso.data_r_1541_sv2v_reg  <= 1'b0;
      \piso.data_r_1540_sv2v_reg  <= 1'b0;
      \piso.data_r_1539_sv2v_reg  <= 1'b0;
      \piso.data_r_1538_sv2v_reg  <= 1'b0;
      \piso.data_r_1537_sv2v_reg  <= 1'b0;
      \piso.data_r_1536_sv2v_reg  <= 1'b0;
      \piso.data_r_1535_sv2v_reg  <= 1'b0;
      \piso.data_r_1534_sv2v_reg  <= 1'b0;
      \piso.data_r_1533_sv2v_reg  <= 1'b0;
      \piso.data_r_1532_sv2v_reg  <= 1'b0;
      \piso.data_r_1531_sv2v_reg  <= 1'b0;
      \piso.data_r_1530_sv2v_reg  <= 1'b0;
      \piso.data_r_1529_sv2v_reg  <= 1'b0;
      \piso.data_r_1528_sv2v_reg  <= 1'b0;
      \piso.data_r_1527_sv2v_reg  <= 1'b0;
      \piso.data_r_1526_sv2v_reg  <= 1'b0;
      \piso.data_r_1525_sv2v_reg  <= 1'b0;
      \piso.data_r_1524_sv2v_reg  <= 1'b0;
      \piso.data_r_1523_sv2v_reg  <= 1'b0;
      \piso.data_r_1522_sv2v_reg  <= 1'b0;
      \piso.data_r_1521_sv2v_reg  <= 1'b0;
      \piso.data_r_1520_sv2v_reg  <= 1'b0;
      \piso.data_r_1519_sv2v_reg  <= 1'b0;
      \piso.data_r_1518_sv2v_reg  <= 1'b0;
      \piso.data_r_1517_sv2v_reg  <= 1'b0;
      \piso.data_r_1516_sv2v_reg  <= 1'b0;
      \piso.data_r_1515_sv2v_reg  <= 1'b0;
      \piso.data_r_1514_sv2v_reg  <= 1'b0;
      \piso.data_r_1513_sv2v_reg  <= 1'b0;
      \piso.data_r_1512_sv2v_reg  <= 1'b0;
      \piso.data_r_1511_sv2v_reg  <= 1'b0;
      \piso.data_r_1510_sv2v_reg  <= 1'b0;
      \piso.data_r_1509_sv2v_reg  <= 1'b0;
      \piso.data_r_1508_sv2v_reg  <= 1'b0;
      \piso.data_r_1507_sv2v_reg  <= 1'b0;
      \piso.data_r_1506_sv2v_reg  <= 1'b0;
      \piso.data_r_1505_sv2v_reg  <= 1'b0;
      \piso.data_r_1504_sv2v_reg  <= 1'b0;
      \piso.data_r_1503_sv2v_reg  <= 1'b0;
      \piso.data_r_1502_sv2v_reg  <= 1'b0;
      \piso.data_r_1501_sv2v_reg  <= 1'b0;
      \piso.data_r_1500_sv2v_reg  <= 1'b0;
      \piso.data_r_1499_sv2v_reg  <= 1'b0;
      \piso.data_r_1498_sv2v_reg  <= 1'b0;
      \piso.data_r_1497_sv2v_reg  <= 1'b0;
      \piso.data_r_1496_sv2v_reg  <= 1'b0;
      \piso.data_r_1495_sv2v_reg  <= 1'b0;
      \piso.data_r_1494_sv2v_reg  <= 1'b0;
      \piso.data_r_1493_sv2v_reg  <= 1'b0;
      \piso.data_r_1492_sv2v_reg  <= 1'b0;
      \piso.data_r_1491_sv2v_reg  <= 1'b0;
      \piso.data_r_1490_sv2v_reg  <= 1'b0;
      \piso.data_r_1489_sv2v_reg  <= 1'b0;
      \piso.data_r_1488_sv2v_reg  <= 1'b0;
      \piso.data_r_1487_sv2v_reg  <= 1'b0;
      \piso.data_r_1486_sv2v_reg  <= 1'b0;
      \piso.data_r_1485_sv2v_reg  <= 1'b0;
      \piso.data_r_1484_sv2v_reg  <= 1'b0;
      \piso.data_r_1483_sv2v_reg  <= 1'b0;
      \piso.data_r_1482_sv2v_reg  <= 1'b0;
      \piso.data_r_1481_sv2v_reg  <= 1'b0;
      \piso.data_r_1480_sv2v_reg  <= 1'b0;
      \piso.data_r_1479_sv2v_reg  <= 1'b0;
      \piso.data_r_1478_sv2v_reg  <= 1'b0;
      \piso.data_r_1477_sv2v_reg  <= 1'b0;
      \piso.data_r_1476_sv2v_reg  <= 1'b0;
      \piso.data_r_1475_sv2v_reg  <= 1'b0;
      \piso.data_r_1474_sv2v_reg  <= 1'b0;
      \piso.data_r_1473_sv2v_reg  <= 1'b0;
      \piso.data_r_1472_sv2v_reg  <= 1'b0;
      \piso.data_r_1471_sv2v_reg  <= 1'b0;
      \piso.data_r_1470_sv2v_reg  <= 1'b0;
      \piso.data_r_1469_sv2v_reg  <= 1'b0;
      \piso.data_r_1468_sv2v_reg  <= 1'b0;
      \piso.data_r_1467_sv2v_reg  <= 1'b0;
      \piso.data_r_1466_sv2v_reg  <= 1'b0;
      \piso.data_r_1465_sv2v_reg  <= 1'b0;
      \piso.data_r_1464_sv2v_reg  <= 1'b0;
      \piso.data_r_1463_sv2v_reg  <= 1'b0;
      \piso.data_r_1462_sv2v_reg  <= 1'b0;
      \piso.data_r_1461_sv2v_reg  <= 1'b0;
      \piso.data_r_1460_sv2v_reg  <= 1'b0;
      \piso.data_r_1459_sv2v_reg  <= 1'b0;
      \piso.data_r_1458_sv2v_reg  <= 1'b0;
      \piso.data_r_1457_sv2v_reg  <= 1'b0;
      \piso.data_r_1456_sv2v_reg  <= 1'b0;
      \piso.data_r_1455_sv2v_reg  <= 1'b0;
      \piso.data_r_1454_sv2v_reg  <= 1'b0;
      \piso.data_r_1453_sv2v_reg  <= 1'b0;
      \piso.data_r_1452_sv2v_reg  <= 1'b0;
      \piso.data_r_1451_sv2v_reg  <= 1'b0;
      \piso.data_r_1450_sv2v_reg  <= 1'b0;
      \piso.data_r_1449_sv2v_reg  <= 1'b0;
      \piso.data_r_1448_sv2v_reg  <= 1'b0;
      \piso.data_r_1447_sv2v_reg  <= 1'b0;
      \piso.data_r_1446_sv2v_reg  <= 1'b0;
      \piso.data_r_1445_sv2v_reg  <= 1'b0;
      \piso.data_r_1444_sv2v_reg  <= 1'b0;
      \piso.data_r_1443_sv2v_reg  <= 1'b0;
      \piso.data_r_1442_sv2v_reg  <= 1'b0;
      \piso.data_r_1441_sv2v_reg  <= 1'b0;
      \piso.data_r_1440_sv2v_reg  <= 1'b0;
      \piso.data_r_1439_sv2v_reg  <= 1'b0;
      \piso.data_r_1438_sv2v_reg  <= 1'b0;
      \piso.data_r_1437_sv2v_reg  <= 1'b0;
      \piso.data_r_1436_sv2v_reg  <= 1'b0;
      \piso.data_r_1435_sv2v_reg  <= 1'b0;
      \piso.data_r_1434_sv2v_reg  <= 1'b0;
      \piso.data_r_1433_sv2v_reg  <= 1'b0;
      \piso.data_r_1432_sv2v_reg  <= 1'b0;
      \piso.data_r_1431_sv2v_reg  <= 1'b0;
      \piso.data_r_1430_sv2v_reg  <= 1'b0;
      \piso.data_r_1429_sv2v_reg  <= 1'b0;
      \piso.data_r_1428_sv2v_reg  <= 1'b0;
      \piso.data_r_1427_sv2v_reg  <= 1'b0;
      \piso.data_r_1426_sv2v_reg  <= 1'b0;
      \piso.data_r_1425_sv2v_reg  <= 1'b0;
      \piso.data_r_1424_sv2v_reg  <= 1'b0;
      \piso.data_r_1423_sv2v_reg  <= 1'b0;
      \piso.data_r_1422_sv2v_reg  <= 1'b0;
      \piso.data_r_1421_sv2v_reg  <= 1'b0;
      \piso.data_r_1420_sv2v_reg  <= 1'b0;
      \piso.data_r_1419_sv2v_reg  <= 1'b0;
      \piso.data_r_1418_sv2v_reg  <= 1'b0;
      \piso.data_r_1417_sv2v_reg  <= 1'b0;
      \piso.data_r_1416_sv2v_reg  <= 1'b0;
      \piso.data_r_1415_sv2v_reg  <= 1'b0;
      \piso.data_r_1414_sv2v_reg  <= 1'b0;
      \piso.data_r_1413_sv2v_reg  <= 1'b0;
      \piso.data_r_1412_sv2v_reg  <= 1'b0;
      \piso.data_r_1411_sv2v_reg  <= 1'b0;
      \piso.data_r_1410_sv2v_reg  <= 1'b0;
      \piso.data_r_1409_sv2v_reg  <= 1'b0;
      \piso.data_r_1408_sv2v_reg  <= 1'b0;
      \piso.data_r_1407_sv2v_reg  <= 1'b0;
      \piso.data_r_1406_sv2v_reg  <= 1'b0;
      \piso.data_r_1405_sv2v_reg  <= 1'b0;
      \piso.data_r_1404_sv2v_reg  <= 1'b0;
      \piso.data_r_1403_sv2v_reg  <= 1'b0;
      \piso.data_r_1402_sv2v_reg  <= 1'b0;
      \piso.data_r_1401_sv2v_reg  <= 1'b0;
      \piso.data_r_1400_sv2v_reg  <= 1'b0;
      \piso.data_r_1399_sv2v_reg  <= 1'b0;
      \piso.data_r_1398_sv2v_reg  <= 1'b0;
      \piso.data_r_1397_sv2v_reg  <= 1'b0;
      \piso.data_r_1396_sv2v_reg  <= 1'b0;
      \piso.data_r_1395_sv2v_reg  <= 1'b0;
      \piso.data_r_1394_sv2v_reg  <= 1'b0;
      \piso.data_r_1393_sv2v_reg  <= 1'b0;
      \piso.data_r_1392_sv2v_reg  <= 1'b0;
      \piso.data_r_1391_sv2v_reg  <= 1'b0;
      \piso.data_r_1390_sv2v_reg  <= 1'b0;
      \piso.data_r_1389_sv2v_reg  <= 1'b0;
      \piso.data_r_1388_sv2v_reg  <= 1'b0;
      \piso.data_r_1387_sv2v_reg  <= 1'b0;
      \piso.data_r_1386_sv2v_reg  <= 1'b0;
      \piso.data_r_1385_sv2v_reg  <= 1'b0;
      \piso.data_r_1384_sv2v_reg  <= 1'b0;
      \piso.data_r_1383_sv2v_reg  <= 1'b0;
      \piso.data_r_1382_sv2v_reg  <= 1'b0;
      \piso.data_r_1381_sv2v_reg  <= 1'b0;
      \piso.data_r_1380_sv2v_reg  <= 1'b0;
      \piso.data_r_1379_sv2v_reg  <= 1'b0;
      \piso.data_r_1378_sv2v_reg  <= 1'b0;
      \piso.data_r_1377_sv2v_reg  <= 1'b0;
      \piso.data_r_1376_sv2v_reg  <= 1'b0;
      \piso.data_r_1375_sv2v_reg  <= 1'b0;
      \piso.data_r_1374_sv2v_reg  <= 1'b0;
      \piso.data_r_1373_sv2v_reg  <= 1'b0;
      \piso.data_r_1372_sv2v_reg  <= 1'b0;
      \piso.data_r_1371_sv2v_reg  <= 1'b0;
      \piso.data_r_1370_sv2v_reg  <= 1'b0;
      \piso.data_r_1369_sv2v_reg  <= 1'b0;
      \piso.data_r_1368_sv2v_reg  <= 1'b0;
      \piso.data_r_1367_sv2v_reg  <= 1'b0;
      \piso.data_r_1366_sv2v_reg  <= 1'b0;
      \piso.data_r_1365_sv2v_reg  <= 1'b0;
      \piso.data_r_1364_sv2v_reg  <= 1'b0;
      \piso.data_r_1363_sv2v_reg  <= 1'b0;
      \piso.data_r_1362_sv2v_reg  <= 1'b0;
      \piso.data_r_1361_sv2v_reg  <= 1'b0;
      \piso.data_r_1360_sv2v_reg  <= 1'b0;
      \piso.data_r_1359_sv2v_reg  <= 1'b0;
      \piso.data_r_1358_sv2v_reg  <= 1'b0;
      \piso.data_r_1357_sv2v_reg  <= 1'b0;
      \piso.data_r_1356_sv2v_reg  <= 1'b0;
      \piso.data_r_1355_sv2v_reg  <= 1'b0;
      \piso.data_r_1354_sv2v_reg  <= 1'b0;
      \piso.data_r_1353_sv2v_reg  <= 1'b0;
      \piso.data_r_1352_sv2v_reg  <= 1'b0;
      \piso.data_r_1351_sv2v_reg  <= 1'b0;
      \piso.data_r_1350_sv2v_reg  <= 1'b0;
      \piso.data_r_1349_sv2v_reg  <= 1'b0;
      \piso.data_r_1348_sv2v_reg  <= 1'b0;
      \piso.data_r_1347_sv2v_reg  <= 1'b0;
      \piso.data_r_1346_sv2v_reg  <= 1'b0;
      \piso.data_r_1345_sv2v_reg  <= 1'b0;
      \piso.data_r_1344_sv2v_reg  <= 1'b0;
      \piso.data_r_1343_sv2v_reg  <= 1'b0;
      \piso.data_r_1342_sv2v_reg  <= 1'b0;
      \piso.data_r_1341_sv2v_reg  <= 1'b0;
      \piso.data_r_1340_sv2v_reg  <= 1'b0;
      \piso.data_r_1339_sv2v_reg  <= 1'b0;
      \piso.data_r_1338_sv2v_reg  <= 1'b0;
      \piso.data_r_1337_sv2v_reg  <= 1'b0;
      \piso.data_r_1336_sv2v_reg  <= 1'b0;
      \piso.data_r_1335_sv2v_reg  <= 1'b0;
      \piso.data_r_1334_sv2v_reg  <= 1'b0;
      \piso.data_r_1333_sv2v_reg  <= 1'b0;
      \piso.data_r_1332_sv2v_reg  <= 1'b0;
      \piso.data_r_1331_sv2v_reg  <= 1'b0;
      \piso.data_r_1330_sv2v_reg  <= 1'b0;
      \piso.data_r_1329_sv2v_reg  <= 1'b0;
      \piso.data_r_1328_sv2v_reg  <= 1'b0;
      \piso.data_r_1327_sv2v_reg  <= 1'b0;
      \piso.data_r_1326_sv2v_reg  <= 1'b0;
      \piso.data_r_1325_sv2v_reg  <= 1'b0;
      \piso.data_r_1324_sv2v_reg  <= 1'b0;
      \piso.data_r_1323_sv2v_reg  <= 1'b0;
      \piso.data_r_1322_sv2v_reg  <= 1'b0;
      \piso.data_r_1321_sv2v_reg  <= 1'b0;
      \piso.data_r_1320_sv2v_reg  <= 1'b0;
      \piso.data_r_1319_sv2v_reg  <= 1'b0;
      \piso.data_r_1318_sv2v_reg  <= 1'b0;
      \piso.data_r_1317_sv2v_reg  <= 1'b0;
      \piso.data_r_1316_sv2v_reg  <= 1'b0;
      \piso.data_r_1315_sv2v_reg  <= 1'b0;
      \piso.data_r_1314_sv2v_reg  <= 1'b0;
      \piso.data_r_1313_sv2v_reg  <= 1'b0;
      \piso.data_r_1312_sv2v_reg  <= 1'b0;
      \piso.data_r_1311_sv2v_reg  <= 1'b0;
      \piso.data_r_1310_sv2v_reg  <= 1'b0;
      \piso.data_r_1309_sv2v_reg  <= 1'b0;
      \piso.data_r_1308_sv2v_reg  <= 1'b0;
      \piso.data_r_1307_sv2v_reg  <= 1'b0;
      \piso.data_r_1306_sv2v_reg  <= 1'b0;
      \piso.data_r_1305_sv2v_reg  <= 1'b0;
      \piso.data_r_1304_sv2v_reg  <= 1'b0;
      \piso.data_r_1303_sv2v_reg  <= 1'b0;
      \piso.data_r_1302_sv2v_reg  <= 1'b0;
      \piso.data_r_1301_sv2v_reg  <= 1'b0;
      \piso.data_r_1300_sv2v_reg  <= 1'b0;
      \piso.data_r_1299_sv2v_reg  <= 1'b0;
      \piso.data_r_1298_sv2v_reg  <= 1'b0;
      \piso.data_r_1297_sv2v_reg  <= 1'b0;
      \piso.data_r_1296_sv2v_reg  <= 1'b0;
      \piso.data_r_1295_sv2v_reg  <= 1'b0;
      \piso.data_r_1294_sv2v_reg  <= 1'b0;
      \piso.data_r_1293_sv2v_reg  <= 1'b0;
      \piso.data_r_1292_sv2v_reg  <= 1'b0;
      \piso.data_r_1291_sv2v_reg  <= 1'b0;
      \piso.data_r_1290_sv2v_reg  <= 1'b0;
      \piso.data_r_1289_sv2v_reg  <= 1'b0;
      \piso.data_r_1288_sv2v_reg  <= 1'b0;
      \piso.data_r_1287_sv2v_reg  <= 1'b0;
      \piso.data_r_1286_sv2v_reg  <= 1'b0;
      \piso.data_r_1285_sv2v_reg  <= 1'b0;
      \piso.data_r_1284_sv2v_reg  <= 1'b0;
      \piso.data_r_1283_sv2v_reg  <= 1'b0;
      \piso.data_r_1282_sv2v_reg  <= 1'b0;
      \piso.data_r_1281_sv2v_reg  <= 1'b0;
      \piso.data_r_1280_sv2v_reg  <= 1'b0;
      \piso.data_r_1279_sv2v_reg  <= 1'b0;
      \piso.data_r_1278_sv2v_reg  <= 1'b0;
      \piso.data_r_1277_sv2v_reg  <= 1'b0;
      \piso.data_r_1276_sv2v_reg  <= 1'b0;
      \piso.data_r_1275_sv2v_reg  <= 1'b0;
      \piso.data_r_1274_sv2v_reg  <= 1'b0;
      \piso.data_r_1273_sv2v_reg  <= 1'b0;
      \piso.data_r_1272_sv2v_reg  <= 1'b0;
      \piso.data_r_1271_sv2v_reg  <= 1'b0;
      \piso.data_r_1270_sv2v_reg  <= 1'b0;
      \piso.data_r_1269_sv2v_reg  <= 1'b0;
      \piso.data_r_1268_sv2v_reg  <= 1'b0;
      \piso.data_r_1267_sv2v_reg  <= 1'b0;
      \piso.data_r_1266_sv2v_reg  <= 1'b0;
      \piso.data_r_1265_sv2v_reg  <= 1'b0;
      \piso.data_r_1264_sv2v_reg  <= 1'b0;
      \piso.data_r_1263_sv2v_reg  <= 1'b0;
      \piso.data_r_1262_sv2v_reg  <= 1'b0;
      \piso.data_r_1261_sv2v_reg  <= 1'b0;
      \piso.data_r_1260_sv2v_reg  <= 1'b0;
      \piso.data_r_1259_sv2v_reg  <= 1'b0;
      \piso.data_r_1258_sv2v_reg  <= 1'b0;
      \piso.data_r_1257_sv2v_reg  <= 1'b0;
      \piso.data_r_1256_sv2v_reg  <= 1'b0;
      \piso.data_r_1255_sv2v_reg  <= 1'b0;
      \piso.data_r_1254_sv2v_reg  <= 1'b0;
      \piso.data_r_1253_sv2v_reg  <= 1'b0;
      \piso.data_r_1252_sv2v_reg  <= 1'b0;
      \piso.data_r_1251_sv2v_reg  <= 1'b0;
      \piso.data_r_1250_sv2v_reg  <= 1'b0;
      \piso.data_r_1249_sv2v_reg  <= 1'b0;
      \piso.data_r_1248_sv2v_reg  <= 1'b0;
      \piso.data_r_1247_sv2v_reg  <= 1'b0;
      \piso.data_r_1246_sv2v_reg  <= 1'b0;
      \piso.data_r_1245_sv2v_reg  <= 1'b0;
      \piso.data_r_1244_sv2v_reg  <= 1'b0;
      \piso.data_r_1243_sv2v_reg  <= 1'b0;
      \piso.data_r_1242_sv2v_reg  <= 1'b0;
      \piso.data_r_1241_sv2v_reg  <= 1'b0;
      \piso.data_r_1240_sv2v_reg  <= 1'b0;
      \piso.data_r_1239_sv2v_reg  <= 1'b0;
      \piso.data_r_1238_sv2v_reg  <= 1'b0;
      \piso.data_r_1237_sv2v_reg  <= 1'b0;
      \piso.data_r_1236_sv2v_reg  <= 1'b0;
      \piso.data_r_1235_sv2v_reg  <= 1'b0;
      \piso.data_r_1234_sv2v_reg  <= 1'b0;
      \piso.data_r_1233_sv2v_reg  <= 1'b0;
      \piso.data_r_1232_sv2v_reg  <= 1'b0;
      \piso.data_r_1231_sv2v_reg  <= 1'b0;
      \piso.data_r_1230_sv2v_reg  <= 1'b0;
      \piso.data_r_1229_sv2v_reg  <= 1'b0;
      \piso.data_r_1228_sv2v_reg  <= 1'b0;
      \piso.data_r_1227_sv2v_reg  <= 1'b0;
      \piso.data_r_1226_sv2v_reg  <= 1'b0;
      \piso.data_r_1225_sv2v_reg  <= 1'b0;
      \piso.data_r_1224_sv2v_reg  <= 1'b0;
      \piso.data_r_1223_sv2v_reg  <= 1'b0;
      \piso.data_r_1222_sv2v_reg  <= 1'b0;
      \piso.data_r_1221_sv2v_reg  <= 1'b0;
      \piso.data_r_1220_sv2v_reg  <= 1'b0;
      \piso.data_r_1219_sv2v_reg  <= 1'b0;
      \piso.data_r_1218_sv2v_reg  <= 1'b0;
      \piso.data_r_1217_sv2v_reg  <= 1'b0;
      \piso.data_r_1216_sv2v_reg  <= 1'b0;
      \piso.data_r_1215_sv2v_reg  <= 1'b0;
      \piso.data_r_1214_sv2v_reg  <= 1'b0;
      \piso.data_r_1213_sv2v_reg  <= 1'b0;
      \piso.data_r_1212_sv2v_reg  <= 1'b0;
      \piso.data_r_1211_sv2v_reg  <= 1'b0;
      \piso.data_r_1210_sv2v_reg  <= 1'b0;
      \piso.data_r_1209_sv2v_reg  <= 1'b0;
      \piso.data_r_1208_sv2v_reg  <= 1'b0;
      \piso.data_r_1207_sv2v_reg  <= 1'b0;
      \piso.data_r_1206_sv2v_reg  <= 1'b0;
      \piso.data_r_1205_sv2v_reg  <= 1'b0;
      \piso.data_r_1204_sv2v_reg  <= 1'b0;
      \piso.data_r_1203_sv2v_reg  <= 1'b0;
      \piso.data_r_1202_sv2v_reg  <= 1'b0;
      \piso.data_r_1201_sv2v_reg  <= 1'b0;
      \piso.data_r_1200_sv2v_reg  <= 1'b0;
      \piso.data_r_1199_sv2v_reg  <= 1'b0;
      \piso.data_r_1198_sv2v_reg  <= 1'b0;
      \piso.data_r_1197_sv2v_reg  <= 1'b0;
      \piso.data_r_1196_sv2v_reg  <= 1'b0;
      \piso.data_r_1195_sv2v_reg  <= 1'b0;
      \piso.data_r_1194_sv2v_reg  <= 1'b0;
      \piso.data_r_1193_sv2v_reg  <= 1'b0;
      \piso.data_r_1192_sv2v_reg  <= 1'b0;
      \piso.data_r_1191_sv2v_reg  <= 1'b0;
      \piso.data_r_1190_sv2v_reg  <= 1'b0;
      \piso.data_r_1189_sv2v_reg  <= 1'b0;
      \piso.data_r_1188_sv2v_reg  <= 1'b0;
      \piso.data_r_1187_sv2v_reg  <= 1'b0;
      \piso.data_r_1186_sv2v_reg  <= 1'b0;
      \piso.data_r_1185_sv2v_reg  <= 1'b0;
      \piso.data_r_1184_sv2v_reg  <= 1'b0;
      \piso.data_r_1183_sv2v_reg  <= 1'b0;
      \piso.data_r_1182_sv2v_reg  <= 1'b0;
      \piso.data_r_1181_sv2v_reg  <= 1'b0;
      \piso.data_r_1180_sv2v_reg  <= 1'b0;
      \piso.data_r_1179_sv2v_reg  <= 1'b0;
      \piso.data_r_1178_sv2v_reg  <= 1'b0;
      \piso.data_r_1177_sv2v_reg  <= 1'b0;
      \piso.data_r_1176_sv2v_reg  <= 1'b0;
      \piso.data_r_1175_sv2v_reg  <= 1'b0;
      \piso.data_r_1174_sv2v_reg  <= 1'b0;
      \piso.data_r_1173_sv2v_reg  <= 1'b0;
      \piso.data_r_1172_sv2v_reg  <= 1'b0;
      \piso.data_r_1171_sv2v_reg  <= 1'b0;
      \piso.data_r_1170_sv2v_reg  <= 1'b0;
      \piso.data_r_1169_sv2v_reg  <= 1'b0;
      \piso.data_r_1168_sv2v_reg  <= 1'b0;
      \piso.data_r_1167_sv2v_reg  <= 1'b0;
      \piso.data_r_1166_sv2v_reg  <= 1'b0;
      \piso.data_r_1165_sv2v_reg  <= 1'b0;
      \piso.data_r_1164_sv2v_reg  <= 1'b0;
      \piso.data_r_1163_sv2v_reg  <= 1'b0;
      \piso.data_r_1162_sv2v_reg  <= 1'b0;
      \piso.data_r_1161_sv2v_reg  <= 1'b0;
      \piso.data_r_1160_sv2v_reg  <= 1'b0;
      \piso.data_r_1159_sv2v_reg  <= 1'b0;
      \piso.data_r_1158_sv2v_reg  <= 1'b0;
      \piso.data_r_1157_sv2v_reg  <= 1'b0;
      \piso.data_r_1156_sv2v_reg  <= 1'b0;
      \piso.data_r_1155_sv2v_reg  <= 1'b0;
      \piso.data_r_1154_sv2v_reg  <= 1'b0;
      \piso.data_r_1153_sv2v_reg  <= 1'b0;
      \piso.data_r_1152_sv2v_reg  <= 1'b0;
      \piso.data_r_1151_sv2v_reg  <= 1'b0;
      \piso.data_r_1150_sv2v_reg  <= 1'b0;
      \piso.data_r_1149_sv2v_reg  <= 1'b0;
      \piso.data_r_1148_sv2v_reg  <= 1'b0;
      \piso.data_r_1147_sv2v_reg  <= 1'b0;
      \piso.data_r_1146_sv2v_reg  <= 1'b0;
      \piso.data_r_1145_sv2v_reg  <= 1'b0;
      \piso.data_r_1144_sv2v_reg  <= 1'b0;
      \piso.data_r_1143_sv2v_reg  <= 1'b0;
      \piso.data_r_1142_sv2v_reg  <= 1'b0;
      \piso.data_r_1141_sv2v_reg  <= 1'b0;
      \piso.data_r_1140_sv2v_reg  <= 1'b0;
      \piso.data_r_1139_sv2v_reg  <= 1'b0;
      \piso.data_r_1138_sv2v_reg  <= 1'b0;
      \piso.data_r_1137_sv2v_reg  <= 1'b0;
      \piso.data_r_1136_sv2v_reg  <= 1'b0;
      \piso.data_r_1135_sv2v_reg  <= 1'b0;
      \piso.data_r_1134_sv2v_reg  <= 1'b0;
      \piso.data_r_1133_sv2v_reg  <= 1'b0;
      \piso.data_r_1132_sv2v_reg  <= 1'b0;
      \piso.data_r_1131_sv2v_reg  <= 1'b0;
      \piso.data_r_1130_sv2v_reg  <= 1'b0;
      \piso.data_r_1129_sv2v_reg  <= 1'b0;
      \piso.data_r_1128_sv2v_reg  <= 1'b0;
      \piso.data_r_1127_sv2v_reg  <= 1'b0;
      \piso.data_r_1126_sv2v_reg  <= 1'b0;
      \piso.data_r_1125_sv2v_reg  <= 1'b0;
      \piso.data_r_1124_sv2v_reg  <= 1'b0;
      \piso.data_r_1123_sv2v_reg  <= 1'b0;
      \piso.data_r_1122_sv2v_reg  <= 1'b0;
      \piso.data_r_1121_sv2v_reg  <= 1'b0;
      \piso.data_r_1120_sv2v_reg  <= 1'b0;
      \piso.data_r_1119_sv2v_reg  <= 1'b0;
      \piso.data_r_1118_sv2v_reg  <= 1'b0;
      \piso.data_r_1117_sv2v_reg  <= 1'b0;
      \piso.data_r_1116_sv2v_reg  <= 1'b0;
      \piso.data_r_1115_sv2v_reg  <= 1'b0;
      \piso.data_r_1114_sv2v_reg  <= 1'b0;
      \piso.data_r_1113_sv2v_reg  <= 1'b0;
      \piso.data_r_1112_sv2v_reg  <= 1'b0;
      \piso.data_r_1111_sv2v_reg  <= 1'b0;
      \piso.data_r_1110_sv2v_reg  <= 1'b0;
      \piso.data_r_1109_sv2v_reg  <= 1'b0;
      \piso.data_r_1108_sv2v_reg  <= 1'b0;
      \piso.data_r_1107_sv2v_reg  <= 1'b0;
      \piso.data_r_1106_sv2v_reg  <= 1'b0;
      \piso.data_r_1105_sv2v_reg  <= 1'b0;
      \piso.data_r_1104_sv2v_reg  <= 1'b0;
      \piso.data_r_1103_sv2v_reg  <= 1'b0;
      \piso.data_r_1102_sv2v_reg  <= 1'b0;
      \piso.data_r_1101_sv2v_reg  <= 1'b0;
      \piso.data_r_1100_sv2v_reg  <= 1'b0;
      \piso.data_r_1099_sv2v_reg  <= 1'b0;
      \piso.data_r_1098_sv2v_reg  <= 1'b0;
      \piso.data_r_1097_sv2v_reg  <= 1'b0;
      \piso.data_r_1096_sv2v_reg  <= 1'b0;
      \piso.data_r_1095_sv2v_reg  <= 1'b0;
      \piso.data_r_1094_sv2v_reg  <= 1'b0;
      \piso.data_r_1093_sv2v_reg  <= 1'b0;
      \piso.data_r_1092_sv2v_reg  <= 1'b0;
      \piso.data_r_1091_sv2v_reg  <= 1'b0;
      \piso.data_r_1090_sv2v_reg  <= 1'b0;
      \piso.data_r_1089_sv2v_reg  <= 1'b0;
      \piso.data_r_1088_sv2v_reg  <= 1'b0;
      \piso.data_r_1087_sv2v_reg  <= 1'b0;
      \piso.data_r_1086_sv2v_reg  <= 1'b0;
      \piso.data_r_1085_sv2v_reg  <= 1'b0;
      \piso.data_r_1084_sv2v_reg  <= 1'b0;
      \piso.data_r_1083_sv2v_reg  <= 1'b0;
      \piso.data_r_1082_sv2v_reg  <= 1'b0;
      \piso.data_r_1081_sv2v_reg  <= 1'b0;
      \piso.data_r_1080_sv2v_reg  <= 1'b0;
      \piso.data_r_1079_sv2v_reg  <= 1'b0;
      \piso.data_r_1078_sv2v_reg  <= 1'b0;
      \piso.data_r_1077_sv2v_reg  <= 1'b0;
      \piso.data_r_1076_sv2v_reg  <= 1'b0;
      \piso.data_r_1075_sv2v_reg  <= 1'b0;
      \piso.data_r_1074_sv2v_reg  <= 1'b0;
      \piso.data_r_1073_sv2v_reg  <= 1'b0;
      \piso.data_r_1072_sv2v_reg  <= 1'b0;
      \piso.data_r_1071_sv2v_reg  <= 1'b0;
      \piso.data_r_1070_sv2v_reg  <= 1'b0;
      \piso.data_r_1069_sv2v_reg  <= 1'b0;
      \piso.data_r_1068_sv2v_reg  <= 1'b0;
      \piso.data_r_1067_sv2v_reg  <= 1'b0;
      \piso.data_r_1066_sv2v_reg  <= 1'b0;
      \piso.data_r_1065_sv2v_reg  <= 1'b0;
      \piso.data_r_1064_sv2v_reg  <= 1'b0;
      \piso.data_r_1063_sv2v_reg  <= 1'b0;
      \piso.data_r_1062_sv2v_reg  <= 1'b0;
      \piso.data_r_1061_sv2v_reg  <= 1'b0;
      \piso.data_r_1060_sv2v_reg  <= 1'b0;
      \piso.data_r_1059_sv2v_reg  <= 1'b0;
      \piso.data_r_1058_sv2v_reg  <= 1'b0;
      \piso.data_r_1057_sv2v_reg  <= 1'b0;
      \piso.data_r_1056_sv2v_reg  <= 1'b0;
      \piso.data_r_1055_sv2v_reg  <= 1'b0;
      \piso.data_r_1054_sv2v_reg  <= 1'b0;
      \piso.data_r_1053_sv2v_reg  <= 1'b0;
      \piso.data_r_1052_sv2v_reg  <= 1'b0;
      \piso.data_r_1051_sv2v_reg  <= 1'b0;
      \piso.data_r_1050_sv2v_reg  <= 1'b0;
      \piso.data_r_1049_sv2v_reg  <= 1'b0;
      \piso.data_r_1048_sv2v_reg  <= 1'b0;
      \piso.data_r_1047_sv2v_reg  <= 1'b0;
      \piso.data_r_1046_sv2v_reg  <= 1'b0;
      \piso.data_r_1045_sv2v_reg  <= 1'b0;
      \piso.data_r_1044_sv2v_reg  <= 1'b0;
      \piso.data_r_1043_sv2v_reg  <= 1'b0;
      \piso.data_r_1042_sv2v_reg  <= 1'b0;
      \piso.data_r_1041_sv2v_reg  <= 1'b0;
      \piso.data_r_1040_sv2v_reg  <= 1'b0;
      \piso.data_r_1039_sv2v_reg  <= 1'b0;
      \piso.data_r_1038_sv2v_reg  <= 1'b0;
      \piso.data_r_1037_sv2v_reg  <= 1'b0;
      \piso.data_r_1036_sv2v_reg  <= 1'b0;
      \piso.data_r_1035_sv2v_reg  <= 1'b0;
      \piso.data_r_1034_sv2v_reg  <= 1'b0;
      \piso.data_r_1033_sv2v_reg  <= 1'b0;
      \piso.data_r_1032_sv2v_reg  <= 1'b0;
      \piso.data_r_1031_sv2v_reg  <= 1'b0;
      \piso.data_r_1030_sv2v_reg  <= 1'b0;
      \piso.data_r_1029_sv2v_reg  <= 1'b0;
      \piso.data_r_1028_sv2v_reg  <= 1'b0;
      \piso.data_r_1027_sv2v_reg  <= 1'b0;
      \piso.data_r_1026_sv2v_reg  <= 1'b0;
      \piso.data_r_1025_sv2v_reg  <= 1'b0;
      \piso.data_r_1024_sv2v_reg  <= 1'b0;
      \piso.data_r_1023_sv2v_reg  <= 1'b0;
      \piso.data_r_1022_sv2v_reg  <= 1'b0;
      \piso.data_r_1021_sv2v_reg  <= 1'b0;
      \piso.data_r_1020_sv2v_reg  <= 1'b0;
      \piso.data_r_1019_sv2v_reg  <= 1'b0;
      \piso.data_r_1018_sv2v_reg  <= 1'b0;
      \piso.data_r_1017_sv2v_reg  <= 1'b0;
      \piso.data_r_1016_sv2v_reg  <= 1'b0;
      \piso.data_r_1015_sv2v_reg  <= 1'b0;
      \piso.data_r_1014_sv2v_reg  <= 1'b0;
      \piso.data_r_1013_sv2v_reg  <= 1'b0;
      \piso.data_r_1012_sv2v_reg  <= 1'b0;
      \piso.data_r_1011_sv2v_reg  <= 1'b0;
      \piso.data_r_1010_sv2v_reg  <= 1'b0;
      \piso.data_r_1009_sv2v_reg  <= 1'b0;
      \piso.data_r_1008_sv2v_reg  <= 1'b0;
      \piso.data_r_1007_sv2v_reg  <= 1'b0;
      \piso.data_r_1006_sv2v_reg  <= 1'b0;
      \piso.data_r_1005_sv2v_reg  <= 1'b0;
      \piso.data_r_1004_sv2v_reg  <= 1'b0;
      \piso.data_r_1003_sv2v_reg  <= 1'b0;
      \piso.data_r_1002_sv2v_reg  <= 1'b0;
      \piso.data_r_1001_sv2v_reg  <= 1'b0;
      \piso.data_r_1000_sv2v_reg  <= 1'b0;
      \piso.data_r_999_sv2v_reg  <= 1'b0;
      \piso.data_r_998_sv2v_reg  <= 1'b0;
      \piso.data_r_997_sv2v_reg  <= 1'b0;
      \piso.data_r_996_sv2v_reg  <= 1'b0;
      \piso.data_r_995_sv2v_reg  <= 1'b0;
      \piso.data_r_994_sv2v_reg  <= 1'b0;
      \piso.data_r_993_sv2v_reg  <= 1'b0;
      \piso.data_r_992_sv2v_reg  <= 1'b0;
      \piso.data_r_991_sv2v_reg  <= 1'b0;
      \piso.data_r_990_sv2v_reg  <= 1'b0;
      \piso.data_r_989_sv2v_reg  <= 1'b0;
      \piso.data_r_988_sv2v_reg  <= 1'b0;
      \piso.data_r_987_sv2v_reg  <= 1'b0;
      \piso.data_r_986_sv2v_reg  <= 1'b0;
      \piso.data_r_985_sv2v_reg  <= 1'b0;
      \piso.data_r_984_sv2v_reg  <= 1'b0;
      \piso.data_r_983_sv2v_reg  <= 1'b0;
      \piso.data_r_982_sv2v_reg  <= 1'b0;
      \piso.data_r_981_sv2v_reg  <= 1'b0;
      \piso.data_r_980_sv2v_reg  <= 1'b0;
      \piso.data_r_979_sv2v_reg  <= 1'b0;
      \piso.data_r_978_sv2v_reg  <= 1'b0;
      \piso.data_r_977_sv2v_reg  <= 1'b0;
      \piso.data_r_976_sv2v_reg  <= 1'b0;
      \piso.data_r_975_sv2v_reg  <= 1'b0;
      \piso.data_r_974_sv2v_reg  <= 1'b0;
      \piso.data_r_973_sv2v_reg  <= 1'b0;
      \piso.data_r_972_sv2v_reg  <= 1'b0;
      \piso.data_r_971_sv2v_reg  <= 1'b0;
      \piso.data_r_970_sv2v_reg  <= 1'b0;
      \piso.data_r_969_sv2v_reg  <= 1'b0;
      \piso.data_r_968_sv2v_reg  <= 1'b0;
      \piso.data_r_967_sv2v_reg  <= 1'b0;
      \piso.data_r_966_sv2v_reg  <= 1'b0;
      \piso.data_r_965_sv2v_reg  <= 1'b0;
      \piso.data_r_964_sv2v_reg  <= 1'b0;
      \piso.data_r_963_sv2v_reg  <= 1'b0;
      \piso.data_r_962_sv2v_reg  <= 1'b0;
      \piso.data_r_961_sv2v_reg  <= 1'b0;
      \piso.data_r_960_sv2v_reg  <= 1'b0;
      \piso.data_r_959_sv2v_reg  <= 1'b0;
      \piso.data_r_958_sv2v_reg  <= 1'b0;
      \piso.data_r_957_sv2v_reg  <= 1'b0;
      \piso.data_r_956_sv2v_reg  <= 1'b0;
      \piso.data_r_955_sv2v_reg  <= 1'b0;
      \piso.data_r_954_sv2v_reg  <= 1'b0;
      \piso.data_r_953_sv2v_reg  <= 1'b0;
      \piso.data_r_952_sv2v_reg  <= 1'b0;
      \piso.data_r_951_sv2v_reg  <= 1'b0;
      \piso.data_r_950_sv2v_reg  <= 1'b0;
      \piso.data_r_949_sv2v_reg  <= 1'b0;
      \piso.data_r_948_sv2v_reg  <= 1'b0;
      \piso.data_r_947_sv2v_reg  <= 1'b0;
      \piso.data_r_946_sv2v_reg  <= 1'b0;
      \piso.data_r_945_sv2v_reg  <= 1'b0;
      \piso.data_r_944_sv2v_reg  <= 1'b0;
      \piso.data_r_943_sv2v_reg  <= 1'b0;
      \piso.data_r_942_sv2v_reg  <= 1'b0;
      \piso.data_r_941_sv2v_reg  <= 1'b0;
      \piso.data_r_940_sv2v_reg  <= 1'b0;
      \piso.data_r_939_sv2v_reg  <= 1'b0;
      \piso.data_r_938_sv2v_reg  <= 1'b0;
      \piso.data_r_937_sv2v_reg  <= 1'b0;
      \piso.data_r_936_sv2v_reg  <= 1'b0;
      \piso.data_r_935_sv2v_reg  <= 1'b0;
      \piso.data_r_934_sv2v_reg  <= 1'b0;
      \piso.data_r_933_sv2v_reg  <= 1'b0;
      \piso.data_r_932_sv2v_reg  <= 1'b0;
      \piso.data_r_931_sv2v_reg  <= 1'b0;
      \piso.data_r_930_sv2v_reg  <= 1'b0;
      \piso.data_r_929_sv2v_reg  <= 1'b0;
      \piso.data_r_928_sv2v_reg  <= 1'b0;
      \piso.data_r_927_sv2v_reg  <= 1'b0;
      \piso.data_r_926_sv2v_reg  <= 1'b0;
      \piso.data_r_925_sv2v_reg  <= 1'b0;
      \piso.data_r_924_sv2v_reg  <= 1'b0;
      \piso.data_r_923_sv2v_reg  <= 1'b0;
      \piso.data_r_922_sv2v_reg  <= 1'b0;
      \piso.data_r_921_sv2v_reg  <= 1'b0;
      \piso.data_r_920_sv2v_reg  <= 1'b0;
      \piso.data_r_919_sv2v_reg  <= 1'b0;
      \piso.data_r_918_sv2v_reg  <= 1'b0;
      \piso.data_r_917_sv2v_reg  <= 1'b0;
      \piso.data_r_916_sv2v_reg  <= 1'b0;
      \piso.data_r_915_sv2v_reg  <= 1'b0;
      \piso.data_r_914_sv2v_reg  <= 1'b0;
      \piso.data_r_913_sv2v_reg  <= 1'b0;
      \piso.data_r_912_sv2v_reg  <= 1'b0;
      \piso.data_r_911_sv2v_reg  <= 1'b0;
      \piso.data_r_910_sv2v_reg  <= 1'b0;
      \piso.data_r_909_sv2v_reg  <= 1'b0;
      \piso.data_r_908_sv2v_reg  <= 1'b0;
      \piso.data_r_907_sv2v_reg  <= 1'b0;
      \piso.data_r_906_sv2v_reg  <= 1'b0;
      \piso.data_r_905_sv2v_reg  <= 1'b0;
      \piso.data_r_904_sv2v_reg  <= 1'b0;
      \piso.data_r_903_sv2v_reg  <= 1'b0;
      \piso.data_r_902_sv2v_reg  <= 1'b0;
      \piso.data_r_901_sv2v_reg  <= 1'b0;
      \piso.data_r_900_sv2v_reg  <= 1'b0;
      \piso.data_r_899_sv2v_reg  <= 1'b0;
      \piso.data_r_898_sv2v_reg  <= 1'b0;
      \piso.data_r_897_sv2v_reg  <= 1'b0;
      \piso.data_r_896_sv2v_reg  <= 1'b0;
      \piso.data_r_895_sv2v_reg  <= 1'b0;
      \piso.data_r_894_sv2v_reg  <= 1'b0;
      \piso.data_r_893_sv2v_reg  <= 1'b0;
      \piso.data_r_892_sv2v_reg  <= 1'b0;
      \piso.data_r_891_sv2v_reg  <= 1'b0;
      \piso.data_r_890_sv2v_reg  <= 1'b0;
      \piso.data_r_889_sv2v_reg  <= 1'b0;
      \piso.data_r_888_sv2v_reg  <= 1'b0;
      \piso.data_r_887_sv2v_reg  <= 1'b0;
      \piso.data_r_886_sv2v_reg  <= 1'b0;
      \piso.data_r_885_sv2v_reg  <= 1'b0;
      \piso.data_r_884_sv2v_reg  <= 1'b0;
      \piso.data_r_883_sv2v_reg  <= 1'b0;
      \piso.data_r_882_sv2v_reg  <= 1'b0;
      \piso.data_r_881_sv2v_reg  <= 1'b0;
      \piso.data_r_880_sv2v_reg  <= 1'b0;
      \piso.data_r_879_sv2v_reg  <= 1'b0;
      \piso.data_r_878_sv2v_reg  <= 1'b0;
      \piso.data_r_877_sv2v_reg  <= 1'b0;
      \piso.data_r_876_sv2v_reg  <= 1'b0;
      \piso.data_r_875_sv2v_reg  <= 1'b0;
      \piso.data_r_874_sv2v_reg  <= 1'b0;
      \piso.data_r_873_sv2v_reg  <= 1'b0;
      \piso.data_r_872_sv2v_reg  <= 1'b0;
      \piso.data_r_871_sv2v_reg  <= 1'b0;
      \piso.data_r_870_sv2v_reg  <= 1'b0;
      \piso.data_r_869_sv2v_reg  <= 1'b0;
      \piso.data_r_868_sv2v_reg  <= 1'b0;
      \piso.data_r_867_sv2v_reg  <= 1'b0;
      \piso.data_r_866_sv2v_reg  <= 1'b0;
      \piso.data_r_865_sv2v_reg  <= 1'b0;
      \piso.data_r_864_sv2v_reg  <= 1'b0;
      \piso.data_r_863_sv2v_reg  <= 1'b0;
      \piso.data_r_862_sv2v_reg  <= 1'b0;
      \piso.data_r_861_sv2v_reg  <= 1'b0;
      \piso.data_r_860_sv2v_reg  <= 1'b0;
      \piso.data_r_859_sv2v_reg  <= 1'b0;
      \piso.data_r_858_sv2v_reg  <= 1'b0;
      \piso.data_r_857_sv2v_reg  <= 1'b0;
      \piso.data_r_856_sv2v_reg  <= 1'b0;
      \piso.data_r_855_sv2v_reg  <= 1'b0;
      \piso.data_r_854_sv2v_reg  <= 1'b0;
      \piso.data_r_853_sv2v_reg  <= 1'b0;
      \piso.data_r_852_sv2v_reg  <= 1'b0;
      \piso.data_r_851_sv2v_reg  <= 1'b0;
      \piso.data_r_850_sv2v_reg  <= 1'b0;
      \piso.data_r_849_sv2v_reg  <= 1'b0;
      \piso.data_r_848_sv2v_reg  <= 1'b0;
      \piso.data_r_847_sv2v_reg  <= 1'b0;
      \piso.data_r_846_sv2v_reg  <= 1'b0;
      \piso.data_r_845_sv2v_reg  <= 1'b0;
      \piso.data_r_844_sv2v_reg  <= 1'b0;
      \piso.data_r_843_sv2v_reg  <= 1'b0;
      \piso.data_r_842_sv2v_reg  <= 1'b0;
      \piso.data_r_841_sv2v_reg  <= 1'b0;
      \piso.data_r_840_sv2v_reg  <= 1'b0;
      \piso.data_r_839_sv2v_reg  <= 1'b0;
      \piso.data_r_838_sv2v_reg  <= 1'b0;
      \piso.data_r_837_sv2v_reg  <= 1'b0;
      \piso.data_r_836_sv2v_reg  <= 1'b0;
      \piso.data_r_835_sv2v_reg  <= 1'b0;
      \piso.data_r_834_sv2v_reg  <= 1'b0;
      \piso.data_r_833_sv2v_reg  <= 1'b0;
      \piso.data_r_832_sv2v_reg  <= 1'b0;
      \piso.data_r_831_sv2v_reg  <= 1'b0;
      \piso.data_r_830_sv2v_reg  <= 1'b0;
      \piso.data_r_829_sv2v_reg  <= 1'b0;
      \piso.data_r_828_sv2v_reg  <= 1'b0;
      \piso.data_r_827_sv2v_reg  <= 1'b0;
      \piso.data_r_826_sv2v_reg  <= 1'b0;
      \piso.data_r_825_sv2v_reg  <= 1'b0;
      \piso.data_r_824_sv2v_reg  <= 1'b0;
      \piso.data_r_823_sv2v_reg  <= 1'b0;
      \piso.data_r_822_sv2v_reg  <= 1'b0;
      \piso.data_r_821_sv2v_reg  <= 1'b0;
      \piso.data_r_820_sv2v_reg  <= 1'b0;
      \piso.data_r_819_sv2v_reg  <= 1'b0;
      \piso.data_r_818_sv2v_reg  <= 1'b0;
      \piso.data_r_817_sv2v_reg  <= 1'b0;
      \piso.data_r_816_sv2v_reg  <= 1'b0;
      \piso.data_r_815_sv2v_reg  <= 1'b0;
      \piso.data_r_814_sv2v_reg  <= 1'b0;
      \piso.data_r_813_sv2v_reg  <= 1'b0;
      \piso.data_r_812_sv2v_reg  <= 1'b0;
      \piso.data_r_811_sv2v_reg  <= 1'b0;
      \piso.data_r_810_sv2v_reg  <= 1'b0;
      \piso.data_r_809_sv2v_reg  <= 1'b0;
      \piso.data_r_808_sv2v_reg  <= 1'b0;
      \piso.data_r_807_sv2v_reg  <= 1'b0;
      \piso.data_r_806_sv2v_reg  <= 1'b0;
      \piso.data_r_805_sv2v_reg  <= 1'b0;
      \piso.data_r_804_sv2v_reg  <= 1'b0;
      \piso.data_r_803_sv2v_reg  <= 1'b0;
      \piso.data_r_802_sv2v_reg  <= 1'b0;
      \piso.data_r_801_sv2v_reg  <= 1'b0;
      \piso.data_r_800_sv2v_reg  <= 1'b0;
      \piso.data_r_799_sv2v_reg  <= 1'b0;
      \piso.data_r_798_sv2v_reg  <= 1'b0;
      \piso.data_r_797_sv2v_reg  <= 1'b0;
      \piso.data_r_796_sv2v_reg  <= 1'b0;
      \piso.data_r_795_sv2v_reg  <= 1'b0;
      \piso.data_r_794_sv2v_reg  <= 1'b0;
      \piso.data_r_793_sv2v_reg  <= 1'b0;
      \piso.data_r_792_sv2v_reg  <= 1'b0;
      \piso.data_r_791_sv2v_reg  <= 1'b0;
      \piso.data_r_790_sv2v_reg  <= 1'b0;
      \piso.data_r_789_sv2v_reg  <= 1'b0;
      \piso.data_r_788_sv2v_reg  <= 1'b0;
      \piso.data_r_787_sv2v_reg  <= 1'b0;
      \piso.data_r_786_sv2v_reg  <= 1'b0;
      \piso.data_r_785_sv2v_reg  <= 1'b0;
      \piso.data_r_784_sv2v_reg  <= 1'b0;
      \piso.data_r_783_sv2v_reg  <= 1'b0;
      \piso.data_r_782_sv2v_reg  <= 1'b0;
      \piso.data_r_781_sv2v_reg  <= 1'b0;
      \piso.data_r_780_sv2v_reg  <= 1'b0;
      \piso.data_r_779_sv2v_reg  <= 1'b0;
      \piso.data_r_778_sv2v_reg  <= 1'b0;
      \piso.data_r_777_sv2v_reg  <= 1'b0;
      \piso.data_r_776_sv2v_reg  <= 1'b0;
      \piso.data_r_775_sv2v_reg  <= 1'b0;
      \piso.data_r_774_sv2v_reg  <= 1'b0;
      \piso.data_r_773_sv2v_reg  <= 1'b0;
      \piso.data_r_772_sv2v_reg  <= 1'b0;
      \piso.data_r_771_sv2v_reg  <= 1'b0;
      \piso.data_r_770_sv2v_reg  <= 1'b0;
      \piso.data_r_769_sv2v_reg  <= 1'b0;
      \piso.data_r_768_sv2v_reg  <= 1'b0;
      \piso.data_r_767_sv2v_reg  <= 1'b0;
      \piso.data_r_766_sv2v_reg  <= 1'b0;
      \piso.data_r_765_sv2v_reg  <= 1'b0;
      \piso.data_r_764_sv2v_reg  <= 1'b0;
      \piso.data_r_763_sv2v_reg  <= 1'b0;
      \piso.data_r_762_sv2v_reg  <= 1'b0;
      \piso.data_r_761_sv2v_reg  <= 1'b0;
      \piso.data_r_760_sv2v_reg  <= 1'b0;
      \piso.data_r_759_sv2v_reg  <= 1'b0;
      \piso.data_r_758_sv2v_reg  <= 1'b0;
      \piso.data_r_757_sv2v_reg  <= 1'b0;
      \piso.data_r_756_sv2v_reg  <= 1'b0;
      \piso.data_r_755_sv2v_reg  <= 1'b0;
      \piso.data_r_754_sv2v_reg  <= 1'b0;
      \piso.data_r_753_sv2v_reg  <= 1'b0;
      \piso.data_r_752_sv2v_reg  <= 1'b0;
      \piso.data_r_751_sv2v_reg  <= 1'b0;
      \piso.data_r_750_sv2v_reg  <= 1'b0;
      \piso.data_r_749_sv2v_reg  <= 1'b0;
      \piso.data_r_748_sv2v_reg  <= 1'b0;
      \piso.data_r_747_sv2v_reg  <= 1'b0;
      \piso.data_r_746_sv2v_reg  <= 1'b0;
      \piso.data_r_745_sv2v_reg  <= 1'b0;
      \piso.data_r_744_sv2v_reg  <= 1'b0;
      \piso.data_r_743_sv2v_reg  <= 1'b0;
      \piso.data_r_742_sv2v_reg  <= 1'b0;
      \piso.data_r_741_sv2v_reg  <= 1'b0;
      \piso.data_r_740_sv2v_reg  <= 1'b0;
      \piso.data_r_739_sv2v_reg  <= 1'b0;
      \piso.data_r_738_sv2v_reg  <= 1'b0;
      \piso.data_r_737_sv2v_reg  <= 1'b0;
      \piso.data_r_736_sv2v_reg  <= 1'b0;
      \piso.data_r_735_sv2v_reg  <= 1'b0;
      \piso.data_r_734_sv2v_reg  <= 1'b0;
      \piso.data_r_733_sv2v_reg  <= 1'b0;
      \piso.data_r_732_sv2v_reg  <= 1'b0;
      \piso.data_r_731_sv2v_reg  <= 1'b0;
      \piso.data_r_730_sv2v_reg  <= 1'b0;
      \piso.data_r_729_sv2v_reg  <= 1'b0;
      \piso.data_r_728_sv2v_reg  <= 1'b0;
      \piso.data_r_727_sv2v_reg  <= 1'b0;
      \piso.data_r_726_sv2v_reg  <= 1'b0;
      \piso.data_r_725_sv2v_reg  <= 1'b0;
      \piso.data_r_724_sv2v_reg  <= 1'b0;
      \piso.data_r_723_sv2v_reg  <= 1'b0;
      \piso.data_r_722_sv2v_reg  <= 1'b0;
      \piso.data_r_721_sv2v_reg  <= 1'b0;
      \piso.data_r_720_sv2v_reg  <= 1'b0;
      \piso.data_r_719_sv2v_reg  <= 1'b0;
      \piso.data_r_718_sv2v_reg  <= 1'b0;
      \piso.data_r_717_sv2v_reg  <= 1'b0;
      \piso.data_r_716_sv2v_reg  <= 1'b0;
      \piso.data_r_715_sv2v_reg  <= 1'b0;
      \piso.data_r_714_sv2v_reg  <= 1'b0;
      \piso.data_r_713_sv2v_reg  <= 1'b0;
      \piso.data_r_712_sv2v_reg  <= 1'b0;
      \piso.data_r_711_sv2v_reg  <= 1'b0;
      \piso.data_r_710_sv2v_reg  <= 1'b0;
      \piso.data_r_709_sv2v_reg  <= 1'b0;
      \piso.data_r_708_sv2v_reg  <= 1'b0;
      \piso.data_r_707_sv2v_reg  <= 1'b0;
      \piso.data_r_706_sv2v_reg  <= 1'b0;
      \piso.data_r_705_sv2v_reg  <= 1'b0;
      \piso.data_r_704_sv2v_reg  <= 1'b0;
      \piso.data_r_703_sv2v_reg  <= 1'b0;
      \piso.data_r_702_sv2v_reg  <= 1'b0;
      \piso.data_r_701_sv2v_reg  <= 1'b0;
      \piso.data_r_700_sv2v_reg  <= 1'b0;
      \piso.data_r_699_sv2v_reg  <= 1'b0;
      \piso.data_r_698_sv2v_reg  <= 1'b0;
      \piso.data_r_697_sv2v_reg  <= 1'b0;
      \piso.data_r_696_sv2v_reg  <= 1'b0;
      \piso.data_r_695_sv2v_reg  <= 1'b0;
      \piso.data_r_694_sv2v_reg  <= 1'b0;
      \piso.data_r_693_sv2v_reg  <= 1'b0;
      \piso.data_r_692_sv2v_reg  <= 1'b0;
      \piso.data_r_691_sv2v_reg  <= 1'b0;
      \piso.data_r_690_sv2v_reg  <= 1'b0;
      \piso.data_r_689_sv2v_reg  <= 1'b0;
      \piso.data_r_688_sv2v_reg  <= 1'b0;
      \piso.data_r_687_sv2v_reg  <= 1'b0;
      \piso.data_r_686_sv2v_reg  <= 1'b0;
      \piso.data_r_685_sv2v_reg  <= 1'b0;
      \piso.data_r_684_sv2v_reg  <= 1'b0;
      \piso.data_r_683_sv2v_reg  <= 1'b0;
      \piso.data_r_682_sv2v_reg  <= 1'b0;
      \piso.data_r_681_sv2v_reg  <= 1'b0;
      \piso.data_r_680_sv2v_reg  <= 1'b0;
      \piso.data_r_679_sv2v_reg  <= 1'b0;
      \piso.data_r_678_sv2v_reg  <= 1'b0;
      \piso.data_r_677_sv2v_reg  <= 1'b0;
      \piso.data_r_676_sv2v_reg  <= 1'b0;
      \piso.data_r_675_sv2v_reg  <= 1'b0;
      \piso.data_r_674_sv2v_reg  <= 1'b0;
      \piso.data_r_673_sv2v_reg  <= 1'b0;
      \piso.data_r_672_sv2v_reg  <= 1'b0;
      \piso.data_r_671_sv2v_reg  <= 1'b0;
      \piso.data_r_670_sv2v_reg  <= 1'b0;
      \piso.data_r_669_sv2v_reg  <= 1'b0;
      \piso.data_r_668_sv2v_reg  <= 1'b0;
      \piso.data_r_667_sv2v_reg  <= 1'b0;
      \piso.data_r_666_sv2v_reg  <= 1'b0;
      \piso.data_r_665_sv2v_reg  <= 1'b0;
      \piso.data_r_664_sv2v_reg  <= 1'b0;
      \piso.data_r_663_sv2v_reg  <= 1'b0;
      \piso.data_r_662_sv2v_reg  <= 1'b0;
      \piso.data_r_661_sv2v_reg  <= 1'b0;
      \piso.data_r_660_sv2v_reg  <= 1'b0;
      \piso.data_r_659_sv2v_reg  <= 1'b0;
      \piso.data_r_658_sv2v_reg  <= 1'b0;
      \piso.data_r_657_sv2v_reg  <= 1'b0;
      \piso.data_r_656_sv2v_reg  <= 1'b0;
      \piso.data_r_655_sv2v_reg  <= 1'b0;
      \piso.data_r_654_sv2v_reg  <= 1'b0;
      \piso.data_r_653_sv2v_reg  <= 1'b0;
      \piso.data_r_652_sv2v_reg  <= 1'b0;
      \piso.data_r_651_sv2v_reg  <= 1'b0;
      \piso.data_r_650_sv2v_reg  <= 1'b0;
      \piso.data_r_649_sv2v_reg  <= 1'b0;
      \piso.data_r_648_sv2v_reg  <= 1'b0;
      \piso.data_r_647_sv2v_reg  <= 1'b0;
      \piso.data_r_646_sv2v_reg  <= 1'b0;
      \piso.data_r_645_sv2v_reg  <= 1'b0;
      \piso.data_r_644_sv2v_reg  <= 1'b0;
      \piso.data_r_643_sv2v_reg  <= 1'b0;
      \piso.data_r_642_sv2v_reg  <= 1'b0;
      \piso.data_r_641_sv2v_reg  <= 1'b0;
      \piso.data_r_640_sv2v_reg  <= 1'b0;
      \piso.data_r_639_sv2v_reg  <= 1'b0;
      \piso.data_r_638_sv2v_reg  <= 1'b0;
      \piso.data_r_637_sv2v_reg  <= 1'b0;
      \piso.data_r_636_sv2v_reg  <= 1'b0;
      \piso.data_r_635_sv2v_reg  <= 1'b0;
      \piso.data_r_634_sv2v_reg  <= 1'b0;
      \piso.data_r_633_sv2v_reg  <= 1'b0;
      \piso.data_r_632_sv2v_reg  <= 1'b0;
      \piso.data_r_631_sv2v_reg  <= 1'b0;
      \piso.data_r_630_sv2v_reg  <= 1'b0;
      \piso.data_r_629_sv2v_reg  <= 1'b0;
      \piso.data_r_628_sv2v_reg  <= 1'b0;
      \piso.data_r_627_sv2v_reg  <= 1'b0;
      \piso.data_r_626_sv2v_reg  <= 1'b0;
      \piso.data_r_625_sv2v_reg  <= 1'b0;
      \piso.data_r_624_sv2v_reg  <= 1'b0;
      \piso.data_r_623_sv2v_reg  <= 1'b0;
      \piso.data_r_622_sv2v_reg  <= 1'b0;
      \piso.data_r_621_sv2v_reg  <= 1'b0;
      \piso.data_r_620_sv2v_reg  <= 1'b0;
      \piso.data_r_619_sv2v_reg  <= 1'b0;
      \piso.data_r_618_sv2v_reg  <= 1'b0;
      \piso.data_r_617_sv2v_reg  <= 1'b0;
      \piso.data_r_616_sv2v_reg  <= 1'b0;
      \piso.data_r_615_sv2v_reg  <= 1'b0;
      \piso.data_r_614_sv2v_reg  <= 1'b0;
      \piso.data_r_613_sv2v_reg  <= 1'b0;
      \piso.data_r_612_sv2v_reg  <= 1'b0;
      \piso.data_r_611_sv2v_reg  <= 1'b0;
      \piso.data_r_610_sv2v_reg  <= 1'b0;
      \piso.data_r_609_sv2v_reg  <= 1'b0;
      \piso.data_r_608_sv2v_reg  <= 1'b0;
      \piso.data_r_607_sv2v_reg  <= 1'b0;
      \piso.data_r_606_sv2v_reg  <= 1'b0;
      \piso.data_r_605_sv2v_reg  <= 1'b0;
      \piso.data_r_604_sv2v_reg  <= 1'b0;
      \piso.data_r_603_sv2v_reg  <= 1'b0;
      \piso.data_r_602_sv2v_reg  <= 1'b0;
      \piso.data_r_601_sv2v_reg  <= 1'b0;
      \piso.data_r_600_sv2v_reg  <= 1'b0;
      \piso.data_r_599_sv2v_reg  <= 1'b0;
      \piso.data_r_598_sv2v_reg  <= 1'b0;
      \piso.data_r_597_sv2v_reg  <= 1'b0;
      \piso.data_r_596_sv2v_reg  <= 1'b0;
      \piso.data_r_595_sv2v_reg  <= 1'b0;
      \piso.data_r_594_sv2v_reg  <= 1'b0;
      \piso.data_r_593_sv2v_reg  <= 1'b0;
      \piso.data_r_592_sv2v_reg  <= 1'b0;
      \piso.data_r_591_sv2v_reg  <= 1'b0;
      \piso.data_r_590_sv2v_reg  <= 1'b0;
      \piso.data_r_589_sv2v_reg  <= 1'b0;
      \piso.data_r_588_sv2v_reg  <= 1'b0;
      \piso.data_r_587_sv2v_reg  <= 1'b0;
      \piso.data_r_586_sv2v_reg  <= 1'b0;
      \piso.data_r_585_sv2v_reg  <= 1'b0;
      \piso.data_r_584_sv2v_reg  <= 1'b0;
      \piso.data_r_583_sv2v_reg  <= 1'b0;
      \piso.data_r_582_sv2v_reg  <= 1'b0;
      \piso.data_r_581_sv2v_reg  <= 1'b0;
      \piso.data_r_580_sv2v_reg  <= 1'b0;
      \piso.data_r_579_sv2v_reg  <= 1'b0;
      \piso.data_r_578_sv2v_reg  <= 1'b0;
      \piso.data_r_577_sv2v_reg  <= 1'b0;
      \piso.data_r_576_sv2v_reg  <= 1'b0;
      \piso.data_r_575_sv2v_reg  <= 1'b0;
      \piso.data_r_574_sv2v_reg  <= 1'b0;
      \piso.data_r_573_sv2v_reg  <= 1'b0;
      \piso.data_r_572_sv2v_reg  <= 1'b0;
      \piso.data_r_571_sv2v_reg  <= 1'b0;
      \piso.data_r_570_sv2v_reg  <= 1'b0;
      \piso.data_r_569_sv2v_reg  <= 1'b0;
      \piso.data_r_568_sv2v_reg  <= 1'b0;
      \piso.data_r_567_sv2v_reg  <= 1'b0;
      \piso.data_r_566_sv2v_reg  <= 1'b0;
      \piso.data_r_565_sv2v_reg  <= 1'b0;
      \piso.data_r_564_sv2v_reg  <= 1'b0;
      \piso.data_r_563_sv2v_reg  <= 1'b0;
      \piso.data_r_562_sv2v_reg  <= 1'b0;
      \piso.data_r_561_sv2v_reg  <= 1'b0;
      \piso.data_r_560_sv2v_reg  <= 1'b0;
      \piso.data_r_559_sv2v_reg  <= 1'b0;
      \piso.data_r_558_sv2v_reg  <= 1'b0;
      \piso.data_r_557_sv2v_reg  <= 1'b0;
      \piso.data_r_556_sv2v_reg  <= 1'b0;
      \piso.data_r_555_sv2v_reg  <= 1'b0;
      \piso.data_r_554_sv2v_reg  <= 1'b0;
      \piso.data_r_553_sv2v_reg  <= 1'b0;
      \piso.data_r_552_sv2v_reg  <= 1'b0;
      \piso.data_r_551_sv2v_reg  <= 1'b0;
      \piso.data_r_550_sv2v_reg  <= 1'b0;
      \piso.data_r_549_sv2v_reg  <= 1'b0;
      \piso.data_r_548_sv2v_reg  <= 1'b0;
      \piso.data_r_547_sv2v_reg  <= 1'b0;
      \piso.data_r_546_sv2v_reg  <= 1'b0;
      \piso.data_r_545_sv2v_reg  <= 1'b0;
      \piso.data_r_544_sv2v_reg  <= 1'b0;
      \piso.data_r_543_sv2v_reg  <= 1'b0;
      \piso.data_r_542_sv2v_reg  <= 1'b0;
      \piso.data_r_541_sv2v_reg  <= 1'b0;
      \piso.data_r_540_sv2v_reg  <= 1'b0;
      \piso.data_r_539_sv2v_reg  <= 1'b0;
      \piso.data_r_538_sv2v_reg  <= 1'b0;
      \piso.data_r_537_sv2v_reg  <= 1'b0;
      \piso.data_r_536_sv2v_reg  <= 1'b0;
      \piso.data_r_535_sv2v_reg  <= 1'b0;
      \piso.data_r_534_sv2v_reg  <= 1'b0;
      \piso.data_r_533_sv2v_reg  <= 1'b0;
      \piso.data_r_532_sv2v_reg  <= 1'b0;
      \piso.data_r_531_sv2v_reg  <= 1'b0;
      \piso.data_r_530_sv2v_reg  <= 1'b0;
      \piso.data_r_529_sv2v_reg  <= 1'b0;
      \piso.data_r_528_sv2v_reg  <= 1'b0;
      \piso.data_r_527_sv2v_reg  <= 1'b0;
      \piso.data_r_526_sv2v_reg  <= 1'b0;
      \piso.data_r_525_sv2v_reg  <= 1'b0;
      \piso.data_r_524_sv2v_reg  <= 1'b0;
      \piso.data_r_523_sv2v_reg  <= 1'b0;
      \piso.data_r_522_sv2v_reg  <= 1'b0;
      \piso.data_r_521_sv2v_reg  <= 1'b0;
      \piso.data_r_520_sv2v_reg  <= 1'b0;
      \piso.data_r_519_sv2v_reg  <= 1'b0;
      \piso.data_r_518_sv2v_reg  <= 1'b0;
      \piso.data_r_517_sv2v_reg  <= 1'b0;
      \piso.data_r_516_sv2v_reg  <= 1'b0;
      \piso.data_r_515_sv2v_reg  <= 1'b0;
      \piso.data_r_514_sv2v_reg  <= 1'b0;
      \piso.data_r_513_sv2v_reg  <= 1'b0;
      \piso.data_r_512_sv2v_reg  <= 1'b0;
      \piso.data_r_511_sv2v_reg  <= 1'b0;
      \piso.data_r_510_sv2v_reg  <= 1'b0;
      \piso.data_r_509_sv2v_reg  <= 1'b0;
      \piso.data_r_508_sv2v_reg  <= 1'b0;
      \piso.data_r_507_sv2v_reg  <= 1'b0;
      \piso.data_r_506_sv2v_reg  <= 1'b0;
      \piso.data_r_505_sv2v_reg  <= 1'b0;
      \piso.data_r_504_sv2v_reg  <= 1'b0;
      \piso.data_r_503_sv2v_reg  <= 1'b0;
      \piso.data_r_502_sv2v_reg  <= 1'b0;
      \piso.data_r_501_sv2v_reg  <= 1'b0;
      \piso.data_r_500_sv2v_reg  <= 1'b0;
      \piso.data_r_499_sv2v_reg  <= 1'b0;
      \piso.data_r_498_sv2v_reg  <= 1'b0;
      \piso.data_r_497_sv2v_reg  <= 1'b0;
      \piso.data_r_496_sv2v_reg  <= 1'b0;
      \piso.data_r_495_sv2v_reg  <= 1'b0;
      \piso.data_r_494_sv2v_reg  <= 1'b0;
      \piso.data_r_493_sv2v_reg  <= 1'b0;
      \piso.data_r_492_sv2v_reg  <= 1'b0;
      \piso.data_r_491_sv2v_reg  <= 1'b0;
      \piso.data_r_490_sv2v_reg  <= 1'b0;
      \piso.data_r_489_sv2v_reg  <= 1'b0;
      \piso.data_r_488_sv2v_reg  <= 1'b0;
      \piso.data_r_487_sv2v_reg  <= 1'b0;
      \piso.data_r_486_sv2v_reg  <= 1'b0;
      \piso.data_r_485_sv2v_reg  <= 1'b0;
      \piso.data_r_484_sv2v_reg  <= 1'b0;
      \piso.data_r_483_sv2v_reg  <= 1'b0;
      \piso.data_r_482_sv2v_reg  <= 1'b0;
      \piso.data_r_481_sv2v_reg  <= 1'b0;
      \piso.data_r_480_sv2v_reg  <= 1'b0;
      \piso.data_r_479_sv2v_reg  <= 1'b0;
      \piso.data_r_478_sv2v_reg  <= 1'b0;
      \piso.data_r_477_sv2v_reg  <= 1'b0;
      \piso.data_r_476_sv2v_reg  <= 1'b0;
      \piso.data_r_475_sv2v_reg  <= 1'b0;
      \piso.data_r_474_sv2v_reg  <= 1'b0;
      \piso.data_r_473_sv2v_reg  <= 1'b0;
      \piso.data_r_472_sv2v_reg  <= 1'b0;
      \piso.data_r_471_sv2v_reg  <= 1'b0;
      \piso.data_r_470_sv2v_reg  <= 1'b0;
      \piso.data_r_469_sv2v_reg  <= 1'b0;
      \piso.data_r_468_sv2v_reg  <= 1'b0;
      \piso.data_r_467_sv2v_reg  <= 1'b0;
      \piso.data_r_466_sv2v_reg  <= 1'b0;
      \piso.data_r_465_sv2v_reg  <= 1'b0;
      \piso.data_r_464_sv2v_reg  <= 1'b0;
      \piso.data_r_463_sv2v_reg  <= 1'b0;
      \piso.data_r_462_sv2v_reg  <= 1'b0;
      \piso.data_r_461_sv2v_reg  <= 1'b0;
      \piso.data_r_460_sv2v_reg  <= 1'b0;
      \piso.data_r_459_sv2v_reg  <= 1'b0;
      \piso.data_r_458_sv2v_reg  <= 1'b0;
      \piso.data_r_457_sv2v_reg  <= 1'b0;
      \piso.data_r_456_sv2v_reg  <= 1'b0;
      \piso.data_r_455_sv2v_reg  <= 1'b0;
      \piso.data_r_454_sv2v_reg  <= 1'b0;
      \piso.data_r_453_sv2v_reg  <= 1'b0;
      \piso.data_r_452_sv2v_reg  <= 1'b0;
      \piso.data_r_451_sv2v_reg  <= 1'b0;
      \piso.data_r_450_sv2v_reg  <= 1'b0;
      \piso.data_r_449_sv2v_reg  <= 1'b0;
      \piso.data_r_448_sv2v_reg  <= 1'b0;
      \piso.data_r_447_sv2v_reg  <= 1'b0;
      \piso.data_r_446_sv2v_reg  <= 1'b0;
      \piso.data_r_445_sv2v_reg  <= 1'b0;
      \piso.data_r_444_sv2v_reg  <= 1'b0;
      \piso.data_r_443_sv2v_reg  <= 1'b0;
      \piso.data_r_442_sv2v_reg  <= 1'b0;
      \piso.data_r_441_sv2v_reg  <= 1'b0;
      \piso.data_r_440_sv2v_reg  <= 1'b0;
      \piso.data_r_439_sv2v_reg  <= 1'b0;
      \piso.data_r_438_sv2v_reg  <= 1'b0;
      \piso.data_r_437_sv2v_reg  <= 1'b0;
      \piso.data_r_436_sv2v_reg  <= 1'b0;
      \piso.data_r_435_sv2v_reg  <= 1'b0;
      \piso.data_r_434_sv2v_reg  <= 1'b0;
      \piso.data_r_433_sv2v_reg  <= 1'b0;
      \piso.data_r_432_sv2v_reg  <= 1'b0;
      \piso.data_r_431_sv2v_reg  <= 1'b0;
      \piso.data_r_430_sv2v_reg  <= 1'b0;
      \piso.data_r_429_sv2v_reg  <= 1'b0;
      \piso.data_r_428_sv2v_reg  <= 1'b0;
      \piso.data_r_427_sv2v_reg  <= 1'b0;
      \piso.data_r_426_sv2v_reg  <= 1'b0;
      \piso.data_r_425_sv2v_reg  <= 1'b0;
      \piso.data_r_424_sv2v_reg  <= 1'b0;
      \piso.data_r_423_sv2v_reg  <= 1'b0;
      \piso.data_r_422_sv2v_reg  <= 1'b0;
      \piso.data_r_421_sv2v_reg  <= 1'b0;
      \piso.data_r_420_sv2v_reg  <= 1'b0;
      \piso.data_r_419_sv2v_reg  <= 1'b0;
      \piso.data_r_418_sv2v_reg  <= 1'b0;
      \piso.data_r_417_sv2v_reg  <= 1'b0;
      \piso.data_r_416_sv2v_reg  <= 1'b0;
      \piso.data_r_415_sv2v_reg  <= 1'b0;
      \piso.data_r_414_sv2v_reg  <= 1'b0;
      \piso.data_r_413_sv2v_reg  <= 1'b0;
      \piso.data_r_412_sv2v_reg  <= 1'b0;
      \piso.data_r_411_sv2v_reg  <= 1'b0;
      \piso.data_r_410_sv2v_reg  <= 1'b0;
      \piso.data_r_409_sv2v_reg  <= 1'b0;
      \piso.data_r_408_sv2v_reg  <= 1'b0;
      \piso.data_r_407_sv2v_reg  <= 1'b0;
      \piso.data_r_406_sv2v_reg  <= 1'b0;
      \piso.data_r_405_sv2v_reg  <= 1'b0;
      \piso.data_r_404_sv2v_reg  <= 1'b0;
      \piso.data_r_403_sv2v_reg  <= 1'b0;
      \piso.data_r_402_sv2v_reg  <= 1'b0;
      \piso.data_r_401_sv2v_reg  <= 1'b0;
      \piso.data_r_400_sv2v_reg  <= 1'b0;
      \piso.data_r_399_sv2v_reg  <= 1'b0;
      \piso.data_r_398_sv2v_reg  <= 1'b0;
      \piso.data_r_397_sv2v_reg  <= 1'b0;
      \piso.data_r_396_sv2v_reg  <= 1'b0;
      \piso.data_r_395_sv2v_reg  <= 1'b0;
      \piso.data_r_394_sv2v_reg  <= 1'b0;
      \piso.data_r_393_sv2v_reg  <= 1'b0;
      \piso.data_r_392_sv2v_reg  <= 1'b0;
      \piso.data_r_391_sv2v_reg  <= 1'b0;
      \piso.data_r_390_sv2v_reg  <= 1'b0;
      \piso.data_r_389_sv2v_reg  <= 1'b0;
      \piso.data_r_388_sv2v_reg  <= 1'b0;
      \piso.data_r_387_sv2v_reg  <= 1'b0;
      \piso.data_r_386_sv2v_reg  <= 1'b0;
      \piso.data_r_385_sv2v_reg  <= 1'b0;
      \piso.data_r_384_sv2v_reg  <= 1'b0;
      \piso.data_r_383_sv2v_reg  <= 1'b0;
      \piso.data_r_382_sv2v_reg  <= 1'b0;
      \piso.data_r_381_sv2v_reg  <= 1'b0;
      \piso.data_r_380_sv2v_reg  <= 1'b0;
      \piso.data_r_379_sv2v_reg  <= 1'b0;
      \piso.data_r_378_sv2v_reg  <= 1'b0;
      \piso.data_r_377_sv2v_reg  <= 1'b0;
      \piso.data_r_376_sv2v_reg  <= 1'b0;
      \piso.data_r_375_sv2v_reg  <= 1'b0;
      \piso.data_r_374_sv2v_reg  <= 1'b0;
      \piso.data_r_373_sv2v_reg  <= 1'b0;
      \piso.data_r_372_sv2v_reg  <= 1'b0;
      \piso.data_r_371_sv2v_reg  <= 1'b0;
      \piso.data_r_370_sv2v_reg  <= 1'b0;
      \piso.data_r_369_sv2v_reg  <= 1'b0;
      \piso.data_r_368_sv2v_reg  <= 1'b0;
      \piso.data_r_367_sv2v_reg  <= 1'b0;
      \piso.data_r_366_sv2v_reg  <= 1'b0;
      \piso.data_r_365_sv2v_reg  <= 1'b0;
      \piso.data_r_364_sv2v_reg  <= 1'b0;
      \piso.data_r_363_sv2v_reg  <= 1'b0;
      \piso.data_r_362_sv2v_reg  <= 1'b0;
      \piso.data_r_361_sv2v_reg  <= 1'b0;
      \piso.data_r_360_sv2v_reg  <= 1'b0;
      \piso.data_r_359_sv2v_reg  <= 1'b0;
      \piso.data_r_358_sv2v_reg  <= 1'b0;
      \piso.data_r_357_sv2v_reg  <= 1'b0;
      \piso.data_r_356_sv2v_reg  <= 1'b0;
      \piso.data_r_355_sv2v_reg  <= 1'b0;
      \piso.data_r_354_sv2v_reg  <= 1'b0;
      \piso.data_r_353_sv2v_reg  <= 1'b0;
      \piso.data_r_352_sv2v_reg  <= 1'b0;
      \piso.data_r_351_sv2v_reg  <= 1'b0;
      \piso.data_r_350_sv2v_reg  <= 1'b0;
      \piso.data_r_349_sv2v_reg  <= 1'b0;
      \piso.data_r_348_sv2v_reg  <= 1'b0;
      \piso.data_r_347_sv2v_reg  <= 1'b0;
      \piso.data_r_346_sv2v_reg  <= 1'b0;
      \piso.data_r_345_sv2v_reg  <= 1'b0;
      \piso.data_r_344_sv2v_reg  <= 1'b0;
      \piso.data_r_343_sv2v_reg  <= 1'b0;
      \piso.data_r_342_sv2v_reg  <= 1'b0;
      \piso.data_r_341_sv2v_reg  <= 1'b0;
      \piso.data_r_340_sv2v_reg  <= 1'b0;
      \piso.data_r_339_sv2v_reg  <= 1'b0;
      \piso.data_r_338_sv2v_reg  <= 1'b0;
      \piso.data_r_337_sv2v_reg  <= 1'b0;
      \piso.data_r_336_sv2v_reg  <= 1'b0;
      \piso.data_r_335_sv2v_reg  <= 1'b0;
      \piso.data_r_334_sv2v_reg  <= 1'b0;
      \piso.data_r_333_sv2v_reg  <= 1'b0;
      \piso.data_r_332_sv2v_reg  <= 1'b0;
      \piso.data_r_331_sv2v_reg  <= 1'b0;
      \piso.data_r_330_sv2v_reg  <= 1'b0;
      \piso.data_r_329_sv2v_reg  <= 1'b0;
      \piso.data_r_328_sv2v_reg  <= 1'b0;
      \piso.data_r_327_sv2v_reg  <= 1'b0;
      \piso.data_r_326_sv2v_reg  <= 1'b0;
      \piso.data_r_325_sv2v_reg  <= 1'b0;
      \piso.data_r_324_sv2v_reg  <= 1'b0;
      \piso.data_r_323_sv2v_reg  <= 1'b0;
      \piso.data_r_322_sv2v_reg  <= 1'b0;
      \piso.data_r_321_sv2v_reg  <= 1'b0;
      \piso.data_r_320_sv2v_reg  <= 1'b0;
      \piso.data_r_319_sv2v_reg  <= 1'b0;
      \piso.data_r_318_sv2v_reg  <= 1'b0;
      \piso.data_r_317_sv2v_reg  <= 1'b0;
      \piso.data_r_316_sv2v_reg  <= 1'b0;
      \piso.data_r_315_sv2v_reg  <= 1'b0;
      \piso.data_r_314_sv2v_reg  <= 1'b0;
      \piso.data_r_313_sv2v_reg  <= 1'b0;
      \piso.data_r_312_sv2v_reg  <= 1'b0;
      \piso.data_r_311_sv2v_reg  <= 1'b0;
      \piso.data_r_310_sv2v_reg  <= 1'b0;
      \piso.data_r_309_sv2v_reg  <= 1'b0;
      \piso.data_r_308_sv2v_reg  <= 1'b0;
      \piso.data_r_307_sv2v_reg  <= 1'b0;
      \piso.data_r_306_sv2v_reg  <= 1'b0;
      \piso.data_r_305_sv2v_reg  <= 1'b0;
      \piso.data_r_304_sv2v_reg  <= 1'b0;
      \piso.data_r_303_sv2v_reg  <= 1'b0;
      \piso.data_r_302_sv2v_reg  <= 1'b0;
      \piso.data_r_301_sv2v_reg  <= 1'b0;
      \piso.data_r_300_sv2v_reg  <= 1'b0;
      \piso.data_r_299_sv2v_reg  <= 1'b0;
      \piso.data_r_298_sv2v_reg  <= 1'b0;
      \piso.data_r_297_sv2v_reg  <= 1'b0;
      \piso.data_r_296_sv2v_reg  <= 1'b0;
      \piso.data_r_295_sv2v_reg  <= 1'b0;
      \piso.data_r_294_sv2v_reg  <= 1'b0;
      \piso.data_r_293_sv2v_reg  <= 1'b0;
      \piso.data_r_292_sv2v_reg  <= 1'b0;
      \piso.data_r_291_sv2v_reg  <= 1'b0;
      \piso.data_r_290_sv2v_reg  <= 1'b0;
      \piso.data_r_289_sv2v_reg  <= 1'b0;
      \piso.data_r_288_sv2v_reg  <= 1'b0;
      \piso.data_r_287_sv2v_reg  <= 1'b0;
      \piso.data_r_286_sv2v_reg  <= 1'b0;
      \piso.data_r_285_sv2v_reg  <= 1'b0;
      \piso.data_r_284_sv2v_reg  <= 1'b0;
      \piso.data_r_283_sv2v_reg  <= 1'b0;
      \piso.data_r_282_sv2v_reg  <= 1'b0;
      \piso.data_r_281_sv2v_reg  <= 1'b0;
      \piso.data_r_280_sv2v_reg  <= 1'b0;
      \piso.data_r_279_sv2v_reg  <= 1'b0;
      \piso.data_r_278_sv2v_reg  <= 1'b0;
      \piso.data_r_277_sv2v_reg  <= 1'b0;
      \piso.data_r_276_sv2v_reg  <= 1'b0;
      \piso.data_r_275_sv2v_reg  <= 1'b0;
      \piso.data_r_274_sv2v_reg  <= 1'b0;
      \piso.data_r_273_sv2v_reg  <= 1'b0;
      \piso.data_r_272_sv2v_reg  <= 1'b0;
      \piso.data_r_271_sv2v_reg  <= 1'b0;
      \piso.data_r_270_sv2v_reg  <= 1'b0;
      \piso.data_r_269_sv2v_reg  <= 1'b0;
      \piso.data_r_268_sv2v_reg  <= 1'b0;
      \piso.data_r_267_sv2v_reg  <= 1'b0;
      \piso.data_r_266_sv2v_reg  <= 1'b0;
      \piso.data_r_265_sv2v_reg  <= 1'b0;
      \piso.data_r_264_sv2v_reg  <= 1'b0;
      \piso.data_r_263_sv2v_reg  <= 1'b0;
      \piso.data_r_262_sv2v_reg  <= 1'b0;
      \piso.data_r_261_sv2v_reg  <= 1'b0;
      \piso.data_r_260_sv2v_reg  <= 1'b0;
      \piso.data_r_259_sv2v_reg  <= 1'b0;
      \piso.data_r_258_sv2v_reg  <= 1'b0;
      \piso.data_r_257_sv2v_reg  <= 1'b0;
      \piso.data_r_256_sv2v_reg  <= 1'b0;
      \piso.data_r_255_sv2v_reg  <= 1'b0;
      \piso.data_r_254_sv2v_reg  <= 1'b0;
      \piso.data_r_253_sv2v_reg  <= 1'b0;
      \piso.data_r_252_sv2v_reg  <= 1'b0;
      \piso.data_r_251_sv2v_reg  <= 1'b0;
      \piso.data_r_250_sv2v_reg  <= 1'b0;
      \piso.data_r_249_sv2v_reg  <= 1'b0;
      \piso.data_r_248_sv2v_reg  <= 1'b0;
      \piso.data_r_247_sv2v_reg  <= 1'b0;
      \piso.data_r_246_sv2v_reg  <= 1'b0;
      \piso.data_r_245_sv2v_reg  <= 1'b0;
      \piso.data_r_244_sv2v_reg  <= 1'b0;
      \piso.data_r_243_sv2v_reg  <= 1'b0;
      \piso.data_r_242_sv2v_reg  <= 1'b0;
      \piso.data_r_241_sv2v_reg  <= 1'b0;
      \piso.data_r_240_sv2v_reg  <= 1'b0;
      \piso.data_r_239_sv2v_reg  <= 1'b0;
      \piso.data_r_238_sv2v_reg  <= 1'b0;
      \piso.data_r_237_sv2v_reg  <= 1'b0;
      \piso.data_r_236_sv2v_reg  <= 1'b0;
      \piso.data_r_235_sv2v_reg  <= 1'b0;
      \piso.data_r_234_sv2v_reg  <= 1'b0;
      \piso.data_r_233_sv2v_reg  <= 1'b0;
      \piso.data_r_232_sv2v_reg  <= 1'b0;
      \piso.data_r_231_sv2v_reg  <= 1'b0;
      \piso.data_r_230_sv2v_reg  <= 1'b0;
      \piso.data_r_229_sv2v_reg  <= 1'b0;
      \piso.data_r_228_sv2v_reg  <= 1'b0;
      \piso.data_r_227_sv2v_reg  <= 1'b0;
      \piso.data_r_226_sv2v_reg  <= 1'b0;
      \piso.data_r_225_sv2v_reg  <= 1'b0;
      \piso.data_r_224_sv2v_reg  <= 1'b0;
      \piso.data_r_223_sv2v_reg  <= 1'b0;
      \piso.data_r_222_sv2v_reg  <= 1'b0;
      \piso.data_r_221_sv2v_reg  <= 1'b0;
      \piso.data_r_220_sv2v_reg  <= 1'b0;
      \piso.data_r_219_sv2v_reg  <= 1'b0;
      \piso.data_r_218_sv2v_reg  <= 1'b0;
      \piso.data_r_217_sv2v_reg  <= 1'b0;
      \piso.data_r_216_sv2v_reg  <= 1'b0;
      \piso.data_r_215_sv2v_reg  <= 1'b0;
      \piso.data_r_214_sv2v_reg  <= 1'b0;
      \piso.data_r_213_sv2v_reg  <= 1'b0;
      \piso.data_r_212_sv2v_reg  <= 1'b0;
      \piso.data_r_211_sv2v_reg  <= 1'b0;
      \piso.data_r_210_sv2v_reg  <= 1'b0;
      \piso.data_r_209_sv2v_reg  <= 1'b0;
      \piso.data_r_208_sv2v_reg  <= 1'b0;
      \piso.data_r_207_sv2v_reg  <= 1'b0;
      \piso.data_r_206_sv2v_reg  <= 1'b0;
      \piso.data_r_205_sv2v_reg  <= 1'b0;
      \piso.data_r_204_sv2v_reg  <= 1'b0;
      \piso.data_r_203_sv2v_reg  <= 1'b0;
      \piso.data_r_202_sv2v_reg  <= 1'b0;
      \piso.data_r_201_sv2v_reg  <= 1'b0;
      \piso.data_r_200_sv2v_reg  <= 1'b0;
      \piso.data_r_199_sv2v_reg  <= 1'b0;
      \piso.data_r_198_sv2v_reg  <= 1'b0;
      \piso.data_r_197_sv2v_reg  <= 1'b0;
      \piso.data_r_196_sv2v_reg  <= 1'b0;
      \piso.data_r_195_sv2v_reg  <= 1'b0;
      \piso.data_r_194_sv2v_reg  <= 1'b0;
      \piso.data_r_193_sv2v_reg  <= 1'b0;
      \piso.data_r_192_sv2v_reg  <= 1'b0;
      \piso.data_r_191_sv2v_reg  <= 1'b0;
      \piso.data_r_190_sv2v_reg  <= 1'b0;
      \piso.data_r_189_sv2v_reg  <= 1'b0;
      \piso.data_r_188_sv2v_reg  <= 1'b0;
      \piso.data_r_187_sv2v_reg  <= 1'b0;
      \piso.data_r_186_sv2v_reg  <= 1'b0;
      \piso.data_r_185_sv2v_reg  <= 1'b0;
      \piso.data_r_184_sv2v_reg  <= 1'b0;
      \piso.data_r_183_sv2v_reg  <= 1'b0;
      \piso.data_r_182_sv2v_reg  <= 1'b0;
      \piso.data_r_181_sv2v_reg  <= 1'b0;
      \piso.data_r_180_sv2v_reg  <= 1'b0;
      \piso.data_r_179_sv2v_reg  <= 1'b0;
      \piso.data_r_178_sv2v_reg  <= 1'b0;
      \piso.data_r_177_sv2v_reg  <= 1'b0;
      \piso.data_r_176_sv2v_reg  <= 1'b0;
      \piso.data_r_175_sv2v_reg  <= 1'b0;
      \piso.data_r_174_sv2v_reg  <= 1'b0;
      \piso.data_r_173_sv2v_reg  <= 1'b0;
      \piso.data_r_172_sv2v_reg  <= 1'b0;
      \piso.data_r_171_sv2v_reg  <= 1'b0;
      \piso.data_r_170_sv2v_reg  <= 1'b0;
      \piso.data_r_169_sv2v_reg  <= 1'b0;
      \piso.data_r_168_sv2v_reg  <= 1'b0;
      \piso.data_r_167_sv2v_reg  <= 1'b0;
      \piso.data_r_166_sv2v_reg  <= 1'b0;
      \piso.data_r_165_sv2v_reg  <= 1'b0;
      \piso.data_r_164_sv2v_reg  <= 1'b0;
      \piso.data_r_163_sv2v_reg  <= 1'b0;
      \piso.data_r_162_sv2v_reg  <= 1'b0;
      \piso.data_r_161_sv2v_reg  <= 1'b0;
      \piso.data_r_160_sv2v_reg  <= 1'b0;
      \piso.data_r_159_sv2v_reg  <= 1'b0;
      \piso.data_r_158_sv2v_reg  <= 1'b0;
      \piso.data_r_157_sv2v_reg  <= 1'b0;
      \piso.data_r_156_sv2v_reg  <= 1'b0;
      \piso.data_r_155_sv2v_reg  <= 1'b0;
      \piso.data_r_154_sv2v_reg  <= 1'b0;
      \piso.data_r_153_sv2v_reg  <= 1'b0;
      \piso.data_r_152_sv2v_reg  <= 1'b0;
      \piso.data_r_151_sv2v_reg  <= 1'b0;
      \piso.data_r_150_sv2v_reg  <= 1'b0;
      \piso.data_r_149_sv2v_reg  <= 1'b0;
      \piso.data_r_148_sv2v_reg  <= 1'b0;
      \piso.data_r_147_sv2v_reg  <= 1'b0;
      \piso.data_r_146_sv2v_reg  <= 1'b0;
      \piso.data_r_145_sv2v_reg  <= 1'b0;
      \piso.data_r_144_sv2v_reg  <= 1'b0;
      \piso.data_r_143_sv2v_reg  <= 1'b0;
      \piso.data_r_142_sv2v_reg  <= 1'b0;
      \piso.data_r_141_sv2v_reg  <= 1'b0;
      \piso.data_r_140_sv2v_reg  <= 1'b0;
      \piso.data_r_139_sv2v_reg  <= 1'b0;
      \piso.data_r_138_sv2v_reg  <= 1'b0;
      \piso.data_r_137_sv2v_reg  <= 1'b0;
      \piso.data_r_136_sv2v_reg  <= 1'b0;
      \piso.data_r_135_sv2v_reg  <= 1'b0;
      \piso.data_r_134_sv2v_reg  <= 1'b0;
      \piso.data_r_133_sv2v_reg  <= 1'b0;
      \piso.data_r_132_sv2v_reg  <= 1'b0;
      \piso.data_r_131_sv2v_reg  <= 1'b0;
      \piso.data_r_130_sv2v_reg  <= 1'b0;
      \piso.data_r_129_sv2v_reg  <= 1'b0;
      \piso.data_r_128_sv2v_reg  <= 1'b0;
      \piso.data_r_127_sv2v_reg  <= 1'b0;
      \piso.data_r_126_sv2v_reg  <= 1'b0;
      \piso.data_r_125_sv2v_reg  <= 1'b0;
      \piso.data_r_124_sv2v_reg  <= 1'b0;
      \piso.data_r_123_sv2v_reg  <= 1'b0;
      \piso.data_r_122_sv2v_reg  <= 1'b0;
      \piso.data_r_121_sv2v_reg  <= 1'b0;
      \piso.data_r_120_sv2v_reg  <= 1'b0;
      \piso.data_r_119_sv2v_reg  <= 1'b0;
      \piso.data_r_118_sv2v_reg  <= 1'b0;
      \piso.data_r_117_sv2v_reg  <= 1'b0;
      \piso.data_r_116_sv2v_reg  <= 1'b0;
      \piso.data_r_115_sv2v_reg  <= 1'b0;
      \piso.data_r_114_sv2v_reg  <= 1'b0;
      \piso.data_r_113_sv2v_reg  <= 1'b0;
      \piso.data_r_112_sv2v_reg  <= 1'b0;
      \piso.data_r_111_sv2v_reg  <= 1'b0;
      \piso.data_r_110_sv2v_reg  <= 1'b0;
      \piso.data_r_109_sv2v_reg  <= 1'b0;
      \piso.data_r_108_sv2v_reg  <= 1'b0;
      \piso.data_r_107_sv2v_reg  <= 1'b0;
      \piso.data_r_106_sv2v_reg  <= 1'b0;
      \piso.data_r_105_sv2v_reg  <= 1'b0;
      \piso.data_r_104_sv2v_reg  <= 1'b0;
      \piso.data_r_103_sv2v_reg  <= 1'b0;
      \piso.data_r_102_sv2v_reg  <= 1'b0;
      \piso.data_r_101_sv2v_reg  <= 1'b0;
      \piso.data_r_100_sv2v_reg  <= 1'b0;
      \piso.data_r_99_sv2v_reg  <= 1'b0;
      \piso.data_r_98_sv2v_reg  <= 1'b0;
      \piso.data_r_97_sv2v_reg  <= 1'b0;
      \piso.data_r_96_sv2v_reg  <= 1'b0;
      \piso.data_r_95_sv2v_reg  <= 1'b0;
      \piso.data_r_94_sv2v_reg  <= 1'b0;
      \piso.data_r_93_sv2v_reg  <= 1'b0;
      \piso.data_r_92_sv2v_reg  <= 1'b0;
      \piso.data_r_91_sv2v_reg  <= 1'b0;
      \piso.data_r_90_sv2v_reg  <= 1'b0;
      \piso.data_r_89_sv2v_reg  <= 1'b0;
      \piso.data_r_88_sv2v_reg  <= 1'b0;
      \piso.data_r_87_sv2v_reg  <= 1'b0;
      \piso.data_r_86_sv2v_reg  <= 1'b0;
      \piso.data_r_85_sv2v_reg  <= 1'b0;
      \piso.data_r_84_sv2v_reg  <= 1'b0;
      \piso.data_r_83_sv2v_reg  <= 1'b0;
      \piso.data_r_82_sv2v_reg  <= 1'b0;
      \piso.data_r_81_sv2v_reg  <= 1'b0;
      \piso.data_r_80_sv2v_reg  <= 1'b0;
      \piso.data_r_79_sv2v_reg  <= 1'b0;
      \piso.data_r_78_sv2v_reg  <= 1'b0;
      \piso.data_r_77_sv2v_reg  <= 1'b0;
      \piso.data_r_76_sv2v_reg  <= 1'b0;
      \piso.data_r_75_sv2v_reg  <= 1'b0;
      \piso.data_r_74_sv2v_reg  <= 1'b0;
      \piso.data_r_73_sv2v_reg  <= 1'b0;
      \piso.data_r_72_sv2v_reg  <= 1'b0;
      \piso.data_r_71_sv2v_reg  <= 1'b0;
      \piso.data_r_70_sv2v_reg  <= 1'b0;
      \piso.data_r_69_sv2v_reg  <= 1'b0;
      \piso.data_r_68_sv2v_reg  <= 1'b0;
      \piso.data_r_67_sv2v_reg  <= 1'b0;
      \piso.data_r_66_sv2v_reg  <= 1'b0;
      \piso.data_r_65_sv2v_reg  <= 1'b0;
      \piso.data_r_64_sv2v_reg  <= 1'b0;
      \piso.data_r_63_sv2v_reg  <= 1'b0;
      \piso.data_r_62_sv2v_reg  <= 1'b0;
      \piso.data_r_61_sv2v_reg  <= 1'b0;
      \piso.data_r_60_sv2v_reg  <= 1'b0;
      \piso.data_r_59_sv2v_reg  <= 1'b0;
      \piso.data_r_58_sv2v_reg  <= 1'b0;
      \piso.data_r_57_sv2v_reg  <= 1'b0;
      \piso.data_r_56_sv2v_reg  <= 1'b0;
      \piso.data_r_55_sv2v_reg  <= 1'b0;
      \piso.data_r_54_sv2v_reg  <= 1'b0;
      \piso.data_r_53_sv2v_reg  <= 1'b0;
      \piso.data_r_52_sv2v_reg  <= 1'b0;
      \piso.data_r_51_sv2v_reg  <= 1'b0;
      \piso.data_r_50_sv2v_reg  <= 1'b0;
      \piso.data_r_49_sv2v_reg  <= 1'b0;
      \piso.data_r_48_sv2v_reg  <= 1'b0;
      \piso.data_r_47_sv2v_reg  <= 1'b0;
      \piso.data_r_46_sv2v_reg  <= 1'b0;
      \piso.data_r_45_sv2v_reg  <= 1'b0;
      \piso.data_r_44_sv2v_reg  <= 1'b0;
      \piso.data_r_43_sv2v_reg  <= 1'b0;
      \piso.data_r_42_sv2v_reg  <= 1'b0;
      \piso.data_r_41_sv2v_reg  <= 1'b0;
      \piso.data_r_40_sv2v_reg  <= 1'b0;
      \piso.data_r_39_sv2v_reg  <= 1'b0;
      \piso.data_r_38_sv2v_reg  <= 1'b0;
      \piso.data_r_37_sv2v_reg  <= 1'b0;
      \piso.data_r_36_sv2v_reg  <= 1'b0;
      \piso.data_r_35_sv2v_reg  <= 1'b0;
      \piso.data_r_34_sv2v_reg  <= 1'b0;
      \piso.data_r_33_sv2v_reg  <= 1'b0;
      \piso.data_r_32_sv2v_reg  <= 1'b0;
      \piso.data_r_31_sv2v_reg  <= 1'b0;
      \piso.data_r_30_sv2v_reg  <= 1'b0;
      \piso.data_r_29_sv2v_reg  <= 1'b0;
      \piso.data_r_28_sv2v_reg  <= 1'b0;
      \piso.data_r_27_sv2v_reg  <= 1'b0;
      \piso.data_r_26_sv2v_reg  <= 1'b0;
      \piso.data_r_25_sv2v_reg  <= 1'b0;
      \piso.data_r_24_sv2v_reg  <= 1'b0;
      \piso.data_r_23_sv2v_reg  <= 1'b0;
      \piso.data_r_22_sv2v_reg  <= 1'b0;
      \piso.data_r_21_sv2v_reg  <= 1'b0;
      \piso.data_r_20_sv2v_reg  <= 1'b0;
      \piso.data_r_19_sv2v_reg  <= 1'b0;
      \piso.data_r_18_sv2v_reg  <= 1'b0;
      \piso.data_r_17_sv2v_reg  <= 1'b0;
      \piso.data_r_16_sv2v_reg  <= 1'b0;
      \piso.data_r_15_sv2v_reg  <= 1'b0;
      \piso.data_r_14_sv2v_reg  <= 1'b0;
      \piso.data_r_13_sv2v_reg  <= 1'b0;
      \piso.data_r_12_sv2v_reg  <= 1'b0;
      \piso.data_r_11_sv2v_reg  <= 1'b0;
      \piso.data_r_10_sv2v_reg  <= 1'b0;
      \piso.data_r_9_sv2v_reg  <= 1'b0;
      \piso.data_r_8_sv2v_reg  <= 1'b0;
      \piso.data_r_7_sv2v_reg  <= 1'b0;
      \piso.data_r_6_sv2v_reg  <= 1'b0;
      \piso.data_r_5_sv2v_reg  <= 1'b0;
      \piso.data_r_4_sv2v_reg  <= 1'b0;
      \piso.data_r_3_sv2v_reg  <= 1'b0;
      \piso.data_r_2_sv2v_reg  <= 1'b0;
      \piso.data_r_1_sv2v_reg  <= 1'b0;
      \piso.data_r_0_sv2v_reg  <= 1'b0;
    end else if(N6) begin
      \piso.data_r_4095_sv2v_reg  <= \piso.data_li [4095];
      \piso.data_r_4094_sv2v_reg  <= \piso.data_li [4094];
      \piso.data_r_4093_sv2v_reg  <= \piso.data_li [4093];
      \piso.data_r_4092_sv2v_reg  <= \piso.data_li [4092];
      \piso.data_r_4091_sv2v_reg  <= \piso.data_li [4091];
      \piso.data_r_4090_sv2v_reg  <= \piso.data_li [4090];
      \piso.data_r_4089_sv2v_reg  <= \piso.data_li [4089];
      \piso.data_r_4088_sv2v_reg  <= \piso.data_li [4088];
      \piso.data_r_4087_sv2v_reg  <= \piso.data_li [4087];
      \piso.data_r_4086_sv2v_reg  <= \piso.data_li [4086];
      \piso.data_r_4085_sv2v_reg  <= \piso.data_li [4085];
      \piso.data_r_4084_sv2v_reg  <= \piso.data_li [4084];
      \piso.data_r_4083_sv2v_reg  <= \piso.data_li [4083];
      \piso.data_r_4082_sv2v_reg  <= \piso.data_li [4082];
      \piso.data_r_4081_sv2v_reg  <= \piso.data_li [4081];
      \piso.data_r_4080_sv2v_reg  <= \piso.data_li [4080];
      \piso.data_r_4079_sv2v_reg  <= \piso.data_li [4079];
      \piso.data_r_4078_sv2v_reg  <= \piso.data_li [4078];
      \piso.data_r_4077_sv2v_reg  <= \piso.data_li [4077];
      \piso.data_r_4076_sv2v_reg  <= \piso.data_li [4076];
      \piso.data_r_4075_sv2v_reg  <= \piso.data_li [4075];
      \piso.data_r_4074_sv2v_reg  <= \piso.data_li [4074];
      \piso.data_r_4073_sv2v_reg  <= \piso.data_li [4073];
      \piso.data_r_4072_sv2v_reg  <= \piso.data_li [4072];
      \piso.data_r_4071_sv2v_reg  <= \piso.data_li [4071];
      \piso.data_r_4070_sv2v_reg  <= \piso.data_li [4070];
      \piso.data_r_4069_sv2v_reg  <= \piso.data_li [4069];
      \piso.data_r_4068_sv2v_reg  <= \piso.data_li [4068];
      \piso.data_r_4067_sv2v_reg  <= \piso.data_li [4067];
      \piso.data_r_4066_sv2v_reg  <= \piso.data_li [4066];
      \piso.data_r_4065_sv2v_reg  <= \piso.data_li [4065];
      \piso.data_r_4064_sv2v_reg  <= \piso.data_li [4064];
      \piso.data_r_4063_sv2v_reg  <= \piso.data_li [4063];
      \piso.data_r_4062_sv2v_reg  <= \piso.data_li [4062];
      \piso.data_r_4061_sv2v_reg  <= \piso.data_li [4061];
      \piso.data_r_4060_sv2v_reg  <= \piso.data_li [4060];
      \piso.data_r_4059_sv2v_reg  <= \piso.data_li [4059];
      \piso.data_r_4058_sv2v_reg  <= \piso.data_li [4058];
      \piso.data_r_4057_sv2v_reg  <= \piso.data_li [4057];
      \piso.data_r_4056_sv2v_reg  <= \piso.data_li [4056];
      \piso.data_r_4055_sv2v_reg  <= \piso.data_li [4055];
      \piso.data_r_4054_sv2v_reg  <= \piso.data_li [4054];
      \piso.data_r_4053_sv2v_reg  <= \piso.data_li [4053];
      \piso.data_r_4052_sv2v_reg  <= \piso.data_li [4052];
      \piso.data_r_4051_sv2v_reg  <= \piso.data_li [4051];
      \piso.data_r_4050_sv2v_reg  <= \piso.data_li [4050];
      \piso.data_r_4049_sv2v_reg  <= \piso.data_li [4049];
      \piso.data_r_4048_sv2v_reg  <= \piso.data_li [4048];
      \piso.data_r_4047_sv2v_reg  <= \piso.data_li [4047];
      \piso.data_r_4046_sv2v_reg  <= \piso.data_li [4046];
      \piso.data_r_4045_sv2v_reg  <= \piso.data_li [4045];
      \piso.data_r_4044_sv2v_reg  <= \piso.data_li [4044];
      \piso.data_r_4043_sv2v_reg  <= \piso.data_li [4043];
      \piso.data_r_4042_sv2v_reg  <= \piso.data_li [4042];
      \piso.data_r_4041_sv2v_reg  <= \piso.data_li [4041];
      \piso.data_r_4040_sv2v_reg  <= \piso.data_li [4040];
      \piso.data_r_4039_sv2v_reg  <= \piso.data_li [4039];
      \piso.data_r_4038_sv2v_reg  <= \piso.data_li [4038];
      \piso.data_r_4037_sv2v_reg  <= \piso.data_li [4037];
      \piso.data_r_4036_sv2v_reg  <= \piso.data_li [4036];
      \piso.data_r_4035_sv2v_reg  <= \piso.data_li [4035];
      \piso.data_r_4034_sv2v_reg  <= \piso.data_li [4034];
      \piso.data_r_4033_sv2v_reg  <= \piso.data_li [4033];
      \piso.data_r_4032_sv2v_reg  <= \piso.data_li [4032];
      \piso.data_r_4031_sv2v_reg  <= \piso.data_li [4031];
      \piso.data_r_4030_sv2v_reg  <= \piso.data_li [4030];
      \piso.data_r_4029_sv2v_reg  <= \piso.data_li [4029];
      \piso.data_r_4028_sv2v_reg  <= \piso.data_li [4028];
      \piso.data_r_4027_sv2v_reg  <= \piso.data_li [4027];
      \piso.data_r_4026_sv2v_reg  <= \piso.data_li [4026];
      \piso.data_r_4025_sv2v_reg  <= \piso.data_li [4025];
      \piso.data_r_4024_sv2v_reg  <= \piso.data_li [4024];
      \piso.data_r_4023_sv2v_reg  <= \piso.data_li [4023];
      \piso.data_r_4022_sv2v_reg  <= \piso.data_li [4022];
      \piso.data_r_4021_sv2v_reg  <= \piso.data_li [4021];
      \piso.data_r_4020_sv2v_reg  <= \piso.data_li [4020];
      \piso.data_r_4019_sv2v_reg  <= \piso.data_li [4019];
      \piso.data_r_4018_sv2v_reg  <= \piso.data_li [4018];
      \piso.data_r_4017_sv2v_reg  <= \piso.data_li [4017];
      \piso.data_r_4016_sv2v_reg  <= \piso.data_li [4016];
      \piso.data_r_4015_sv2v_reg  <= \piso.data_li [4015];
      \piso.data_r_4014_sv2v_reg  <= \piso.data_li [4014];
      \piso.data_r_4013_sv2v_reg  <= \piso.data_li [4013];
      \piso.data_r_4012_sv2v_reg  <= \piso.data_li [4012];
      \piso.data_r_4011_sv2v_reg  <= \piso.data_li [4011];
      \piso.data_r_4010_sv2v_reg  <= \piso.data_li [4010];
      \piso.data_r_4009_sv2v_reg  <= \piso.data_li [4009];
      \piso.data_r_4008_sv2v_reg  <= \piso.data_li [4008];
      \piso.data_r_4007_sv2v_reg  <= \piso.data_li [4007];
      \piso.data_r_4006_sv2v_reg  <= \piso.data_li [4006];
      \piso.data_r_4005_sv2v_reg  <= \piso.data_li [4005];
      \piso.data_r_4004_sv2v_reg  <= \piso.data_li [4004];
      \piso.data_r_4003_sv2v_reg  <= \piso.data_li [4003];
      \piso.data_r_4002_sv2v_reg  <= \piso.data_li [4002];
      \piso.data_r_4001_sv2v_reg  <= \piso.data_li [4001];
      \piso.data_r_4000_sv2v_reg  <= \piso.data_li [4000];
      \piso.data_r_3999_sv2v_reg  <= \piso.data_li [3999];
      \piso.data_r_3998_sv2v_reg  <= \piso.data_li [3998];
      \piso.data_r_3997_sv2v_reg  <= \piso.data_li [3997];
      \piso.data_r_3996_sv2v_reg  <= \piso.data_li [3996];
      \piso.data_r_3995_sv2v_reg  <= \piso.data_li [3995];
      \piso.data_r_3994_sv2v_reg  <= \piso.data_li [3994];
      \piso.data_r_3993_sv2v_reg  <= \piso.data_li [3993];
      \piso.data_r_3992_sv2v_reg  <= \piso.data_li [3992];
      \piso.data_r_3991_sv2v_reg  <= \piso.data_li [3991];
      \piso.data_r_3990_sv2v_reg  <= \piso.data_li [3990];
      \piso.data_r_3989_sv2v_reg  <= \piso.data_li [3989];
      \piso.data_r_3988_sv2v_reg  <= \piso.data_li [3988];
      \piso.data_r_3987_sv2v_reg  <= \piso.data_li [3987];
      \piso.data_r_3986_sv2v_reg  <= \piso.data_li [3986];
      \piso.data_r_3985_sv2v_reg  <= \piso.data_li [3985];
      \piso.data_r_3984_sv2v_reg  <= \piso.data_li [3984];
      \piso.data_r_3983_sv2v_reg  <= \piso.data_li [3983];
      \piso.data_r_3982_sv2v_reg  <= \piso.data_li [3982];
      \piso.data_r_3981_sv2v_reg  <= \piso.data_li [3981];
      \piso.data_r_3980_sv2v_reg  <= \piso.data_li [3980];
      \piso.data_r_3979_sv2v_reg  <= \piso.data_li [3979];
      \piso.data_r_3978_sv2v_reg  <= \piso.data_li [3978];
      \piso.data_r_3977_sv2v_reg  <= \piso.data_li [3977];
      \piso.data_r_3976_sv2v_reg  <= \piso.data_li [3976];
      \piso.data_r_3975_sv2v_reg  <= \piso.data_li [3975];
      \piso.data_r_3974_sv2v_reg  <= \piso.data_li [3974];
      \piso.data_r_3973_sv2v_reg  <= \piso.data_li [3973];
      \piso.data_r_3972_sv2v_reg  <= \piso.data_li [3972];
      \piso.data_r_3971_sv2v_reg  <= \piso.data_li [3971];
      \piso.data_r_3970_sv2v_reg  <= \piso.data_li [3970];
      \piso.data_r_3969_sv2v_reg  <= \piso.data_li [3969];
      \piso.data_r_3968_sv2v_reg  <= \piso.data_li [3968];
      \piso.data_r_3967_sv2v_reg  <= \piso.data_li [3967];
      \piso.data_r_3966_sv2v_reg  <= \piso.data_li [3966];
      \piso.data_r_3965_sv2v_reg  <= \piso.data_li [3965];
      \piso.data_r_3964_sv2v_reg  <= \piso.data_li [3964];
      \piso.data_r_3963_sv2v_reg  <= \piso.data_li [3963];
      \piso.data_r_3962_sv2v_reg  <= \piso.data_li [3962];
      \piso.data_r_3961_sv2v_reg  <= \piso.data_li [3961];
      \piso.data_r_3960_sv2v_reg  <= \piso.data_li [3960];
      \piso.data_r_3959_sv2v_reg  <= \piso.data_li [3959];
      \piso.data_r_3958_sv2v_reg  <= \piso.data_li [3958];
      \piso.data_r_3957_sv2v_reg  <= \piso.data_li [3957];
      \piso.data_r_3956_sv2v_reg  <= \piso.data_li [3956];
      \piso.data_r_3955_sv2v_reg  <= \piso.data_li [3955];
      \piso.data_r_3954_sv2v_reg  <= \piso.data_li [3954];
      \piso.data_r_3953_sv2v_reg  <= \piso.data_li [3953];
      \piso.data_r_3952_sv2v_reg  <= \piso.data_li [3952];
      \piso.data_r_3951_sv2v_reg  <= \piso.data_li [3951];
      \piso.data_r_3950_sv2v_reg  <= \piso.data_li [3950];
      \piso.data_r_3949_sv2v_reg  <= \piso.data_li [3949];
      \piso.data_r_3948_sv2v_reg  <= \piso.data_li [3948];
      \piso.data_r_3947_sv2v_reg  <= \piso.data_li [3947];
      \piso.data_r_3946_sv2v_reg  <= \piso.data_li [3946];
      \piso.data_r_3945_sv2v_reg  <= \piso.data_li [3945];
      \piso.data_r_3944_sv2v_reg  <= \piso.data_li [3944];
      \piso.data_r_3943_sv2v_reg  <= \piso.data_li [3943];
      \piso.data_r_3942_sv2v_reg  <= \piso.data_li [3942];
      \piso.data_r_3941_sv2v_reg  <= \piso.data_li [3941];
      \piso.data_r_3940_sv2v_reg  <= \piso.data_li [3940];
      \piso.data_r_3939_sv2v_reg  <= \piso.data_li [3939];
      \piso.data_r_3938_sv2v_reg  <= \piso.data_li [3938];
      \piso.data_r_3937_sv2v_reg  <= \piso.data_li [3937];
      \piso.data_r_3936_sv2v_reg  <= \piso.data_li [3936];
      \piso.data_r_3935_sv2v_reg  <= \piso.data_li [3935];
      \piso.data_r_3934_sv2v_reg  <= \piso.data_li [3934];
      \piso.data_r_3933_sv2v_reg  <= \piso.data_li [3933];
      \piso.data_r_3932_sv2v_reg  <= \piso.data_li [3932];
      \piso.data_r_3931_sv2v_reg  <= \piso.data_li [3931];
      \piso.data_r_3930_sv2v_reg  <= \piso.data_li [3930];
      \piso.data_r_3929_sv2v_reg  <= \piso.data_li [3929];
      \piso.data_r_3928_sv2v_reg  <= \piso.data_li [3928];
      \piso.data_r_3927_sv2v_reg  <= \piso.data_li [3927];
      \piso.data_r_3926_sv2v_reg  <= \piso.data_li [3926];
      \piso.data_r_3925_sv2v_reg  <= \piso.data_li [3925];
      \piso.data_r_3924_sv2v_reg  <= \piso.data_li [3924];
      \piso.data_r_3923_sv2v_reg  <= \piso.data_li [3923];
      \piso.data_r_3922_sv2v_reg  <= \piso.data_li [3922];
      \piso.data_r_3921_sv2v_reg  <= \piso.data_li [3921];
      \piso.data_r_3920_sv2v_reg  <= \piso.data_li [3920];
      \piso.data_r_3919_sv2v_reg  <= \piso.data_li [3919];
      \piso.data_r_3918_sv2v_reg  <= \piso.data_li [3918];
      \piso.data_r_3917_sv2v_reg  <= \piso.data_li [3917];
      \piso.data_r_3916_sv2v_reg  <= \piso.data_li [3916];
      \piso.data_r_3915_sv2v_reg  <= \piso.data_li [3915];
      \piso.data_r_3914_sv2v_reg  <= \piso.data_li [3914];
      \piso.data_r_3913_sv2v_reg  <= \piso.data_li [3913];
      \piso.data_r_3912_sv2v_reg  <= \piso.data_li [3912];
      \piso.data_r_3911_sv2v_reg  <= \piso.data_li [3911];
      \piso.data_r_3910_sv2v_reg  <= \piso.data_li [3910];
      \piso.data_r_3909_sv2v_reg  <= \piso.data_li [3909];
      \piso.data_r_3908_sv2v_reg  <= \piso.data_li [3908];
      \piso.data_r_3907_sv2v_reg  <= \piso.data_li [3907];
      \piso.data_r_3906_sv2v_reg  <= \piso.data_li [3906];
      \piso.data_r_3905_sv2v_reg  <= \piso.data_li [3905];
      \piso.data_r_3904_sv2v_reg  <= \piso.data_li [3904];
      \piso.data_r_3903_sv2v_reg  <= \piso.data_li [3903];
      \piso.data_r_3902_sv2v_reg  <= \piso.data_li [3902];
      \piso.data_r_3901_sv2v_reg  <= \piso.data_li [3901];
      \piso.data_r_3900_sv2v_reg  <= \piso.data_li [3900];
      \piso.data_r_3899_sv2v_reg  <= \piso.data_li [3899];
      \piso.data_r_3898_sv2v_reg  <= \piso.data_li [3898];
      \piso.data_r_3897_sv2v_reg  <= \piso.data_li [3897];
      \piso.data_r_3896_sv2v_reg  <= \piso.data_li [3896];
      \piso.data_r_3895_sv2v_reg  <= \piso.data_li [3895];
      \piso.data_r_3894_sv2v_reg  <= \piso.data_li [3894];
      \piso.data_r_3893_sv2v_reg  <= \piso.data_li [3893];
      \piso.data_r_3892_sv2v_reg  <= \piso.data_li [3892];
      \piso.data_r_3891_sv2v_reg  <= \piso.data_li [3891];
      \piso.data_r_3890_sv2v_reg  <= \piso.data_li [3890];
      \piso.data_r_3889_sv2v_reg  <= \piso.data_li [3889];
      \piso.data_r_3888_sv2v_reg  <= \piso.data_li [3888];
      \piso.data_r_3887_sv2v_reg  <= \piso.data_li [3887];
      \piso.data_r_3886_sv2v_reg  <= \piso.data_li [3886];
      \piso.data_r_3885_sv2v_reg  <= \piso.data_li [3885];
      \piso.data_r_3884_sv2v_reg  <= \piso.data_li [3884];
      \piso.data_r_3883_sv2v_reg  <= \piso.data_li [3883];
      \piso.data_r_3882_sv2v_reg  <= \piso.data_li [3882];
      \piso.data_r_3881_sv2v_reg  <= \piso.data_li [3881];
      \piso.data_r_3880_sv2v_reg  <= \piso.data_li [3880];
      \piso.data_r_3879_sv2v_reg  <= \piso.data_li [3879];
      \piso.data_r_3878_sv2v_reg  <= \piso.data_li [3878];
      \piso.data_r_3877_sv2v_reg  <= \piso.data_li [3877];
      \piso.data_r_3876_sv2v_reg  <= \piso.data_li [3876];
      \piso.data_r_3875_sv2v_reg  <= \piso.data_li [3875];
      \piso.data_r_3874_sv2v_reg  <= \piso.data_li [3874];
      \piso.data_r_3873_sv2v_reg  <= \piso.data_li [3873];
      \piso.data_r_3872_sv2v_reg  <= \piso.data_li [3872];
      \piso.data_r_3871_sv2v_reg  <= \piso.data_li [3871];
      \piso.data_r_3870_sv2v_reg  <= \piso.data_li [3870];
      \piso.data_r_3869_sv2v_reg  <= \piso.data_li [3869];
      \piso.data_r_3868_sv2v_reg  <= \piso.data_li [3868];
      \piso.data_r_3867_sv2v_reg  <= \piso.data_li [3867];
      \piso.data_r_3866_sv2v_reg  <= \piso.data_li [3866];
      \piso.data_r_3865_sv2v_reg  <= \piso.data_li [3865];
      \piso.data_r_3864_sv2v_reg  <= \piso.data_li [3864];
      \piso.data_r_3863_sv2v_reg  <= \piso.data_li [3863];
      \piso.data_r_3862_sv2v_reg  <= \piso.data_li [3862];
      \piso.data_r_3861_sv2v_reg  <= \piso.data_li [3861];
      \piso.data_r_3860_sv2v_reg  <= \piso.data_li [3860];
      \piso.data_r_3859_sv2v_reg  <= \piso.data_li [3859];
      \piso.data_r_3858_sv2v_reg  <= \piso.data_li [3858];
      \piso.data_r_3857_sv2v_reg  <= \piso.data_li [3857];
      \piso.data_r_3856_sv2v_reg  <= \piso.data_li [3856];
      \piso.data_r_3855_sv2v_reg  <= \piso.data_li [3855];
      \piso.data_r_3854_sv2v_reg  <= \piso.data_li [3854];
      \piso.data_r_3853_sv2v_reg  <= \piso.data_li [3853];
      \piso.data_r_3852_sv2v_reg  <= \piso.data_li [3852];
      \piso.data_r_3851_sv2v_reg  <= \piso.data_li [3851];
      \piso.data_r_3850_sv2v_reg  <= \piso.data_li [3850];
      \piso.data_r_3849_sv2v_reg  <= \piso.data_li [3849];
      \piso.data_r_3848_sv2v_reg  <= \piso.data_li [3848];
      \piso.data_r_3847_sv2v_reg  <= \piso.data_li [3847];
      \piso.data_r_3846_sv2v_reg  <= \piso.data_li [3846];
      \piso.data_r_3845_sv2v_reg  <= \piso.data_li [3845];
      \piso.data_r_3844_sv2v_reg  <= \piso.data_li [3844];
      \piso.data_r_3843_sv2v_reg  <= \piso.data_li [3843];
      \piso.data_r_3842_sv2v_reg  <= \piso.data_li [3842];
      \piso.data_r_3841_sv2v_reg  <= \piso.data_li [3841];
      \piso.data_r_3840_sv2v_reg  <= \piso.data_li [3840];
      \piso.data_r_3839_sv2v_reg  <= \piso.data_li [3839];
      \piso.data_r_3838_sv2v_reg  <= \piso.data_li [3838];
      \piso.data_r_3837_sv2v_reg  <= \piso.data_li [3837];
      \piso.data_r_3836_sv2v_reg  <= \piso.data_li [3836];
      \piso.data_r_3835_sv2v_reg  <= \piso.data_li [3835];
      \piso.data_r_3834_sv2v_reg  <= \piso.data_li [3834];
      \piso.data_r_3833_sv2v_reg  <= \piso.data_li [3833];
      \piso.data_r_3832_sv2v_reg  <= \piso.data_li [3832];
      \piso.data_r_3831_sv2v_reg  <= \piso.data_li [3831];
      \piso.data_r_3830_sv2v_reg  <= \piso.data_li [3830];
      \piso.data_r_3829_sv2v_reg  <= \piso.data_li [3829];
      \piso.data_r_3828_sv2v_reg  <= \piso.data_li [3828];
      \piso.data_r_3827_sv2v_reg  <= \piso.data_li [3827];
      \piso.data_r_3826_sv2v_reg  <= \piso.data_li [3826];
      \piso.data_r_3825_sv2v_reg  <= \piso.data_li [3825];
      \piso.data_r_3824_sv2v_reg  <= \piso.data_li [3824];
      \piso.data_r_3823_sv2v_reg  <= \piso.data_li [3823];
      \piso.data_r_3822_sv2v_reg  <= \piso.data_li [3822];
      \piso.data_r_3821_sv2v_reg  <= \piso.data_li [3821];
      \piso.data_r_3820_sv2v_reg  <= \piso.data_li [3820];
      \piso.data_r_3819_sv2v_reg  <= \piso.data_li [3819];
      \piso.data_r_3818_sv2v_reg  <= \piso.data_li [3818];
      \piso.data_r_3817_sv2v_reg  <= \piso.data_li [3817];
      \piso.data_r_3816_sv2v_reg  <= \piso.data_li [3816];
      \piso.data_r_3815_sv2v_reg  <= \piso.data_li [3815];
      \piso.data_r_3814_sv2v_reg  <= \piso.data_li [3814];
      \piso.data_r_3813_sv2v_reg  <= \piso.data_li [3813];
      \piso.data_r_3812_sv2v_reg  <= \piso.data_li [3812];
      \piso.data_r_3811_sv2v_reg  <= \piso.data_li [3811];
      \piso.data_r_3810_sv2v_reg  <= \piso.data_li [3810];
      \piso.data_r_3809_sv2v_reg  <= \piso.data_li [3809];
      \piso.data_r_3808_sv2v_reg  <= \piso.data_li [3808];
      \piso.data_r_3807_sv2v_reg  <= \piso.data_li [3807];
      \piso.data_r_3806_sv2v_reg  <= \piso.data_li [3806];
      \piso.data_r_3805_sv2v_reg  <= \piso.data_li [3805];
      \piso.data_r_3804_sv2v_reg  <= \piso.data_li [3804];
      \piso.data_r_3803_sv2v_reg  <= \piso.data_li [3803];
      \piso.data_r_3802_sv2v_reg  <= \piso.data_li [3802];
      \piso.data_r_3801_sv2v_reg  <= \piso.data_li [3801];
      \piso.data_r_3800_sv2v_reg  <= \piso.data_li [3800];
      \piso.data_r_3799_sv2v_reg  <= \piso.data_li [3799];
      \piso.data_r_3798_sv2v_reg  <= \piso.data_li [3798];
      \piso.data_r_3797_sv2v_reg  <= \piso.data_li [3797];
      \piso.data_r_3796_sv2v_reg  <= \piso.data_li [3796];
      \piso.data_r_3795_sv2v_reg  <= \piso.data_li [3795];
      \piso.data_r_3794_sv2v_reg  <= \piso.data_li [3794];
      \piso.data_r_3793_sv2v_reg  <= \piso.data_li [3793];
      \piso.data_r_3792_sv2v_reg  <= \piso.data_li [3792];
      \piso.data_r_3791_sv2v_reg  <= \piso.data_li [3791];
      \piso.data_r_3790_sv2v_reg  <= \piso.data_li [3790];
      \piso.data_r_3789_sv2v_reg  <= \piso.data_li [3789];
      \piso.data_r_3788_sv2v_reg  <= \piso.data_li [3788];
      \piso.data_r_3787_sv2v_reg  <= \piso.data_li [3787];
      \piso.data_r_3786_sv2v_reg  <= \piso.data_li [3786];
      \piso.data_r_3785_sv2v_reg  <= \piso.data_li [3785];
      \piso.data_r_3784_sv2v_reg  <= \piso.data_li [3784];
      \piso.data_r_3783_sv2v_reg  <= \piso.data_li [3783];
      \piso.data_r_3782_sv2v_reg  <= \piso.data_li [3782];
      \piso.data_r_3781_sv2v_reg  <= \piso.data_li [3781];
      \piso.data_r_3780_sv2v_reg  <= \piso.data_li [3780];
      \piso.data_r_3779_sv2v_reg  <= \piso.data_li [3779];
      \piso.data_r_3778_sv2v_reg  <= \piso.data_li [3778];
      \piso.data_r_3777_sv2v_reg  <= \piso.data_li [3777];
      \piso.data_r_3776_sv2v_reg  <= \piso.data_li [3776];
      \piso.data_r_3775_sv2v_reg  <= \piso.data_li [3775];
      \piso.data_r_3774_sv2v_reg  <= \piso.data_li [3774];
      \piso.data_r_3773_sv2v_reg  <= \piso.data_li [3773];
      \piso.data_r_3772_sv2v_reg  <= \piso.data_li [3772];
      \piso.data_r_3771_sv2v_reg  <= \piso.data_li [3771];
      \piso.data_r_3770_sv2v_reg  <= \piso.data_li [3770];
      \piso.data_r_3769_sv2v_reg  <= \piso.data_li [3769];
      \piso.data_r_3768_sv2v_reg  <= \piso.data_li [3768];
      \piso.data_r_3767_sv2v_reg  <= \piso.data_li [3767];
      \piso.data_r_3766_sv2v_reg  <= \piso.data_li [3766];
      \piso.data_r_3765_sv2v_reg  <= \piso.data_li [3765];
      \piso.data_r_3764_sv2v_reg  <= \piso.data_li [3764];
      \piso.data_r_3763_sv2v_reg  <= \piso.data_li [3763];
      \piso.data_r_3762_sv2v_reg  <= \piso.data_li [3762];
      \piso.data_r_3761_sv2v_reg  <= \piso.data_li [3761];
      \piso.data_r_3760_sv2v_reg  <= \piso.data_li [3760];
      \piso.data_r_3759_sv2v_reg  <= \piso.data_li [3759];
      \piso.data_r_3758_sv2v_reg  <= \piso.data_li [3758];
      \piso.data_r_3757_sv2v_reg  <= \piso.data_li [3757];
      \piso.data_r_3756_sv2v_reg  <= \piso.data_li [3756];
      \piso.data_r_3755_sv2v_reg  <= \piso.data_li [3755];
      \piso.data_r_3754_sv2v_reg  <= \piso.data_li [3754];
      \piso.data_r_3753_sv2v_reg  <= \piso.data_li [3753];
      \piso.data_r_3752_sv2v_reg  <= \piso.data_li [3752];
      \piso.data_r_3751_sv2v_reg  <= \piso.data_li [3751];
      \piso.data_r_3750_sv2v_reg  <= \piso.data_li [3750];
      \piso.data_r_3749_sv2v_reg  <= \piso.data_li [3749];
      \piso.data_r_3748_sv2v_reg  <= \piso.data_li [3748];
      \piso.data_r_3747_sv2v_reg  <= \piso.data_li [3747];
      \piso.data_r_3746_sv2v_reg  <= \piso.data_li [3746];
      \piso.data_r_3745_sv2v_reg  <= \piso.data_li [3745];
      \piso.data_r_3744_sv2v_reg  <= \piso.data_li [3744];
      \piso.data_r_3743_sv2v_reg  <= \piso.data_li [3743];
      \piso.data_r_3742_sv2v_reg  <= \piso.data_li [3742];
      \piso.data_r_3741_sv2v_reg  <= \piso.data_li [3741];
      \piso.data_r_3740_sv2v_reg  <= \piso.data_li [3740];
      \piso.data_r_3739_sv2v_reg  <= \piso.data_li [3739];
      \piso.data_r_3738_sv2v_reg  <= \piso.data_li [3738];
      \piso.data_r_3737_sv2v_reg  <= \piso.data_li [3737];
      \piso.data_r_3736_sv2v_reg  <= \piso.data_li [3736];
      \piso.data_r_3735_sv2v_reg  <= \piso.data_li [3735];
      \piso.data_r_3734_sv2v_reg  <= \piso.data_li [3734];
      \piso.data_r_3733_sv2v_reg  <= \piso.data_li [3733];
      \piso.data_r_3732_sv2v_reg  <= \piso.data_li [3732];
      \piso.data_r_3731_sv2v_reg  <= \piso.data_li [3731];
      \piso.data_r_3730_sv2v_reg  <= \piso.data_li [3730];
      \piso.data_r_3729_sv2v_reg  <= \piso.data_li [3729];
      \piso.data_r_3728_sv2v_reg  <= \piso.data_li [3728];
      \piso.data_r_3727_sv2v_reg  <= \piso.data_li [3727];
      \piso.data_r_3726_sv2v_reg  <= \piso.data_li [3726];
      \piso.data_r_3725_sv2v_reg  <= \piso.data_li [3725];
      \piso.data_r_3724_sv2v_reg  <= \piso.data_li [3724];
      \piso.data_r_3723_sv2v_reg  <= \piso.data_li [3723];
      \piso.data_r_3722_sv2v_reg  <= \piso.data_li [3722];
      \piso.data_r_3721_sv2v_reg  <= \piso.data_li [3721];
      \piso.data_r_3720_sv2v_reg  <= \piso.data_li [3720];
      \piso.data_r_3719_sv2v_reg  <= \piso.data_li [3719];
      \piso.data_r_3718_sv2v_reg  <= \piso.data_li [3718];
      \piso.data_r_3717_sv2v_reg  <= \piso.data_li [3717];
      \piso.data_r_3716_sv2v_reg  <= \piso.data_li [3716];
      \piso.data_r_3715_sv2v_reg  <= \piso.data_li [3715];
      \piso.data_r_3714_sv2v_reg  <= \piso.data_li [3714];
      \piso.data_r_3713_sv2v_reg  <= \piso.data_li [3713];
      \piso.data_r_3712_sv2v_reg  <= \piso.data_li [3712];
      \piso.data_r_3711_sv2v_reg  <= \piso.data_li [3711];
      \piso.data_r_3710_sv2v_reg  <= \piso.data_li [3710];
      \piso.data_r_3709_sv2v_reg  <= \piso.data_li [3709];
      \piso.data_r_3708_sv2v_reg  <= \piso.data_li [3708];
      \piso.data_r_3707_sv2v_reg  <= \piso.data_li [3707];
      \piso.data_r_3706_sv2v_reg  <= \piso.data_li [3706];
      \piso.data_r_3705_sv2v_reg  <= \piso.data_li [3705];
      \piso.data_r_3704_sv2v_reg  <= \piso.data_li [3704];
      \piso.data_r_3703_sv2v_reg  <= \piso.data_li [3703];
      \piso.data_r_3702_sv2v_reg  <= \piso.data_li [3702];
      \piso.data_r_3701_sv2v_reg  <= \piso.data_li [3701];
      \piso.data_r_3700_sv2v_reg  <= \piso.data_li [3700];
      \piso.data_r_3699_sv2v_reg  <= \piso.data_li [3699];
      \piso.data_r_3698_sv2v_reg  <= \piso.data_li [3698];
      \piso.data_r_3697_sv2v_reg  <= \piso.data_li [3697];
      \piso.data_r_3696_sv2v_reg  <= \piso.data_li [3696];
      \piso.data_r_3695_sv2v_reg  <= \piso.data_li [3695];
      \piso.data_r_3694_sv2v_reg  <= \piso.data_li [3694];
      \piso.data_r_3693_sv2v_reg  <= \piso.data_li [3693];
      \piso.data_r_3692_sv2v_reg  <= \piso.data_li [3692];
      \piso.data_r_3691_sv2v_reg  <= \piso.data_li [3691];
      \piso.data_r_3690_sv2v_reg  <= \piso.data_li [3690];
      \piso.data_r_3689_sv2v_reg  <= \piso.data_li [3689];
      \piso.data_r_3688_sv2v_reg  <= \piso.data_li [3688];
      \piso.data_r_3687_sv2v_reg  <= \piso.data_li [3687];
      \piso.data_r_3686_sv2v_reg  <= \piso.data_li [3686];
      \piso.data_r_3685_sv2v_reg  <= \piso.data_li [3685];
      \piso.data_r_3684_sv2v_reg  <= \piso.data_li [3684];
      \piso.data_r_3683_sv2v_reg  <= \piso.data_li [3683];
      \piso.data_r_3682_sv2v_reg  <= \piso.data_li [3682];
      \piso.data_r_3681_sv2v_reg  <= \piso.data_li [3681];
      \piso.data_r_3680_sv2v_reg  <= \piso.data_li [3680];
      \piso.data_r_3679_sv2v_reg  <= \piso.data_li [3679];
      \piso.data_r_3678_sv2v_reg  <= \piso.data_li [3678];
      \piso.data_r_3677_sv2v_reg  <= \piso.data_li [3677];
      \piso.data_r_3676_sv2v_reg  <= \piso.data_li [3676];
      \piso.data_r_3675_sv2v_reg  <= \piso.data_li [3675];
      \piso.data_r_3674_sv2v_reg  <= \piso.data_li [3674];
      \piso.data_r_3673_sv2v_reg  <= \piso.data_li [3673];
      \piso.data_r_3672_sv2v_reg  <= \piso.data_li [3672];
      \piso.data_r_3671_sv2v_reg  <= \piso.data_li [3671];
      \piso.data_r_3670_sv2v_reg  <= \piso.data_li [3670];
      \piso.data_r_3669_sv2v_reg  <= \piso.data_li [3669];
      \piso.data_r_3668_sv2v_reg  <= \piso.data_li [3668];
      \piso.data_r_3667_sv2v_reg  <= \piso.data_li [3667];
      \piso.data_r_3666_sv2v_reg  <= \piso.data_li [3666];
      \piso.data_r_3665_sv2v_reg  <= \piso.data_li [3665];
      \piso.data_r_3664_sv2v_reg  <= \piso.data_li [3664];
      \piso.data_r_3663_sv2v_reg  <= \piso.data_li [3663];
      \piso.data_r_3662_sv2v_reg  <= \piso.data_li [3662];
      \piso.data_r_3661_sv2v_reg  <= \piso.data_li [3661];
      \piso.data_r_3660_sv2v_reg  <= \piso.data_li [3660];
      \piso.data_r_3659_sv2v_reg  <= \piso.data_li [3659];
      \piso.data_r_3658_sv2v_reg  <= \piso.data_li [3658];
      \piso.data_r_3657_sv2v_reg  <= \piso.data_li [3657];
      \piso.data_r_3656_sv2v_reg  <= \piso.data_li [3656];
      \piso.data_r_3655_sv2v_reg  <= \piso.data_li [3655];
      \piso.data_r_3654_sv2v_reg  <= \piso.data_li [3654];
      \piso.data_r_3653_sv2v_reg  <= \piso.data_li [3653];
      \piso.data_r_3652_sv2v_reg  <= \piso.data_li [3652];
      \piso.data_r_3651_sv2v_reg  <= \piso.data_li [3651];
      \piso.data_r_3650_sv2v_reg  <= \piso.data_li [3650];
      \piso.data_r_3649_sv2v_reg  <= \piso.data_li [3649];
      \piso.data_r_3648_sv2v_reg  <= \piso.data_li [3648];
      \piso.data_r_3647_sv2v_reg  <= \piso.data_li [3647];
      \piso.data_r_3646_sv2v_reg  <= \piso.data_li [3646];
      \piso.data_r_3645_sv2v_reg  <= \piso.data_li [3645];
      \piso.data_r_3644_sv2v_reg  <= \piso.data_li [3644];
      \piso.data_r_3643_sv2v_reg  <= \piso.data_li [3643];
      \piso.data_r_3642_sv2v_reg  <= \piso.data_li [3642];
      \piso.data_r_3641_sv2v_reg  <= \piso.data_li [3641];
      \piso.data_r_3640_sv2v_reg  <= \piso.data_li [3640];
      \piso.data_r_3639_sv2v_reg  <= \piso.data_li [3639];
      \piso.data_r_3638_sv2v_reg  <= \piso.data_li [3638];
      \piso.data_r_3637_sv2v_reg  <= \piso.data_li [3637];
      \piso.data_r_3636_sv2v_reg  <= \piso.data_li [3636];
      \piso.data_r_3635_sv2v_reg  <= \piso.data_li [3635];
      \piso.data_r_3634_sv2v_reg  <= \piso.data_li [3634];
      \piso.data_r_3633_sv2v_reg  <= \piso.data_li [3633];
      \piso.data_r_3632_sv2v_reg  <= \piso.data_li [3632];
      \piso.data_r_3631_sv2v_reg  <= \piso.data_li [3631];
      \piso.data_r_3630_sv2v_reg  <= \piso.data_li [3630];
      \piso.data_r_3629_sv2v_reg  <= \piso.data_li [3629];
      \piso.data_r_3628_sv2v_reg  <= \piso.data_li [3628];
      \piso.data_r_3627_sv2v_reg  <= \piso.data_li [3627];
      \piso.data_r_3626_sv2v_reg  <= \piso.data_li [3626];
      \piso.data_r_3625_sv2v_reg  <= \piso.data_li [3625];
      \piso.data_r_3624_sv2v_reg  <= \piso.data_li [3624];
      \piso.data_r_3623_sv2v_reg  <= \piso.data_li [3623];
      \piso.data_r_3622_sv2v_reg  <= \piso.data_li [3622];
      \piso.data_r_3621_sv2v_reg  <= \piso.data_li [3621];
      \piso.data_r_3620_sv2v_reg  <= \piso.data_li [3620];
      \piso.data_r_3619_sv2v_reg  <= \piso.data_li [3619];
      \piso.data_r_3618_sv2v_reg  <= \piso.data_li [3618];
      \piso.data_r_3617_sv2v_reg  <= \piso.data_li [3617];
      \piso.data_r_3616_sv2v_reg  <= \piso.data_li [3616];
      \piso.data_r_3615_sv2v_reg  <= \piso.data_li [3615];
      \piso.data_r_3614_sv2v_reg  <= \piso.data_li [3614];
      \piso.data_r_3613_sv2v_reg  <= \piso.data_li [3613];
      \piso.data_r_3612_sv2v_reg  <= \piso.data_li [3612];
      \piso.data_r_3611_sv2v_reg  <= \piso.data_li [3611];
      \piso.data_r_3610_sv2v_reg  <= \piso.data_li [3610];
      \piso.data_r_3609_sv2v_reg  <= \piso.data_li [3609];
      \piso.data_r_3608_sv2v_reg  <= \piso.data_li [3608];
      \piso.data_r_3607_sv2v_reg  <= \piso.data_li [3607];
      \piso.data_r_3606_sv2v_reg  <= \piso.data_li [3606];
      \piso.data_r_3605_sv2v_reg  <= \piso.data_li [3605];
      \piso.data_r_3604_sv2v_reg  <= \piso.data_li [3604];
      \piso.data_r_3603_sv2v_reg  <= \piso.data_li [3603];
      \piso.data_r_3602_sv2v_reg  <= \piso.data_li [3602];
      \piso.data_r_3601_sv2v_reg  <= \piso.data_li [3601];
      \piso.data_r_3600_sv2v_reg  <= \piso.data_li [3600];
      \piso.data_r_3599_sv2v_reg  <= \piso.data_li [3599];
      \piso.data_r_3598_sv2v_reg  <= \piso.data_li [3598];
      \piso.data_r_3597_sv2v_reg  <= \piso.data_li [3597];
      \piso.data_r_3596_sv2v_reg  <= \piso.data_li [3596];
      \piso.data_r_3595_sv2v_reg  <= \piso.data_li [3595];
      \piso.data_r_3594_sv2v_reg  <= \piso.data_li [3594];
      \piso.data_r_3593_sv2v_reg  <= \piso.data_li [3593];
      \piso.data_r_3592_sv2v_reg  <= \piso.data_li [3592];
      \piso.data_r_3591_sv2v_reg  <= \piso.data_li [3591];
      \piso.data_r_3590_sv2v_reg  <= \piso.data_li [3590];
      \piso.data_r_3589_sv2v_reg  <= \piso.data_li [3589];
      \piso.data_r_3588_sv2v_reg  <= \piso.data_li [3588];
      \piso.data_r_3587_sv2v_reg  <= \piso.data_li [3587];
      \piso.data_r_3586_sv2v_reg  <= \piso.data_li [3586];
      \piso.data_r_3585_sv2v_reg  <= \piso.data_li [3585];
      \piso.data_r_3584_sv2v_reg  <= \piso.data_li [3584];
      \piso.data_r_3583_sv2v_reg  <= \piso.data_li [3583];
      \piso.data_r_3582_sv2v_reg  <= \piso.data_li [3582];
      \piso.data_r_3581_sv2v_reg  <= \piso.data_li [3581];
      \piso.data_r_3580_sv2v_reg  <= \piso.data_li [3580];
      \piso.data_r_3579_sv2v_reg  <= \piso.data_li [3579];
      \piso.data_r_3578_sv2v_reg  <= \piso.data_li [3578];
      \piso.data_r_3577_sv2v_reg  <= \piso.data_li [3577];
      \piso.data_r_3576_sv2v_reg  <= \piso.data_li [3576];
      \piso.data_r_3575_sv2v_reg  <= \piso.data_li [3575];
      \piso.data_r_3574_sv2v_reg  <= \piso.data_li [3574];
      \piso.data_r_3573_sv2v_reg  <= \piso.data_li [3573];
      \piso.data_r_3572_sv2v_reg  <= \piso.data_li [3572];
      \piso.data_r_3571_sv2v_reg  <= \piso.data_li [3571];
      \piso.data_r_3570_sv2v_reg  <= \piso.data_li [3570];
      \piso.data_r_3569_sv2v_reg  <= \piso.data_li [3569];
      \piso.data_r_3568_sv2v_reg  <= \piso.data_li [3568];
      \piso.data_r_3567_sv2v_reg  <= \piso.data_li [3567];
      \piso.data_r_3566_sv2v_reg  <= \piso.data_li [3566];
      \piso.data_r_3565_sv2v_reg  <= \piso.data_li [3565];
      \piso.data_r_3564_sv2v_reg  <= \piso.data_li [3564];
      \piso.data_r_3563_sv2v_reg  <= \piso.data_li [3563];
      \piso.data_r_3562_sv2v_reg  <= \piso.data_li [3562];
      \piso.data_r_3561_sv2v_reg  <= \piso.data_li [3561];
      \piso.data_r_3560_sv2v_reg  <= \piso.data_li [3560];
      \piso.data_r_3559_sv2v_reg  <= \piso.data_li [3559];
      \piso.data_r_3558_sv2v_reg  <= \piso.data_li [3558];
      \piso.data_r_3557_sv2v_reg  <= \piso.data_li [3557];
      \piso.data_r_3556_sv2v_reg  <= \piso.data_li [3556];
      \piso.data_r_3555_sv2v_reg  <= \piso.data_li [3555];
      \piso.data_r_3554_sv2v_reg  <= \piso.data_li [3554];
      \piso.data_r_3553_sv2v_reg  <= \piso.data_li [3553];
      \piso.data_r_3552_sv2v_reg  <= \piso.data_li [3552];
      \piso.data_r_3551_sv2v_reg  <= \piso.data_li [3551];
      \piso.data_r_3550_sv2v_reg  <= \piso.data_li [3550];
      \piso.data_r_3549_sv2v_reg  <= \piso.data_li [3549];
      \piso.data_r_3548_sv2v_reg  <= \piso.data_li [3548];
      \piso.data_r_3547_sv2v_reg  <= \piso.data_li [3547];
      \piso.data_r_3546_sv2v_reg  <= \piso.data_li [3546];
      \piso.data_r_3545_sv2v_reg  <= \piso.data_li [3545];
      \piso.data_r_3544_sv2v_reg  <= \piso.data_li [3544];
      \piso.data_r_3543_sv2v_reg  <= \piso.data_li [3543];
      \piso.data_r_3542_sv2v_reg  <= \piso.data_li [3542];
      \piso.data_r_3541_sv2v_reg  <= \piso.data_li [3541];
      \piso.data_r_3540_sv2v_reg  <= \piso.data_li [3540];
      \piso.data_r_3539_sv2v_reg  <= \piso.data_li [3539];
      \piso.data_r_3538_sv2v_reg  <= \piso.data_li [3538];
      \piso.data_r_3537_sv2v_reg  <= \piso.data_li [3537];
      \piso.data_r_3536_sv2v_reg  <= \piso.data_li [3536];
      \piso.data_r_3535_sv2v_reg  <= \piso.data_li [3535];
      \piso.data_r_3534_sv2v_reg  <= \piso.data_li [3534];
      \piso.data_r_3533_sv2v_reg  <= \piso.data_li [3533];
      \piso.data_r_3532_sv2v_reg  <= \piso.data_li [3532];
      \piso.data_r_3531_sv2v_reg  <= \piso.data_li [3531];
      \piso.data_r_3530_sv2v_reg  <= \piso.data_li [3530];
      \piso.data_r_3529_sv2v_reg  <= \piso.data_li [3529];
      \piso.data_r_3528_sv2v_reg  <= \piso.data_li [3528];
      \piso.data_r_3527_sv2v_reg  <= \piso.data_li [3527];
      \piso.data_r_3526_sv2v_reg  <= \piso.data_li [3526];
      \piso.data_r_3525_sv2v_reg  <= \piso.data_li [3525];
      \piso.data_r_3524_sv2v_reg  <= \piso.data_li [3524];
      \piso.data_r_3523_sv2v_reg  <= \piso.data_li [3523];
      \piso.data_r_3522_sv2v_reg  <= \piso.data_li [3522];
      \piso.data_r_3521_sv2v_reg  <= \piso.data_li [3521];
      \piso.data_r_3520_sv2v_reg  <= \piso.data_li [3520];
      \piso.data_r_3519_sv2v_reg  <= \piso.data_li [3519];
      \piso.data_r_3518_sv2v_reg  <= \piso.data_li [3518];
      \piso.data_r_3517_sv2v_reg  <= \piso.data_li [3517];
      \piso.data_r_3516_sv2v_reg  <= \piso.data_li [3516];
      \piso.data_r_3515_sv2v_reg  <= \piso.data_li [3515];
      \piso.data_r_3514_sv2v_reg  <= \piso.data_li [3514];
      \piso.data_r_3513_sv2v_reg  <= \piso.data_li [3513];
      \piso.data_r_3512_sv2v_reg  <= \piso.data_li [3512];
      \piso.data_r_3511_sv2v_reg  <= \piso.data_li [3511];
      \piso.data_r_3510_sv2v_reg  <= \piso.data_li [3510];
      \piso.data_r_3509_sv2v_reg  <= \piso.data_li [3509];
      \piso.data_r_3508_sv2v_reg  <= \piso.data_li [3508];
      \piso.data_r_3507_sv2v_reg  <= \piso.data_li [3507];
      \piso.data_r_3506_sv2v_reg  <= \piso.data_li [3506];
      \piso.data_r_3505_sv2v_reg  <= \piso.data_li [3505];
      \piso.data_r_3504_sv2v_reg  <= \piso.data_li [3504];
      \piso.data_r_3503_sv2v_reg  <= \piso.data_li [3503];
      \piso.data_r_3502_sv2v_reg  <= \piso.data_li [3502];
      \piso.data_r_3501_sv2v_reg  <= \piso.data_li [3501];
      \piso.data_r_3500_sv2v_reg  <= \piso.data_li [3500];
      \piso.data_r_3499_sv2v_reg  <= \piso.data_li [3499];
      \piso.data_r_3498_sv2v_reg  <= \piso.data_li [3498];
      \piso.data_r_3497_sv2v_reg  <= \piso.data_li [3497];
      \piso.data_r_3496_sv2v_reg  <= \piso.data_li [3496];
      \piso.data_r_3495_sv2v_reg  <= \piso.data_li [3495];
      \piso.data_r_3494_sv2v_reg  <= \piso.data_li [3494];
      \piso.data_r_3493_sv2v_reg  <= \piso.data_li [3493];
      \piso.data_r_3492_sv2v_reg  <= \piso.data_li [3492];
      \piso.data_r_3491_sv2v_reg  <= \piso.data_li [3491];
      \piso.data_r_3490_sv2v_reg  <= \piso.data_li [3490];
      \piso.data_r_3489_sv2v_reg  <= \piso.data_li [3489];
      \piso.data_r_3488_sv2v_reg  <= \piso.data_li [3488];
      \piso.data_r_3487_sv2v_reg  <= \piso.data_li [3487];
      \piso.data_r_3486_sv2v_reg  <= \piso.data_li [3486];
      \piso.data_r_3485_sv2v_reg  <= \piso.data_li [3485];
      \piso.data_r_3484_sv2v_reg  <= \piso.data_li [3484];
      \piso.data_r_3483_sv2v_reg  <= \piso.data_li [3483];
      \piso.data_r_3482_sv2v_reg  <= \piso.data_li [3482];
      \piso.data_r_3481_sv2v_reg  <= \piso.data_li [3481];
      \piso.data_r_3480_sv2v_reg  <= \piso.data_li [3480];
      \piso.data_r_3479_sv2v_reg  <= \piso.data_li [3479];
      \piso.data_r_3478_sv2v_reg  <= \piso.data_li [3478];
      \piso.data_r_3477_sv2v_reg  <= \piso.data_li [3477];
      \piso.data_r_3476_sv2v_reg  <= \piso.data_li [3476];
      \piso.data_r_3475_sv2v_reg  <= \piso.data_li [3475];
      \piso.data_r_3474_sv2v_reg  <= \piso.data_li [3474];
      \piso.data_r_3473_sv2v_reg  <= \piso.data_li [3473];
      \piso.data_r_3472_sv2v_reg  <= \piso.data_li [3472];
      \piso.data_r_3471_sv2v_reg  <= \piso.data_li [3471];
      \piso.data_r_3470_sv2v_reg  <= \piso.data_li [3470];
      \piso.data_r_3469_sv2v_reg  <= \piso.data_li [3469];
      \piso.data_r_3468_sv2v_reg  <= \piso.data_li [3468];
      \piso.data_r_3467_sv2v_reg  <= \piso.data_li [3467];
      \piso.data_r_3466_sv2v_reg  <= \piso.data_li [3466];
      \piso.data_r_3465_sv2v_reg  <= \piso.data_li [3465];
      \piso.data_r_3464_sv2v_reg  <= \piso.data_li [3464];
      \piso.data_r_3463_sv2v_reg  <= \piso.data_li [3463];
      \piso.data_r_3462_sv2v_reg  <= \piso.data_li [3462];
      \piso.data_r_3461_sv2v_reg  <= \piso.data_li [3461];
      \piso.data_r_3460_sv2v_reg  <= \piso.data_li [3460];
      \piso.data_r_3459_sv2v_reg  <= \piso.data_li [3459];
      \piso.data_r_3458_sv2v_reg  <= \piso.data_li [3458];
      \piso.data_r_3457_sv2v_reg  <= \piso.data_li [3457];
      \piso.data_r_3456_sv2v_reg  <= \piso.data_li [3456];
      \piso.data_r_3455_sv2v_reg  <= \piso.data_li [3455];
      \piso.data_r_3454_sv2v_reg  <= \piso.data_li [3454];
      \piso.data_r_3453_sv2v_reg  <= \piso.data_li [3453];
      \piso.data_r_3452_sv2v_reg  <= \piso.data_li [3452];
      \piso.data_r_3451_sv2v_reg  <= \piso.data_li [3451];
      \piso.data_r_3450_sv2v_reg  <= \piso.data_li [3450];
      \piso.data_r_3449_sv2v_reg  <= \piso.data_li [3449];
      \piso.data_r_3448_sv2v_reg  <= \piso.data_li [3448];
      \piso.data_r_3447_sv2v_reg  <= \piso.data_li [3447];
      \piso.data_r_3446_sv2v_reg  <= \piso.data_li [3446];
      \piso.data_r_3445_sv2v_reg  <= \piso.data_li [3445];
      \piso.data_r_3444_sv2v_reg  <= \piso.data_li [3444];
      \piso.data_r_3443_sv2v_reg  <= \piso.data_li [3443];
      \piso.data_r_3442_sv2v_reg  <= \piso.data_li [3442];
      \piso.data_r_3441_sv2v_reg  <= \piso.data_li [3441];
      \piso.data_r_3440_sv2v_reg  <= \piso.data_li [3440];
      \piso.data_r_3439_sv2v_reg  <= \piso.data_li [3439];
      \piso.data_r_3438_sv2v_reg  <= \piso.data_li [3438];
      \piso.data_r_3437_sv2v_reg  <= \piso.data_li [3437];
      \piso.data_r_3436_sv2v_reg  <= \piso.data_li [3436];
      \piso.data_r_3435_sv2v_reg  <= \piso.data_li [3435];
      \piso.data_r_3434_sv2v_reg  <= \piso.data_li [3434];
      \piso.data_r_3433_sv2v_reg  <= \piso.data_li [3433];
      \piso.data_r_3432_sv2v_reg  <= \piso.data_li [3432];
      \piso.data_r_3431_sv2v_reg  <= \piso.data_li [3431];
      \piso.data_r_3430_sv2v_reg  <= \piso.data_li [3430];
      \piso.data_r_3429_sv2v_reg  <= \piso.data_li [3429];
      \piso.data_r_3428_sv2v_reg  <= \piso.data_li [3428];
      \piso.data_r_3427_sv2v_reg  <= \piso.data_li [3427];
      \piso.data_r_3426_sv2v_reg  <= \piso.data_li [3426];
      \piso.data_r_3425_sv2v_reg  <= \piso.data_li [3425];
      \piso.data_r_3424_sv2v_reg  <= \piso.data_li [3424];
      \piso.data_r_3423_sv2v_reg  <= \piso.data_li [3423];
      \piso.data_r_3422_sv2v_reg  <= \piso.data_li [3422];
      \piso.data_r_3421_sv2v_reg  <= \piso.data_li [3421];
      \piso.data_r_3420_sv2v_reg  <= \piso.data_li [3420];
      \piso.data_r_3419_sv2v_reg  <= \piso.data_li [3419];
      \piso.data_r_3418_sv2v_reg  <= \piso.data_li [3418];
      \piso.data_r_3417_sv2v_reg  <= \piso.data_li [3417];
      \piso.data_r_3416_sv2v_reg  <= \piso.data_li [3416];
      \piso.data_r_3415_sv2v_reg  <= \piso.data_li [3415];
      \piso.data_r_3414_sv2v_reg  <= \piso.data_li [3414];
      \piso.data_r_3413_sv2v_reg  <= \piso.data_li [3413];
      \piso.data_r_3412_sv2v_reg  <= \piso.data_li [3412];
      \piso.data_r_3411_sv2v_reg  <= \piso.data_li [3411];
      \piso.data_r_3410_sv2v_reg  <= \piso.data_li [3410];
      \piso.data_r_3409_sv2v_reg  <= \piso.data_li [3409];
      \piso.data_r_3408_sv2v_reg  <= \piso.data_li [3408];
      \piso.data_r_3407_sv2v_reg  <= \piso.data_li [3407];
      \piso.data_r_3406_sv2v_reg  <= \piso.data_li [3406];
      \piso.data_r_3405_sv2v_reg  <= \piso.data_li [3405];
      \piso.data_r_3404_sv2v_reg  <= \piso.data_li [3404];
      \piso.data_r_3403_sv2v_reg  <= \piso.data_li [3403];
      \piso.data_r_3402_sv2v_reg  <= \piso.data_li [3402];
      \piso.data_r_3401_sv2v_reg  <= \piso.data_li [3401];
      \piso.data_r_3400_sv2v_reg  <= \piso.data_li [3400];
      \piso.data_r_3399_sv2v_reg  <= \piso.data_li [3399];
      \piso.data_r_3398_sv2v_reg  <= \piso.data_li [3398];
      \piso.data_r_3397_sv2v_reg  <= \piso.data_li [3397];
      \piso.data_r_3396_sv2v_reg  <= \piso.data_li [3396];
      \piso.data_r_3395_sv2v_reg  <= \piso.data_li [3395];
      \piso.data_r_3394_sv2v_reg  <= \piso.data_li [3394];
      \piso.data_r_3393_sv2v_reg  <= \piso.data_li [3393];
      \piso.data_r_3392_sv2v_reg  <= \piso.data_li [3392];
      \piso.data_r_3391_sv2v_reg  <= \piso.data_li [3391];
      \piso.data_r_3390_sv2v_reg  <= \piso.data_li [3390];
      \piso.data_r_3389_sv2v_reg  <= \piso.data_li [3389];
      \piso.data_r_3388_sv2v_reg  <= \piso.data_li [3388];
      \piso.data_r_3387_sv2v_reg  <= \piso.data_li [3387];
      \piso.data_r_3386_sv2v_reg  <= \piso.data_li [3386];
      \piso.data_r_3385_sv2v_reg  <= \piso.data_li [3385];
      \piso.data_r_3384_sv2v_reg  <= \piso.data_li [3384];
      \piso.data_r_3383_sv2v_reg  <= \piso.data_li [3383];
      \piso.data_r_3382_sv2v_reg  <= \piso.data_li [3382];
      \piso.data_r_3381_sv2v_reg  <= \piso.data_li [3381];
      \piso.data_r_3380_sv2v_reg  <= \piso.data_li [3380];
      \piso.data_r_3379_sv2v_reg  <= \piso.data_li [3379];
      \piso.data_r_3378_sv2v_reg  <= \piso.data_li [3378];
      \piso.data_r_3377_sv2v_reg  <= \piso.data_li [3377];
      \piso.data_r_3376_sv2v_reg  <= \piso.data_li [3376];
      \piso.data_r_3375_sv2v_reg  <= \piso.data_li [3375];
      \piso.data_r_3374_sv2v_reg  <= \piso.data_li [3374];
      \piso.data_r_3373_sv2v_reg  <= \piso.data_li [3373];
      \piso.data_r_3372_sv2v_reg  <= \piso.data_li [3372];
      \piso.data_r_3371_sv2v_reg  <= \piso.data_li [3371];
      \piso.data_r_3370_sv2v_reg  <= \piso.data_li [3370];
      \piso.data_r_3369_sv2v_reg  <= \piso.data_li [3369];
      \piso.data_r_3368_sv2v_reg  <= \piso.data_li [3368];
      \piso.data_r_3367_sv2v_reg  <= \piso.data_li [3367];
      \piso.data_r_3366_sv2v_reg  <= \piso.data_li [3366];
      \piso.data_r_3365_sv2v_reg  <= \piso.data_li [3365];
      \piso.data_r_3364_sv2v_reg  <= \piso.data_li [3364];
      \piso.data_r_3363_sv2v_reg  <= \piso.data_li [3363];
      \piso.data_r_3362_sv2v_reg  <= \piso.data_li [3362];
      \piso.data_r_3361_sv2v_reg  <= \piso.data_li [3361];
      \piso.data_r_3360_sv2v_reg  <= \piso.data_li [3360];
      \piso.data_r_3359_sv2v_reg  <= \piso.data_li [3359];
      \piso.data_r_3358_sv2v_reg  <= \piso.data_li [3358];
      \piso.data_r_3357_sv2v_reg  <= \piso.data_li [3357];
      \piso.data_r_3356_sv2v_reg  <= \piso.data_li [3356];
      \piso.data_r_3355_sv2v_reg  <= \piso.data_li [3355];
      \piso.data_r_3354_sv2v_reg  <= \piso.data_li [3354];
      \piso.data_r_3353_sv2v_reg  <= \piso.data_li [3353];
      \piso.data_r_3352_sv2v_reg  <= \piso.data_li [3352];
      \piso.data_r_3351_sv2v_reg  <= \piso.data_li [3351];
      \piso.data_r_3350_sv2v_reg  <= \piso.data_li [3350];
      \piso.data_r_3349_sv2v_reg  <= \piso.data_li [3349];
      \piso.data_r_3348_sv2v_reg  <= \piso.data_li [3348];
      \piso.data_r_3347_sv2v_reg  <= \piso.data_li [3347];
      \piso.data_r_3346_sv2v_reg  <= \piso.data_li [3346];
      \piso.data_r_3345_sv2v_reg  <= \piso.data_li [3345];
      \piso.data_r_3344_sv2v_reg  <= \piso.data_li [3344];
      \piso.data_r_3343_sv2v_reg  <= \piso.data_li [3343];
      \piso.data_r_3342_sv2v_reg  <= \piso.data_li [3342];
      \piso.data_r_3341_sv2v_reg  <= \piso.data_li [3341];
      \piso.data_r_3340_sv2v_reg  <= \piso.data_li [3340];
      \piso.data_r_3339_sv2v_reg  <= \piso.data_li [3339];
      \piso.data_r_3338_sv2v_reg  <= \piso.data_li [3338];
      \piso.data_r_3337_sv2v_reg  <= \piso.data_li [3337];
      \piso.data_r_3336_sv2v_reg  <= \piso.data_li [3336];
      \piso.data_r_3335_sv2v_reg  <= \piso.data_li [3335];
      \piso.data_r_3334_sv2v_reg  <= \piso.data_li [3334];
      \piso.data_r_3333_sv2v_reg  <= \piso.data_li [3333];
      \piso.data_r_3332_sv2v_reg  <= \piso.data_li [3332];
      \piso.data_r_3331_sv2v_reg  <= \piso.data_li [3331];
      \piso.data_r_3330_sv2v_reg  <= \piso.data_li [3330];
      \piso.data_r_3329_sv2v_reg  <= \piso.data_li [3329];
      \piso.data_r_3328_sv2v_reg  <= \piso.data_li [3328];
      \piso.data_r_3327_sv2v_reg  <= \piso.data_li [3327];
      \piso.data_r_3326_sv2v_reg  <= \piso.data_li [3326];
      \piso.data_r_3325_sv2v_reg  <= \piso.data_li [3325];
      \piso.data_r_3324_sv2v_reg  <= \piso.data_li [3324];
      \piso.data_r_3323_sv2v_reg  <= \piso.data_li [3323];
      \piso.data_r_3322_sv2v_reg  <= \piso.data_li [3322];
      \piso.data_r_3321_sv2v_reg  <= \piso.data_li [3321];
      \piso.data_r_3320_sv2v_reg  <= \piso.data_li [3320];
      \piso.data_r_3319_sv2v_reg  <= \piso.data_li [3319];
      \piso.data_r_3318_sv2v_reg  <= \piso.data_li [3318];
      \piso.data_r_3317_sv2v_reg  <= \piso.data_li [3317];
      \piso.data_r_3316_sv2v_reg  <= \piso.data_li [3316];
      \piso.data_r_3315_sv2v_reg  <= \piso.data_li [3315];
      \piso.data_r_3314_sv2v_reg  <= \piso.data_li [3314];
      \piso.data_r_3313_sv2v_reg  <= \piso.data_li [3313];
      \piso.data_r_3312_sv2v_reg  <= \piso.data_li [3312];
      \piso.data_r_3311_sv2v_reg  <= \piso.data_li [3311];
      \piso.data_r_3310_sv2v_reg  <= \piso.data_li [3310];
      \piso.data_r_3309_sv2v_reg  <= \piso.data_li [3309];
      \piso.data_r_3308_sv2v_reg  <= \piso.data_li [3308];
      \piso.data_r_3307_sv2v_reg  <= \piso.data_li [3307];
      \piso.data_r_3306_sv2v_reg  <= \piso.data_li [3306];
      \piso.data_r_3305_sv2v_reg  <= \piso.data_li [3305];
      \piso.data_r_3304_sv2v_reg  <= \piso.data_li [3304];
      \piso.data_r_3303_sv2v_reg  <= \piso.data_li [3303];
      \piso.data_r_3302_sv2v_reg  <= \piso.data_li [3302];
      \piso.data_r_3301_sv2v_reg  <= \piso.data_li [3301];
      \piso.data_r_3300_sv2v_reg  <= \piso.data_li [3300];
      \piso.data_r_3299_sv2v_reg  <= \piso.data_li [3299];
      \piso.data_r_3298_sv2v_reg  <= \piso.data_li [3298];
      \piso.data_r_3297_sv2v_reg  <= \piso.data_li [3297];
      \piso.data_r_3296_sv2v_reg  <= \piso.data_li [3296];
      \piso.data_r_3295_sv2v_reg  <= \piso.data_li [3295];
      \piso.data_r_3294_sv2v_reg  <= \piso.data_li [3294];
      \piso.data_r_3293_sv2v_reg  <= \piso.data_li [3293];
      \piso.data_r_3292_sv2v_reg  <= \piso.data_li [3292];
      \piso.data_r_3291_sv2v_reg  <= \piso.data_li [3291];
      \piso.data_r_3290_sv2v_reg  <= \piso.data_li [3290];
      \piso.data_r_3289_sv2v_reg  <= \piso.data_li [3289];
      \piso.data_r_3288_sv2v_reg  <= \piso.data_li [3288];
      \piso.data_r_3287_sv2v_reg  <= \piso.data_li [3287];
      \piso.data_r_3286_sv2v_reg  <= \piso.data_li [3286];
      \piso.data_r_3285_sv2v_reg  <= \piso.data_li [3285];
      \piso.data_r_3284_sv2v_reg  <= \piso.data_li [3284];
      \piso.data_r_3283_sv2v_reg  <= \piso.data_li [3283];
      \piso.data_r_3282_sv2v_reg  <= \piso.data_li [3282];
      \piso.data_r_3281_sv2v_reg  <= \piso.data_li [3281];
      \piso.data_r_3280_sv2v_reg  <= \piso.data_li [3280];
      \piso.data_r_3279_sv2v_reg  <= \piso.data_li [3279];
      \piso.data_r_3278_sv2v_reg  <= \piso.data_li [3278];
      \piso.data_r_3277_sv2v_reg  <= \piso.data_li [3277];
      \piso.data_r_3276_sv2v_reg  <= \piso.data_li [3276];
      \piso.data_r_3275_sv2v_reg  <= \piso.data_li [3275];
      \piso.data_r_3274_sv2v_reg  <= \piso.data_li [3274];
      \piso.data_r_3273_sv2v_reg  <= \piso.data_li [3273];
      \piso.data_r_3272_sv2v_reg  <= \piso.data_li [3272];
      \piso.data_r_3271_sv2v_reg  <= \piso.data_li [3271];
      \piso.data_r_3270_sv2v_reg  <= \piso.data_li [3270];
      \piso.data_r_3269_sv2v_reg  <= \piso.data_li [3269];
      \piso.data_r_3268_sv2v_reg  <= \piso.data_li [3268];
      \piso.data_r_3267_sv2v_reg  <= \piso.data_li [3267];
      \piso.data_r_3266_sv2v_reg  <= \piso.data_li [3266];
      \piso.data_r_3265_sv2v_reg  <= \piso.data_li [3265];
      \piso.data_r_3264_sv2v_reg  <= \piso.data_li [3264];
      \piso.data_r_3263_sv2v_reg  <= \piso.data_li [3263];
      \piso.data_r_3262_sv2v_reg  <= \piso.data_li [3262];
      \piso.data_r_3261_sv2v_reg  <= \piso.data_li [3261];
      \piso.data_r_3260_sv2v_reg  <= \piso.data_li [3260];
      \piso.data_r_3259_sv2v_reg  <= \piso.data_li [3259];
      \piso.data_r_3258_sv2v_reg  <= \piso.data_li [3258];
      \piso.data_r_3257_sv2v_reg  <= \piso.data_li [3257];
      \piso.data_r_3256_sv2v_reg  <= \piso.data_li [3256];
      \piso.data_r_3255_sv2v_reg  <= \piso.data_li [3255];
      \piso.data_r_3254_sv2v_reg  <= \piso.data_li [3254];
      \piso.data_r_3253_sv2v_reg  <= \piso.data_li [3253];
      \piso.data_r_3252_sv2v_reg  <= \piso.data_li [3252];
      \piso.data_r_3251_sv2v_reg  <= \piso.data_li [3251];
      \piso.data_r_3250_sv2v_reg  <= \piso.data_li [3250];
      \piso.data_r_3249_sv2v_reg  <= \piso.data_li [3249];
      \piso.data_r_3248_sv2v_reg  <= \piso.data_li [3248];
      \piso.data_r_3247_sv2v_reg  <= \piso.data_li [3247];
      \piso.data_r_3246_sv2v_reg  <= \piso.data_li [3246];
      \piso.data_r_3245_sv2v_reg  <= \piso.data_li [3245];
      \piso.data_r_3244_sv2v_reg  <= \piso.data_li [3244];
      \piso.data_r_3243_sv2v_reg  <= \piso.data_li [3243];
      \piso.data_r_3242_sv2v_reg  <= \piso.data_li [3242];
      \piso.data_r_3241_sv2v_reg  <= \piso.data_li [3241];
      \piso.data_r_3240_sv2v_reg  <= \piso.data_li [3240];
      \piso.data_r_3239_sv2v_reg  <= \piso.data_li [3239];
      \piso.data_r_3238_sv2v_reg  <= \piso.data_li [3238];
      \piso.data_r_3237_sv2v_reg  <= \piso.data_li [3237];
      \piso.data_r_3236_sv2v_reg  <= \piso.data_li [3236];
      \piso.data_r_3235_sv2v_reg  <= \piso.data_li [3235];
      \piso.data_r_3234_sv2v_reg  <= \piso.data_li [3234];
      \piso.data_r_3233_sv2v_reg  <= \piso.data_li [3233];
      \piso.data_r_3232_sv2v_reg  <= \piso.data_li [3232];
      \piso.data_r_3231_sv2v_reg  <= \piso.data_li [3231];
      \piso.data_r_3230_sv2v_reg  <= \piso.data_li [3230];
      \piso.data_r_3229_sv2v_reg  <= \piso.data_li [3229];
      \piso.data_r_3228_sv2v_reg  <= \piso.data_li [3228];
      \piso.data_r_3227_sv2v_reg  <= \piso.data_li [3227];
      \piso.data_r_3226_sv2v_reg  <= \piso.data_li [3226];
      \piso.data_r_3225_sv2v_reg  <= \piso.data_li [3225];
      \piso.data_r_3224_sv2v_reg  <= \piso.data_li [3224];
      \piso.data_r_3223_sv2v_reg  <= \piso.data_li [3223];
      \piso.data_r_3222_sv2v_reg  <= \piso.data_li [3222];
      \piso.data_r_3221_sv2v_reg  <= \piso.data_li [3221];
      \piso.data_r_3220_sv2v_reg  <= \piso.data_li [3220];
      \piso.data_r_3219_sv2v_reg  <= \piso.data_li [3219];
      \piso.data_r_3218_sv2v_reg  <= \piso.data_li [3218];
      \piso.data_r_3217_sv2v_reg  <= \piso.data_li [3217];
      \piso.data_r_3216_sv2v_reg  <= \piso.data_li [3216];
      \piso.data_r_3215_sv2v_reg  <= \piso.data_li [3215];
      \piso.data_r_3214_sv2v_reg  <= \piso.data_li [3214];
      \piso.data_r_3213_sv2v_reg  <= \piso.data_li [3213];
      \piso.data_r_3212_sv2v_reg  <= \piso.data_li [3212];
      \piso.data_r_3211_sv2v_reg  <= \piso.data_li [3211];
      \piso.data_r_3210_sv2v_reg  <= \piso.data_li [3210];
      \piso.data_r_3209_sv2v_reg  <= \piso.data_li [3209];
      \piso.data_r_3208_sv2v_reg  <= \piso.data_li [3208];
      \piso.data_r_3207_sv2v_reg  <= \piso.data_li [3207];
      \piso.data_r_3206_sv2v_reg  <= \piso.data_li [3206];
      \piso.data_r_3205_sv2v_reg  <= \piso.data_li [3205];
      \piso.data_r_3204_sv2v_reg  <= \piso.data_li [3204];
      \piso.data_r_3203_sv2v_reg  <= \piso.data_li [3203];
      \piso.data_r_3202_sv2v_reg  <= \piso.data_li [3202];
      \piso.data_r_3201_sv2v_reg  <= \piso.data_li [3201];
      \piso.data_r_3200_sv2v_reg  <= \piso.data_li [3200];
      \piso.data_r_3199_sv2v_reg  <= \piso.data_li [3199];
      \piso.data_r_3198_sv2v_reg  <= \piso.data_li [3198];
      \piso.data_r_3197_sv2v_reg  <= \piso.data_li [3197];
      \piso.data_r_3196_sv2v_reg  <= \piso.data_li [3196];
      \piso.data_r_3195_sv2v_reg  <= \piso.data_li [3195];
      \piso.data_r_3194_sv2v_reg  <= \piso.data_li [3194];
      \piso.data_r_3193_sv2v_reg  <= \piso.data_li [3193];
      \piso.data_r_3192_sv2v_reg  <= \piso.data_li [3192];
      \piso.data_r_3191_sv2v_reg  <= \piso.data_li [3191];
      \piso.data_r_3190_sv2v_reg  <= \piso.data_li [3190];
      \piso.data_r_3189_sv2v_reg  <= \piso.data_li [3189];
      \piso.data_r_3188_sv2v_reg  <= \piso.data_li [3188];
      \piso.data_r_3187_sv2v_reg  <= \piso.data_li [3187];
      \piso.data_r_3186_sv2v_reg  <= \piso.data_li [3186];
      \piso.data_r_3185_sv2v_reg  <= \piso.data_li [3185];
      \piso.data_r_3184_sv2v_reg  <= \piso.data_li [3184];
      \piso.data_r_3183_sv2v_reg  <= \piso.data_li [3183];
      \piso.data_r_3182_sv2v_reg  <= \piso.data_li [3182];
      \piso.data_r_3181_sv2v_reg  <= \piso.data_li [3181];
      \piso.data_r_3180_sv2v_reg  <= \piso.data_li [3180];
      \piso.data_r_3179_sv2v_reg  <= \piso.data_li [3179];
      \piso.data_r_3178_sv2v_reg  <= \piso.data_li [3178];
      \piso.data_r_3177_sv2v_reg  <= \piso.data_li [3177];
      \piso.data_r_3176_sv2v_reg  <= \piso.data_li [3176];
      \piso.data_r_3175_sv2v_reg  <= \piso.data_li [3175];
      \piso.data_r_3174_sv2v_reg  <= \piso.data_li [3174];
      \piso.data_r_3173_sv2v_reg  <= \piso.data_li [3173];
      \piso.data_r_3172_sv2v_reg  <= \piso.data_li [3172];
      \piso.data_r_3171_sv2v_reg  <= \piso.data_li [3171];
      \piso.data_r_3170_sv2v_reg  <= \piso.data_li [3170];
      \piso.data_r_3169_sv2v_reg  <= \piso.data_li [3169];
      \piso.data_r_3168_sv2v_reg  <= \piso.data_li [3168];
      \piso.data_r_3167_sv2v_reg  <= \piso.data_li [3167];
      \piso.data_r_3166_sv2v_reg  <= \piso.data_li [3166];
      \piso.data_r_3165_sv2v_reg  <= \piso.data_li [3165];
      \piso.data_r_3164_sv2v_reg  <= \piso.data_li [3164];
      \piso.data_r_3163_sv2v_reg  <= \piso.data_li [3163];
      \piso.data_r_3162_sv2v_reg  <= \piso.data_li [3162];
      \piso.data_r_3161_sv2v_reg  <= \piso.data_li [3161];
      \piso.data_r_3160_sv2v_reg  <= \piso.data_li [3160];
      \piso.data_r_3159_sv2v_reg  <= \piso.data_li [3159];
      \piso.data_r_3158_sv2v_reg  <= \piso.data_li [3158];
      \piso.data_r_3157_sv2v_reg  <= \piso.data_li [3157];
      \piso.data_r_3156_sv2v_reg  <= \piso.data_li [3156];
      \piso.data_r_3155_sv2v_reg  <= \piso.data_li [3155];
      \piso.data_r_3154_sv2v_reg  <= \piso.data_li [3154];
      \piso.data_r_3153_sv2v_reg  <= \piso.data_li [3153];
      \piso.data_r_3152_sv2v_reg  <= \piso.data_li [3152];
      \piso.data_r_3151_sv2v_reg  <= \piso.data_li [3151];
      \piso.data_r_3150_sv2v_reg  <= \piso.data_li [3150];
      \piso.data_r_3149_sv2v_reg  <= \piso.data_li [3149];
      \piso.data_r_3148_sv2v_reg  <= \piso.data_li [3148];
      \piso.data_r_3147_sv2v_reg  <= \piso.data_li [3147];
      \piso.data_r_3146_sv2v_reg  <= \piso.data_li [3146];
      \piso.data_r_3145_sv2v_reg  <= \piso.data_li [3145];
      \piso.data_r_3144_sv2v_reg  <= \piso.data_li [3144];
      \piso.data_r_3143_sv2v_reg  <= \piso.data_li [3143];
      \piso.data_r_3142_sv2v_reg  <= \piso.data_li [3142];
      \piso.data_r_3141_sv2v_reg  <= \piso.data_li [3141];
      \piso.data_r_3140_sv2v_reg  <= \piso.data_li [3140];
      \piso.data_r_3139_sv2v_reg  <= \piso.data_li [3139];
      \piso.data_r_3138_sv2v_reg  <= \piso.data_li [3138];
      \piso.data_r_3137_sv2v_reg  <= \piso.data_li [3137];
      \piso.data_r_3136_sv2v_reg  <= \piso.data_li [3136];
      \piso.data_r_3135_sv2v_reg  <= \piso.data_li [3135];
      \piso.data_r_3134_sv2v_reg  <= \piso.data_li [3134];
      \piso.data_r_3133_sv2v_reg  <= \piso.data_li [3133];
      \piso.data_r_3132_sv2v_reg  <= \piso.data_li [3132];
      \piso.data_r_3131_sv2v_reg  <= \piso.data_li [3131];
      \piso.data_r_3130_sv2v_reg  <= \piso.data_li [3130];
      \piso.data_r_3129_sv2v_reg  <= \piso.data_li [3129];
      \piso.data_r_3128_sv2v_reg  <= \piso.data_li [3128];
      \piso.data_r_3127_sv2v_reg  <= \piso.data_li [3127];
      \piso.data_r_3126_sv2v_reg  <= \piso.data_li [3126];
      \piso.data_r_3125_sv2v_reg  <= \piso.data_li [3125];
      \piso.data_r_3124_sv2v_reg  <= \piso.data_li [3124];
      \piso.data_r_3123_sv2v_reg  <= \piso.data_li [3123];
      \piso.data_r_3122_sv2v_reg  <= \piso.data_li [3122];
      \piso.data_r_3121_sv2v_reg  <= \piso.data_li [3121];
      \piso.data_r_3120_sv2v_reg  <= \piso.data_li [3120];
      \piso.data_r_3119_sv2v_reg  <= \piso.data_li [3119];
      \piso.data_r_3118_sv2v_reg  <= \piso.data_li [3118];
      \piso.data_r_3117_sv2v_reg  <= \piso.data_li [3117];
      \piso.data_r_3116_sv2v_reg  <= \piso.data_li [3116];
      \piso.data_r_3115_sv2v_reg  <= \piso.data_li [3115];
      \piso.data_r_3114_sv2v_reg  <= \piso.data_li [3114];
      \piso.data_r_3113_sv2v_reg  <= \piso.data_li [3113];
      \piso.data_r_3112_sv2v_reg  <= \piso.data_li [3112];
      \piso.data_r_3111_sv2v_reg  <= \piso.data_li [3111];
      \piso.data_r_3110_sv2v_reg  <= \piso.data_li [3110];
      \piso.data_r_3109_sv2v_reg  <= \piso.data_li [3109];
      \piso.data_r_3108_sv2v_reg  <= \piso.data_li [3108];
      \piso.data_r_3107_sv2v_reg  <= \piso.data_li [3107];
      \piso.data_r_3106_sv2v_reg  <= \piso.data_li [3106];
      \piso.data_r_3105_sv2v_reg  <= \piso.data_li [3105];
      \piso.data_r_3104_sv2v_reg  <= \piso.data_li [3104];
      \piso.data_r_3103_sv2v_reg  <= \piso.data_li [3103];
      \piso.data_r_3102_sv2v_reg  <= \piso.data_li [3102];
      \piso.data_r_3101_sv2v_reg  <= \piso.data_li [3101];
      \piso.data_r_3100_sv2v_reg  <= \piso.data_li [3100];
      \piso.data_r_3099_sv2v_reg  <= \piso.data_li [3099];
      \piso.data_r_3098_sv2v_reg  <= \piso.data_li [3098];
      \piso.data_r_3097_sv2v_reg  <= \piso.data_li [3097];
      \piso.data_r_3096_sv2v_reg  <= \piso.data_li [3096];
      \piso.data_r_3095_sv2v_reg  <= \piso.data_li [3095];
      \piso.data_r_3094_sv2v_reg  <= \piso.data_li [3094];
      \piso.data_r_3093_sv2v_reg  <= \piso.data_li [3093];
      \piso.data_r_3092_sv2v_reg  <= \piso.data_li [3092];
      \piso.data_r_3091_sv2v_reg  <= \piso.data_li [3091];
      \piso.data_r_3090_sv2v_reg  <= \piso.data_li [3090];
      \piso.data_r_3089_sv2v_reg  <= \piso.data_li [3089];
      \piso.data_r_3088_sv2v_reg  <= \piso.data_li [3088];
      \piso.data_r_3087_sv2v_reg  <= \piso.data_li [3087];
      \piso.data_r_3086_sv2v_reg  <= \piso.data_li [3086];
      \piso.data_r_3085_sv2v_reg  <= \piso.data_li [3085];
      \piso.data_r_3084_sv2v_reg  <= \piso.data_li [3084];
      \piso.data_r_3083_sv2v_reg  <= \piso.data_li [3083];
      \piso.data_r_3082_sv2v_reg  <= \piso.data_li [3082];
      \piso.data_r_3081_sv2v_reg  <= \piso.data_li [3081];
      \piso.data_r_3080_sv2v_reg  <= \piso.data_li [3080];
      \piso.data_r_3079_sv2v_reg  <= \piso.data_li [3079];
      \piso.data_r_3078_sv2v_reg  <= \piso.data_li [3078];
      \piso.data_r_3077_sv2v_reg  <= \piso.data_li [3077];
      \piso.data_r_3076_sv2v_reg  <= \piso.data_li [3076];
      \piso.data_r_3075_sv2v_reg  <= \piso.data_li [3075];
      \piso.data_r_3074_sv2v_reg  <= \piso.data_li [3074];
      \piso.data_r_3073_sv2v_reg  <= \piso.data_li [3073];
      \piso.data_r_3072_sv2v_reg  <= \piso.data_li [3072];
      \piso.data_r_3071_sv2v_reg  <= \piso.data_li [3071];
      \piso.data_r_3070_sv2v_reg  <= \piso.data_li [3070];
      \piso.data_r_3069_sv2v_reg  <= \piso.data_li [3069];
      \piso.data_r_3068_sv2v_reg  <= \piso.data_li [3068];
      \piso.data_r_3067_sv2v_reg  <= \piso.data_li [3067];
      \piso.data_r_3066_sv2v_reg  <= \piso.data_li [3066];
      \piso.data_r_3065_sv2v_reg  <= \piso.data_li [3065];
      \piso.data_r_3064_sv2v_reg  <= \piso.data_li [3064];
      \piso.data_r_3063_sv2v_reg  <= \piso.data_li [3063];
      \piso.data_r_3062_sv2v_reg  <= \piso.data_li [3062];
      \piso.data_r_3061_sv2v_reg  <= \piso.data_li [3061];
      \piso.data_r_3060_sv2v_reg  <= \piso.data_li [3060];
      \piso.data_r_3059_sv2v_reg  <= \piso.data_li [3059];
      \piso.data_r_3058_sv2v_reg  <= \piso.data_li [3058];
      \piso.data_r_3057_sv2v_reg  <= \piso.data_li [3057];
      \piso.data_r_3056_sv2v_reg  <= \piso.data_li [3056];
      \piso.data_r_3055_sv2v_reg  <= \piso.data_li [3055];
      \piso.data_r_3054_sv2v_reg  <= \piso.data_li [3054];
      \piso.data_r_3053_sv2v_reg  <= \piso.data_li [3053];
      \piso.data_r_3052_sv2v_reg  <= \piso.data_li [3052];
      \piso.data_r_3051_sv2v_reg  <= \piso.data_li [3051];
      \piso.data_r_3050_sv2v_reg  <= \piso.data_li [3050];
      \piso.data_r_3049_sv2v_reg  <= \piso.data_li [3049];
      \piso.data_r_3048_sv2v_reg  <= \piso.data_li [3048];
      \piso.data_r_3047_sv2v_reg  <= \piso.data_li [3047];
      \piso.data_r_3046_sv2v_reg  <= \piso.data_li [3046];
      \piso.data_r_3045_sv2v_reg  <= \piso.data_li [3045];
      \piso.data_r_3044_sv2v_reg  <= \piso.data_li [3044];
      \piso.data_r_3043_sv2v_reg  <= \piso.data_li [3043];
      \piso.data_r_3042_sv2v_reg  <= \piso.data_li [3042];
      \piso.data_r_3041_sv2v_reg  <= \piso.data_li [3041];
      \piso.data_r_3040_sv2v_reg  <= \piso.data_li [3040];
      \piso.data_r_3039_sv2v_reg  <= \piso.data_li [3039];
      \piso.data_r_3038_sv2v_reg  <= \piso.data_li [3038];
      \piso.data_r_3037_sv2v_reg  <= \piso.data_li [3037];
      \piso.data_r_3036_sv2v_reg  <= \piso.data_li [3036];
      \piso.data_r_3035_sv2v_reg  <= \piso.data_li [3035];
      \piso.data_r_3034_sv2v_reg  <= \piso.data_li [3034];
      \piso.data_r_3033_sv2v_reg  <= \piso.data_li [3033];
      \piso.data_r_3032_sv2v_reg  <= \piso.data_li [3032];
      \piso.data_r_3031_sv2v_reg  <= \piso.data_li [3031];
      \piso.data_r_3030_sv2v_reg  <= \piso.data_li [3030];
      \piso.data_r_3029_sv2v_reg  <= \piso.data_li [3029];
      \piso.data_r_3028_sv2v_reg  <= \piso.data_li [3028];
      \piso.data_r_3027_sv2v_reg  <= \piso.data_li [3027];
      \piso.data_r_3026_sv2v_reg  <= \piso.data_li [3026];
      \piso.data_r_3025_sv2v_reg  <= \piso.data_li [3025];
      \piso.data_r_3024_sv2v_reg  <= \piso.data_li [3024];
      \piso.data_r_3023_sv2v_reg  <= \piso.data_li [3023];
      \piso.data_r_3022_sv2v_reg  <= \piso.data_li [3022];
      \piso.data_r_3021_sv2v_reg  <= \piso.data_li [3021];
      \piso.data_r_3020_sv2v_reg  <= \piso.data_li [3020];
      \piso.data_r_3019_sv2v_reg  <= \piso.data_li [3019];
      \piso.data_r_3018_sv2v_reg  <= \piso.data_li [3018];
      \piso.data_r_3017_sv2v_reg  <= \piso.data_li [3017];
      \piso.data_r_3016_sv2v_reg  <= \piso.data_li [3016];
      \piso.data_r_3015_sv2v_reg  <= \piso.data_li [3015];
      \piso.data_r_3014_sv2v_reg  <= \piso.data_li [3014];
      \piso.data_r_3013_sv2v_reg  <= \piso.data_li [3013];
      \piso.data_r_3012_sv2v_reg  <= \piso.data_li [3012];
      \piso.data_r_3011_sv2v_reg  <= \piso.data_li [3011];
      \piso.data_r_3010_sv2v_reg  <= \piso.data_li [3010];
      \piso.data_r_3009_sv2v_reg  <= \piso.data_li [3009];
      \piso.data_r_3008_sv2v_reg  <= \piso.data_li [3008];
      \piso.data_r_3007_sv2v_reg  <= \piso.data_li [3007];
      \piso.data_r_3006_sv2v_reg  <= \piso.data_li [3006];
      \piso.data_r_3005_sv2v_reg  <= \piso.data_li [3005];
      \piso.data_r_3004_sv2v_reg  <= \piso.data_li [3004];
      \piso.data_r_3003_sv2v_reg  <= \piso.data_li [3003];
      \piso.data_r_3002_sv2v_reg  <= \piso.data_li [3002];
      \piso.data_r_3001_sv2v_reg  <= \piso.data_li [3001];
      \piso.data_r_3000_sv2v_reg  <= \piso.data_li [3000];
      \piso.data_r_2999_sv2v_reg  <= \piso.data_li [2999];
      \piso.data_r_2998_sv2v_reg  <= \piso.data_li [2998];
      \piso.data_r_2997_sv2v_reg  <= \piso.data_li [2997];
      \piso.data_r_2996_sv2v_reg  <= \piso.data_li [2996];
      \piso.data_r_2995_sv2v_reg  <= \piso.data_li [2995];
      \piso.data_r_2994_sv2v_reg  <= \piso.data_li [2994];
      \piso.data_r_2993_sv2v_reg  <= \piso.data_li [2993];
      \piso.data_r_2992_sv2v_reg  <= \piso.data_li [2992];
      \piso.data_r_2991_sv2v_reg  <= \piso.data_li [2991];
      \piso.data_r_2990_sv2v_reg  <= \piso.data_li [2990];
      \piso.data_r_2989_sv2v_reg  <= \piso.data_li [2989];
      \piso.data_r_2988_sv2v_reg  <= \piso.data_li [2988];
      \piso.data_r_2987_sv2v_reg  <= \piso.data_li [2987];
      \piso.data_r_2986_sv2v_reg  <= \piso.data_li [2986];
      \piso.data_r_2985_sv2v_reg  <= \piso.data_li [2985];
      \piso.data_r_2984_sv2v_reg  <= \piso.data_li [2984];
      \piso.data_r_2983_sv2v_reg  <= \piso.data_li [2983];
      \piso.data_r_2982_sv2v_reg  <= \piso.data_li [2982];
      \piso.data_r_2981_sv2v_reg  <= \piso.data_li [2981];
      \piso.data_r_2980_sv2v_reg  <= \piso.data_li [2980];
      \piso.data_r_2979_sv2v_reg  <= \piso.data_li [2979];
      \piso.data_r_2978_sv2v_reg  <= \piso.data_li [2978];
      \piso.data_r_2977_sv2v_reg  <= \piso.data_li [2977];
      \piso.data_r_2976_sv2v_reg  <= \piso.data_li [2976];
      \piso.data_r_2975_sv2v_reg  <= \piso.data_li [2975];
      \piso.data_r_2974_sv2v_reg  <= \piso.data_li [2974];
      \piso.data_r_2973_sv2v_reg  <= \piso.data_li [2973];
      \piso.data_r_2972_sv2v_reg  <= \piso.data_li [2972];
      \piso.data_r_2971_sv2v_reg  <= \piso.data_li [2971];
      \piso.data_r_2970_sv2v_reg  <= \piso.data_li [2970];
      \piso.data_r_2969_sv2v_reg  <= \piso.data_li [2969];
      \piso.data_r_2968_sv2v_reg  <= \piso.data_li [2968];
      \piso.data_r_2967_sv2v_reg  <= \piso.data_li [2967];
      \piso.data_r_2966_sv2v_reg  <= \piso.data_li [2966];
      \piso.data_r_2965_sv2v_reg  <= \piso.data_li [2965];
      \piso.data_r_2964_sv2v_reg  <= \piso.data_li [2964];
      \piso.data_r_2963_sv2v_reg  <= \piso.data_li [2963];
      \piso.data_r_2962_sv2v_reg  <= \piso.data_li [2962];
      \piso.data_r_2961_sv2v_reg  <= \piso.data_li [2961];
      \piso.data_r_2960_sv2v_reg  <= \piso.data_li [2960];
      \piso.data_r_2959_sv2v_reg  <= \piso.data_li [2959];
      \piso.data_r_2958_sv2v_reg  <= \piso.data_li [2958];
      \piso.data_r_2957_sv2v_reg  <= \piso.data_li [2957];
      \piso.data_r_2956_sv2v_reg  <= \piso.data_li [2956];
      \piso.data_r_2955_sv2v_reg  <= \piso.data_li [2955];
      \piso.data_r_2954_sv2v_reg  <= \piso.data_li [2954];
      \piso.data_r_2953_sv2v_reg  <= \piso.data_li [2953];
      \piso.data_r_2952_sv2v_reg  <= \piso.data_li [2952];
      \piso.data_r_2951_sv2v_reg  <= \piso.data_li [2951];
      \piso.data_r_2950_sv2v_reg  <= \piso.data_li [2950];
      \piso.data_r_2949_sv2v_reg  <= \piso.data_li [2949];
      \piso.data_r_2948_sv2v_reg  <= \piso.data_li [2948];
      \piso.data_r_2947_sv2v_reg  <= \piso.data_li [2947];
      \piso.data_r_2946_sv2v_reg  <= \piso.data_li [2946];
      \piso.data_r_2945_sv2v_reg  <= \piso.data_li [2945];
      \piso.data_r_2944_sv2v_reg  <= \piso.data_li [2944];
      \piso.data_r_2943_sv2v_reg  <= \piso.data_li [2943];
      \piso.data_r_2942_sv2v_reg  <= \piso.data_li [2942];
      \piso.data_r_2941_sv2v_reg  <= \piso.data_li [2941];
      \piso.data_r_2940_sv2v_reg  <= \piso.data_li [2940];
      \piso.data_r_2939_sv2v_reg  <= \piso.data_li [2939];
      \piso.data_r_2938_sv2v_reg  <= \piso.data_li [2938];
      \piso.data_r_2937_sv2v_reg  <= \piso.data_li [2937];
      \piso.data_r_2936_sv2v_reg  <= \piso.data_li [2936];
      \piso.data_r_2935_sv2v_reg  <= \piso.data_li [2935];
      \piso.data_r_2934_sv2v_reg  <= \piso.data_li [2934];
      \piso.data_r_2933_sv2v_reg  <= \piso.data_li [2933];
      \piso.data_r_2932_sv2v_reg  <= \piso.data_li [2932];
      \piso.data_r_2931_sv2v_reg  <= \piso.data_li [2931];
      \piso.data_r_2930_sv2v_reg  <= \piso.data_li [2930];
      \piso.data_r_2929_sv2v_reg  <= \piso.data_li [2929];
      \piso.data_r_2928_sv2v_reg  <= \piso.data_li [2928];
      \piso.data_r_2927_sv2v_reg  <= \piso.data_li [2927];
      \piso.data_r_2926_sv2v_reg  <= \piso.data_li [2926];
      \piso.data_r_2925_sv2v_reg  <= \piso.data_li [2925];
      \piso.data_r_2924_sv2v_reg  <= \piso.data_li [2924];
      \piso.data_r_2923_sv2v_reg  <= \piso.data_li [2923];
      \piso.data_r_2922_sv2v_reg  <= \piso.data_li [2922];
      \piso.data_r_2921_sv2v_reg  <= \piso.data_li [2921];
      \piso.data_r_2920_sv2v_reg  <= \piso.data_li [2920];
      \piso.data_r_2919_sv2v_reg  <= \piso.data_li [2919];
      \piso.data_r_2918_sv2v_reg  <= \piso.data_li [2918];
      \piso.data_r_2917_sv2v_reg  <= \piso.data_li [2917];
      \piso.data_r_2916_sv2v_reg  <= \piso.data_li [2916];
      \piso.data_r_2915_sv2v_reg  <= \piso.data_li [2915];
      \piso.data_r_2914_sv2v_reg  <= \piso.data_li [2914];
      \piso.data_r_2913_sv2v_reg  <= \piso.data_li [2913];
      \piso.data_r_2912_sv2v_reg  <= \piso.data_li [2912];
      \piso.data_r_2911_sv2v_reg  <= \piso.data_li [2911];
      \piso.data_r_2910_sv2v_reg  <= \piso.data_li [2910];
      \piso.data_r_2909_sv2v_reg  <= \piso.data_li [2909];
      \piso.data_r_2908_sv2v_reg  <= \piso.data_li [2908];
      \piso.data_r_2907_sv2v_reg  <= \piso.data_li [2907];
      \piso.data_r_2906_sv2v_reg  <= \piso.data_li [2906];
      \piso.data_r_2905_sv2v_reg  <= \piso.data_li [2905];
      \piso.data_r_2904_sv2v_reg  <= \piso.data_li [2904];
      \piso.data_r_2903_sv2v_reg  <= \piso.data_li [2903];
      \piso.data_r_2902_sv2v_reg  <= \piso.data_li [2902];
      \piso.data_r_2901_sv2v_reg  <= \piso.data_li [2901];
      \piso.data_r_2900_sv2v_reg  <= \piso.data_li [2900];
      \piso.data_r_2899_sv2v_reg  <= \piso.data_li [2899];
      \piso.data_r_2898_sv2v_reg  <= \piso.data_li [2898];
      \piso.data_r_2897_sv2v_reg  <= \piso.data_li [2897];
      \piso.data_r_2896_sv2v_reg  <= \piso.data_li [2896];
      \piso.data_r_2895_sv2v_reg  <= \piso.data_li [2895];
      \piso.data_r_2894_sv2v_reg  <= \piso.data_li [2894];
      \piso.data_r_2893_sv2v_reg  <= \piso.data_li [2893];
      \piso.data_r_2892_sv2v_reg  <= \piso.data_li [2892];
      \piso.data_r_2891_sv2v_reg  <= \piso.data_li [2891];
      \piso.data_r_2890_sv2v_reg  <= \piso.data_li [2890];
      \piso.data_r_2889_sv2v_reg  <= \piso.data_li [2889];
      \piso.data_r_2888_sv2v_reg  <= \piso.data_li [2888];
      \piso.data_r_2887_sv2v_reg  <= \piso.data_li [2887];
      \piso.data_r_2886_sv2v_reg  <= \piso.data_li [2886];
      \piso.data_r_2885_sv2v_reg  <= \piso.data_li [2885];
      \piso.data_r_2884_sv2v_reg  <= \piso.data_li [2884];
      \piso.data_r_2883_sv2v_reg  <= \piso.data_li [2883];
      \piso.data_r_2882_sv2v_reg  <= \piso.data_li [2882];
      \piso.data_r_2881_sv2v_reg  <= \piso.data_li [2881];
      \piso.data_r_2880_sv2v_reg  <= \piso.data_li [2880];
      \piso.data_r_2879_sv2v_reg  <= \piso.data_li [2879];
      \piso.data_r_2878_sv2v_reg  <= \piso.data_li [2878];
      \piso.data_r_2877_sv2v_reg  <= \piso.data_li [2877];
      \piso.data_r_2876_sv2v_reg  <= \piso.data_li [2876];
      \piso.data_r_2875_sv2v_reg  <= \piso.data_li [2875];
      \piso.data_r_2874_sv2v_reg  <= \piso.data_li [2874];
      \piso.data_r_2873_sv2v_reg  <= \piso.data_li [2873];
      \piso.data_r_2872_sv2v_reg  <= \piso.data_li [2872];
      \piso.data_r_2871_sv2v_reg  <= \piso.data_li [2871];
      \piso.data_r_2870_sv2v_reg  <= \piso.data_li [2870];
      \piso.data_r_2869_sv2v_reg  <= \piso.data_li [2869];
      \piso.data_r_2868_sv2v_reg  <= \piso.data_li [2868];
      \piso.data_r_2867_sv2v_reg  <= \piso.data_li [2867];
      \piso.data_r_2866_sv2v_reg  <= \piso.data_li [2866];
      \piso.data_r_2865_sv2v_reg  <= \piso.data_li [2865];
      \piso.data_r_2864_sv2v_reg  <= \piso.data_li [2864];
      \piso.data_r_2863_sv2v_reg  <= \piso.data_li [2863];
      \piso.data_r_2862_sv2v_reg  <= \piso.data_li [2862];
      \piso.data_r_2861_sv2v_reg  <= \piso.data_li [2861];
      \piso.data_r_2860_sv2v_reg  <= \piso.data_li [2860];
      \piso.data_r_2859_sv2v_reg  <= \piso.data_li [2859];
      \piso.data_r_2858_sv2v_reg  <= \piso.data_li [2858];
      \piso.data_r_2857_sv2v_reg  <= \piso.data_li [2857];
      \piso.data_r_2856_sv2v_reg  <= \piso.data_li [2856];
      \piso.data_r_2855_sv2v_reg  <= \piso.data_li [2855];
      \piso.data_r_2854_sv2v_reg  <= \piso.data_li [2854];
      \piso.data_r_2853_sv2v_reg  <= \piso.data_li [2853];
      \piso.data_r_2852_sv2v_reg  <= \piso.data_li [2852];
      \piso.data_r_2851_sv2v_reg  <= \piso.data_li [2851];
      \piso.data_r_2850_sv2v_reg  <= \piso.data_li [2850];
      \piso.data_r_2849_sv2v_reg  <= \piso.data_li [2849];
      \piso.data_r_2848_sv2v_reg  <= \piso.data_li [2848];
      \piso.data_r_2847_sv2v_reg  <= \piso.data_li [2847];
      \piso.data_r_2846_sv2v_reg  <= \piso.data_li [2846];
      \piso.data_r_2845_sv2v_reg  <= \piso.data_li [2845];
      \piso.data_r_2844_sv2v_reg  <= \piso.data_li [2844];
      \piso.data_r_2843_sv2v_reg  <= \piso.data_li [2843];
      \piso.data_r_2842_sv2v_reg  <= \piso.data_li [2842];
      \piso.data_r_2841_sv2v_reg  <= \piso.data_li [2841];
      \piso.data_r_2840_sv2v_reg  <= \piso.data_li [2840];
      \piso.data_r_2839_sv2v_reg  <= \piso.data_li [2839];
      \piso.data_r_2838_sv2v_reg  <= \piso.data_li [2838];
      \piso.data_r_2837_sv2v_reg  <= \piso.data_li [2837];
      \piso.data_r_2836_sv2v_reg  <= \piso.data_li [2836];
      \piso.data_r_2835_sv2v_reg  <= \piso.data_li [2835];
      \piso.data_r_2834_sv2v_reg  <= \piso.data_li [2834];
      \piso.data_r_2833_sv2v_reg  <= \piso.data_li [2833];
      \piso.data_r_2832_sv2v_reg  <= \piso.data_li [2832];
      \piso.data_r_2831_sv2v_reg  <= \piso.data_li [2831];
      \piso.data_r_2830_sv2v_reg  <= \piso.data_li [2830];
      \piso.data_r_2829_sv2v_reg  <= \piso.data_li [2829];
      \piso.data_r_2828_sv2v_reg  <= \piso.data_li [2828];
      \piso.data_r_2827_sv2v_reg  <= \piso.data_li [2827];
      \piso.data_r_2826_sv2v_reg  <= \piso.data_li [2826];
      \piso.data_r_2825_sv2v_reg  <= \piso.data_li [2825];
      \piso.data_r_2824_sv2v_reg  <= \piso.data_li [2824];
      \piso.data_r_2823_sv2v_reg  <= \piso.data_li [2823];
      \piso.data_r_2822_sv2v_reg  <= \piso.data_li [2822];
      \piso.data_r_2821_sv2v_reg  <= \piso.data_li [2821];
      \piso.data_r_2820_sv2v_reg  <= \piso.data_li [2820];
      \piso.data_r_2819_sv2v_reg  <= \piso.data_li [2819];
      \piso.data_r_2818_sv2v_reg  <= \piso.data_li [2818];
      \piso.data_r_2817_sv2v_reg  <= \piso.data_li [2817];
      \piso.data_r_2816_sv2v_reg  <= \piso.data_li [2816];
      \piso.data_r_2815_sv2v_reg  <= \piso.data_li [2815];
      \piso.data_r_2814_sv2v_reg  <= \piso.data_li [2814];
      \piso.data_r_2813_sv2v_reg  <= \piso.data_li [2813];
      \piso.data_r_2812_sv2v_reg  <= \piso.data_li [2812];
      \piso.data_r_2811_sv2v_reg  <= \piso.data_li [2811];
      \piso.data_r_2810_sv2v_reg  <= \piso.data_li [2810];
      \piso.data_r_2809_sv2v_reg  <= \piso.data_li [2809];
      \piso.data_r_2808_sv2v_reg  <= \piso.data_li [2808];
      \piso.data_r_2807_sv2v_reg  <= \piso.data_li [2807];
      \piso.data_r_2806_sv2v_reg  <= \piso.data_li [2806];
      \piso.data_r_2805_sv2v_reg  <= \piso.data_li [2805];
      \piso.data_r_2804_sv2v_reg  <= \piso.data_li [2804];
      \piso.data_r_2803_sv2v_reg  <= \piso.data_li [2803];
      \piso.data_r_2802_sv2v_reg  <= \piso.data_li [2802];
      \piso.data_r_2801_sv2v_reg  <= \piso.data_li [2801];
      \piso.data_r_2800_sv2v_reg  <= \piso.data_li [2800];
      \piso.data_r_2799_sv2v_reg  <= \piso.data_li [2799];
      \piso.data_r_2798_sv2v_reg  <= \piso.data_li [2798];
      \piso.data_r_2797_sv2v_reg  <= \piso.data_li [2797];
      \piso.data_r_2796_sv2v_reg  <= \piso.data_li [2796];
      \piso.data_r_2795_sv2v_reg  <= \piso.data_li [2795];
      \piso.data_r_2794_sv2v_reg  <= \piso.data_li [2794];
      \piso.data_r_2793_sv2v_reg  <= \piso.data_li [2793];
      \piso.data_r_2792_sv2v_reg  <= \piso.data_li [2792];
      \piso.data_r_2791_sv2v_reg  <= \piso.data_li [2791];
      \piso.data_r_2790_sv2v_reg  <= \piso.data_li [2790];
      \piso.data_r_2789_sv2v_reg  <= \piso.data_li [2789];
      \piso.data_r_2788_sv2v_reg  <= \piso.data_li [2788];
      \piso.data_r_2787_sv2v_reg  <= \piso.data_li [2787];
      \piso.data_r_2786_sv2v_reg  <= \piso.data_li [2786];
      \piso.data_r_2785_sv2v_reg  <= \piso.data_li [2785];
      \piso.data_r_2784_sv2v_reg  <= \piso.data_li [2784];
      \piso.data_r_2783_sv2v_reg  <= \piso.data_li [2783];
      \piso.data_r_2782_sv2v_reg  <= \piso.data_li [2782];
      \piso.data_r_2781_sv2v_reg  <= \piso.data_li [2781];
      \piso.data_r_2780_sv2v_reg  <= \piso.data_li [2780];
      \piso.data_r_2779_sv2v_reg  <= \piso.data_li [2779];
      \piso.data_r_2778_sv2v_reg  <= \piso.data_li [2778];
      \piso.data_r_2777_sv2v_reg  <= \piso.data_li [2777];
      \piso.data_r_2776_sv2v_reg  <= \piso.data_li [2776];
      \piso.data_r_2775_sv2v_reg  <= \piso.data_li [2775];
      \piso.data_r_2774_sv2v_reg  <= \piso.data_li [2774];
      \piso.data_r_2773_sv2v_reg  <= \piso.data_li [2773];
      \piso.data_r_2772_sv2v_reg  <= \piso.data_li [2772];
      \piso.data_r_2771_sv2v_reg  <= \piso.data_li [2771];
      \piso.data_r_2770_sv2v_reg  <= \piso.data_li [2770];
      \piso.data_r_2769_sv2v_reg  <= \piso.data_li [2769];
      \piso.data_r_2768_sv2v_reg  <= \piso.data_li [2768];
      \piso.data_r_2767_sv2v_reg  <= \piso.data_li [2767];
      \piso.data_r_2766_sv2v_reg  <= \piso.data_li [2766];
      \piso.data_r_2765_sv2v_reg  <= \piso.data_li [2765];
      \piso.data_r_2764_sv2v_reg  <= \piso.data_li [2764];
      \piso.data_r_2763_sv2v_reg  <= \piso.data_li [2763];
      \piso.data_r_2762_sv2v_reg  <= \piso.data_li [2762];
      \piso.data_r_2761_sv2v_reg  <= \piso.data_li [2761];
      \piso.data_r_2760_sv2v_reg  <= \piso.data_li [2760];
      \piso.data_r_2759_sv2v_reg  <= \piso.data_li [2759];
      \piso.data_r_2758_sv2v_reg  <= \piso.data_li [2758];
      \piso.data_r_2757_sv2v_reg  <= \piso.data_li [2757];
      \piso.data_r_2756_sv2v_reg  <= \piso.data_li [2756];
      \piso.data_r_2755_sv2v_reg  <= \piso.data_li [2755];
      \piso.data_r_2754_sv2v_reg  <= \piso.data_li [2754];
      \piso.data_r_2753_sv2v_reg  <= \piso.data_li [2753];
      \piso.data_r_2752_sv2v_reg  <= \piso.data_li [2752];
      \piso.data_r_2751_sv2v_reg  <= \piso.data_li [2751];
      \piso.data_r_2750_sv2v_reg  <= \piso.data_li [2750];
      \piso.data_r_2749_sv2v_reg  <= \piso.data_li [2749];
      \piso.data_r_2748_sv2v_reg  <= \piso.data_li [2748];
      \piso.data_r_2747_sv2v_reg  <= \piso.data_li [2747];
      \piso.data_r_2746_sv2v_reg  <= \piso.data_li [2746];
      \piso.data_r_2745_sv2v_reg  <= \piso.data_li [2745];
      \piso.data_r_2744_sv2v_reg  <= \piso.data_li [2744];
      \piso.data_r_2743_sv2v_reg  <= \piso.data_li [2743];
      \piso.data_r_2742_sv2v_reg  <= \piso.data_li [2742];
      \piso.data_r_2741_sv2v_reg  <= \piso.data_li [2741];
      \piso.data_r_2740_sv2v_reg  <= \piso.data_li [2740];
      \piso.data_r_2739_sv2v_reg  <= \piso.data_li [2739];
      \piso.data_r_2738_sv2v_reg  <= \piso.data_li [2738];
      \piso.data_r_2737_sv2v_reg  <= \piso.data_li [2737];
      \piso.data_r_2736_sv2v_reg  <= \piso.data_li [2736];
      \piso.data_r_2735_sv2v_reg  <= \piso.data_li [2735];
      \piso.data_r_2734_sv2v_reg  <= \piso.data_li [2734];
      \piso.data_r_2733_sv2v_reg  <= \piso.data_li [2733];
      \piso.data_r_2732_sv2v_reg  <= \piso.data_li [2732];
      \piso.data_r_2731_sv2v_reg  <= \piso.data_li [2731];
      \piso.data_r_2730_sv2v_reg  <= \piso.data_li [2730];
      \piso.data_r_2729_sv2v_reg  <= \piso.data_li [2729];
      \piso.data_r_2728_sv2v_reg  <= \piso.data_li [2728];
      \piso.data_r_2727_sv2v_reg  <= \piso.data_li [2727];
      \piso.data_r_2726_sv2v_reg  <= \piso.data_li [2726];
      \piso.data_r_2725_sv2v_reg  <= \piso.data_li [2725];
      \piso.data_r_2724_sv2v_reg  <= \piso.data_li [2724];
      \piso.data_r_2723_sv2v_reg  <= \piso.data_li [2723];
      \piso.data_r_2722_sv2v_reg  <= \piso.data_li [2722];
      \piso.data_r_2721_sv2v_reg  <= \piso.data_li [2721];
      \piso.data_r_2720_sv2v_reg  <= \piso.data_li [2720];
      \piso.data_r_2719_sv2v_reg  <= \piso.data_li [2719];
      \piso.data_r_2718_sv2v_reg  <= \piso.data_li [2718];
      \piso.data_r_2717_sv2v_reg  <= \piso.data_li [2717];
      \piso.data_r_2716_sv2v_reg  <= \piso.data_li [2716];
      \piso.data_r_2715_sv2v_reg  <= \piso.data_li [2715];
      \piso.data_r_2714_sv2v_reg  <= \piso.data_li [2714];
      \piso.data_r_2713_sv2v_reg  <= \piso.data_li [2713];
      \piso.data_r_2712_sv2v_reg  <= \piso.data_li [2712];
      \piso.data_r_2711_sv2v_reg  <= \piso.data_li [2711];
      \piso.data_r_2710_sv2v_reg  <= \piso.data_li [2710];
      \piso.data_r_2709_sv2v_reg  <= \piso.data_li [2709];
      \piso.data_r_2708_sv2v_reg  <= \piso.data_li [2708];
      \piso.data_r_2707_sv2v_reg  <= \piso.data_li [2707];
      \piso.data_r_2706_sv2v_reg  <= \piso.data_li [2706];
      \piso.data_r_2705_sv2v_reg  <= \piso.data_li [2705];
      \piso.data_r_2704_sv2v_reg  <= \piso.data_li [2704];
      \piso.data_r_2703_sv2v_reg  <= \piso.data_li [2703];
      \piso.data_r_2702_sv2v_reg  <= \piso.data_li [2702];
      \piso.data_r_2701_sv2v_reg  <= \piso.data_li [2701];
      \piso.data_r_2700_sv2v_reg  <= \piso.data_li [2700];
      \piso.data_r_2699_sv2v_reg  <= \piso.data_li [2699];
      \piso.data_r_2698_sv2v_reg  <= \piso.data_li [2698];
      \piso.data_r_2697_sv2v_reg  <= \piso.data_li [2697];
      \piso.data_r_2696_sv2v_reg  <= \piso.data_li [2696];
      \piso.data_r_2695_sv2v_reg  <= \piso.data_li [2695];
      \piso.data_r_2694_sv2v_reg  <= \piso.data_li [2694];
      \piso.data_r_2693_sv2v_reg  <= \piso.data_li [2693];
      \piso.data_r_2692_sv2v_reg  <= \piso.data_li [2692];
      \piso.data_r_2691_sv2v_reg  <= \piso.data_li [2691];
      \piso.data_r_2690_sv2v_reg  <= \piso.data_li [2690];
      \piso.data_r_2689_sv2v_reg  <= \piso.data_li [2689];
      \piso.data_r_2688_sv2v_reg  <= \piso.data_li [2688];
      \piso.data_r_2687_sv2v_reg  <= \piso.data_li [2687];
      \piso.data_r_2686_sv2v_reg  <= \piso.data_li [2686];
      \piso.data_r_2685_sv2v_reg  <= \piso.data_li [2685];
      \piso.data_r_2684_sv2v_reg  <= \piso.data_li [2684];
      \piso.data_r_2683_sv2v_reg  <= \piso.data_li [2683];
      \piso.data_r_2682_sv2v_reg  <= \piso.data_li [2682];
      \piso.data_r_2681_sv2v_reg  <= \piso.data_li [2681];
      \piso.data_r_2680_sv2v_reg  <= \piso.data_li [2680];
      \piso.data_r_2679_sv2v_reg  <= \piso.data_li [2679];
      \piso.data_r_2678_sv2v_reg  <= \piso.data_li [2678];
      \piso.data_r_2677_sv2v_reg  <= \piso.data_li [2677];
      \piso.data_r_2676_sv2v_reg  <= \piso.data_li [2676];
      \piso.data_r_2675_sv2v_reg  <= \piso.data_li [2675];
      \piso.data_r_2674_sv2v_reg  <= \piso.data_li [2674];
      \piso.data_r_2673_sv2v_reg  <= \piso.data_li [2673];
      \piso.data_r_2672_sv2v_reg  <= \piso.data_li [2672];
      \piso.data_r_2671_sv2v_reg  <= \piso.data_li [2671];
      \piso.data_r_2670_sv2v_reg  <= \piso.data_li [2670];
      \piso.data_r_2669_sv2v_reg  <= \piso.data_li [2669];
      \piso.data_r_2668_sv2v_reg  <= \piso.data_li [2668];
      \piso.data_r_2667_sv2v_reg  <= \piso.data_li [2667];
      \piso.data_r_2666_sv2v_reg  <= \piso.data_li [2666];
      \piso.data_r_2665_sv2v_reg  <= \piso.data_li [2665];
      \piso.data_r_2664_sv2v_reg  <= \piso.data_li [2664];
      \piso.data_r_2663_sv2v_reg  <= \piso.data_li [2663];
      \piso.data_r_2662_sv2v_reg  <= \piso.data_li [2662];
      \piso.data_r_2661_sv2v_reg  <= \piso.data_li [2661];
      \piso.data_r_2660_sv2v_reg  <= \piso.data_li [2660];
      \piso.data_r_2659_sv2v_reg  <= \piso.data_li [2659];
      \piso.data_r_2658_sv2v_reg  <= \piso.data_li [2658];
      \piso.data_r_2657_sv2v_reg  <= \piso.data_li [2657];
      \piso.data_r_2656_sv2v_reg  <= \piso.data_li [2656];
      \piso.data_r_2655_sv2v_reg  <= \piso.data_li [2655];
      \piso.data_r_2654_sv2v_reg  <= \piso.data_li [2654];
      \piso.data_r_2653_sv2v_reg  <= \piso.data_li [2653];
      \piso.data_r_2652_sv2v_reg  <= \piso.data_li [2652];
      \piso.data_r_2651_sv2v_reg  <= \piso.data_li [2651];
      \piso.data_r_2650_sv2v_reg  <= \piso.data_li [2650];
      \piso.data_r_2649_sv2v_reg  <= \piso.data_li [2649];
      \piso.data_r_2648_sv2v_reg  <= \piso.data_li [2648];
      \piso.data_r_2647_sv2v_reg  <= \piso.data_li [2647];
      \piso.data_r_2646_sv2v_reg  <= \piso.data_li [2646];
      \piso.data_r_2645_sv2v_reg  <= \piso.data_li [2645];
      \piso.data_r_2644_sv2v_reg  <= \piso.data_li [2644];
      \piso.data_r_2643_sv2v_reg  <= \piso.data_li [2643];
      \piso.data_r_2642_sv2v_reg  <= \piso.data_li [2642];
      \piso.data_r_2641_sv2v_reg  <= \piso.data_li [2641];
      \piso.data_r_2640_sv2v_reg  <= \piso.data_li [2640];
      \piso.data_r_2639_sv2v_reg  <= \piso.data_li [2639];
      \piso.data_r_2638_sv2v_reg  <= \piso.data_li [2638];
      \piso.data_r_2637_sv2v_reg  <= \piso.data_li [2637];
      \piso.data_r_2636_sv2v_reg  <= \piso.data_li [2636];
      \piso.data_r_2635_sv2v_reg  <= \piso.data_li [2635];
      \piso.data_r_2634_sv2v_reg  <= \piso.data_li [2634];
      \piso.data_r_2633_sv2v_reg  <= \piso.data_li [2633];
      \piso.data_r_2632_sv2v_reg  <= \piso.data_li [2632];
      \piso.data_r_2631_sv2v_reg  <= \piso.data_li [2631];
      \piso.data_r_2630_sv2v_reg  <= \piso.data_li [2630];
      \piso.data_r_2629_sv2v_reg  <= \piso.data_li [2629];
      \piso.data_r_2628_sv2v_reg  <= \piso.data_li [2628];
      \piso.data_r_2627_sv2v_reg  <= \piso.data_li [2627];
      \piso.data_r_2626_sv2v_reg  <= \piso.data_li [2626];
      \piso.data_r_2625_sv2v_reg  <= \piso.data_li [2625];
      \piso.data_r_2624_sv2v_reg  <= \piso.data_li [2624];
      \piso.data_r_2623_sv2v_reg  <= \piso.data_li [2623];
      \piso.data_r_2622_sv2v_reg  <= \piso.data_li [2622];
      \piso.data_r_2621_sv2v_reg  <= \piso.data_li [2621];
      \piso.data_r_2620_sv2v_reg  <= \piso.data_li [2620];
      \piso.data_r_2619_sv2v_reg  <= \piso.data_li [2619];
      \piso.data_r_2618_sv2v_reg  <= \piso.data_li [2618];
      \piso.data_r_2617_sv2v_reg  <= \piso.data_li [2617];
      \piso.data_r_2616_sv2v_reg  <= \piso.data_li [2616];
      \piso.data_r_2615_sv2v_reg  <= \piso.data_li [2615];
      \piso.data_r_2614_sv2v_reg  <= \piso.data_li [2614];
      \piso.data_r_2613_sv2v_reg  <= \piso.data_li [2613];
      \piso.data_r_2612_sv2v_reg  <= \piso.data_li [2612];
      \piso.data_r_2611_sv2v_reg  <= \piso.data_li [2611];
      \piso.data_r_2610_sv2v_reg  <= \piso.data_li [2610];
      \piso.data_r_2609_sv2v_reg  <= \piso.data_li [2609];
      \piso.data_r_2608_sv2v_reg  <= \piso.data_li [2608];
      \piso.data_r_2607_sv2v_reg  <= \piso.data_li [2607];
      \piso.data_r_2606_sv2v_reg  <= \piso.data_li [2606];
      \piso.data_r_2605_sv2v_reg  <= \piso.data_li [2605];
      \piso.data_r_2604_sv2v_reg  <= \piso.data_li [2604];
      \piso.data_r_2603_sv2v_reg  <= \piso.data_li [2603];
      \piso.data_r_2602_sv2v_reg  <= \piso.data_li [2602];
      \piso.data_r_2601_sv2v_reg  <= \piso.data_li [2601];
      \piso.data_r_2600_sv2v_reg  <= \piso.data_li [2600];
      \piso.data_r_2599_sv2v_reg  <= \piso.data_li [2599];
      \piso.data_r_2598_sv2v_reg  <= \piso.data_li [2598];
      \piso.data_r_2597_sv2v_reg  <= \piso.data_li [2597];
      \piso.data_r_2596_sv2v_reg  <= \piso.data_li [2596];
      \piso.data_r_2595_sv2v_reg  <= \piso.data_li [2595];
      \piso.data_r_2594_sv2v_reg  <= \piso.data_li [2594];
      \piso.data_r_2593_sv2v_reg  <= \piso.data_li [2593];
      \piso.data_r_2592_sv2v_reg  <= \piso.data_li [2592];
      \piso.data_r_2591_sv2v_reg  <= \piso.data_li [2591];
      \piso.data_r_2590_sv2v_reg  <= \piso.data_li [2590];
      \piso.data_r_2589_sv2v_reg  <= \piso.data_li [2589];
      \piso.data_r_2588_sv2v_reg  <= \piso.data_li [2588];
      \piso.data_r_2587_sv2v_reg  <= \piso.data_li [2587];
      \piso.data_r_2586_sv2v_reg  <= \piso.data_li [2586];
      \piso.data_r_2585_sv2v_reg  <= \piso.data_li [2585];
      \piso.data_r_2584_sv2v_reg  <= \piso.data_li [2584];
      \piso.data_r_2583_sv2v_reg  <= \piso.data_li [2583];
      \piso.data_r_2582_sv2v_reg  <= \piso.data_li [2582];
      \piso.data_r_2581_sv2v_reg  <= \piso.data_li [2581];
      \piso.data_r_2580_sv2v_reg  <= \piso.data_li [2580];
      \piso.data_r_2579_sv2v_reg  <= \piso.data_li [2579];
      \piso.data_r_2578_sv2v_reg  <= \piso.data_li [2578];
      \piso.data_r_2577_sv2v_reg  <= \piso.data_li [2577];
      \piso.data_r_2576_sv2v_reg  <= \piso.data_li [2576];
      \piso.data_r_2575_sv2v_reg  <= \piso.data_li [2575];
      \piso.data_r_2574_sv2v_reg  <= \piso.data_li [2574];
      \piso.data_r_2573_sv2v_reg  <= \piso.data_li [2573];
      \piso.data_r_2572_sv2v_reg  <= \piso.data_li [2572];
      \piso.data_r_2571_sv2v_reg  <= \piso.data_li [2571];
      \piso.data_r_2570_sv2v_reg  <= \piso.data_li [2570];
      \piso.data_r_2569_sv2v_reg  <= \piso.data_li [2569];
      \piso.data_r_2568_sv2v_reg  <= \piso.data_li [2568];
      \piso.data_r_2567_sv2v_reg  <= \piso.data_li [2567];
      \piso.data_r_2566_sv2v_reg  <= \piso.data_li [2566];
      \piso.data_r_2565_sv2v_reg  <= \piso.data_li [2565];
      \piso.data_r_2564_sv2v_reg  <= \piso.data_li [2564];
      \piso.data_r_2563_sv2v_reg  <= \piso.data_li [2563];
      \piso.data_r_2562_sv2v_reg  <= \piso.data_li [2562];
      \piso.data_r_2561_sv2v_reg  <= \piso.data_li [2561];
      \piso.data_r_2560_sv2v_reg  <= \piso.data_li [2560];
      \piso.data_r_2559_sv2v_reg  <= \piso.data_li [2559];
      \piso.data_r_2558_sv2v_reg  <= \piso.data_li [2558];
      \piso.data_r_2557_sv2v_reg  <= \piso.data_li [2557];
      \piso.data_r_2556_sv2v_reg  <= \piso.data_li [2556];
      \piso.data_r_2555_sv2v_reg  <= \piso.data_li [2555];
      \piso.data_r_2554_sv2v_reg  <= \piso.data_li [2554];
      \piso.data_r_2553_sv2v_reg  <= \piso.data_li [2553];
      \piso.data_r_2552_sv2v_reg  <= \piso.data_li [2552];
      \piso.data_r_2551_sv2v_reg  <= \piso.data_li [2551];
      \piso.data_r_2550_sv2v_reg  <= \piso.data_li [2550];
      \piso.data_r_2549_sv2v_reg  <= \piso.data_li [2549];
      \piso.data_r_2548_sv2v_reg  <= \piso.data_li [2548];
      \piso.data_r_2547_sv2v_reg  <= \piso.data_li [2547];
      \piso.data_r_2546_sv2v_reg  <= \piso.data_li [2546];
      \piso.data_r_2545_sv2v_reg  <= \piso.data_li [2545];
      \piso.data_r_2544_sv2v_reg  <= \piso.data_li [2544];
      \piso.data_r_2543_sv2v_reg  <= \piso.data_li [2543];
      \piso.data_r_2542_sv2v_reg  <= \piso.data_li [2542];
      \piso.data_r_2541_sv2v_reg  <= \piso.data_li [2541];
      \piso.data_r_2540_sv2v_reg  <= \piso.data_li [2540];
      \piso.data_r_2539_sv2v_reg  <= \piso.data_li [2539];
      \piso.data_r_2538_sv2v_reg  <= \piso.data_li [2538];
      \piso.data_r_2537_sv2v_reg  <= \piso.data_li [2537];
      \piso.data_r_2536_sv2v_reg  <= \piso.data_li [2536];
      \piso.data_r_2535_sv2v_reg  <= \piso.data_li [2535];
      \piso.data_r_2534_sv2v_reg  <= \piso.data_li [2534];
      \piso.data_r_2533_sv2v_reg  <= \piso.data_li [2533];
      \piso.data_r_2532_sv2v_reg  <= \piso.data_li [2532];
      \piso.data_r_2531_sv2v_reg  <= \piso.data_li [2531];
      \piso.data_r_2530_sv2v_reg  <= \piso.data_li [2530];
      \piso.data_r_2529_sv2v_reg  <= \piso.data_li [2529];
      \piso.data_r_2528_sv2v_reg  <= \piso.data_li [2528];
      \piso.data_r_2527_sv2v_reg  <= \piso.data_li [2527];
      \piso.data_r_2526_sv2v_reg  <= \piso.data_li [2526];
      \piso.data_r_2525_sv2v_reg  <= \piso.data_li [2525];
      \piso.data_r_2524_sv2v_reg  <= \piso.data_li [2524];
      \piso.data_r_2523_sv2v_reg  <= \piso.data_li [2523];
      \piso.data_r_2522_sv2v_reg  <= \piso.data_li [2522];
      \piso.data_r_2521_sv2v_reg  <= \piso.data_li [2521];
      \piso.data_r_2520_sv2v_reg  <= \piso.data_li [2520];
      \piso.data_r_2519_sv2v_reg  <= \piso.data_li [2519];
      \piso.data_r_2518_sv2v_reg  <= \piso.data_li [2518];
      \piso.data_r_2517_sv2v_reg  <= \piso.data_li [2517];
      \piso.data_r_2516_sv2v_reg  <= \piso.data_li [2516];
      \piso.data_r_2515_sv2v_reg  <= \piso.data_li [2515];
      \piso.data_r_2514_sv2v_reg  <= \piso.data_li [2514];
      \piso.data_r_2513_sv2v_reg  <= \piso.data_li [2513];
      \piso.data_r_2512_sv2v_reg  <= \piso.data_li [2512];
      \piso.data_r_2511_sv2v_reg  <= \piso.data_li [2511];
      \piso.data_r_2510_sv2v_reg  <= \piso.data_li [2510];
      \piso.data_r_2509_sv2v_reg  <= \piso.data_li [2509];
      \piso.data_r_2508_sv2v_reg  <= \piso.data_li [2508];
      \piso.data_r_2507_sv2v_reg  <= \piso.data_li [2507];
      \piso.data_r_2506_sv2v_reg  <= \piso.data_li [2506];
      \piso.data_r_2505_sv2v_reg  <= \piso.data_li [2505];
      \piso.data_r_2504_sv2v_reg  <= \piso.data_li [2504];
      \piso.data_r_2503_sv2v_reg  <= \piso.data_li [2503];
      \piso.data_r_2502_sv2v_reg  <= \piso.data_li [2502];
      \piso.data_r_2501_sv2v_reg  <= \piso.data_li [2501];
      \piso.data_r_2500_sv2v_reg  <= \piso.data_li [2500];
      \piso.data_r_2499_sv2v_reg  <= \piso.data_li [2499];
      \piso.data_r_2498_sv2v_reg  <= \piso.data_li [2498];
      \piso.data_r_2497_sv2v_reg  <= \piso.data_li [2497];
      \piso.data_r_2496_sv2v_reg  <= \piso.data_li [2496];
      \piso.data_r_2495_sv2v_reg  <= \piso.data_li [2495];
      \piso.data_r_2494_sv2v_reg  <= \piso.data_li [2494];
      \piso.data_r_2493_sv2v_reg  <= \piso.data_li [2493];
      \piso.data_r_2492_sv2v_reg  <= \piso.data_li [2492];
      \piso.data_r_2491_sv2v_reg  <= \piso.data_li [2491];
      \piso.data_r_2490_sv2v_reg  <= \piso.data_li [2490];
      \piso.data_r_2489_sv2v_reg  <= \piso.data_li [2489];
      \piso.data_r_2488_sv2v_reg  <= \piso.data_li [2488];
      \piso.data_r_2487_sv2v_reg  <= \piso.data_li [2487];
      \piso.data_r_2486_sv2v_reg  <= \piso.data_li [2486];
      \piso.data_r_2485_sv2v_reg  <= \piso.data_li [2485];
      \piso.data_r_2484_sv2v_reg  <= \piso.data_li [2484];
      \piso.data_r_2483_sv2v_reg  <= \piso.data_li [2483];
      \piso.data_r_2482_sv2v_reg  <= \piso.data_li [2482];
      \piso.data_r_2481_sv2v_reg  <= \piso.data_li [2481];
      \piso.data_r_2480_sv2v_reg  <= \piso.data_li [2480];
      \piso.data_r_2479_sv2v_reg  <= \piso.data_li [2479];
      \piso.data_r_2478_sv2v_reg  <= \piso.data_li [2478];
      \piso.data_r_2477_sv2v_reg  <= \piso.data_li [2477];
      \piso.data_r_2476_sv2v_reg  <= \piso.data_li [2476];
      \piso.data_r_2475_sv2v_reg  <= \piso.data_li [2475];
      \piso.data_r_2474_sv2v_reg  <= \piso.data_li [2474];
      \piso.data_r_2473_sv2v_reg  <= \piso.data_li [2473];
      \piso.data_r_2472_sv2v_reg  <= \piso.data_li [2472];
      \piso.data_r_2471_sv2v_reg  <= \piso.data_li [2471];
      \piso.data_r_2470_sv2v_reg  <= \piso.data_li [2470];
      \piso.data_r_2469_sv2v_reg  <= \piso.data_li [2469];
      \piso.data_r_2468_sv2v_reg  <= \piso.data_li [2468];
      \piso.data_r_2467_sv2v_reg  <= \piso.data_li [2467];
      \piso.data_r_2466_sv2v_reg  <= \piso.data_li [2466];
      \piso.data_r_2465_sv2v_reg  <= \piso.data_li [2465];
      \piso.data_r_2464_sv2v_reg  <= \piso.data_li [2464];
      \piso.data_r_2463_sv2v_reg  <= \piso.data_li [2463];
      \piso.data_r_2462_sv2v_reg  <= \piso.data_li [2462];
      \piso.data_r_2461_sv2v_reg  <= \piso.data_li [2461];
      \piso.data_r_2460_sv2v_reg  <= \piso.data_li [2460];
      \piso.data_r_2459_sv2v_reg  <= \piso.data_li [2459];
      \piso.data_r_2458_sv2v_reg  <= \piso.data_li [2458];
      \piso.data_r_2457_sv2v_reg  <= \piso.data_li [2457];
      \piso.data_r_2456_sv2v_reg  <= \piso.data_li [2456];
      \piso.data_r_2455_sv2v_reg  <= \piso.data_li [2455];
      \piso.data_r_2454_sv2v_reg  <= \piso.data_li [2454];
      \piso.data_r_2453_sv2v_reg  <= \piso.data_li [2453];
      \piso.data_r_2452_sv2v_reg  <= \piso.data_li [2452];
      \piso.data_r_2451_sv2v_reg  <= \piso.data_li [2451];
      \piso.data_r_2450_sv2v_reg  <= \piso.data_li [2450];
      \piso.data_r_2449_sv2v_reg  <= \piso.data_li [2449];
      \piso.data_r_2448_sv2v_reg  <= \piso.data_li [2448];
      \piso.data_r_2447_sv2v_reg  <= \piso.data_li [2447];
      \piso.data_r_2446_sv2v_reg  <= \piso.data_li [2446];
      \piso.data_r_2445_sv2v_reg  <= \piso.data_li [2445];
      \piso.data_r_2444_sv2v_reg  <= \piso.data_li [2444];
      \piso.data_r_2443_sv2v_reg  <= \piso.data_li [2443];
      \piso.data_r_2442_sv2v_reg  <= \piso.data_li [2442];
      \piso.data_r_2441_sv2v_reg  <= \piso.data_li [2441];
      \piso.data_r_2440_sv2v_reg  <= \piso.data_li [2440];
      \piso.data_r_2439_sv2v_reg  <= \piso.data_li [2439];
      \piso.data_r_2438_sv2v_reg  <= \piso.data_li [2438];
      \piso.data_r_2437_sv2v_reg  <= \piso.data_li [2437];
      \piso.data_r_2436_sv2v_reg  <= \piso.data_li [2436];
      \piso.data_r_2435_sv2v_reg  <= \piso.data_li [2435];
      \piso.data_r_2434_sv2v_reg  <= \piso.data_li [2434];
      \piso.data_r_2433_sv2v_reg  <= \piso.data_li [2433];
      \piso.data_r_2432_sv2v_reg  <= \piso.data_li [2432];
      \piso.data_r_2431_sv2v_reg  <= \piso.data_li [2431];
      \piso.data_r_2430_sv2v_reg  <= \piso.data_li [2430];
      \piso.data_r_2429_sv2v_reg  <= \piso.data_li [2429];
      \piso.data_r_2428_sv2v_reg  <= \piso.data_li [2428];
      \piso.data_r_2427_sv2v_reg  <= \piso.data_li [2427];
      \piso.data_r_2426_sv2v_reg  <= \piso.data_li [2426];
      \piso.data_r_2425_sv2v_reg  <= \piso.data_li [2425];
      \piso.data_r_2424_sv2v_reg  <= \piso.data_li [2424];
      \piso.data_r_2423_sv2v_reg  <= \piso.data_li [2423];
      \piso.data_r_2422_sv2v_reg  <= \piso.data_li [2422];
      \piso.data_r_2421_sv2v_reg  <= \piso.data_li [2421];
      \piso.data_r_2420_sv2v_reg  <= \piso.data_li [2420];
      \piso.data_r_2419_sv2v_reg  <= \piso.data_li [2419];
      \piso.data_r_2418_sv2v_reg  <= \piso.data_li [2418];
      \piso.data_r_2417_sv2v_reg  <= \piso.data_li [2417];
      \piso.data_r_2416_sv2v_reg  <= \piso.data_li [2416];
      \piso.data_r_2415_sv2v_reg  <= \piso.data_li [2415];
      \piso.data_r_2414_sv2v_reg  <= \piso.data_li [2414];
      \piso.data_r_2413_sv2v_reg  <= \piso.data_li [2413];
      \piso.data_r_2412_sv2v_reg  <= \piso.data_li [2412];
      \piso.data_r_2411_sv2v_reg  <= \piso.data_li [2411];
      \piso.data_r_2410_sv2v_reg  <= \piso.data_li [2410];
      \piso.data_r_2409_sv2v_reg  <= \piso.data_li [2409];
      \piso.data_r_2408_sv2v_reg  <= \piso.data_li [2408];
      \piso.data_r_2407_sv2v_reg  <= \piso.data_li [2407];
      \piso.data_r_2406_sv2v_reg  <= \piso.data_li [2406];
      \piso.data_r_2405_sv2v_reg  <= \piso.data_li [2405];
      \piso.data_r_2404_sv2v_reg  <= \piso.data_li [2404];
      \piso.data_r_2403_sv2v_reg  <= \piso.data_li [2403];
      \piso.data_r_2402_sv2v_reg  <= \piso.data_li [2402];
      \piso.data_r_2401_sv2v_reg  <= \piso.data_li [2401];
      \piso.data_r_2400_sv2v_reg  <= \piso.data_li [2400];
      \piso.data_r_2399_sv2v_reg  <= \piso.data_li [2399];
      \piso.data_r_2398_sv2v_reg  <= \piso.data_li [2398];
      \piso.data_r_2397_sv2v_reg  <= \piso.data_li [2397];
      \piso.data_r_2396_sv2v_reg  <= \piso.data_li [2396];
      \piso.data_r_2395_sv2v_reg  <= \piso.data_li [2395];
      \piso.data_r_2394_sv2v_reg  <= \piso.data_li [2394];
      \piso.data_r_2393_sv2v_reg  <= \piso.data_li [2393];
      \piso.data_r_2392_sv2v_reg  <= \piso.data_li [2392];
      \piso.data_r_2391_sv2v_reg  <= \piso.data_li [2391];
      \piso.data_r_2390_sv2v_reg  <= \piso.data_li [2390];
      \piso.data_r_2389_sv2v_reg  <= \piso.data_li [2389];
      \piso.data_r_2388_sv2v_reg  <= \piso.data_li [2388];
      \piso.data_r_2387_sv2v_reg  <= \piso.data_li [2387];
      \piso.data_r_2386_sv2v_reg  <= \piso.data_li [2386];
      \piso.data_r_2385_sv2v_reg  <= \piso.data_li [2385];
      \piso.data_r_2384_sv2v_reg  <= \piso.data_li [2384];
      \piso.data_r_2383_sv2v_reg  <= \piso.data_li [2383];
      \piso.data_r_2382_sv2v_reg  <= \piso.data_li [2382];
      \piso.data_r_2381_sv2v_reg  <= \piso.data_li [2381];
      \piso.data_r_2380_sv2v_reg  <= \piso.data_li [2380];
      \piso.data_r_2379_sv2v_reg  <= \piso.data_li [2379];
      \piso.data_r_2378_sv2v_reg  <= \piso.data_li [2378];
      \piso.data_r_2377_sv2v_reg  <= \piso.data_li [2377];
      \piso.data_r_2376_sv2v_reg  <= \piso.data_li [2376];
      \piso.data_r_2375_sv2v_reg  <= \piso.data_li [2375];
      \piso.data_r_2374_sv2v_reg  <= \piso.data_li [2374];
      \piso.data_r_2373_sv2v_reg  <= \piso.data_li [2373];
      \piso.data_r_2372_sv2v_reg  <= \piso.data_li [2372];
      \piso.data_r_2371_sv2v_reg  <= \piso.data_li [2371];
      \piso.data_r_2370_sv2v_reg  <= \piso.data_li [2370];
      \piso.data_r_2369_sv2v_reg  <= \piso.data_li [2369];
      \piso.data_r_2368_sv2v_reg  <= \piso.data_li [2368];
      \piso.data_r_2367_sv2v_reg  <= \piso.data_li [2367];
      \piso.data_r_2366_sv2v_reg  <= \piso.data_li [2366];
      \piso.data_r_2365_sv2v_reg  <= \piso.data_li [2365];
      \piso.data_r_2364_sv2v_reg  <= \piso.data_li [2364];
      \piso.data_r_2363_sv2v_reg  <= \piso.data_li [2363];
      \piso.data_r_2362_sv2v_reg  <= \piso.data_li [2362];
      \piso.data_r_2361_sv2v_reg  <= \piso.data_li [2361];
      \piso.data_r_2360_sv2v_reg  <= \piso.data_li [2360];
      \piso.data_r_2359_sv2v_reg  <= \piso.data_li [2359];
      \piso.data_r_2358_sv2v_reg  <= \piso.data_li [2358];
      \piso.data_r_2357_sv2v_reg  <= \piso.data_li [2357];
      \piso.data_r_2356_sv2v_reg  <= \piso.data_li [2356];
      \piso.data_r_2355_sv2v_reg  <= \piso.data_li [2355];
      \piso.data_r_2354_sv2v_reg  <= \piso.data_li [2354];
      \piso.data_r_2353_sv2v_reg  <= \piso.data_li [2353];
      \piso.data_r_2352_sv2v_reg  <= \piso.data_li [2352];
      \piso.data_r_2351_sv2v_reg  <= \piso.data_li [2351];
      \piso.data_r_2350_sv2v_reg  <= \piso.data_li [2350];
      \piso.data_r_2349_sv2v_reg  <= \piso.data_li [2349];
      \piso.data_r_2348_sv2v_reg  <= \piso.data_li [2348];
      \piso.data_r_2347_sv2v_reg  <= \piso.data_li [2347];
      \piso.data_r_2346_sv2v_reg  <= \piso.data_li [2346];
      \piso.data_r_2345_sv2v_reg  <= \piso.data_li [2345];
      \piso.data_r_2344_sv2v_reg  <= \piso.data_li [2344];
      \piso.data_r_2343_sv2v_reg  <= \piso.data_li [2343];
      \piso.data_r_2342_sv2v_reg  <= \piso.data_li [2342];
      \piso.data_r_2341_sv2v_reg  <= \piso.data_li [2341];
      \piso.data_r_2340_sv2v_reg  <= \piso.data_li [2340];
      \piso.data_r_2339_sv2v_reg  <= \piso.data_li [2339];
      \piso.data_r_2338_sv2v_reg  <= \piso.data_li [2338];
      \piso.data_r_2337_sv2v_reg  <= \piso.data_li [2337];
      \piso.data_r_2336_sv2v_reg  <= \piso.data_li [2336];
      \piso.data_r_2335_sv2v_reg  <= \piso.data_li [2335];
      \piso.data_r_2334_sv2v_reg  <= \piso.data_li [2334];
      \piso.data_r_2333_sv2v_reg  <= \piso.data_li [2333];
      \piso.data_r_2332_sv2v_reg  <= \piso.data_li [2332];
      \piso.data_r_2331_sv2v_reg  <= \piso.data_li [2331];
      \piso.data_r_2330_sv2v_reg  <= \piso.data_li [2330];
      \piso.data_r_2329_sv2v_reg  <= \piso.data_li [2329];
      \piso.data_r_2328_sv2v_reg  <= \piso.data_li [2328];
      \piso.data_r_2327_sv2v_reg  <= \piso.data_li [2327];
      \piso.data_r_2326_sv2v_reg  <= \piso.data_li [2326];
      \piso.data_r_2325_sv2v_reg  <= \piso.data_li [2325];
      \piso.data_r_2324_sv2v_reg  <= \piso.data_li [2324];
      \piso.data_r_2323_sv2v_reg  <= \piso.data_li [2323];
      \piso.data_r_2322_sv2v_reg  <= \piso.data_li [2322];
      \piso.data_r_2321_sv2v_reg  <= \piso.data_li [2321];
      \piso.data_r_2320_sv2v_reg  <= \piso.data_li [2320];
      \piso.data_r_2319_sv2v_reg  <= \piso.data_li [2319];
      \piso.data_r_2318_sv2v_reg  <= \piso.data_li [2318];
      \piso.data_r_2317_sv2v_reg  <= \piso.data_li [2317];
      \piso.data_r_2316_sv2v_reg  <= \piso.data_li [2316];
      \piso.data_r_2315_sv2v_reg  <= \piso.data_li [2315];
      \piso.data_r_2314_sv2v_reg  <= \piso.data_li [2314];
      \piso.data_r_2313_sv2v_reg  <= \piso.data_li [2313];
      \piso.data_r_2312_sv2v_reg  <= \piso.data_li [2312];
      \piso.data_r_2311_sv2v_reg  <= \piso.data_li [2311];
      \piso.data_r_2310_sv2v_reg  <= \piso.data_li [2310];
      \piso.data_r_2309_sv2v_reg  <= \piso.data_li [2309];
      \piso.data_r_2308_sv2v_reg  <= \piso.data_li [2308];
      \piso.data_r_2307_sv2v_reg  <= \piso.data_li [2307];
      \piso.data_r_2306_sv2v_reg  <= \piso.data_li [2306];
      \piso.data_r_2305_sv2v_reg  <= \piso.data_li [2305];
      \piso.data_r_2304_sv2v_reg  <= \piso.data_li [2304];
      \piso.data_r_2303_sv2v_reg  <= \piso.data_li [2303];
      \piso.data_r_2302_sv2v_reg  <= \piso.data_li [2302];
      \piso.data_r_2301_sv2v_reg  <= \piso.data_li [2301];
      \piso.data_r_2300_sv2v_reg  <= \piso.data_li [2300];
      \piso.data_r_2299_sv2v_reg  <= \piso.data_li [2299];
      \piso.data_r_2298_sv2v_reg  <= \piso.data_li [2298];
      \piso.data_r_2297_sv2v_reg  <= \piso.data_li [2297];
      \piso.data_r_2296_sv2v_reg  <= \piso.data_li [2296];
      \piso.data_r_2295_sv2v_reg  <= \piso.data_li [2295];
      \piso.data_r_2294_sv2v_reg  <= \piso.data_li [2294];
      \piso.data_r_2293_sv2v_reg  <= \piso.data_li [2293];
      \piso.data_r_2292_sv2v_reg  <= \piso.data_li [2292];
      \piso.data_r_2291_sv2v_reg  <= \piso.data_li [2291];
      \piso.data_r_2290_sv2v_reg  <= \piso.data_li [2290];
      \piso.data_r_2289_sv2v_reg  <= \piso.data_li [2289];
      \piso.data_r_2288_sv2v_reg  <= \piso.data_li [2288];
      \piso.data_r_2287_sv2v_reg  <= \piso.data_li [2287];
      \piso.data_r_2286_sv2v_reg  <= \piso.data_li [2286];
      \piso.data_r_2285_sv2v_reg  <= \piso.data_li [2285];
      \piso.data_r_2284_sv2v_reg  <= \piso.data_li [2284];
      \piso.data_r_2283_sv2v_reg  <= \piso.data_li [2283];
      \piso.data_r_2282_sv2v_reg  <= \piso.data_li [2282];
      \piso.data_r_2281_sv2v_reg  <= \piso.data_li [2281];
      \piso.data_r_2280_sv2v_reg  <= \piso.data_li [2280];
      \piso.data_r_2279_sv2v_reg  <= \piso.data_li [2279];
      \piso.data_r_2278_sv2v_reg  <= \piso.data_li [2278];
      \piso.data_r_2277_sv2v_reg  <= \piso.data_li [2277];
      \piso.data_r_2276_sv2v_reg  <= \piso.data_li [2276];
      \piso.data_r_2275_sv2v_reg  <= \piso.data_li [2275];
      \piso.data_r_2274_sv2v_reg  <= \piso.data_li [2274];
      \piso.data_r_2273_sv2v_reg  <= \piso.data_li [2273];
      \piso.data_r_2272_sv2v_reg  <= \piso.data_li [2272];
      \piso.data_r_2271_sv2v_reg  <= \piso.data_li [2271];
      \piso.data_r_2270_sv2v_reg  <= \piso.data_li [2270];
      \piso.data_r_2269_sv2v_reg  <= \piso.data_li [2269];
      \piso.data_r_2268_sv2v_reg  <= \piso.data_li [2268];
      \piso.data_r_2267_sv2v_reg  <= \piso.data_li [2267];
      \piso.data_r_2266_sv2v_reg  <= \piso.data_li [2266];
      \piso.data_r_2265_sv2v_reg  <= \piso.data_li [2265];
      \piso.data_r_2264_sv2v_reg  <= \piso.data_li [2264];
      \piso.data_r_2263_sv2v_reg  <= \piso.data_li [2263];
      \piso.data_r_2262_sv2v_reg  <= \piso.data_li [2262];
      \piso.data_r_2261_sv2v_reg  <= \piso.data_li [2261];
      \piso.data_r_2260_sv2v_reg  <= \piso.data_li [2260];
      \piso.data_r_2259_sv2v_reg  <= \piso.data_li [2259];
      \piso.data_r_2258_sv2v_reg  <= \piso.data_li [2258];
      \piso.data_r_2257_sv2v_reg  <= \piso.data_li [2257];
      \piso.data_r_2256_sv2v_reg  <= \piso.data_li [2256];
      \piso.data_r_2255_sv2v_reg  <= \piso.data_li [2255];
      \piso.data_r_2254_sv2v_reg  <= \piso.data_li [2254];
      \piso.data_r_2253_sv2v_reg  <= \piso.data_li [2253];
      \piso.data_r_2252_sv2v_reg  <= \piso.data_li [2252];
      \piso.data_r_2251_sv2v_reg  <= \piso.data_li [2251];
      \piso.data_r_2250_sv2v_reg  <= \piso.data_li [2250];
      \piso.data_r_2249_sv2v_reg  <= \piso.data_li [2249];
      \piso.data_r_2248_sv2v_reg  <= \piso.data_li [2248];
      \piso.data_r_2247_sv2v_reg  <= \piso.data_li [2247];
      \piso.data_r_2246_sv2v_reg  <= \piso.data_li [2246];
      \piso.data_r_2245_sv2v_reg  <= \piso.data_li [2245];
      \piso.data_r_2244_sv2v_reg  <= \piso.data_li [2244];
      \piso.data_r_2243_sv2v_reg  <= \piso.data_li [2243];
      \piso.data_r_2242_sv2v_reg  <= \piso.data_li [2242];
      \piso.data_r_2241_sv2v_reg  <= \piso.data_li [2241];
      \piso.data_r_2240_sv2v_reg  <= \piso.data_li [2240];
      \piso.data_r_2239_sv2v_reg  <= \piso.data_li [2239];
      \piso.data_r_2238_sv2v_reg  <= \piso.data_li [2238];
      \piso.data_r_2237_sv2v_reg  <= \piso.data_li [2237];
      \piso.data_r_2236_sv2v_reg  <= \piso.data_li [2236];
      \piso.data_r_2235_sv2v_reg  <= \piso.data_li [2235];
      \piso.data_r_2234_sv2v_reg  <= \piso.data_li [2234];
      \piso.data_r_2233_sv2v_reg  <= \piso.data_li [2233];
      \piso.data_r_2232_sv2v_reg  <= \piso.data_li [2232];
      \piso.data_r_2231_sv2v_reg  <= \piso.data_li [2231];
      \piso.data_r_2230_sv2v_reg  <= \piso.data_li [2230];
      \piso.data_r_2229_sv2v_reg  <= \piso.data_li [2229];
      \piso.data_r_2228_sv2v_reg  <= \piso.data_li [2228];
      \piso.data_r_2227_sv2v_reg  <= \piso.data_li [2227];
      \piso.data_r_2226_sv2v_reg  <= \piso.data_li [2226];
      \piso.data_r_2225_sv2v_reg  <= \piso.data_li [2225];
      \piso.data_r_2224_sv2v_reg  <= \piso.data_li [2224];
      \piso.data_r_2223_sv2v_reg  <= \piso.data_li [2223];
      \piso.data_r_2222_sv2v_reg  <= \piso.data_li [2222];
      \piso.data_r_2221_sv2v_reg  <= \piso.data_li [2221];
      \piso.data_r_2220_sv2v_reg  <= \piso.data_li [2220];
      \piso.data_r_2219_sv2v_reg  <= \piso.data_li [2219];
      \piso.data_r_2218_sv2v_reg  <= \piso.data_li [2218];
      \piso.data_r_2217_sv2v_reg  <= \piso.data_li [2217];
      \piso.data_r_2216_sv2v_reg  <= \piso.data_li [2216];
      \piso.data_r_2215_sv2v_reg  <= \piso.data_li [2215];
      \piso.data_r_2214_sv2v_reg  <= \piso.data_li [2214];
      \piso.data_r_2213_sv2v_reg  <= \piso.data_li [2213];
      \piso.data_r_2212_sv2v_reg  <= \piso.data_li [2212];
      \piso.data_r_2211_sv2v_reg  <= \piso.data_li [2211];
      \piso.data_r_2210_sv2v_reg  <= \piso.data_li [2210];
      \piso.data_r_2209_sv2v_reg  <= \piso.data_li [2209];
      \piso.data_r_2208_sv2v_reg  <= \piso.data_li [2208];
      \piso.data_r_2207_sv2v_reg  <= \piso.data_li [2207];
      \piso.data_r_2206_sv2v_reg  <= \piso.data_li [2206];
      \piso.data_r_2205_sv2v_reg  <= \piso.data_li [2205];
      \piso.data_r_2204_sv2v_reg  <= \piso.data_li [2204];
      \piso.data_r_2203_sv2v_reg  <= \piso.data_li [2203];
      \piso.data_r_2202_sv2v_reg  <= \piso.data_li [2202];
      \piso.data_r_2201_sv2v_reg  <= \piso.data_li [2201];
      \piso.data_r_2200_sv2v_reg  <= \piso.data_li [2200];
      \piso.data_r_2199_sv2v_reg  <= \piso.data_li [2199];
      \piso.data_r_2198_sv2v_reg  <= \piso.data_li [2198];
      \piso.data_r_2197_sv2v_reg  <= \piso.data_li [2197];
      \piso.data_r_2196_sv2v_reg  <= \piso.data_li [2196];
      \piso.data_r_2195_sv2v_reg  <= \piso.data_li [2195];
      \piso.data_r_2194_sv2v_reg  <= \piso.data_li [2194];
      \piso.data_r_2193_sv2v_reg  <= \piso.data_li [2193];
      \piso.data_r_2192_sv2v_reg  <= \piso.data_li [2192];
      \piso.data_r_2191_sv2v_reg  <= \piso.data_li [2191];
      \piso.data_r_2190_sv2v_reg  <= \piso.data_li [2190];
      \piso.data_r_2189_sv2v_reg  <= \piso.data_li [2189];
      \piso.data_r_2188_sv2v_reg  <= \piso.data_li [2188];
      \piso.data_r_2187_sv2v_reg  <= \piso.data_li [2187];
      \piso.data_r_2186_sv2v_reg  <= \piso.data_li [2186];
      \piso.data_r_2185_sv2v_reg  <= \piso.data_li [2185];
      \piso.data_r_2184_sv2v_reg  <= \piso.data_li [2184];
      \piso.data_r_2183_sv2v_reg  <= \piso.data_li [2183];
      \piso.data_r_2182_sv2v_reg  <= \piso.data_li [2182];
      \piso.data_r_2181_sv2v_reg  <= \piso.data_li [2181];
      \piso.data_r_2180_sv2v_reg  <= \piso.data_li [2180];
      \piso.data_r_2179_sv2v_reg  <= \piso.data_li [2179];
      \piso.data_r_2178_sv2v_reg  <= \piso.data_li [2178];
      \piso.data_r_2177_sv2v_reg  <= \piso.data_li [2177];
      \piso.data_r_2176_sv2v_reg  <= \piso.data_li [2176];
      \piso.data_r_2175_sv2v_reg  <= \piso.data_li [2175];
      \piso.data_r_2174_sv2v_reg  <= \piso.data_li [2174];
      \piso.data_r_2173_sv2v_reg  <= \piso.data_li [2173];
      \piso.data_r_2172_sv2v_reg  <= \piso.data_li [2172];
      \piso.data_r_2171_sv2v_reg  <= \piso.data_li [2171];
      \piso.data_r_2170_sv2v_reg  <= \piso.data_li [2170];
      \piso.data_r_2169_sv2v_reg  <= \piso.data_li [2169];
      \piso.data_r_2168_sv2v_reg  <= \piso.data_li [2168];
      \piso.data_r_2167_sv2v_reg  <= \piso.data_li [2167];
      \piso.data_r_2166_sv2v_reg  <= \piso.data_li [2166];
      \piso.data_r_2165_sv2v_reg  <= \piso.data_li [2165];
      \piso.data_r_2164_sv2v_reg  <= \piso.data_li [2164];
      \piso.data_r_2163_sv2v_reg  <= \piso.data_li [2163];
      \piso.data_r_2162_sv2v_reg  <= \piso.data_li [2162];
      \piso.data_r_2161_sv2v_reg  <= \piso.data_li [2161];
      \piso.data_r_2160_sv2v_reg  <= \piso.data_li [2160];
      \piso.data_r_2159_sv2v_reg  <= \piso.data_li [2159];
      \piso.data_r_2158_sv2v_reg  <= \piso.data_li [2158];
      \piso.data_r_2157_sv2v_reg  <= \piso.data_li [2157];
      \piso.data_r_2156_sv2v_reg  <= \piso.data_li [2156];
      \piso.data_r_2155_sv2v_reg  <= \piso.data_li [2155];
      \piso.data_r_2154_sv2v_reg  <= \piso.data_li [2154];
      \piso.data_r_2153_sv2v_reg  <= \piso.data_li [2153];
      \piso.data_r_2152_sv2v_reg  <= \piso.data_li [2152];
      \piso.data_r_2151_sv2v_reg  <= \piso.data_li [2151];
      \piso.data_r_2150_sv2v_reg  <= \piso.data_li [2150];
      \piso.data_r_2149_sv2v_reg  <= \piso.data_li [2149];
      \piso.data_r_2148_sv2v_reg  <= \piso.data_li [2148];
      \piso.data_r_2147_sv2v_reg  <= \piso.data_li [2147];
      \piso.data_r_2146_sv2v_reg  <= \piso.data_li [2146];
      \piso.data_r_2145_sv2v_reg  <= \piso.data_li [2145];
      \piso.data_r_2144_sv2v_reg  <= \piso.data_li [2144];
      \piso.data_r_2143_sv2v_reg  <= \piso.data_li [2143];
      \piso.data_r_2142_sv2v_reg  <= \piso.data_li [2142];
      \piso.data_r_2141_sv2v_reg  <= \piso.data_li [2141];
      \piso.data_r_2140_sv2v_reg  <= \piso.data_li [2140];
      \piso.data_r_2139_sv2v_reg  <= \piso.data_li [2139];
      \piso.data_r_2138_sv2v_reg  <= \piso.data_li [2138];
      \piso.data_r_2137_sv2v_reg  <= \piso.data_li [2137];
      \piso.data_r_2136_sv2v_reg  <= \piso.data_li [2136];
      \piso.data_r_2135_sv2v_reg  <= \piso.data_li [2135];
      \piso.data_r_2134_sv2v_reg  <= \piso.data_li [2134];
      \piso.data_r_2133_sv2v_reg  <= \piso.data_li [2133];
      \piso.data_r_2132_sv2v_reg  <= \piso.data_li [2132];
      \piso.data_r_2131_sv2v_reg  <= \piso.data_li [2131];
      \piso.data_r_2130_sv2v_reg  <= \piso.data_li [2130];
      \piso.data_r_2129_sv2v_reg  <= \piso.data_li [2129];
      \piso.data_r_2128_sv2v_reg  <= \piso.data_li [2128];
      \piso.data_r_2127_sv2v_reg  <= \piso.data_li [2127];
      \piso.data_r_2126_sv2v_reg  <= \piso.data_li [2126];
      \piso.data_r_2125_sv2v_reg  <= \piso.data_li [2125];
      \piso.data_r_2124_sv2v_reg  <= \piso.data_li [2124];
      \piso.data_r_2123_sv2v_reg  <= \piso.data_li [2123];
      \piso.data_r_2122_sv2v_reg  <= \piso.data_li [2122];
      \piso.data_r_2121_sv2v_reg  <= \piso.data_li [2121];
      \piso.data_r_2120_sv2v_reg  <= \piso.data_li [2120];
      \piso.data_r_2119_sv2v_reg  <= \piso.data_li [2119];
      \piso.data_r_2118_sv2v_reg  <= \piso.data_li [2118];
      \piso.data_r_2117_sv2v_reg  <= \piso.data_li [2117];
      \piso.data_r_2116_sv2v_reg  <= \piso.data_li [2116];
      \piso.data_r_2115_sv2v_reg  <= \piso.data_li [2115];
      \piso.data_r_2114_sv2v_reg  <= \piso.data_li [2114];
      \piso.data_r_2113_sv2v_reg  <= \piso.data_li [2113];
      \piso.data_r_2112_sv2v_reg  <= \piso.data_li [2112];
      \piso.data_r_2111_sv2v_reg  <= \piso.data_li [2111];
      \piso.data_r_2110_sv2v_reg  <= \piso.data_li [2110];
      \piso.data_r_2109_sv2v_reg  <= \piso.data_li [2109];
      \piso.data_r_2108_sv2v_reg  <= \piso.data_li [2108];
      \piso.data_r_2107_sv2v_reg  <= \piso.data_li [2107];
      \piso.data_r_2106_sv2v_reg  <= \piso.data_li [2106];
      \piso.data_r_2105_sv2v_reg  <= \piso.data_li [2105];
      \piso.data_r_2104_sv2v_reg  <= \piso.data_li [2104];
      \piso.data_r_2103_sv2v_reg  <= \piso.data_li [2103];
      \piso.data_r_2102_sv2v_reg  <= \piso.data_li [2102];
      \piso.data_r_2101_sv2v_reg  <= \piso.data_li [2101];
      \piso.data_r_2100_sv2v_reg  <= \piso.data_li [2100];
      \piso.data_r_2099_sv2v_reg  <= \piso.data_li [2099];
      \piso.data_r_2098_sv2v_reg  <= \piso.data_li [2098];
      \piso.data_r_2097_sv2v_reg  <= \piso.data_li [2097];
      \piso.data_r_2096_sv2v_reg  <= \piso.data_li [2096];
      \piso.data_r_2095_sv2v_reg  <= \piso.data_li [2095];
      \piso.data_r_2094_sv2v_reg  <= \piso.data_li [2094];
      \piso.data_r_2093_sv2v_reg  <= \piso.data_li [2093];
      \piso.data_r_2092_sv2v_reg  <= \piso.data_li [2092];
      \piso.data_r_2091_sv2v_reg  <= \piso.data_li [2091];
      \piso.data_r_2090_sv2v_reg  <= \piso.data_li [2090];
      \piso.data_r_2089_sv2v_reg  <= \piso.data_li [2089];
      \piso.data_r_2088_sv2v_reg  <= \piso.data_li [2088];
      \piso.data_r_2087_sv2v_reg  <= \piso.data_li [2087];
      \piso.data_r_2086_sv2v_reg  <= \piso.data_li [2086];
      \piso.data_r_2085_sv2v_reg  <= \piso.data_li [2085];
      \piso.data_r_2084_sv2v_reg  <= \piso.data_li [2084];
      \piso.data_r_2083_sv2v_reg  <= \piso.data_li [2083];
      \piso.data_r_2082_sv2v_reg  <= \piso.data_li [2082];
      \piso.data_r_2081_sv2v_reg  <= \piso.data_li [2081];
      \piso.data_r_2080_sv2v_reg  <= \piso.data_li [2080];
      \piso.data_r_2079_sv2v_reg  <= \piso.data_li [2079];
      \piso.data_r_2078_sv2v_reg  <= \piso.data_li [2078];
      \piso.data_r_2077_sv2v_reg  <= \piso.data_li [2077];
      \piso.data_r_2076_sv2v_reg  <= \piso.data_li [2076];
      \piso.data_r_2075_sv2v_reg  <= \piso.data_li [2075];
      \piso.data_r_2074_sv2v_reg  <= \piso.data_li [2074];
      \piso.data_r_2073_sv2v_reg  <= \piso.data_li [2073];
      \piso.data_r_2072_sv2v_reg  <= \piso.data_li [2072];
      \piso.data_r_2071_sv2v_reg  <= \piso.data_li [2071];
      \piso.data_r_2070_sv2v_reg  <= \piso.data_li [2070];
      \piso.data_r_2069_sv2v_reg  <= \piso.data_li [2069];
      \piso.data_r_2068_sv2v_reg  <= \piso.data_li [2068];
      \piso.data_r_2067_sv2v_reg  <= \piso.data_li [2067];
      \piso.data_r_2066_sv2v_reg  <= \piso.data_li [2066];
      \piso.data_r_2065_sv2v_reg  <= \piso.data_li [2065];
      \piso.data_r_2064_sv2v_reg  <= \piso.data_li [2064];
      \piso.data_r_2063_sv2v_reg  <= \piso.data_li [2063];
      \piso.data_r_2062_sv2v_reg  <= \piso.data_li [2062];
      \piso.data_r_2061_sv2v_reg  <= \piso.data_li [2061];
      \piso.data_r_2060_sv2v_reg  <= \piso.data_li [2060];
      \piso.data_r_2059_sv2v_reg  <= \piso.data_li [2059];
      \piso.data_r_2058_sv2v_reg  <= \piso.data_li [2058];
      \piso.data_r_2057_sv2v_reg  <= \piso.data_li [2057];
      \piso.data_r_2056_sv2v_reg  <= \piso.data_li [2056];
      \piso.data_r_2055_sv2v_reg  <= \piso.data_li [2055];
      \piso.data_r_2054_sv2v_reg  <= \piso.data_li [2054];
      \piso.data_r_2053_sv2v_reg  <= \piso.data_li [2053];
      \piso.data_r_2052_sv2v_reg  <= \piso.data_li [2052];
      \piso.data_r_2051_sv2v_reg  <= \piso.data_li [2051];
      \piso.data_r_2050_sv2v_reg  <= \piso.data_li [2050];
      \piso.data_r_2049_sv2v_reg  <= \piso.data_li [2049];
      \piso.data_r_2048_sv2v_reg  <= \piso.data_li [2048];
      \piso.data_r_2047_sv2v_reg  <= \piso.data_li [2047];
      \piso.data_r_2046_sv2v_reg  <= \piso.data_li [2046];
      \piso.data_r_2045_sv2v_reg  <= \piso.data_li [2045];
      \piso.data_r_2044_sv2v_reg  <= \piso.data_li [2044];
      \piso.data_r_2043_sv2v_reg  <= \piso.data_li [2043];
      \piso.data_r_2042_sv2v_reg  <= \piso.data_li [2042];
      \piso.data_r_2041_sv2v_reg  <= \piso.data_li [2041];
      \piso.data_r_2040_sv2v_reg  <= \piso.data_li [2040];
      \piso.data_r_2039_sv2v_reg  <= \piso.data_li [2039];
      \piso.data_r_2038_sv2v_reg  <= \piso.data_li [2038];
      \piso.data_r_2037_sv2v_reg  <= \piso.data_li [2037];
      \piso.data_r_2036_sv2v_reg  <= \piso.data_li [2036];
      \piso.data_r_2035_sv2v_reg  <= \piso.data_li [2035];
      \piso.data_r_2034_sv2v_reg  <= \piso.data_li [2034];
      \piso.data_r_2033_sv2v_reg  <= \piso.data_li [2033];
      \piso.data_r_2032_sv2v_reg  <= \piso.data_li [2032];
      \piso.data_r_2031_sv2v_reg  <= \piso.data_li [2031];
      \piso.data_r_2030_sv2v_reg  <= \piso.data_li [2030];
      \piso.data_r_2029_sv2v_reg  <= \piso.data_li [2029];
      \piso.data_r_2028_sv2v_reg  <= \piso.data_li [2028];
      \piso.data_r_2027_sv2v_reg  <= \piso.data_li [2027];
      \piso.data_r_2026_sv2v_reg  <= \piso.data_li [2026];
      \piso.data_r_2025_sv2v_reg  <= \piso.data_li [2025];
      \piso.data_r_2024_sv2v_reg  <= \piso.data_li [2024];
      \piso.data_r_2023_sv2v_reg  <= \piso.data_li [2023];
      \piso.data_r_2022_sv2v_reg  <= \piso.data_li [2022];
      \piso.data_r_2021_sv2v_reg  <= \piso.data_li [2021];
      \piso.data_r_2020_sv2v_reg  <= \piso.data_li [2020];
      \piso.data_r_2019_sv2v_reg  <= \piso.data_li [2019];
      \piso.data_r_2018_sv2v_reg  <= \piso.data_li [2018];
      \piso.data_r_2017_sv2v_reg  <= \piso.data_li [2017];
      \piso.data_r_2016_sv2v_reg  <= \piso.data_li [2016];
      \piso.data_r_2015_sv2v_reg  <= \piso.data_li [2015];
      \piso.data_r_2014_sv2v_reg  <= \piso.data_li [2014];
      \piso.data_r_2013_sv2v_reg  <= \piso.data_li [2013];
      \piso.data_r_2012_sv2v_reg  <= \piso.data_li [2012];
      \piso.data_r_2011_sv2v_reg  <= \piso.data_li [2011];
      \piso.data_r_2010_sv2v_reg  <= \piso.data_li [2010];
      \piso.data_r_2009_sv2v_reg  <= \piso.data_li [2009];
      \piso.data_r_2008_sv2v_reg  <= \piso.data_li [2008];
      \piso.data_r_2007_sv2v_reg  <= \piso.data_li [2007];
      \piso.data_r_2006_sv2v_reg  <= \piso.data_li [2006];
      \piso.data_r_2005_sv2v_reg  <= \piso.data_li [2005];
      \piso.data_r_2004_sv2v_reg  <= \piso.data_li [2004];
      \piso.data_r_2003_sv2v_reg  <= \piso.data_li [2003];
      \piso.data_r_2002_sv2v_reg  <= \piso.data_li [2002];
      \piso.data_r_2001_sv2v_reg  <= \piso.data_li [2001];
      \piso.data_r_2000_sv2v_reg  <= \piso.data_li [2000];
      \piso.data_r_1999_sv2v_reg  <= \piso.data_li [1999];
      \piso.data_r_1998_sv2v_reg  <= \piso.data_li [1998];
      \piso.data_r_1997_sv2v_reg  <= \piso.data_li [1997];
      \piso.data_r_1996_sv2v_reg  <= \piso.data_li [1996];
      \piso.data_r_1995_sv2v_reg  <= \piso.data_li [1995];
      \piso.data_r_1994_sv2v_reg  <= \piso.data_li [1994];
      \piso.data_r_1993_sv2v_reg  <= \piso.data_li [1993];
      \piso.data_r_1992_sv2v_reg  <= \piso.data_li [1992];
      \piso.data_r_1991_sv2v_reg  <= \piso.data_li [1991];
      \piso.data_r_1990_sv2v_reg  <= \piso.data_li [1990];
      \piso.data_r_1989_sv2v_reg  <= \piso.data_li [1989];
      \piso.data_r_1988_sv2v_reg  <= \piso.data_li [1988];
      \piso.data_r_1987_sv2v_reg  <= \piso.data_li [1987];
      \piso.data_r_1986_sv2v_reg  <= \piso.data_li [1986];
      \piso.data_r_1985_sv2v_reg  <= \piso.data_li [1985];
      \piso.data_r_1984_sv2v_reg  <= \piso.data_li [1984];
      \piso.data_r_1983_sv2v_reg  <= \piso.data_li [1983];
      \piso.data_r_1982_sv2v_reg  <= \piso.data_li [1982];
      \piso.data_r_1981_sv2v_reg  <= \piso.data_li [1981];
      \piso.data_r_1980_sv2v_reg  <= \piso.data_li [1980];
      \piso.data_r_1979_sv2v_reg  <= \piso.data_li [1979];
      \piso.data_r_1978_sv2v_reg  <= \piso.data_li [1978];
      \piso.data_r_1977_sv2v_reg  <= \piso.data_li [1977];
      \piso.data_r_1976_sv2v_reg  <= \piso.data_li [1976];
      \piso.data_r_1975_sv2v_reg  <= \piso.data_li [1975];
      \piso.data_r_1974_sv2v_reg  <= \piso.data_li [1974];
      \piso.data_r_1973_sv2v_reg  <= \piso.data_li [1973];
      \piso.data_r_1972_sv2v_reg  <= \piso.data_li [1972];
      \piso.data_r_1971_sv2v_reg  <= \piso.data_li [1971];
      \piso.data_r_1970_sv2v_reg  <= \piso.data_li [1970];
      \piso.data_r_1969_sv2v_reg  <= \piso.data_li [1969];
      \piso.data_r_1968_sv2v_reg  <= \piso.data_li [1968];
      \piso.data_r_1967_sv2v_reg  <= \piso.data_li [1967];
      \piso.data_r_1966_sv2v_reg  <= \piso.data_li [1966];
      \piso.data_r_1965_sv2v_reg  <= \piso.data_li [1965];
      \piso.data_r_1964_sv2v_reg  <= \piso.data_li [1964];
      \piso.data_r_1963_sv2v_reg  <= \piso.data_li [1963];
      \piso.data_r_1962_sv2v_reg  <= \piso.data_li [1962];
      \piso.data_r_1961_sv2v_reg  <= \piso.data_li [1961];
      \piso.data_r_1960_sv2v_reg  <= \piso.data_li [1960];
      \piso.data_r_1959_sv2v_reg  <= \piso.data_li [1959];
      \piso.data_r_1958_sv2v_reg  <= \piso.data_li [1958];
      \piso.data_r_1957_sv2v_reg  <= \piso.data_li [1957];
      \piso.data_r_1956_sv2v_reg  <= \piso.data_li [1956];
      \piso.data_r_1955_sv2v_reg  <= \piso.data_li [1955];
      \piso.data_r_1954_sv2v_reg  <= \piso.data_li [1954];
      \piso.data_r_1953_sv2v_reg  <= \piso.data_li [1953];
      \piso.data_r_1952_sv2v_reg  <= \piso.data_li [1952];
      \piso.data_r_1951_sv2v_reg  <= \piso.data_li [1951];
      \piso.data_r_1950_sv2v_reg  <= \piso.data_li [1950];
      \piso.data_r_1949_sv2v_reg  <= \piso.data_li [1949];
      \piso.data_r_1948_sv2v_reg  <= \piso.data_li [1948];
      \piso.data_r_1947_sv2v_reg  <= \piso.data_li [1947];
      \piso.data_r_1946_sv2v_reg  <= \piso.data_li [1946];
      \piso.data_r_1945_sv2v_reg  <= \piso.data_li [1945];
      \piso.data_r_1944_sv2v_reg  <= \piso.data_li [1944];
      \piso.data_r_1943_sv2v_reg  <= \piso.data_li [1943];
      \piso.data_r_1942_sv2v_reg  <= \piso.data_li [1942];
      \piso.data_r_1941_sv2v_reg  <= \piso.data_li [1941];
      \piso.data_r_1940_sv2v_reg  <= \piso.data_li [1940];
      \piso.data_r_1939_sv2v_reg  <= \piso.data_li [1939];
      \piso.data_r_1938_sv2v_reg  <= \piso.data_li [1938];
      \piso.data_r_1937_sv2v_reg  <= \piso.data_li [1937];
      \piso.data_r_1936_sv2v_reg  <= \piso.data_li [1936];
      \piso.data_r_1935_sv2v_reg  <= \piso.data_li [1935];
      \piso.data_r_1934_sv2v_reg  <= \piso.data_li [1934];
      \piso.data_r_1933_sv2v_reg  <= \piso.data_li [1933];
      \piso.data_r_1932_sv2v_reg  <= \piso.data_li [1932];
      \piso.data_r_1931_sv2v_reg  <= \piso.data_li [1931];
      \piso.data_r_1930_sv2v_reg  <= \piso.data_li [1930];
      \piso.data_r_1929_sv2v_reg  <= \piso.data_li [1929];
      \piso.data_r_1928_sv2v_reg  <= \piso.data_li [1928];
      \piso.data_r_1927_sv2v_reg  <= \piso.data_li [1927];
      \piso.data_r_1926_sv2v_reg  <= \piso.data_li [1926];
      \piso.data_r_1925_sv2v_reg  <= \piso.data_li [1925];
      \piso.data_r_1924_sv2v_reg  <= \piso.data_li [1924];
      \piso.data_r_1923_sv2v_reg  <= \piso.data_li [1923];
      \piso.data_r_1922_sv2v_reg  <= \piso.data_li [1922];
      \piso.data_r_1921_sv2v_reg  <= \piso.data_li [1921];
      \piso.data_r_1920_sv2v_reg  <= \piso.data_li [1920];
      \piso.data_r_1919_sv2v_reg  <= \piso.data_li [1919];
      \piso.data_r_1918_sv2v_reg  <= \piso.data_li [1918];
      \piso.data_r_1917_sv2v_reg  <= \piso.data_li [1917];
      \piso.data_r_1916_sv2v_reg  <= \piso.data_li [1916];
      \piso.data_r_1915_sv2v_reg  <= \piso.data_li [1915];
      \piso.data_r_1914_sv2v_reg  <= \piso.data_li [1914];
      \piso.data_r_1913_sv2v_reg  <= \piso.data_li [1913];
      \piso.data_r_1912_sv2v_reg  <= \piso.data_li [1912];
      \piso.data_r_1911_sv2v_reg  <= \piso.data_li [1911];
      \piso.data_r_1910_sv2v_reg  <= \piso.data_li [1910];
      \piso.data_r_1909_sv2v_reg  <= \piso.data_li [1909];
      \piso.data_r_1908_sv2v_reg  <= \piso.data_li [1908];
      \piso.data_r_1907_sv2v_reg  <= \piso.data_li [1907];
      \piso.data_r_1906_sv2v_reg  <= \piso.data_li [1906];
      \piso.data_r_1905_sv2v_reg  <= \piso.data_li [1905];
      \piso.data_r_1904_sv2v_reg  <= \piso.data_li [1904];
      \piso.data_r_1903_sv2v_reg  <= \piso.data_li [1903];
      \piso.data_r_1902_sv2v_reg  <= \piso.data_li [1902];
      \piso.data_r_1901_sv2v_reg  <= \piso.data_li [1901];
      \piso.data_r_1900_sv2v_reg  <= \piso.data_li [1900];
      \piso.data_r_1899_sv2v_reg  <= \piso.data_li [1899];
      \piso.data_r_1898_sv2v_reg  <= \piso.data_li [1898];
      \piso.data_r_1897_sv2v_reg  <= \piso.data_li [1897];
      \piso.data_r_1896_sv2v_reg  <= \piso.data_li [1896];
      \piso.data_r_1895_sv2v_reg  <= \piso.data_li [1895];
      \piso.data_r_1894_sv2v_reg  <= \piso.data_li [1894];
      \piso.data_r_1893_sv2v_reg  <= \piso.data_li [1893];
      \piso.data_r_1892_sv2v_reg  <= \piso.data_li [1892];
      \piso.data_r_1891_sv2v_reg  <= \piso.data_li [1891];
      \piso.data_r_1890_sv2v_reg  <= \piso.data_li [1890];
      \piso.data_r_1889_sv2v_reg  <= \piso.data_li [1889];
      \piso.data_r_1888_sv2v_reg  <= \piso.data_li [1888];
      \piso.data_r_1887_sv2v_reg  <= \piso.data_li [1887];
      \piso.data_r_1886_sv2v_reg  <= \piso.data_li [1886];
      \piso.data_r_1885_sv2v_reg  <= \piso.data_li [1885];
      \piso.data_r_1884_sv2v_reg  <= \piso.data_li [1884];
      \piso.data_r_1883_sv2v_reg  <= \piso.data_li [1883];
      \piso.data_r_1882_sv2v_reg  <= \piso.data_li [1882];
      \piso.data_r_1881_sv2v_reg  <= \piso.data_li [1881];
      \piso.data_r_1880_sv2v_reg  <= \piso.data_li [1880];
      \piso.data_r_1879_sv2v_reg  <= \piso.data_li [1879];
      \piso.data_r_1878_sv2v_reg  <= \piso.data_li [1878];
      \piso.data_r_1877_sv2v_reg  <= \piso.data_li [1877];
      \piso.data_r_1876_sv2v_reg  <= \piso.data_li [1876];
      \piso.data_r_1875_sv2v_reg  <= \piso.data_li [1875];
      \piso.data_r_1874_sv2v_reg  <= \piso.data_li [1874];
      \piso.data_r_1873_sv2v_reg  <= \piso.data_li [1873];
      \piso.data_r_1872_sv2v_reg  <= \piso.data_li [1872];
      \piso.data_r_1871_sv2v_reg  <= \piso.data_li [1871];
      \piso.data_r_1870_sv2v_reg  <= \piso.data_li [1870];
      \piso.data_r_1869_sv2v_reg  <= \piso.data_li [1869];
      \piso.data_r_1868_sv2v_reg  <= \piso.data_li [1868];
      \piso.data_r_1867_sv2v_reg  <= \piso.data_li [1867];
      \piso.data_r_1866_sv2v_reg  <= \piso.data_li [1866];
      \piso.data_r_1865_sv2v_reg  <= \piso.data_li [1865];
      \piso.data_r_1864_sv2v_reg  <= \piso.data_li [1864];
      \piso.data_r_1863_sv2v_reg  <= \piso.data_li [1863];
      \piso.data_r_1862_sv2v_reg  <= \piso.data_li [1862];
      \piso.data_r_1861_sv2v_reg  <= \piso.data_li [1861];
      \piso.data_r_1860_sv2v_reg  <= \piso.data_li [1860];
      \piso.data_r_1859_sv2v_reg  <= \piso.data_li [1859];
      \piso.data_r_1858_sv2v_reg  <= \piso.data_li [1858];
      \piso.data_r_1857_sv2v_reg  <= \piso.data_li [1857];
      \piso.data_r_1856_sv2v_reg  <= \piso.data_li [1856];
      \piso.data_r_1855_sv2v_reg  <= \piso.data_li [1855];
      \piso.data_r_1854_sv2v_reg  <= \piso.data_li [1854];
      \piso.data_r_1853_sv2v_reg  <= \piso.data_li [1853];
      \piso.data_r_1852_sv2v_reg  <= \piso.data_li [1852];
      \piso.data_r_1851_sv2v_reg  <= \piso.data_li [1851];
      \piso.data_r_1850_sv2v_reg  <= \piso.data_li [1850];
      \piso.data_r_1849_sv2v_reg  <= \piso.data_li [1849];
      \piso.data_r_1848_sv2v_reg  <= \piso.data_li [1848];
      \piso.data_r_1847_sv2v_reg  <= \piso.data_li [1847];
      \piso.data_r_1846_sv2v_reg  <= \piso.data_li [1846];
      \piso.data_r_1845_sv2v_reg  <= \piso.data_li [1845];
      \piso.data_r_1844_sv2v_reg  <= \piso.data_li [1844];
      \piso.data_r_1843_sv2v_reg  <= \piso.data_li [1843];
      \piso.data_r_1842_sv2v_reg  <= \piso.data_li [1842];
      \piso.data_r_1841_sv2v_reg  <= \piso.data_li [1841];
      \piso.data_r_1840_sv2v_reg  <= \piso.data_li [1840];
      \piso.data_r_1839_sv2v_reg  <= \piso.data_li [1839];
      \piso.data_r_1838_sv2v_reg  <= \piso.data_li [1838];
      \piso.data_r_1837_sv2v_reg  <= \piso.data_li [1837];
      \piso.data_r_1836_sv2v_reg  <= \piso.data_li [1836];
      \piso.data_r_1835_sv2v_reg  <= \piso.data_li [1835];
      \piso.data_r_1834_sv2v_reg  <= \piso.data_li [1834];
      \piso.data_r_1833_sv2v_reg  <= \piso.data_li [1833];
      \piso.data_r_1832_sv2v_reg  <= \piso.data_li [1832];
      \piso.data_r_1831_sv2v_reg  <= \piso.data_li [1831];
      \piso.data_r_1830_sv2v_reg  <= \piso.data_li [1830];
      \piso.data_r_1829_sv2v_reg  <= \piso.data_li [1829];
      \piso.data_r_1828_sv2v_reg  <= \piso.data_li [1828];
      \piso.data_r_1827_sv2v_reg  <= \piso.data_li [1827];
      \piso.data_r_1826_sv2v_reg  <= \piso.data_li [1826];
      \piso.data_r_1825_sv2v_reg  <= \piso.data_li [1825];
      \piso.data_r_1824_sv2v_reg  <= \piso.data_li [1824];
      \piso.data_r_1823_sv2v_reg  <= \piso.data_li [1823];
      \piso.data_r_1822_sv2v_reg  <= \piso.data_li [1822];
      \piso.data_r_1821_sv2v_reg  <= \piso.data_li [1821];
      \piso.data_r_1820_sv2v_reg  <= \piso.data_li [1820];
      \piso.data_r_1819_sv2v_reg  <= \piso.data_li [1819];
      \piso.data_r_1818_sv2v_reg  <= \piso.data_li [1818];
      \piso.data_r_1817_sv2v_reg  <= \piso.data_li [1817];
      \piso.data_r_1816_sv2v_reg  <= \piso.data_li [1816];
      \piso.data_r_1815_sv2v_reg  <= \piso.data_li [1815];
      \piso.data_r_1814_sv2v_reg  <= \piso.data_li [1814];
      \piso.data_r_1813_sv2v_reg  <= \piso.data_li [1813];
      \piso.data_r_1812_sv2v_reg  <= \piso.data_li [1812];
      \piso.data_r_1811_sv2v_reg  <= \piso.data_li [1811];
      \piso.data_r_1810_sv2v_reg  <= \piso.data_li [1810];
      \piso.data_r_1809_sv2v_reg  <= \piso.data_li [1809];
      \piso.data_r_1808_sv2v_reg  <= \piso.data_li [1808];
      \piso.data_r_1807_sv2v_reg  <= \piso.data_li [1807];
      \piso.data_r_1806_sv2v_reg  <= \piso.data_li [1806];
      \piso.data_r_1805_sv2v_reg  <= \piso.data_li [1805];
      \piso.data_r_1804_sv2v_reg  <= \piso.data_li [1804];
      \piso.data_r_1803_sv2v_reg  <= \piso.data_li [1803];
      \piso.data_r_1802_sv2v_reg  <= \piso.data_li [1802];
      \piso.data_r_1801_sv2v_reg  <= \piso.data_li [1801];
      \piso.data_r_1800_sv2v_reg  <= \piso.data_li [1800];
      \piso.data_r_1799_sv2v_reg  <= \piso.data_li [1799];
      \piso.data_r_1798_sv2v_reg  <= \piso.data_li [1798];
      \piso.data_r_1797_sv2v_reg  <= \piso.data_li [1797];
      \piso.data_r_1796_sv2v_reg  <= \piso.data_li [1796];
      \piso.data_r_1795_sv2v_reg  <= \piso.data_li [1795];
      \piso.data_r_1794_sv2v_reg  <= \piso.data_li [1794];
      \piso.data_r_1793_sv2v_reg  <= \piso.data_li [1793];
      \piso.data_r_1792_sv2v_reg  <= \piso.data_li [1792];
      \piso.data_r_1791_sv2v_reg  <= \piso.data_li [1791];
      \piso.data_r_1790_sv2v_reg  <= \piso.data_li [1790];
      \piso.data_r_1789_sv2v_reg  <= \piso.data_li [1789];
      \piso.data_r_1788_sv2v_reg  <= \piso.data_li [1788];
      \piso.data_r_1787_sv2v_reg  <= \piso.data_li [1787];
      \piso.data_r_1786_sv2v_reg  <= \piso.data_li [1786];
      \piso.data_r_1785_sv2v_reg  <= \piso.data_li [1785];
      \piso.data_r_1784_sv2v_reg  <= \piso.data_li [1784];
      \piso.data_r_1783_sv2v_reg  <= \piso.data_li [1783];
      \piso.data_r_1782_sv2v_reg  <= \piso.data_li [1782];
      \piso.data_r_1781_sv2v_reg  <= \piso.data_li [1781];
      \piso.data_r_1780_sv2v_reg  <= \piso.data_li [1780];
      \piso.data_r_1779_sv2v_reg  <= \piso.data_li [1779];
      \piso.data_r_1778_sv2v_reg  <= \piso.data_li [1778];
      \piso.data_r_1777_sv2v_reg  <= \piso.data_li [1777];
      \piso.data_r_1776_sv2v_reg  <= \piso.data_li [1776];
      \piso.data_r_1775_sv2v_reg  <= \piso.data_li [1775];
      \piso.data_r_1774_sv2v_reg  <= \piso.data_li [1774];
      \piso.data_r_1773_sv2v_reg  <= \piso.data_li [1773];
      \piso.data_r_1772_sv2v_reg  <= \piso.data_li [1772];
      \piso.data_r_1771_sv2v_reg  <= \piso.data_li [1771];
      \piso.data_r_1770_sv2v_reg  <= \piso.data_li [1770];
      \piso.data_r_1769_sv2v_reg  <= \piso.data_li [1769];
      \piso.data_r_1768_sv2v_reg  <= \piso.data_li [1768];
      \piso.data_r_1767_sv2v_reg  <= \piso.data_li [1767];
      \piso.data_r_1766_sv2v_reg  <= \piso.data_li [1766];
      \piso.data_r_1765_sv2v_reg  <= \piso.data_li [1765];
      \piso.data_r_1764_sv2v_reg  <= \piso.data_li [1764];
      \piso.data_r_1763_sv2v_reg  <= \piso.data_li [1763];
      \piso.data_r_1762_sv2v_reg  <= \piso.data_li [1762];
      \piso.data_r_1761_sv2v_reg  <= \piso.data_li [1761];
      \piso.data_r_1760_sv2v_reg  <= \piso.data_li [1760];
      \piso.data_r_1759_sv2v_reg  <= \piso.data_li [1759];
      \piso.data_r_1758_sv2v_reg  <= \piso.data_li [1758];
      \piso.data_r_1757_sv2v_reg  <= \piso.data_li [1757];
      \piso.data_r_1756_sv2v_reg  <= \piso.data_li [1756];
      \piso.data_r_1755_sv2v_reg  <= \piso.data_li [1755];
      \piso.data_r_1754_sv2v_reg  <= \piso.data_li [1754];
      \piso.data_r_1753_sv2v_reg  <= \piso.data_li [1753];
      \piso.data_r_1752_sv2v_reg  <= \piso.data_li [1752];
      \piso.data_r_1751_sv2v_reg  <= \piso.data_li [1751];
      \piso.data_r_1750_sv2v_reg  <= \piso.data_li [1750];
      \piso.data_r_1749_sv2v_reg  <= \piso.data_li [1749];
      \piso.data_r_1748_sv2v_reg  <= \piso.data_li [1748];
      \piso.data_r_1747_sv2v_reg  <= \piso.data_li [1747];
      \piso.data_r_1746_sv2v_reg  <= \piso.data_li [1746];
      \piso.data_r_1745_sv2v_reg  <= \piso.data_li [1745];
      \piso.data_r_1744_sv2v_reg  <= \piso.data_li [1744];
      \piso.data_r_1743_sv2v_reg  <= \piso.data_li [1743];
      \piso.data_r_1742_sv2v_reg  <= \piso.data_li [1742];
      \piso.data_r_1741_sv2v_reg  <= \piso.data_li [1741];
      \piso.data_r_1740_sv2v_reg  <= \piso.data_li [1740];
      \piso.data_r_1739_sv2v_reg  <= \piso.data_li [1739];
      \piso.data_r_1738_sv2v_reg  <= \piso.data_li [1738];
      \piso.data_r_1737_sv2v_reg  <= \piso.data_li [1737];
      \piso.data_r_1736_sv2v_reg  <= \piso.data_li [1736];
      \piso.data_r_1735_sv2v_reg  <= \piso.data_li [1735];
      \piso.data_r_1734_sv2v_reg  <= \piso.data_li [1734];
      \piso.data_r_1733_sv2v_reg  <= \piso.data_li [1733];
      \piso.data_r_1732_sv2v_reg  <= \piso.data_li [1732];
      \piso.data_r_1731_sv2v_reg  <= \piso.data_li [1731];
      \piso.data_r_1730_sv2v_reg  <= \piso.data_li [1730];
      \piso.data_r_1729_sv2v_reg  <= \piso.data_li [1729];
      \piso.data_r_1728_sv2v_reg  <= \piso.data_li [1728];
      \piso.data_r_1727_sv2v_reg  <= \piso.data_li [1727];
      \piso.data_r_1726_sv2v_reg  <= \piso.data_li [1726];
      \piso.data_r_1725_sv2v_reg  <= \piso.data_li [1725];
      \piso.data_r_1724_sv2v_reg  <= \piso.data_li [1724];
      \piso.data_r_1723_sv2v_reg  <= \piso.data_li [1723];
      \piso.data_r_1722_sv2v_reg  <= \piso.data_li [1722];
      \piso.data_r_1721_sv2v_reg  <= \piso.data_li [1721];
      \piso.data_r_1720_sv2v_reg  <= \piso.data_li [1720];
      \piso.data_r_1719_sv2v_reg  <= \piso.data_li [1719];
      \piso.data_r_1718_sv2v_reg  <= \piso.data_li [1718];
      \piso.data_r_1717_sv2v_reg  <= \piso.data_li [1717];
      \piso.data_r_1716_sv2v_reg  <= \piso.data_li [1716];
      \piso.data_r_1715_sv2v_reg  <= \piso.data_li [1715];
      \piso.data_r_1714_sv2v_reg  <= \piso.data_li [1714];
      \piso.data_r_1713_sv2v_reg  <= \piso.data_li [1713];
      \piso.data_r_1712_sv2v_reg  <= \piso.data_li [1712];
      \piso.data_r_1711_sv2v_reg  <= \piso.data_li [1711];
      \piso.data_r_1710_sv2v_reg  <= \piso.data_li [1710];
      \piso.data_r_1709_sv2v_reg  <= \piso.data_li [1709];
      \piso.data_r_1708_sv2v_reg  <= \piso.data_li [1708];
      \piso.data_r_1707_sv2v_reg  <= \piso.data_li [1707];
      \piso.data_r_1706_sv2v_reg  <= \piso.data_li [1706];
      \piso.data_r_1705_sv2v_reg  <= \piso.data_li [1705];
      \piso.data_r_1704_sv2v_reg  <= \piso.data_li [1704];
      \piso.data_r_1703_sv2v_reg  <= \piso.data_li [1703];
      \piso.data_r_1702_sv2v_reg  <= \piso.data_li [1702];
      \piso.data_r_1701_sv2v_reg  <= \piso.data_li [1701];
      \piso.data_r_1700_sv2v_reg  <= \piso.data_li [1700];
      \piso.data_r_1699_sv2v_reg  <= \piso.data_li [1699];
      \piso.data_r_1698_sv2v_reg  <= \piso.data_li [1698];
      \piso.data_r_1697_sv2v_reg  <= \piso.data_li [1697];
      \piso.data_r_1696_sv2v_reg  <= \piso.data_li [1696];
      \piso.data_r_1695_sv2v_reg  <= \piso.data_li [1695];
      \piso.data_r_1694_sv2v_reg  <= \piso.data_li [1694];
      \piso.data_r_1693_sv2v_reg  <= \piso.data_li [1693];
      \piso.data_r_1692_sv2v_reg  <= \piso.data_li [1692];
      \piso.data_r_1691_sv2v_reg  <= \piso.data_li [1691];
      \piso.data_r_1690_sv2v_reg  <= \piso.data_li [1690];
      \piso.data_r_1689_sv2v_reg  <= \piso.data_li [1689];
      \piso.data_r_1688_sv2v_reg  <= \piso.data_li [1688];
      \piso.data_r_1687_sv2v_reg  <= \piso.data_li [1687];
      \piso.data_r_1686_sv2v_reg  <= \piso.data_li [1686];
      \piso.data_r_1685_sv2v_reg  <= \piso.data_li [1685];
      \piso.data_r_1684_sv2v_reg  <= \piso.data_li [1684];
      \piso.data_r_1683_sv2v_reg  <= \piso.data_li [1683];
      \piso.data_r_1682_sv2v_reg  <= \piso.data_li [1682];
      \piso.data_r_1681_sv2v_reg  <= \piso.data_li [1681];
      \piso.data_r_1680_sv2v_reg  <= \piso.data_li [1680];
      \piso.data_r_1679_sv2v_reg  <= \piso.data_li [1679];
      \piso.data_r_1678_sv2v_reg  <= \piso.data_li [1678];
      \piso.data_r_1677_sv2v_reg  <= \piso.data_li [1677];
      \piso.data_r_1676_sv2v_reg  <= \piso.data_li [1676];
      \piso.data_r_1675_sv2v_reg  <= \piso.data_li [1675];
      \piso.data_r_1674_sv2v_reg  <= \piso.data_li [1674];
      \piso.data_r_1673_sv2v_reg  <= \piso.data_li [1673];
      \piso.data_r_1672_sv2v_reg  <= \piso.data_li [1672];
      \piso.data_r_1671_sv2v_reg  <= \piso.data_li [1671];
      \piso.data_r_1670_sv2v_reg  <= \piso.data_li [1670];
      \piso.data_r_1669_sv2v_reg  <= \piso.data_li [1669];
      \piso.data_r_1668_sv2v_reg  <= \piso.data_li [1668];
      \piso.data_r_1667_sv2v_reg  <= \piso.data_li [1667];
      \piso.data_r_1666_sv2v_reg  <= \piso.data_li [1666];
      \piso.data_r_1665_sv2v_reg  <= \piso.data_li [1665];
      \piso.data_r_1664_sv2v_reg  <= \piso.data_li [1664];
      \piso.data_r_1663_sv2v_reg  <= \piso.data_li [1663];
      \piso.data_r_1662_sv2v_reg  <= \piso.data_li [1662];
      \piso.data_r_1661_sv2v_reg  <= \piso.data_li [1661];
      \piso.data_r_1660_sv2v_reg  <= \piso.data_li [1660];
      \piso.data_r_1659_sv2v_reg  <= \piso.data_li [1659];
      \piso.data_r_1658_sv2v_reg  <= \piso.data_li [1658];
      \piso.data_r_1657_sv2v_reg  <= \piso.data_li [1657];
      \piso.data_r_1656_sv2v_reg  <= \piso.data_li [1656];
      \piso.data_r_1655_sv2v_reg  <= \piso.data_li [1655];
      \piso.data_r_1654_sv2v_reg  <= \piso.data_li [1654];
      \piso.data_r_1653_sv2v_reg  <= \piso.data_li [1653];
      \piso.data_r_1652_sv2v_reg  <= \piso.data_li [1652];
      \piso.data_r_1651_sv2v_reg  <= \piso.data_li [1651];
      \piso.data_r_1650_sv2v_reg  <= \piso.data_li [1650];
      \piso.data_r_1649_sv2v_reg  <= \piso.data_li [1649];
      \piso.data_r_1648_sv2v_reg  <= \piso.data_li [1648];
      \piso.data_r_1647_sv2v_reg  <= \piso.data_li [1647];
      \piso.data_r_1646_sv2v_reg  <= \piso.data_li [1646];
      \piso.data_r_1645_sv2v_reg  <= \piso.data_li [1645];
      \piso.data_r_1644_sv2v_reg  <= \piso.data_li [1644];
      \piso.data_r_1643_sv2v_reg  <= \piso.data_li [1643];
      \piso.data_r_1642_sv2v_reg  <= \piso.data_li [1642];
      \piso.data_r_1641_sv2v_reg  <= \piso.data_li [1641];
      \piso.data_r_1640_sv2v_reg  <= \piso.data_li [1640];
      \piso.data_r_1639_sv2v_reg  <= \piso.data_li [1639];
      \piso.data_r_1638_sv2v_reg  <= \piso.data_li [1638];
      \piso.data_r_1637_sv2v_reg  <= \piso.data_li [1637];
      \piso.data_r_1636_sv2v_reg  <= \piso.data_li [1636];
      \piso.data_r_1635_sv2v_reg  <= \piso.data_li [1635];
      \piso.data_r_1634_sv2v_reg  <= \piso.data_li [1634];
      \piso.data_r_1633_sv2v_reg  <= \piso.data_li [1633];
      \piso.data_r_1632_sv2v_reg  <= \piso.data_li [1632];
      \piso.data_r_1631_sv2v_reg  <= \piso.data_li [1631];
      \piso.data_r_1630_sv2v_reg  <= \piso.data_li [1630];
      \piso.data_r_1629_sv2v_reg  <= \piso.data_li [1629];
      \piso.data_r_1628_sv2v_reg  <= \piso.data_li [1628];
      \piso.data_r_1627_sv2v_reg  <= \piso.data_li [1627];
      \piso.data_r_1626_sv2v_reg  <= \piso.data_li [1626];
      \piso.data_r_1625_sv2v_reg  <= \piso.data_li [1625];
      \piso.data_r_1624_sv2v_reg  <= \piso.data_li [1624];
      \piso.data_r_1623_sv2v_reg  <= \piso.data_li [1623];
      \piso.data_r_1622_sv2v_reg  <= \piso.data_li [1622];
      \piso.data_r_1621_sv2v_reg  <= \piso.data_li [1621];
      \piso.data_r_1620_sv2v_reg  <= \piso.data_li [1620];
      \piso.data_r_1619_sv2v_reg  <= \piso.data_li [1619];
      \piso.data_r_1618_sv2v_reg  <= \piso.data_li [1618];
      \piso.data_r_1617_sv2v_reg  <= \piso.data_li [1617];
      \piso.data_r_1616_sv2v_reg  <= \piso.data_li [1616];
      \piso.data_r_1615_sv2v_reg  <= \piso.data_li [1615];
      \piso.data_r_1614_sv2v_reg  <= \piso.data_li [1614];
      \piso.data_r_1613_sv2v_reg  <= \piso.data_li [1613];
      \piso.data_r_1612_sv2v_reg  <= \piso.data_li [1612];
      \piso.data_r_1611_sv2v_reg  <= \piso.data_li [1611];
      \piso.data_r_1610_sv2v_reg  <= \piso.data_li [1610];
      \piso.data_r_1609_sv2v_reg  <= \piso.data_li [1609];
      \piso.data_r_1608_sv2v_reg  <= \piso.data_li [1608];
      \piso.data_r_1607_sv2v_reg  <= \piso.data_li [1607];
      \piso.data_r_1606_sv2v_reg  <= \piso.data_li [1606];
      \piso.data_r_1605_sv2v_reg  <= \piso.data_li [1605];
      \piso.data_r_1604_sv2v_reg  <= \piso.data_li [1604];
      \piso.data_r_1603_sv2v_reg  <= \piso.data_li [1603];
      \piso.data_r_1602_sv2v_reg  <= \piso.data_li [1602];
      \piso.data_r_1601_sv2v_reg  <= \piso.data_li [1601];
      \piso.data_r_1600_sv2v_reg  <= \piso.data_li [1600];
      \piso.data_r_1599_sv2v_reg  <= \piso.data_li [1599];
      \piso.data_r_1598_sv2v_reg  <= \piso.data_li [1598];
      \piso.data_r_1597_sv2v_reg  <= \piso.data_li [1597];
      \piso.data_r_1596_sv2v_reg  <= \piso.data_li [1596];
      \piso.data_r_1595_sv2v_reg  <= \piso.data_li [1595];
      \piso.data_r_1594_sv2v_reg  <= \piso.data_li [1594];
      \piso.data_r_1593_sv2v_reg  <= \piso.data_li [1593];
      \piso.data_r_1592_sv2v_reg  <= \piso.data_li [1592];
      \piso.data_r_1591_sv2v_reg  <= \piso.data_li [1591];
      \piso.data_r_1590_sv2v_reg  <= \piso.data_li [1590];
      \piso.data_r_1589_sv2v_reg  <= \piso.data_li [1589];
      \piso.data_r_1588_sv2v_reg  <= \piso.data_li [1588];
      \piso.data_r_1587_sv2v_reg  <= \piso.data_li [1587];
      \piso.data_r_1586_sv2v_reg  <= \piso.data_li [1586];
      \piso.data_r_1585_sv2v_reg  <= \piso.data_li [1585];
      \piso.data_r_1584_sv2v_reg  <= \piso.data_li [1584];
      \piso.data_r_1583_sv2v_reg  <= \piso.data_li [1583];
      \piso.data_r_1582_sv2v_reg  <= \piso.data_li [1582];
      \piso.data_r_1581_sv2v_reg  <= \piso.data_li [1581];
      \piso.data_r_1580_sv2v_reg  <= \piso.data_li [1580];
      \piso.data_r_1579_sv2v_reg  <= \piso.data_li [1579];
      \piso.data_r_1578_sv2v_reg  <= \piso.data_li [1578];
      \piso.data_r_1577_sv2v_reg  <= \piso.data_li [1577];
      \piso.data_r_1576_sv2v_reg  <= \piso.data_li [1576];
      \piso.data_r_1575_sv2v_reg  <= \piso.data_li [1575];
      \piso.data_r_1574_sv2v_reg  <= \piso.data_li [1574];
      \piso.data_r_1573_sv2v_reg  <= \piso.data_li [1573];
      \piso.data_r_1572_sv2v_reg  <= \piso.data_li [1572];
      \piso.data_r_1571_sv2v_reg  <= \piso.data_li [1571];
      \piso.data_r_1570_sv2v_reg  <= \piso.data_li [1570];
      \piso.data_r_1569_sv2v_reg  <= \piso.data_li [1569];
      \piso.data_r_1568_sv2v_reg  <= \piso.data_li [1568];
      \piso.data_r_1567_sv2v_reg  <= \piso.data_li [1567];
      \piso.data_r_1566_sv2v_reg  <= \piso.data_li [1566];
      \piso.data_r_1565_sv2v_reg  <= \piso.data_li [1565];
      \piso.data_r_1564_sv2v_reg  <= \piso.data_li [1564];
      \piso.data_r_1563_sv2v_reg  <= \piso.data_li [1563];
      \piso.data_r_1562_sv2v_reg  <= \piso.data_li [1562];
      \piso.data_r_1561_sv2v_reg  <= \piso.data_li [1561];
      \piso.data_r_1560_sv2v_reg  <= \piso.data_li [1560];
      \piso.data_r_1559_sv2v_reg  <= \piso.data_li [1559];
      \piso.data_r_1558_sv2v_reg  <= \piso.data_li [1558];
      \piso.data_r_1557_sv2v_reg  <= \piso.data_li [1557];
      \piso.data_r_1556_sv2v_reg  <= \piso.data_li [1556];
      \piso.data_r_1555_sv2v_reg  <= \piso.data_li [1555];
      \piso.data_r_1554_sv2v_reg  <= \piso.data_li [1554];
      \piso.data_r_1553_sv2v_reg  <= \piso.data_li [1553];
      \piso.data_r_1552_sv2v_reg  <= \piso.data_li [1552];
      \piso.data_r_1551_sv2v_reg  <= \piso.data_li [1551];
      \piso.data_r_1550_sv2v_reg  <= \piso.data_li [1550];
      \piso.data_r_1549_sv2v_reg  <= \piso.data_li [1549];
      \piso.data_r_1548_sv2v_reg  <= \piso.data_li [1548];
      \piso.data_r_1547_sv2v_reg  <= \piso.data_li [1547];
      \piso.data_r_1546_sv2v_reg  <= \piso.data_li [1546];
      \piso.data_r_1545_sv2v_reg  <= \piso.data_li [1545];
      \piso.data_r_1544_sv2v_reg  <= \piso.data_li [1544];
      \piso.data_r_1543_sv2v_reg  <= \piso.data_li [1543];
      \piso.data_r_1542_sv2v_reg  <= \piso.data_li [1542];
      \piso.data_r_1541_sv2v_reg  <= \piso.data_li [1541];
      \piso.data_r_1540_sv2v_reg  <= \piso.data_li [1540];
      \piso.data_r_1539_sv2v_reg  <= \piso.data_li [1539];
      \piso.data_r_1538_sv2v_reg  <= \piso.data_li [1538];
      \piso.data_r_1537_sv2v_reg  <= \piso.data_li [1537];
      \piso.data_r_1536_sv2v_reg  <= \piso.data_li [1536];
      \piso.data_r_1535_sv2v_reg  <= \piso.data_li [1535];
      \piso.data_r_1534_sv2v_reg  <= \piso.data_li [1534];
      \piso.data_r_1533_sv2v_reg  <= \piso.data_li [1533];
      \piso.data_r_1532_sv2v_reg  <= \piso.data_li [1532];
      \piso.data_r_1531_sv2v_reg  <= \piso.data_li [1531];
      \piso.data_r_1530_sv2v_reg  <= \piso.data_li [1530];
      \piso.data_r_1529_sv2v_reg  <= \piso.data_li [1529];
      \piso.data_r_1528_sv2v_reg  <= \piso.data_li [1528];
      \piso.data_r_1527_sv2v_reg  <= \piso.data_li [1527];
      \piso.data_r_1526_sv2v_reg  <= \piso.data_li [1526];
      \piso.data_r_1525_sv2v_reg  <= \piso.data_li [1525];
      \piso.data_r_1524_sv2v_reg  <= \piso.data_li [1524];
      \piso.data_r_1523_sv2v_reg  <= \piso.data_li [1523];
      \piso.data_r_1522_sv2v_reg  <= \piso.data_li [1522];
      \piso.data_r_1521_sv2v_reg  <= \piso.data_li [1521];
      \piso.data_r_1520_sv2v_reg  <= \piso.data_li [1520];
      \piso.data_r_1519_sv2v_reg  <= \piso.data_li [1519];
      \piso.data_r_1518_sv2v_reg  <= \piso.data_li [1518];
      \piso.data_r_1517_sv2v_reg  <= \piso.data_li [1517];
      \piso.data_r_1516_sv2v_reg  <= \piso.data_li [1516];
      \piso.data_r_1515_sv2v_reg  <= \piso.data_li [1515];
      \piso.data_r_1514_sv2v_reg  <= \piso.data_li [1514];
      \piso.data_r_1513_sv2v_reg  <= \piso.data_li [1513];
      \piso.data_r_1512_sv2v_reg  <= \piso.data_li [1512];
      \piso.data_r_1511_sv2v_reg  <= \piso.data_li [1511];
      \piso.data_r_1510_sv2v_reg  <= \piso.data_li [1510];
      \piso.data_r_1509_sv2v_reg  <= \piso.data_li [1509];
      \piso.data_r_1508_sv2v_reg  <= \piso.data_li [1508];
      \piso.data_r_1507_sv2v_reg  <= \piso.data_li [1507];
      \piso.data_r_1506_sv2v_reg  <= \piso.data_li [1506];
      \piso.data_r_1505_sv2v_reg  <= \piso.data_li [1505];
      \piso.data_r_1504_sv2v_reg  <= \piso.data_li [1504];
      \piso.data_r_1503_sv2v_reg  <= \piso.data_li [1503];
      \piso.data_r_1502_sv2v_reg  <= \piso.data_li [1502];
      \piso.data_r_1501_sv2v_reg  <= \piso.data_li [1501];
      \piso.data_r_1500_sv2v_reg  <= \piso.data_li [1500];
      \piso.data_r_1499_sv2v_reg  <= \piso.data_li [1499];
      \piso.data_r_1498_sv2v_reg  <= \piso.data_li [1498];
      \piso.data_r_1497_sv2v_reg  <= \piso.data_li [1497];
      \piso.data_r_1496_sv2v_reg  <= \piso.data_li [1496];
      \piso.data_r_1495_sv2v_reg  <= \piso.data_li [1495];
      \piso.data_r_1494_sv2v_reg  <= \piso.data_li [1494];
      \piso.data_r_1493_sv2v_reg  <= \piso.data_li [1493];
      \piso.data_r_1492_sv2v_reg  <= \piso.data_li [1492];
      \piso.data_r_1491_sv2v_reg  <= \piso.data_li [1491];
      \piso.data_r_1490_sv2v_reg  <= \piso.data_li [1490];
      \piso.data_r_1489_sv2v_reg  <= \piso.data_li [1489];
      \piso.data_r_1488_sv2v_reg  <= \piso.data_li [1488];
      \piso.data_r_1487_sv2v_reg  <= \piso.data_li [1487];
      \piso.data_r_1486_sv2v_reg  <= \piso.data_li [1486];
      \piso.data_r_1485_sv2v_reg  <= \piso.data_li [1485];
      \piso.data_r_1484_sv2v_reg  <= \piso.data_li [1484];
      \piso.data_r_1483_sv2v_reg  <= \piso.data_li [1483];
      \piso.data_r_1482_sv2v_reg  <= \piso.data_li [1482];
      \piso.data_r_1481_sv2v_reg  <= \piso.data_li [1481];
      \piso.data_r_1480_sv2v_reg  <= \piso.data_li [1480];
      \piso.data_r_1479_sv2v_reg  <= \piso.data_li [1479];
      \piso.data_r_1478_sv2v_reg  <= \piso.data_li [1478];
      \piso.data_r_1477_sv2v_reg  <= \piso.data_li [1477];
      \piso.data_r_1476_sv2v_reg  <= \piso.data_li [1476];
      \piso.data_r_1475_sv2v_reg  <= \piso.data_li [1475];
      \piso.data_r_1474_sv2v_reg  <= \piso.data_li [1474];
      \piso.data_r_1473_sv2v_reg  <= \piso.data_li [1473];
      \piso.data_r_1472_sv2v_reg  <= \piso.data_li [1472];
      \piso.data_r_1471_sv2v_reg  <= \piso.data_li [1471];
      \piso.data_r_1470_sv2v_reg  <= \piso.data_li [1470];
      \piso.data_r_1469_sv2v_reg  <= \piso.data_li [1469];
      \piso.data_r_1468_sv2v_reg  <= \piso.data_li [1468];
      \piso.data_r_1467_sv2v_reg  <= \piso.data_li [1467];
      \piso.data_r_1466_sv2v_reg  <= \piso.data_li [1466];
      \piso.data_r_1465_sv2v_reg  <= \piso.data_li [1465];
      \piso.data_r_1464_sv2v_reg  <= \piso.data_li [1464];
      \piso.data_r_1463_sv2v_reg  <= \piso.data_li [1463];
      \piso.data_r_1462_sv2v_reg  <= \piso.data_li [1462];
      \piso.data_r_1461_sv2v_reg  <= \piso.data_li [1461];
      \piso.data_r_1460_sv2v_reg  <= \piso.data_li [1460];
      \piso.data_r_1459_sv2v_reg  <= \piso.data_li [1459];
      \piso.data_r_1458_sv2v_reg  <= \piso.data_li [1458];
      \piso.data_r_1457_sv2v_reg  <= \piso.data_li [1457];
      \piso.data_r_1456_sv2v_reg  <= \piso.data_li [1456];
      \piso.data_r_1455_sv2v_reg  <= \piso.data_li [1455];
      \piso.data_r_1454_sv2v_reg  <= \piso.data_li [1454];
      \piso.data_r_1453_sv2v_reg  <= \piso.data_li [1453];
      \piso.data_r_1452_sv2v_reg  <= \piso.data_li [1452];
      \piso.data_r_1451_sv2v_reg  <= \piso.data_li [1451];
      \piso.data_r_1450_sv2v_reg  <= \piso.data_li [1450];
      \piso.data_r_1449_sv2v_reg  <= \piso.data_li [1449];
      \piso.data_r_1448_sv2v_reg  <= \piso.data_li [1448];
      \piso.data_r_1447_sv2v_reg  <= \piso.data_li [1447];
      \piso.data_r_1446_sv2v_reg  <= \piso.data_li [1446];
      \piso.data_r_1445_sv2v_reg  <= \piso.data_li [1445];
      \piso.data_r_1444_sv2v_reg  <= \piso.data_li [1444];
      \piso.data_r_1443_sv2v_reg  <= \piso.data_li [1443];
      \piso.data_r_1442_sv2v_reg  <= \piso.data_li [1442];
      \piso.data_r_1441_sv2v_reg  <= \piso.data_li [1441];
      \piso.data_r_1440_sv2v_reg  <= \piso.data_li [1440];
      \piso.data_r_1439_sv2v_reg  <= \piso.data_li [1439];
      \piso.data_r_1438_sv2v_reg  <= \piso.data_li [1438];
      \piso.data_r_1437_sv2v_reg  <= \piso.data_li [1437];
      \piso.data_r_1436_sv2v_reg  <= \piso.data_li [1436];
      \piso.data_r_1435_sv2v_reg  <= \piso.data_li [1435];
      \piso.data_r_1434_sv2v_reg  <= \piso.data_li [1434];
      \piso.data_r_1433_sv2v_reg  <= \piso.data_li [1433];
      \piso.data_r_1432_sv2v_reg  <= \piso.data_li [1432];
      \piso.data_r_1431_sv2v_reg  <= \piso.data_li [1431];
      \piso.data_r_1430_sv2v_reg  <= \piso.data_li [1430];
      \piso.data_r_1429_sv2v_reg  <= \piso.data_li [1429];
      \piso.data_r_1428_sv2v_reg  <= \piso.data_li [1428];
      \piso.data_r_1427_sv2v_reg  <= \piso.data_li [1427];
      \piso.data_r_1426_sv2v_reg  <= \piso.data_li [1426];
      \piso.data_r_1425_sv2v_reg  <= \piso.data_li [1425];
      \piso.data_r_1424_sv2v_reg  <= \piso.data_li [1424];
      \piso.data_r_1423_sv2v_reg  <= \piso.data_li [1423];
      \piso.data_r_1422_sv2v_reg  <= \piso.data_li [1422];
      \piso.data_r_1421_sv2v_reg  <= \piso.data_li [1421];
      \piso.data_r_1420_sv2v_reg  <= \piso.data_li [1420];
      \piso.data_r_1419_sv2v_reg  <= \piso.data_li [1419];
      \piso.data_r_1418_sv2v_reg  <= \piso.data_li [1418];
      \piso.data_r_1417_sv2v_reg  <= \piso.data_li [1417];
      \piso.data_r_1416_sv2v_reg  <= \piso.data_li [1416];
      \piso.data_r_1415_sv2v_reg  <= \piso.data_li [1415];
      \piso.data_r_1414_sv2v_reg  <= \piso.data_li [1414];
      \piso.data_r_1413_sv2v_reg  <= \piso.data_li [1413];
      \piso.data_r_1412_sv2v_reg  <= \piso.data_li [1412];
      \piso.data_r_1411_sv2v_reg  <= \piso.data_li [1411];
      \piso.data_r_1410_sv2v_reg  <= \piso.data_li [1410];
      \piso.data_r_1409_sv2v_reg  <= \piso.data_li [1409];
      \piso.data_r_1408_sv2v_reg  <= \piso.data_li [1408];
      \piso.data_r_1407_sv2v_reg  <= \piso.data_li [1407];
      \piso.data_r_1406_sv2v_reg  <= \piso.data_li [1406];
      \piso.data_r_1405_sv2v_reg  <= \piso.data_li [1405];
      \piso.data_r_1404_sv2v_reg  <= \piso.data_li [1404];
      \piso.data_r_1403_sv2v_reg  <= \piso.data_li [1403];
      \piso.data_r_1402_sv2v_reg  <= \piso.data_li [1402];
      \piso.data_r_1401_sv2v_reg  <= \piso.data_li [1401];
      \piso.data_r_1400_sv2v_reg  <= \piso.data_li [1400];
      \piso.data_r_1399_sv2v_reg  <= \piso.data_li [1399];
      \piso.data_r_1398_sv2v_reg  <= \piso.data_li [1398];
      \piso.data_r_1397_sv2v_reg  <= \piso.data_li [1397];
      \piso.data_r_1396_sv2v_reg  <= \piso.data_li [1396];
      \piso.data_r_1395_sv2v_reg  <= \piso.data_li [1395];
      \piso.data_r_1394_sv2v_reg  <= \piso.data_li [1394];
      \piso.data_r_1393_sv2v_reg  <= \piso.data_li [1393];
      \piso.data_r_1392_sv2v_reg  <= \piso.data_li [1392];
      \piso.data_r_1391_sv2v_reg  <= \piso.data_li [1391];
      \piso.data_r_1390_sv2v_reg  <= \piso.data_li [1390];
      \piso.data_r_1389_sv2v_reg  <= \piso.data_li [1389];
      \piso.data_r_1388_sv2v_reg  <= \piso.data_li [1388];
      \piso.data_r_1387_sv2v_reg  <= \piso.data_li [1387];
      \piso.data_r_1386_sv2v_reg  <= \piso.data_li [1386];
      \piso.data_r_1385_sv2v_reg  <= \piso.data_li [1385];
      \piso.data_r_1384_sv2v_reg  <= \piso.data_li [1384];
      \piso.data_r_1383_sv2v_reg  <= \piso.data_li [1383];
      \piso.data_r_1382_sv2v_reg  <= \piso.data_li [1382];
      \piso.data_r_1381_sv2v_reg  <= \piso.data_li [1381];
      \piso.data_r_1380_sv2v_reg  <= \piso.data_li [1380];
      \piso.data_r_1379_sv2v_reg  <= \piso.data_li [1379];
      \piso.data_r_1378_sv2v_reg  <= \piso.data_li [1378];
      \piso.data_r_1377_sv2v_reg  <= \piso.data_li [1377];
      \piso.data_r_1376_sv2v_reg  <= \piso.data_li [1376];
      \piso.data_r_1375_sv2v_reg  <= \piso.data_li [1375];
      \piso.data_r_1374_sv2v_reg  <= \piso.data_li [1374];
      \piso.data_r_1373_sv2v_reg  <= \piso.data_li [1373];
      \piso.data_r_1372_sv2v_reg  <= \piso.data_li [1372];
      \piso.data_r_1371_sv2v_reg  <= \piso.data_li [1371];
      \piso.data_r_1370_sv2v_reg  <= \piso.data_li [1370];
      \piso.data_r_1369_sv2v_reg  <= \piso.data_li [1369];
      \piso.data_r_1368_sv2v_reg  <= \piso.data_li [1368];
      \piso.data_r_1367_sv2v_reg  <= \piso.data_li [1367];
      \piso.data_r_1366_sv2v_reg  <= \piso.data_li [1366];
      \piso.data_r_1365_sv2v_reg  <= \piso.data_li [1365];
      \piso.data_r_1364_sv2v_reg  <= \piso.data_li [1364];
      \piso.data_r_1363_sv2v_reg  <= \piso.data_li [1363];
      \piso.data_r_1362_sv2v_reg  <= \piso.data_li [1362];
      \piso.data_r_1361_sv2v_reg  <= \piso.data_li [1361];
      \piso.data_r_1360_sv2v_reg  <= \piso.data_li [1360];
      \piso.data_r_1359_sv2v_reg  <= \piso.data_li [1359];
      \piso.data_r_1358_sv2v_reg  <= \piso.data_li [1358];
      \piso.data_r_1357_sv2v_reg  <= \piso.data_li [1357];
      \piso.data_r_1356_sv2v_reg  <= \piso.data_li [1356];
      \piso.data_r_1355_sv2v_reg  <= \piso.data_li [1355];
      \piso.data_r_1354_sv2v_reg  <= \piso.data_li [1354];
      \piso.data_r_1353_sv2v_reg  <= \piso.data_li [1353];
      \piso.data_r_1352_sv2v_reg  <= \piso.data_li [1352];
      \piso.data_r_1351_sv2v_reg  <= \piso.data_li [1351];
      \piso.data_r_1350_sv2v_reg  <= \piso.data_li [1350];
      \piso.data_r_1349_sv2v_reg  <= \piso.data_li [1349];
      \piso.data_r_1348_sv2v_reg  <= \piso.data_li [1348];
      \piso.data_r_1347_sv2v_reg  <= \piso.data_li [1347];
      \piso.data_r_1346_sv2v_reg  <= \piso.data_li [1346];
      \piso.data_r_1345_sv2v_reg  <= \piso.data_li [1345];
      \piso.data_r_1344_sv2v_reg  <= \piso.data_li [1344];
      \piso.data_r_1343_sv2v_reg  <= \piso.data_li [1343];
      \piso.data_r_1342_sv2v_reg  <= \piso.data_li [1342];
      \piso.data_r_1341_sv2v_reg  <= \piso.data_li [1341];
      \piso.data_r_1340_sv2v_reg  <= \piso.data_li [1340];
      \piso.data_r_1339_sv2v_reg  <= \piso.data_li [1339];
      \piso.data_r_1338_sv2v_reg  <= \piso.data_li [1338];
      \piso.data_r_1337_sv2v_reg  <= \piso.data_li [1337];
      \piso.data_r_1336_sv2v_reg  <= \piso.data_li [1336];
      \piso.data_r_1335_sv2v_reg  <= \piso.data_li [1335];
      \piso.data_r_1334_sv2v_reg  <= \piso.data_li [1334];
      \piso.data_r_1333_sv2v_reg  <= \piso.data_li [1333];
      \piso.data_r_1332_sv2v_reg  <= \piso.data_li [1332];
      \piso.data_r_1331_sv2v_reg  <= \piso.data_li [1331];
      \piso.data_r_1330_sv2v_reg  <= \piso.data_li [1330];
      \piso.data_r_1329_sv2v_reg  <= \piso.data_li [1329];
      \piso.data_r_1328_sv2v_reg  <= \piso.data_li [1328];
      \piso.data_r_1327_sv2v_reg  <= \piso.data_li [1327];
      \piso.data_r_1326_sv2v_reg  <= \piso.data_li [1326];
      \piso.data_r_1325_sv2v_reg  <= \piso.data_li [1325];
      \piso.data_r_1324_sv2v_reg  <= \piso.data_li [1324];
      \piso.data_r_1323_sv2v_reg  <= \piso.data_li [1323];
      \piso.data_r_1322_sv2v_reg  <= \piso.data_li [1322];
      \piso.data_r_1321_sv2v_reg  <= \piso.data_li [1321];
      \piso.data_r_1320_sv2v_reg  <= \piso.data_li [1320];
      \piso.data_r_1319_sv2v_reg  <= \piso.data_li [1319];
      \piso.data_r_1318_sv2v_reg  <= \piso.data_li [1318];
      \piso.data_r_1317_sv2v_reg  <= \piso.data_li [1317];
      \piso.data_r_1316_sv2v_reg  <= \piso.data_li [1316];
      \piso.data_r_1315_sv2v_reg  <= \piso.data_li [1315];
      \piso.data_r_1314_sv2v_reg  <= \piso.data_li [1314];
      \piso.data_r_1313_sv2v_reg  <= \piso.data_li [1313];
      \piso.data_r_1312_sv2v_reg  <= \piso.data_li [1312];
      \piso.data_r_1311_sv2v_reg  <= \piso.data_li [1311];
      \piso.data_r_1310_sv2v_reg  <= \piso.data_li [1310];
      \piso.data_r_1309_sv2v_reg  <= \piso.data_li [1309];
      \piso.data_r_1308_sv2v_reg  <= \piso.data_li [1308];
      \piso.data_r_1307_sv2v_reg  <= \piso.data_li [1307];
      \piso.data_r_1306_sv2v_reg  <= \piso.data_li [1306];
      \piso.data_r_1305_sv2v_reg  <= \piso.data_li [1305];
      \piso.data_r_1304_sv2v_reg  <= \piso.data_li [1304];
      \piso.data_r_1303_sv2v_reg  <= \piso.data_li [1303];
      \piso.data_r_1302_sv2v_reg  <= \piso.data_li [1302];
      \piso.data_r_1301_sv2v_reg  <= \piso.data_li [1301];
      \piso.data_r_1300_sv2v_reg  <= \piso.data_li [1300];
      \piso.data_r_1299_sv2v_reg  <= \piso.data_li [1299];
      \piso.data_r_1298_sv2v_reg  <= \piso.data_li [1298];
      \piso.data_r_1297_sv2v_reg  <= \piso.data_li [1297];
      \piso.data_r_1296_sv2v_reg  <= \piso.data_li [1296];
      \piso.data_r_1295_sv2v_reg  <= \piso.data_li [1295];
      \piso.data_r_1294_sv2v_reg  <= \piso.data_li [1294];
      \piso.data_r_1293_sv2v_reg  <= \piso.data_li [1293];
      \piso.data_r_1292_sv2v_reg  <= \piso.data_li [1292];
      \piso.data_r_1291_sv2v_reg  <= \piso.data_li [1291];
      \piso.data_r_1290_sv2v_reg  <= \piso.data_li [1290];
      \piso.data_r_1289_sv2v_reg  <= \piso.data_li [1289];
      \piso.data_r_1288_sv2v_reg  <= \piso.data_li [1288];
      \piso.data_r_1287_sv2v_reg  <= \piso.data_li [1287];
      \piso.data_r_1286_sv2v_reg  <= \piso.data_li [1286];
      \piso.data_r_1285_sv2v_reg  <= \piso.data_li [1285];
      \piso.data_r_1284_sv2v_reg  <= \piso.data_li [1284];
      \piso.data_r_1283_sv2v_reg  <= \piso.data_li [1283];
      \piso.data_r_1282_sv2v_reg  <= \piso.data_li [1282];
      \piso.data_r_1281_sv2v_reg  <= \piso.data_li [1281];
      \piso.data_r_1280_sv2v_reg  <= \piso.data_li [1280];
      \piso.data_r_1279_sv2v_reg  <= \piso.data_li [1279];
      \piso.data_r_1278_sv2v_reg  <= \piso.data_li [1278];
      \piso.data_r_1277_sv2v_reg  <= \piso.data_li [1277];
      \piso.data_r_1276_sv2v_reg  <= \piso.data_li [1276];
      \piso.data_r_1275_sv2v_reg  <= \piso.data_li [1275];
      \piso.data_r_1274_sv2v_reg  <= \piso.data_li [1274];
      \piso.data_r_1273_sv2v_reg  <= \piso.data_li [1273];
      \piso.data_r_1272_sv2v_reg  <= \piso.data_li [1272];
      \piso.data_r_1271_sv2v_reg  <= \piso.data_li [1271];
      \piso.data_r_1270_sv2v_reg  <= \piso.data_li [1270];
      \piso.data_r_1269_sv2v_reg  <= \piso.data_li [1269];
      \piso.data_r_1268_sv2v_reg  <= \piso.data_li [1268];
      \piso.data_r_1267_sv2v_reg  <= \piso.data_li [1267];
      \piso.data_r_1266_sv2v_reg  <= \piso.data_li [1266];
      \piso.data_r_1265_sv2v_reg  <= \piso.data_li [1265];
      \piso.data_r_1264_sv2v_reg  <= \piso.data_li [1264];
      \piso.data_r_1263_sv2v_reg  <= \piso.data_li [1263];
      \piso.data_r_1262_sv2v_reg  <= \piso.data_li [1262];
      \piso.data_r_1261_sv2v_reg  <= \piso.data_li [1261];
      \piso.data_r_1260_sv2v_reg  <= \piso.data_li [1260];
      \piso.data_r_1259_sv2v_reg  <= \piso.data_li [1259];
      \piso.data_r_1258_sv2v_reg  <= \piso.data_li [1258];
      \piso.data_r_1257_sv2v_reg  <= \piso.data_li [1257];
      \piso.data_r_1256_sv2v_reg  <= \piso.data_li [1256];
      \piso.data_r_1255_sv2v_reg  <= \piso.data_li [1255];
      \piso.data_r_1254_sv2v_reg  <= \piso.data_li [1254];
      \piso.data_r_1253_sv2v_reg  <= \piso.data_li [1253];
      \piso.data_r_1252_sv2v_reg  <= \piso.data_li [1252];
      \piso.data_r_1251_sv2v_reg  <= \piso.data_li [1251];
      \piso.data_r_1250_sv2v_reg  <= \piso.data_li [1250];
      \piso.data_r_1249_sv2v_reg  <= \piso.data_li [1249];
      \piso.data_r_1248_sv2v_reg  <= \piso.data_li [1248];
      \piso.data_r_1247_sv2v_reg  <= \piso.data_li [1247];
      \piso.data_r_1246_sv2v_reg  <= \piso.data_li [1246];
      \piso.data_r_1245_sv2v_reg  <= \piso.data_li [1245];
      \piso.data_r_1244_sv2v_reg  <= \piso.data_li [1244];
      \piso.data_r_1243_sv2v_reg  <= \piso.data_li [1243];
      \piso.data_r_1242_sv2v_reg  <= \piso.data_li [1242];
      \piso.data_r_1241_sv2v_reg  <= \piso.data_li [1241];
      \piso.data_r_1240_sv2v_reg  <= \piso.data_li [1240];
      \piso.data_r_1239_sv2v_reg  <= \piso.data_li [1239];
      \piso.data_r_1238_sv2v_reg  <= \piso.data_li [1238];
      \piso.data_r_1237_sv2v_reg  <= \piso.data_li [1237];
      \piso.data_r_1236_sv2v_reg  <= \piso.data_li [1236];
      \piso.data_r_1235_sv2v_reg  <= \piso.data_li [1235];
      \piso.data_r_1234_sv2v_reg  <= \piso.data_li [1234];
      \piso.data_r_1233_sv2v_reg  <= \piso.data_li [1233];
      \piso.data_r_1232_sv2v_reg  <= \piso.data_li [1232];
      \piso.data_r_1231_sv2v_reg  <= \piso.data_li [1231];
      \piso.data_r_1230_sv2v_reg  <= \piso.data_li [1230];
      \piso.data_r_1229_sv2v_reg  <= \piso.data_li [1229];
      \piso.data_r_1228_sv2v_reg  <= \piso.data_li [1228];
      \piso.data_r_1227_sv2v_reg  <= \piso.data_li [1227];
      \piso.data_r_1226_sv2v_reg  <= \piso.data_li [1226];
      \piso.data_r_1225_sv2v_reg  <= \piso.data_li [1225];
      \piso.data_r_1224_sv2v_reg  <= \piso.data_li [1224];
      \piso.data_r_1223_sv2v_reg  <= \piso.data_li [1223];
      \piso.data_r_1222_sv2v_reg  <= \piso.data_li [1222];
      \piso.data_r_1221_sv2v_reg  <= \piso.data_li [1221];
      \piso.data_r_1220_sv2v_reg  <= \piso.data_li [1220];
      \piso.data_r_1219_sv2v_reg  <= \piso.data_li [1219];
      \piso.data_r_1218_sv2v_reg  <= \piso.data_li [1218];
      \piso.data_r_1217_sv2v_reg  <= \piso.data_li [1217];
      \piso.data_r_1216_sv2v_reg  <= \piso.data_li [1216];
      \piso.data_r_1215_sv2v_reg  <= \piso.data_li [1215];
      \piso.data_r_1214_sv2v_reg  <= \piso.data_li [1214];
      \piso.data_r_1213_sv2v_reg  <= \piso.data_li [1213];
      \piso.data_r_1212_sv2v_reg  <= \piso.data_li [1212];
      \piso.data_r_1211_sv2v_reg  <= \piso.data_li [1211];
      \piso.data_r_1210_sv2v_reg  <= \piso.data_li [1210];
      \piso.data_r_1209_sv2v_reg  <= \piso.data_li [1209];
      \piso.data_r_1208_sv2v_reg  <= \piso.data_li [1208];
      \piso.data_r_1207_sv2v_reg  <= \piso.data_li [1207];
      \piso.data_r_1206_sv2v_reg  <= \piso.data_li [1206];
      \piso.data_r_1205_sv2v_reg  <= \piso.data_li [1205];
      \piso.data_r_1204_sv2v_reg  <= \piso.data_li [1204];
      \piso.data_r_1203_sv2v_reg  <= \piso.data_li [1203];
      \piso.data_r_1202_sv2v_reg  <= \piso.data_li [1202];
      \piso.data_r_1201_sv2v_reg  <= \piso.data_li [1201];
      \piso.data_r_1200_sv2v_reg  <= \piso.data_li [1200];
      \piso.data_r_1199_sv2v_reg  <= \piso.data_li [1199];
      \piso.data_r_1198_sv2v_reg  <= \piso.data_li [1198];
      \piso.data_r_1197_sv2v_reg  <= \piso.data_li [1197];
      \piso.data_r_1196_sv2v_reg  <= \piso.data_li [1196];
      \piso.data_r_1195_sv2v_reg  <= \piso.data_li [1195];
      \piso.data_r_1194_sv2v_reg  <= \piso.data_li [1194];
      \piso.data_r_1193_sv2v_reg  <= \piso.data_li [1193];
      \piso.data_r_1192_sv2v_reg  <= \piso.data_li [1192];
      \piso.data_r_1191_sv2v_reg  <= \piso.data_li [1191];
      \piso.data_r_1190_sv2v_reg  <= \piso.data_li [1190];
      \piso.data_r_1189_sv2v_reg  <= \piso.data_li [1189];
      \piso.data_r_1188_sv2v_reg  <= \piso.data_li [1188];
      \piso.data_r_1187_sv2v_reg  <= \piso.data_li [1187];
      \piso.data_r_1186_sv2v_reg  <= \piso.data_li [1186];
      \piso.data_r_1185_sv2v_reg  <= \piso.data_li [1185];
      \piso.data_r_1184_sv2v_reg  <= \piso.data_li [1184];
      \piso.data_r_1183_sv2v_reg  <= \piso.data_li [1183];
      \piso.data_r_1182_sv2v_reg  <= \piso.data_li [1182];
      \piso.data_r_1181_sv2v_reg  <= \piso.data_li [1181];
      \piso.data_r_1180_sv2v_reg  <= \piso.data_li [1180];
      \piso.data_r_1179_sv2v_reg  <= \piso.data_li [1179];
      \piso.data_r_1178_sv2v_reg  <= \piso.data_li [1178];
      \piso.data_r_1177_sv2v_reg  <= \piso.data_li [1177];
      \piso.data_r_1176_sv2v_reg  <= \piso.data_li [1176];
      \piso.data_r_1175_sv2v_reg  <= \piso.data_li [1175];
      \piso.data_r_1174_sv2v_reg  <= \piso.data_li [1174];
      \piso.data_r_1173_sv2v_reg  <= \piso.data_li [1173];
      \piso.data_r_1172_sv2v_reg  <= \piso.data_li [1172];
      \piso.data_r_1171_sv2v_reg  <= \piso.data_li [1171];
      \piso.data_r_1170_sv2v_reg  <= \piso.data_li [1170];
      \piso.data_r_1169_sv2v_reg  <= \piso.data_li [1169];
      \piso.data_r_1168_sv2v_reg  <= \piso.data_li [1168];
      \piso.data_r_1167_sv2v_reg  <= \piso.data_li [1167];
      \piso.data_r_1166_sv2v_reg  <= \piso.data_li [1166];
      \piso.data_r_1165_sv2v_reg  <= \piso.data_li [1165];
      \piso.data_r_1164_sv2v_reg  <= \piso.data_li [1164];
      \piso.data_r_1163_sv2v_reg  <= \piso.data_li [1163];
      \piso.data_r_1162_sv2v_reg  <= \piso.data_li [1162];
      \piso.data_r_1161_sv2v_reg  <= \piso.data_li [1161];
      \piso.data_r_1160_sv2v_reg  <= \piso.data_li [1160];
      \piso.data_r_1159_sv2v_reg  <= \piso.data_li [1159];
      \piso.data_r_1158_sv2v_reg  <= \piso.data_li [1158];
      \piso.data_r_1157_sv2v_reg  <= \piso.data_li [1157];
      \piso.data_r_1156_sv2v_reg  <= \piso.data_li [1156];
      \piso.data_r_1155_sv2v_reg  <= \piso.data_li [1155];
      \piso.data_r_1154_sv2v_reg  <= \piso.data_li [1154];
      \piso.data_r_1153_sv2v_reg  <= \piso.data_li [1153];
      \piso.data_r_1152_sv2v_reg  <= \piso.data_li [1152];
      \piso.data_r_1151_sv2v_reg  <= \piso.data_li [1151];
      \piso.data_r_1150_sv2v_reg  <= \piso.data_li [1150];
      \piso.data_r_1149_sv2v_reg  <= \piso.data_li [1149];
      \piso.data_r_1148_sv2v_reg  <= \piso.data_li [1148];
      \piso.data_r_1147_sv2v_reg  <= \piso.data_li [1147];
      \piso.data_r_1146_sv2v_reg  <= \piso.data_li [1146];
      \piso.data_r_1145_sv2v_reg  <= \piso.data_li [1145];
      \piso.data_r_1144_sv2v_reg  <= \piso.data_li [1144];
      \piso.data_r_1143_sv2v_reg  <= \piso.data_li [1143];
      \piso.data_r_1142_sv2v_reg  <= \piso.data_li [1142];
      \piso.data_r_1141_sv2v_reg  <= \piso.data_li [1141];
      \piso.data_r_1140_sv2v_reg  <= \piso.data_li [1140];
      \piso.data_r_1139_sv2v_reg  <= \piso.data_li [1139];
      \piso.data_r_1138_sv2v_reg  <= \piso.data_li [1138];
      \piso.data_r_1137_sv2v_reg  <= \piso.data_li [1137];
      \piso.data_r_1136_sv2v_reg  <= \piso.data_li [1136];
      \piso.data_r_1135_sv2v_reg  <= \piso.data_li [1135];
      \piso.data_r_1134_sv2v_reg  <= \piso.data_li [1134];
      \piso.data_r_1133_sv2v_reg  <= \piso.data_li [1133];
      \piso.data_r_1132_sv2v_reg  <= \piso.data_li [1132];
      \piso.data_r_1131_sv2v_reg  <= \piso.data_li [1131];
      \piso.data_r_1130_sv2v_reg  <= \piso.data_li [1130];
      \piso.data_r_1129_sv2v_reg  <= \piso.data_li [1129];
      \piso.data_r_1128_sv2v_reg  <= \piso.data_li [1128];
      \piso.data_r_1127_sv2v_reg  <= \piso.data_li [1127];
      \piso.data_r_1126_sv2v_reg  <= \piso.data_li [1126];
      \piso.data_r_1125_sv2v_reg  <= \piso.data_li [1125];
      \piso.data_r_1124_sv2v_reg  <= \piso.data_li [1124];
      \piso.data_r_1123_sv2v_reg  <= \piso.data_li [1123];
      \piso.data_r_1122_sv2v_reg  <= \piso.data_li [1122];
      \piso.data_r_1121_sv2v_reg  <= \piso.data_li [1121];
      \piso.data_r_1120_sv2v_reg  <= \piso.data_li [1120];
      \piso.data_r_1119_sv2v_reg  <= \piso.data_li [1119];
      \piso.data_r_1118_sv2v_reg  <= \piso.data_li [1118];
      \piso.data_r_1117_sv2v_reg  <= \piso.data_li [1117];
      \piso.data_r_1116_sv2v_reg  <= \piso.data_li [1116];
      \piso.data_r_1115_sv2v_reg  <= \piso.data_li [1115];
      \piso.data_r_1114_sv2v_reg  <= \piso.data_li [1114];
      \piso.data_r_1113_sv2v_reg  <= \piso.data_li [1113];
      \piso.data_r_1112_sv2v_reg  <= \piso.data_li [1112];
      \piso.data_r_1111_sv2v_reg  <= \piso.data_li [1111];
      \piso.data_r_1110_sv2v_reg  <= \piso.data_li [1110];
      \piso.data_r_1109_sv2v_reg  <= \piso.data_li [1109];
      \piso.data_r_1108_sv2v_reg  <= \piso.data_li [1108];
      \piso.data_r_1107_sv2v_reg  <= \piso.data_li [1107];
      \piso.data_r_1106_sv2v_reg  <= \piso.data_li [1106];
      \piso.data_r_1105_sv2v_reg  <= \piso.data_li [1105];
      \piso.data_r_1104_sv2v_reg  <= \piso.data_li [1104];
      \piso.data_r_1103_sv2v_reg  <= \piso.data_li [1103];
      \piso.data_r_1102_sv2v_reg  <= \piso.data_li [1102];
      \piso.data_r_1101_sv2v_reg  <= \piso.data_li [1101];
      \piso.data_r_1100_sv2v_reg  <= \piso.data_li [1100];
      \piso.data_r_1099_sv2v_reg  <= \piso.data_li [1099];
      \piso.data_r_1098_sv2v_reg  <= \piso.data_li [1098];
      \piso.data_r_1097_sv2v_reg  <= \piso.data_li [1097];
      \piso.data_r_1096_sv2v_reg  <= \piso.data_li [1096];
      \piso.data_r_1095_sv2v_reg  <= \piso.data_li [1095];
      \piso.data_r_1094_sv2v_reg  <= \piso.data_li [1094];
      \piso.data_r_1093_sv2v_reg  <= \piso.data_li [1093];
      \piso.data_r_1092_sv2v_reg  <= \piso.data_li [1092];
      \piso.data_r_1091_sv2v_reg  <= \piso.data_li [1091];
      \piso.data_r_1090_sv2v_reg  <= \piso.data_li [1090];
      \piso.data_r_1089_sv2v_reg  <= \piso.data_li [1089];
      \piso.data_r_1088_sv2v_reg  <= \piso.data_li [1088];
      \piso.data_r_1087_sv2v_reg  <= \piso.data_li [1087];
      \piso.data_r_1086_sv2v_reg  <= \piso.data_li [1086];
      \piso.data_r_1085_sv2v_reg  <= \piso.data_li [1085];
      \piso.data_r_1084_sv2v_reg  <= \piso.data_li [1084];
      \piso.data_r_1083_sv2v_reg  <= \piso.data_li [1083];
      \piso.data_r_1082_sv2v_reg  <= \piso.data_li [1082];
      \piso.data_r_1081_sv2v_reg  <= \piso.data_li [1081];
      \piso.data_r_1080_sv2v_reg  <= \piso.data_li [1080];
      \piso.data_r_1079_sv2v_reg  <= \piso.data_li [1079];
      \piso.data_r_1078_sv2v_reg  <= \piso.data_li [1078];
      \piso.data_r_1077_sv2v_reg  <= \piso.data_li [1077];
      \piso.data_r_1076_sv2v_reg  <= \piso.data_li [1076];
      \piso.data_r_1075_sv2v_reg  <= \piso.data_li [1075];
      \piso.data_r_1074_sv2v_reg  <= \piso.data_li [1074];
      \piso.data_r_1073_sv2v_reg  <= \piso.data_li [1073];
      \piso.data_r_1072_sv2v_reg  <= \piso.data_li [1072];
      \piso.data_r_1071_sv2v_reg  <= \piso.data_li [1071];
      \piso.data_r_1070_sv2v_reg  <= \piso.data_li [1070];
      \piso.data_r_1069_sv2v_reg  <= \piso.data_li [1069];
      \piso.data_r_1068_sv2v_reg  <= \piso.data_li [1068];
      \piso.data_r_1067_sv2v_reg  <= \piso.data_li [1067];
      \piso.data_r_1066_sv2v_reg  <= \piso.data_li [1066];
      \piso.data_r_1065_sv2v_reg  <= \piso.data_li [1065];
      \piso.data_r_1064_sv2v_reg  <= \piso.data_li [1064];
      \piso.data_r_1063_sv2v_reg  <= \piso.data_li [1063];
      \piso.data_r_1062_sv2v_reg  <= \piso.data_li [1062];
      \piso.data_r_1061_sv2v_reg  <= \piso.data_li [1061];
      \piso.data_r_1060_sv2v_reg  <= \piso.data_li [1060];
      \piso.data_r_1059_sv2v_reg  <= \piso.data_li [1059];
      \piso.data_r_1058_sv2v_reg  <= \piso.data_li [1058];
      \piso.data_r_1057_sv2v_reg  <= \piso.data_li [1057];
      \piso.data_r_1056_sv2v_reg  <= \piso.data_li [1056];
      \piso.data_r_1055_sv2v_reg  <= \piso.data_li [1055];
      \piso.data_r_1054_sv2v_reg  <= \piso.data_li [1054];
      \piso.data_r_1053_sv2v_reg  <= \piso.data_li [1053];
      \piso.data_r_1052_sv2v_reg  <= \piso.data_li [1052];
      \piso.data_r_1051_sv2v_reg  <= \piso.data_li [1051];
      \piso.data_r_1050_sv2v_reg  <= \piso.data_li [1050];
      \piso.data_r_1049_sv2v_reg  <= \piso.data_li [1049];
      \piso.data_r_1048_sv2v_reg  <= \piso.data_li [1048];
      \piso.data_r_1047_sv2v_reg  <= \piso.data_li [1047];
      \piso.data_r_1046_sv2v_reg  <= \piso.data_li [1046];
      \piso.data_r_1045_sv2v_reg  <= \piso.data_li [1045];
      \piso.data_r_1044_sv2v_reg  <= \piso.data_li [1044];
      \piso.data_r_1043_sv2v_reg  <= \piso.data_li [1043];
      \piso.data_r_1042_sv2v_reg  <= \piso.data_li [1042];
      \piso.data_r_1041_sv2v_reg  <= \piso.data_li [1041];
      \piso.data_r_1040_sv2v_reg  <= \piso.data_li [1040];
      \piso.data_r_1039_sv2v_reg  <= \piso.data_li [1039];
      \piso.data_r_1038_sv2v_reg  <= \piso.data_li [1038];
      \piso.data_r_1037_sv2v_reg  <= \piso.data_li [1037];
      \piso.data_r_1036_sv2v_reg  <= \piso.data_li [1036];
      \piso.data_r_1035_sv2v_reg  <= \piso.data_li [1035];
      \piso.data_r_1034_sv2v_reg  <= \piso.data_li [1034];
      \piso.data_r_1033_sv2v_reg  <= \piso.data_li [1033];
      \piso.data_r_1032_sv2v_reg  <= \piso.data_li [1032];
      \piso.data_r_1031_sv2v_reg  <= \piso.data_li [1031];
      \piso.data_r_1030_sv2v_reg  <= \piso.data_li [1030];
      \piso.data_r_1029_sv2v_reg  <= \piso.data_li [1029];
      \piso.data_r_1028_sv2v_reg  <= \piso.data_li [1028];
      \piso.data_r_1027_sv2v_reg  <= \piso.data_li [1027];
      \piso.data_r_1026_sv2v_reg  <= \piso.data_li [1026];
      \piso.data_r_1025_sv2v_reg  <= \piso.data_li [1025];
      \piso.data_r_1024_sv2v_reg  <= \piso.data_li [1024];
      \piso.data_r_1023_sv2v_reg  <= \piso.data_li [1023];
      \piso.data_r_1022_sv2v_reg  <= \piso.data_li [1022];
      \piso.data_r_1021_sv2v_reg  <= \piso.data_li [1021];
      \piso.data_r_1020_sv2v_reg  <= \piso.data_li [1020];
      \piso.data_r_1019_sv2v_reg  <= \piso.data_li [1019];
      \piso.data_r_1018_sv2v_reg  <= \piso.data_li [1018];
      \piso.data_r_1017_sv2v_reg  <= \piso.data_li [1017];
      \piso.data_r_1016_sv2v_reg  <= \piso.data_li [1016];
      \piso.data_r_1015_sv2v_reg  <= \piso.data_li [1015];
      \piso.data_r_1014_sv2v_reg  <= \piso.data_li [1014];
      \piso.data_r_1013_sv2v_reg  <= \piso.data_li [1013];
      \piso.data_r_1012_sv2v_reg  <= \piso.data_li [1012];
      \piso.data_r_1011_sv2v_reg  <= \piso.data_li [1011];
      \piso.data_r_1010_sv2v_reg  <= \piso.data_li [1010];
      \piso.data_r_1009_sv2v_reg  <= \piso.data_li [1009];
      \piso.data_r_1008_sv2v_reg  <= \piso.data_li [1008];
      \piso.data_r_1007_sv2v_reg  <= \piso.data_li [1007];
      \piso.data_r_1006_sv2v_reg  <= \piso.data_li [1006];
      \piso.data_r_1005_sv2v_reg  <= \piso.data_li [1005];
      \piso.data_r_1004_sv2v_reg  <= \piso.data_li [1004];
      \piso.data_r_1003_sv2v_reg  <= \piso.data_li [1003];
      \piso.data_r_1002_sv2v_reg  <= \piso.data_li [1002];
      \piso.data_r_1001_sv2v_reg  <= \piso.data_li [1001];
      \piso.data_r_1000_sv2v_reg  <= \piso.data_li [1000];
      \piso.data_r_999_sv2v_reg  <= \piso.data_li [999];
      \piso.data_r_998_sv2v_reg  <= \piso.data_li [998];
      \piso.data_r_997_sv2v_reg  <= \piso.data_li [997];
      \piso.data_r_996_sv2v_reg  <= \piso.data_li [996];
      \piso.data_r_995_sv2v_reg  <= \piso.data_li [995];
      \piso.data_r_994_sv2v_reg  <= \piso.data_li [994];
      \piso.data_r_993_sv2v_reg  <= \piso.data_li [993];
      \piso.data_r_992_sv2v_reg  <= \piso.data_li [992];
      \piso.data_r_991_sv2v_reg  <= \piso.data_li [991];
      \piso.data_r_990_sv2v_reg  <= \piso.data_li [990];
      \piso.data_r_989_sv2v_reg  <= \piso.data_li [989];
      \piso.data_r_988_sv2v_reg  <= \piso.data_li [988];
      \piso.data_r_987_sv2v_reg  <= \piso.data_li [987];
      \piso.data_r_986_sv2v_reg  <= \piso.data_li [986];
      \piso.data_r_985_sv2v_reg  <= \piso.data_li [985];
      \piso.data_r_984_sv2v_reg  <= \piso.data_li [984];
      \piso.data_r_983_sv2v_reg  <= \piso.data_li [983];
      \piso.data_r_982_sv2v_reg  <= \piso.data_li [982];
      \piso.data_r_981_sv2v_reg  <= \piso.data_li [981];
      \piso.data_r_980_sv2v_reg  <= \piso.data_li [980];
      \piso.data_r_979_sv2v_reg  <= \piso.data_li [979];
      \piso.data_r_978_sv2v_reg  <= \piso.data_li [978];
      \piso.data_r_977_sv2v_reg  <= \piso.data_li [977];
      \piso.data_r_976_sv2v_reg  <= \piso.data_li [976];
      \piso.data_r_975_sv2v_reg  <= \piso.data_li [975];
      \piso.data_r_974_sv2v_reg  <= \piso.data_li [974];
      \piso.data_r_973_sv2v_reg  <= \piso.data_li [973];
      \piso.data_r_972_sv2v_reg  <= \piso.data_li [972];
      \piso.data_r_971_sv2v_reg  <= \piso.data_li [971];
      \piso.data_r_970_sv2v_reg  <= \piso.data_li [970];
      \piso.data_r_969_sv2v_reg  <= \piso.data_li [969];
      \piso.data_r_968_sv2v_reg  <= \piso.data_li [968];
      \piso.data_r_967_sv2v_reg  <= \piso.data_li [967];
      \piso.data_r_966_sv2v_reg  <= \piso.data_li [966];
      \piso.data_r_965_sv2v_reg  <= \piso.data_li [965];
      \piso.data_r_964_sv2v_reg  <= \piso.data_li [964];
      \piso.data_r_963_sv2v_reg  <= \piso.data_li [963];
      \piso.data_r_962_sv2v_reg  <= \piso.data_li [962];
      \piso.data_r_961_sv2v_reg  <= \piso.data_li [961];
      \piso.data_r_960_sv2v_reg  <= \piso.data_li [960];
      \piso.data_r_959_sv2v_reg  <= \piso.data_li [959];
      \piso.data_r_958_sv2v_reg  <= \piso.data_li [958];
      \piso.data_r_957_sv2v_reg  <= \piso.data_li [957];
      \piso.data_r_956_sv2v_reg  <= \piso.data_li [956];
      \piso.data_r_955_sv2v_reg  <= \piso.data_li [955];
      \piso.data_r_954_sv2v_reg  <= \piso.data_li [954];
      \piso.data_r_953_sv2v_reg  <= \piso.data_li [953];
      \piso.data_r_952_sv2v_reg  <= \piso.data_li [952];
      \piso.data_r_951_sv2v_reg  <= \piso.data_li [951];
      \piso.data_r_950_sv2v_reg  <= \piso.data_li [950];
      \piso.data_r_949_sv2v_reg  <= \piso.data_li [949];
      \piso.data_r_948_sv2v_reg  <= \piso.data_li [948];
      \piso.data_r_947_sv2v_reg  <= \piso.data_li [947];
      \piso.data_r_946_sv2v_reg  <= \piso.data_li [946];
      \piso.data_r_945_sv2v_reg  <= \piso.data_li [945];
      \piso.data_r_944_sv2v_reg  <= \piso.data_li [944];
      \piso.data_r_943_sv2v_reg  <= \piso.data_li [943];
      \piso.data_r_942_sv2v_reg  <= \piso.data_li [942];
      \piso.data_r_941_sv2v_reg  <= \piso.data_li [941];
      \piso.data_r_940_sv2v_reg  <= \piso.data_li [940];
      \piso.data_r_939_sv2v_reg  <= \piso.data_li [939];
      \piso.data_r_938_sv2v_reg  <= \piso.data_li [938];
      \piso.data_r_937_sv2v_reg  <= \piso.data_li [937];
      \piso.data_r_936_sv2v_reg  <= \piso.data_li [936];
      \piso.data_r_935_sv2v_reg  <= \piso.data_li [935];
      \piso.data_r_934_sv2v_reg  <= \piso.data_li [934];
      \piso.data_r_933_sv2v_reg  <= \piso.data_li [933];
      \piso.data_r_932_sv2v_reg  <= \piso.data_li [932];
      \piso.data_r_931_sv2v_reg  <= \piso.data_li [931];
      \piso.data_r_930_sv2v_reg  <= \piso.data_li [930];
      \piso.data_r_929_sv2v_reg  <= \piso.data_li [929];
      \piso.data_r_928_sv2v_reg  <= \piso.data_li [928];
      \piso.data_r_927_sv2v_reg  <= \piso.data_li [927];
      \piso.data_r_926_sv2v_reg  <= \piso.data_li [926];
      \piso.data_r_925_sv2v_reg  <= \piso.data_li [925];
      \piso.data_r_924_sv2v_reg  <= \piso.data_li [924];
      \piso.data_r_923_sv2v_reg  <= \piso.data_li [923];
      \piso.data_r_922_sv2v_reg  <= \piso.data_li [922];
      \piso.data_r_921_sv2v_reg  <= \piso.data_li [921];
      \piso.data_r_920_sv2v_reg  <= \piso.data_li [920];
      \piso.data_r_919_sv2v_reg  <= \piso.data_li [919];
      \piso.data_r_918_sv2v_reg  <= \piso.data_li [918];
      \piso.data_r_917_sv2v_reg  <= \piso.data_li [917];
      \piso.data_r_916_sv2v_reg  <= \piso.data_li [916];
      \piso.data_r_915_sv2v_reg  <= \piso.data_li [915];
      \piso.data_r_914_sv2v_reg  <= \piso.data_li [914];
      \piso.data_r_913_sv2v_reg  <= \piso.data_li [913];
      \piso.data_r_912_sv2v_reg  <= \piso.data_li [912];
      \piso.data_r_911_sv2v_reg  <= \piso.data_li [911];
      \piso.data_r_910_sv2v_reg  <= \piso.data_li [910];
      \piso.data_r_909_sv2v_reg  <= \piso.data_li [909];
      \piso.data_r_908_sv2v_reg  <= \piso.data_li [908];
      \piso.data_r_907_sv2v_reg  <= \piso.data_li [907];
      \piso.data_r_906_sv2v_reg  <= \piso.data_li [906];
      \piso.data_r_905_sv2v_reg  <= \piso.data_li [905];
      \piso.data_r_904_sv2v_reg  <= \piso.data_li [904];
      \piso.data_r_903_sv2v_reg  <= \piso.data_li [903];
      \piso.data_r_902_sv2v_reg  <= \piso.data_li [902];
      \piso.data_r_901_sv2v_reg  <= \piso.data_li [901];
      \piso.data_r_900_sv2v_reg  <= \piso.data_li [900];
      \piso.data_r_899_sv2v_reg  <= \piso.data_li [899];
      \piso.data_r_898_sv2v_reg  <= \piso.data_li [898];
      \piso.data_r_897_sv2v_reg  <= \piso.data_li [897];
      \piso.data_r_896_sv2v_reg  <= \piso.data_li [896];
      \piso.data_r_895_sv2v_reg  <= \piso.data_li [895];
      \piso.data_r_894_sv2v_reg  <= \piso.data_li [894];
      \piso.data_r_893_sv2v_reg  <= \piso.data_li [893];
      \piso.data_r_892_sv2v_reg  <= \piso.data_li [892];
      \piso.data_r_891_sv2v_reg  <= \piso.data_li [891];
      \piso.data_r_890_sv2v_reg  <= \piso.data_li [890];
      \piso.data_r_889_sv2v_reg  <= \piso.data_li [889];
      \piso.data_r_888_sv2v_reg  <= \piso.data_li [888];
      \piso.data_r_887_sv2v_reg  <= \piso.data_li [887];
      \piso.data_r_886_sv2v_reg  <= \piso.data_li [886];
      \piso.data_r_885_sv2v_reg  <= \piso.data_li [885];
      \piso.data_r_884_sv2v_reg  <= \piso.data_li [884];
      \piso.data_r_883_sv2v_reg  <= \piso.data_li [883];
      \piso.data_r_882_sv2v_reg  <= \piso.data_li [882];
      \piso.data_r_881_sv2v_reg  <= \piso.data_li [881];
      \piso.data_r_880_sv2v_reg  <= \piso.data_li [880];
      \piso.data_r_879_sv2v_reg  <= \piso.data_li [879];
      \piso.data_r_878_sv2v_reg  <= \piso.data_li [878];
      \piso.data_r_877_sv2v_reg  <= \piso.data_li [877];
      \piso.data_r_876_sv2v_reg  <= \piso.data_li [876];
      \piso.data_r_875_sv2v_reg  <= \piso.data_li [875];
      \piso.data_r_874_sv2v_reg  <= \piso.data_li [874];
      \piso.data_r_873_sv2v_reg  <= \piso.data_li [873];
      \piso.data_r_872_sv2v_reg  <= \piso.data_li [872];
      \piso.data_r_871_sv2v_reg  <= \piso.data_li [871];
      \piso.data_r_870_sv2v_reg  <= \piso.data_li [870];
      \piso.data_r_869_sv2v_reg  <= \piso.data_li [869];
      \piso.data_r_868_sv2v_reg  <= \piso.data_li [868];
      \piso.data_r_867_sv2v_reg  <= \piso.data_li [867];
      \piso.data_r_866_sv2v_reg  <= \piso.data_li [866];
      \piso.data_r_865_sv2v_reg  <= \piso.data_li [865];
      \piso.data_r_864_sv2v_reg  <= \piso.data_li [864];
      \piso.data_r_863_sv2v_reg  <= \piso.data_li [863];
      \piso.data_r_862_sv2v_reg  <= \piso.data_li [862];
      \piso.data_r_861_sv2v_reg  <= \piso.data_li [861];
      \piso.data_r_860_sv2v_reg  <= \piso.data_li [860];
      \piso.data_r_859_sv2v_reg  <= \piso.data_li [859];
      \piso.data_r_858_sv2v_reg  <= \piso.data_li [858];
      \piso.data_r_857_sv2v_reg  <= \piso.data_li [857];
      \piso.data_r_856_sv2v_reg  <= \piso.data_li [856];
      \piso.data_r_855_sv2v_reg  <= \piso.data_li [855];
      \piso.data_r_854_sv2v_reg  <= \piso.data_li [854];
      \piso.data_r_853_sv2v_reg  <= \piso.data_li [853];
      \piso.data_r_852_sv2v_reg  <= \piso.data_li [852];
      \piso.data_r_851_sv2v_reg  <= \piso.data_li [851];
      \piso.data_r_850_sv2v_reg  <= \piso.data_li [850];
      \piso.data_r_849_sv2v_reg  <= \piso.data_li [849];
      \piso.data_r_848_sv2v_reg  <= \piso.data_li [848];
      \piso.data_r_847_sv2v_reg  <= \piso.data_li [847];
      \piso.data_r_846_sv2v_reg  <= \piso.data_li [846];
      \piso.data_r_845_sv2v_reg  <= \piso.data_li [845];
      \piso.data_r_844_sv2v_reg  <= \piso.data_li [844];
      \piso.data_r_843_sv2v_reg  <= \piso.data_li [843];
      \piso.data_r_842_sv2v_reg  <= \piso.data_li [842];
      \piso.data_r_841_sv2v_reg  <= \piso.data_li [841];
      \piso.data_r_840_sv2v_reg  <= \piso.data_li [840];
      \piso.data_r_839_sv2v_reg  <= \piso.data_li [839];
      \piso.data_r_838_sv2v_reg  <= \piso.data_li [838];
      \piso.data_r_837_sv2v_reg  <= \piso.data_li [837];
      \piso.data_r_836_sv2v_reg  <= \piso.data_li [836];
      \piso.data_r_835_sv2v_reg  <= \piso.data_li [835];
      \piso.data_r_834_sv2v_reg  <= \piso.data_li [834];
      \piso.data_r_833_sv2v_reg  <= \piso.data_li [833];
      \piso.data_r_832_sv2v_reg  <= \piso.data_li [832];
      \piso.data_r_831_sv2v_reg  <= \piso.data_li [831];
      \piso.data_r_830_sv2v_reg  <= \piso.data_li [830];
      \piso.data_r_829_sv2v_reg  <= \piso.data_li [829];
      \piso.data_r_828_sv2v_reg  <= \piso.data_li [828];
      \piso.data_r_827_sv2v_reg  <= \piso.data_li [827];
      \piso.data_r_826_sv2v_reg  <= \piso.data_li [826];
      \piso.data_r_825_sv2v_reg  <= \piso.data_li [825];
      \piso.data_r_824_sv2v_reg  <= \piso.data_li [824];
      \piso.data_r_823_sv2v_reg  <= \piso.data_li [823];
      \piso.data_r_822_sv2v_reg  <= \piso.data_li [822];
      \piso.data_r_821_sv2v_reg  <= \piso.data_li [821];
      \piso.data_r_820_sv2v_reg  <= \piso.data_li [820];
      \piso.data_r_819_sv2v_reg  <= \piso.data_li [819];
      \piso.data_r_818_sv2v_reg  <= \piso.data_li [818];
      \piso.data_r_817_sv2v_reg  <= \piso.data_li [817];
      \piso.data_r_816_sv2v_reg  <= \piso.data_li [816];
      \piso.data_r_815_sv2v_reg  <= \piso.data_li [815];
      \piso.data_r_814_sv2v_reg  <= \piso.data_li [814];
      \piso.data_r_813_sv2v_reg  <= \piso.data_li [813];
      \piso.data_r_812_sv2v_reg  <= \piso.data_li [812];
      \piso.data_r_811_sv2v_reg  <= \piso.data_li [811];
      \piso.data_r_810_sv2v_reg  <= \piso.data_li [810];
      \piso.data_r_809_sv2v_reg  <= \piso.data_li [809];
      \piso.data_r_808_sv2v_reg  <= \piso.data_li [808];
      \piso.data_r_807_sv2v_reg  <= \piso.data_li [807];
      \piso.data_r_806_sv2v_reg  <= \piso.data_li [806];
      \piso.data_r_805_sv2v_reg  <= \piso.data_li [805];
      \piso.data_r_804_sv2v_reg  <= \piso.data_li [804];
      \piso.data_r_803_sv2v_reg  <= \piso.data_li [803];
      \piso.data_r_802_sv2v_reg  <= \piso.data_li [802];
      \piso.data_r_801_sv2v_reg  <= \piso.data_li [801];
      \piso.data_r_800_sv2v_reg  <= \piso.data_li [800];
      \piso.data_r_799_sv2v_reg  <= \piso.data_li [799];
      \piso.data_r_798_sv2v_reg  <= \piso.data_li [798];
      \piso.data_r_797_sv2v_reg  <= \piso.data_li [797];
      \piso.data_r_796_sv2v_reg  <= \piso.data_li [796];
      \piso.data_r_795_sv2v_reg  <= \piso.data_li [795];
      \piso.data_r_794_sv2v_reg  <= \piso.data_li [794];
      \piso.data_r_793_sv2v_reg  <= \piso.data_li [793];
      \piso.data_r_792_sv2v_reg  <= \piso.data_li [792];
      \piso.data_r_791_sv2v_reg  <= \piso.data_li [791];
      \piso.data_r_790_sv2v_reg  <= \piso.data_li [790];
      \piso.data_r_789_sv2v_reg  <= \piso.data_li [789];
      \piso.data_r_788_sv2v_reg  <= \piso.data_li [788];
      \piso.data_r_787_sv2v_reg  <= \piso.data_li [787];
      \piso.data_r_786_sv2v_reg  <= \piso.data_li [786];
      \piso.data_r_785_sv2v_reg  <= \piso.data_li [785];
      \piso.data_r_784_sv2v_reg  <= \piso.data_li [784];
      \piso.data_r_783_sv2v_reg  <= \piso.data_li [783];
      \piso.data_r_782_sv2v_reg  <= \piso.data_li [782];
      \piso.data_r_781_sv2v_reg  <= \piso.data_li [781];
      \piso.data_r_780_sv2v_reg  <= \piso.data_li [780];
      \piso.data_r_779_sv2v_reg  <= \piso.data_li [779];
      \piso.data_r_778_sv2v_reg  <= \piso.data_li [778];
      \piso.data_r_777_sv2v_reg  <= \piso.data_li [777];
      \piso.data_r_776_sv2v_reg  <= \piso.data_li [776];
      \piso.data_r_775_sv2v_reg  <= \piso.data_li [775];
      \piso.data_r_774_sv2v_reg  <= \piso.data_li [774];
      \piso.data_r_773_sv2v_reg  <= \piso.data_li [773];
      \piso.data_r_772_sv2v_reg  <= \piso.data_li [772];
      \piso.data_r_771_sv2v_reg  <= \piso.data_li [771];
      \piso.data_r_770_sv2v_reg  <= \piso.data_li [770];
      \piso.data_r_769_sv2v_reg  <= \piso.data_li [769];
      \piso.data_r_768_sv2v_reg  <= \piso.data_li [768];
      \piso.data_r_767_sv2v_reg  <= \piso.data_li [767];
      \piso.data_r_766_sv2v_reg  <= \piso.data_li [766];
      \piso.data_r_765_sv2v_reg  <= \piso.data_li [765];
      \piso.data_r_764_sv2v_reg  <= \piso.data_li [764];
      \piso.data_r_763_sv2v_reg  <= \piso.data_li [763];
      \piso.data_r_762_sv2v_reg  <= \piso.data_li [762];
      \piso.data_r_761_sv2v_reg  <= \piso.data_li [761];
      \piso.data_r_760_sv2v_reg  <= \piso.data_li [760];
      \piso.data_r_759_sv2v_reg  <= \piso.data_li [759];
      \piso.data_r_758_sv2v_reg  <= \piso.data_li [758];
      \piso.data_r_757_sv2v_reg  <= \piso.data_li [757];
      \piso.data_r_756_sv2v_reg  <= \piso.data_li [756];
      \piso.data_r_755_sv2v_reg  <= \piso.data_li [755];
      \piso.data_r_754_sv2v_reg  <= \piso.data_li [754];
      \piso.data_r_753_sv2v_reg  <= \piso.data_li [753];
      \piso.data_r_752_sv2v_reg  <= \piso.data_li [752];
      \piso.data_r_751_sv2v_reg  <= \piso.data_li [751];
      \piso.data_r_750_sv2v_reg  <= \piso.data_li [750];
      \piso.data_r_749_sv2v_reg  <= \piso.data_li [749];
      \piso.data_r_748_sv2v_reg  <= \piso.data_li [748];
      \piso.data_r_747_sv2v_reg  <= \piso.data_li [747];
      \piso.data_r_746_sv2v_reg  <= \piso.data_li [746];
      \piso.data_r_745_sv2v_reg  <= \piso.data_li [745];
      \piso.data_r_744_sv2v_reg  <= \piso.data_li [744];
      \piso.data_r_743_sv2v_reg  <= \piso.data_li [743];
      \piso.data_r_742_sv2v_reg  <= \piso.data_li [742];
      \piso.data_r_741_sv2v_reg  <= \piso.data_li [741];
      \piso.data_r_740_sv2v_reg  <= \piso.data_li [740];
      \piso.data_r_739_sv2v_reg  <= \piso.data_li [739];
      \piso.data_r_738_sv2v_reg  <= \piso.data_li [738];
      \piso.data_r_737_sv2v_reg  <= \piso.data_li [737];
      \piso.data_r_736_sv2v_reg  <= \piso.data_li [736];
      \piso.data_r_735_sv2v_reg  <= \piso.data_li [735];
      \piso.data_r_734_sv2v_reg  <= \piso.data_li [734];
      \piso.data_r_733_sv2v_reg  <= \piso.data_li [733];
      \piso.data_r_732_sv2v_reg  <= \piso.data_li [732];
      \piso.data_r_731_sv2v_reg  <= \piso.data_li [731];
      \piso.data_r_730_sv2v_reg  <= \piso.data_li [730];
      \piso.data_r_729_sv2v_reg  <= \piso.data_li [729];
      \piso.data_r_728_sv2v_reg  <= \piso.data_li [728];
      \piso.data_r_727_sv2v_reg  <= \piso.data_li [727];
      \piso.data_r_726_sv2v_reg  <= \piso.data_li [726];
      \piso.data_r_725_sv2v_reg  <= \piso.data_li [725];
      \piso.data_r_724_sv2v_reg  <= \piso.data_li [724];
      \piso.data_r_723_sv2v_reg  <= \piso.data_li [723];
      \piso.data_r_722_sv2v_reg  <= \piso.data_li [722];
      \piso.data_r_721_sv2v_reg  <= \piso.data_li [721];
      \piso.data_r_720_sv2v_reg  <= \piso.data_li [720];
      \piso.data_r_719_sv2v_reg  <= \piso.data_li [719];
      \piso.data_r_718_sv2v_reg  <= \piso.data_li [718];
      \piso.data_r_717_sv2v_reg  <= \piso.data_li [717];
      \piso.data_r_716_sv2v_reg  <= \piso.data_li [716];
      \piso.data_r_715_sv2v_reg  <= \piso.data_li [715];
      \piso.data_r_714_sv2v_reg  <= \piso.data_li [714];
      \piso.data_r_713_sv2v_reg  <= \piso.data_li [713];
      \piso.data_r_712_sv2v_reg  <= \piso.data_li [712];
      \piso.data_r_711_sv2v_reg  <= \piso.data_li [711];
      \piso.data_r_710_sv2v_reg  <= \piso.data_li [710];
      \piso.data_r_709_sv2v_reg  <= \piso.data_li [709];
      \piso.data_r_708_sv2v_reg  <= \piso.data_li [708];
      \piso.data_r_707_sv2v_reg  <= \piso.data_li [707];
      \piso.data_r_706_sv2v_reg  <= \piso.data_li [706];
      \piso.data_r_705_sv2v_reg  <= \piso.data_li [705];
      \piso.data_r_704_sv2v_reg  <= \piso.data_li [704];
      \piso.data_r_703_sv2v_reg  <= \piso.data_li [703];
      \piso.data_r_702_sv2v_reg  <= \piso.data_li [702];
      \piso.data_r_701_sv2v_reg  <= \piso.data_li [701];
      \piso.data_r_700_sv2v_reg  <= \piso.data_li [700];
      \piso.data_r_699_sv2v_reg  <= \piso.data_li [699];
      \piso.data_r_698_sv2v_reg  <= \piso.data_li [698];
      \piso.data_r_697_sv2v_reg  <= \piso.data_li [697];
      \piso.data_r_696_sv2v_reg  <= \piso.data_li [696];
      \piso.data_r_695_sv2v_reg  <= \piso.data_li [695];
      \piso.data_r_694_sv2v_reg  <= \piso.data_li [694];
      \piso.data_r_693_sv2v_reg  <= \piso.data_li [693];
      \piso.data_r_692_sv2v_reg  <= \piso.data_li [692];
      \piso.data_r_691_sv2v_reg  <= \piso.data_li [691];
      \piso.data_r_690_sv2v_reg  <= \piso.data_li [690];
      \piso.data_r_689_sv2v_reg  <= \piso.data_li [689];
      \piso.data_r_688_sv2v_reg  <= \piso.data_li [688];
      \piso.data_r_687_sv2v_reg  <= \piso.data_li [687];
      \piso.data_r_686_sv2v_reg  <= \piso.data_li [686];
      \piso.data_r_685_sv2v_reg  <= \piso.data_li [685];
      \piso.data_r_684_sv2v_reg  <= \piso.data_li [684];
      \piso.data_r_683_sv2v_reg  <= \piso.data_li [683];
      \piso.data_r_682_sv2v_reg  <= \piso.data_li [682];
      \piso.data_r_681_sv2v_reg  <= \piso.data_li [681];
      \piso.data_r_680_sv2v_reg  <= \piso.data_li [680];
      \piso.data_r_679_sv2v_reg  <= \piso.data_li [679];
      \piso.data_r_678_sv2v_reg  <= \piso.data_li [678];
      \piso.data_r_677_sv2v_reg  <= \piso.data_li [677];
      \piso.data_r_676_sv2v_reg  <= \piso.data_li [676];
      \piso.data_r_675_sv2v_reg  <= \piso.data_li [675];
      \piso.data_r_674_sv2v_reg  <= \piso.data_li [674];
      \piso.data_r_673_sv2v_reg  <= \piso.data_li [673];
      \piso.data_r_672_sv2v_reg  <= \piso.data_li [672];
      \piso.data_r_671_sv2v_reg  <= \piso.data_li [671];
      \piso.data_r_670_sv2v_reg  <= \piso.data_li [670];
      \piso.data_r_669_sv2v_reg  <= \piso.data_li [669];
      \piso.data_r_668_sv2v_reg  <= \piso.data_li [668];
      \piso.data_r_667_sv2v_reg  <= \piso.data_li [667];
      \piso.data_r_666_sv2v_reg  <= \piso.data_li [666];
      \piso.data_r_665_sv2v_reg  <= \piso.data_li [665];
      \piso.data_r_664_sv2v_reg  <= \piso.data_li [664];
      \piso.data_r_663_sv2v_reg  <= \piso.data_li [663];
      \piso.data_r_662_sv2v_reg  <= \piso.data_li [662];
      \piso.data_r_661_sv2v_reg  <= \piso.data_li [661];
      \piso.data_r_660_sv2v_reg  <= \piso.data_li [660];
      \piso.data_r_659_sv2v_reg  <= \piso.data_li [659];
      \piso.data_r_658_sv2v_reg  <= \piso.data_li [658];
      \piso.data_r_657_sv2v_reg  <= \piso.data_li [657];
      \piso.data_r_656_sv2v_reg  <= \piso.data_li [656];
      \piso.data_r_655_sv2v_reg  <= \piso.data_li [655];
      \piso.data_r_654_sv2v_reg  <= \piso.data_li [654];
      \piso.data_r_653_sv2v_reg  <= \piso.data_li [653];
      \piso.data_r_652_sv2v_reg  <= \piso.data_li [652];
      \piso.data_r_651_sv2v_reg  <= \piso.data_li [651];
      \piso.data_r_650_sv2v_reg  <= \piso.data_li [650];
      \piso.data_r_649_sv2v_reg  <= \piso.data_li [649];
      \piso.data_r_648_sv2v_reg  <= \piso.data_li [648];
      \piso.data_r_647_sv2v_reg  <= \piso.data_li [647];
      \piso.data_r_646_sv2v_reg  <= \piso.data_li [646];
      \piso.data_r_645_sv2v_reg  <= \piso.data_li [645];
      \piso.data_r_644_sv2v_reg  <= \piso.data_li [644];
      \piso.data_r_643_sv2v_reg  <= \piso.data_li [643];
      \piso.data_r_642_sv2v_reg  <= \piso.data_li [642];
      \piso.data_r_641_sv2v_reg  <= \piso.data_li [641];
      \piso.data_r_640_sv2v_reg  <= \piso.data_li [640];
      \piso.data_r_639_sv2v_reg  <= \piso.data_li [639];
      \piso.data_r_638_sv2v_reg  <= \piso.data_li [638];
      \piso.data_r_637_sv2v_reg  <= \piso.data_li [637];
      \piso.data_r_636_sv2v_reg  <= \piso.data_li [636];
      \piso.data_r_635_sv2v_reg  <= \piso.data_li [635];
      \piso.data_r_634_sv2v_reg  <= \piso.data_li [634];
      \piso.data_r_633_sv2v_reg  <= \piso.data_li [633];
      \piso.data_r_632_sv2v_reg  <= \piso.data_li [632];
      \piso.data_r_631_sv2v_reg  <= \piso.data_li [631];
      \piso.data_r_630_sv2v_reg  <= \piso.data_li [630];
      \piso.data_r_629_sv2v_reg  <= \piso.data_li [629];
      \piso.data_r_628_sv2v_reg  <= \piso.data_li [628];
      \piso.data_r_627_sv2v_reg  <= \piso.data_li [627];
      \piso.data_r_626_sv2v_reg  <= \piso.data_li [626];
      \piso.data_r_625_sv2v_reg  <= \piso.data_li [625];
      \piso.data_r_624_sv2v_reg  <= \piso.data_li [624];
      \piso.data_r_623_sv2v_reg  <= \piso.data_li [623];
      \piso.data_r_622_sv2v_reg  <= \piso.data_li [622];
      \piso.data_r_621_sv2v_reg  <= \piso.data_li [621];
      \piso.data_r_620_sv2v_reg  <= \piso.data_li [620];
      \piso.data_r_619_sv2v_reg  <= \piso.data_li [619];
      \piso.data_r_618_sv2v_reg  <= \piso.data_li [618];
      \piso.data_r_617_sv2v_reg  <= \piso.data_li [617];
      \piso.data_r_616_sv2v_reg  <= \piso.data_li [616];
      \piso.data_r_615_sv2v_reg  <= \piso.data_li [615];
      \piso.data_r_614_sv2v_reg  <= \piso.data_li [614];
      \piso.data_r_613_sv2v_reg  <= \piso.data_li [613];
      \piso.data_r_612_sv2v_reg  <= \piso.data_li [612];
      \piso.data_r_611_sv2v_reg  <= \piso.data_li [611];
      \piso.data_r_610_sv2v_reg  <= \piso.data_li [610];
      \piso.data_r_609_sv2v_reg  <= \piso.data_li [609];
      \piso.data_r_608_sv2v_reg  <= \piso.data_li [608];
      \piso.data_r_607_sv2v_reg  <= \piso.data_li [607];
      \piso.data_r_606_sv2v_reg  <= \piso.data_li [606];
      \piso.data_r_605_sv2v_reg  <= \piso.data_li [605];
      \piso.data_r_604_sv2v_reg  <= \piso.data_li [604];
      \piso.data_r_603_sv2v_reg  <= \piso.data_li [603];
      \piso.data_r_602_sv2v_reg  <= \piso.data_li [602];
      \piso.data_r_601_sv2v_reg  <= \piso.data_li [601];
      \piso.data_r_600_sv2v_reg  <= \piso.data_li [600];
      \piso.data_r_599_sv2v_reg  <= \piso.data_li [599];
      \piso.data_r_598_sv2v_reg  <= \piso.data_li [598];
      \piso.data_r_597_sv2v_reg  <= \piso.data_li [597];
      \piso.data_r_596_sv2v_reg  <= \piso.data_li [596];
      \piso.data_r_595_sv2v_reg  <= \piso.data_li [595];
      \piso.data_r_594_sv2v_reg  <= \piso.data_li [594];
      \piso.data_r_593_sv2v_reg  <= \piso.data_li [593];
      \piso.data_r_592_sv2v_reg  <= \piso.data_li [592];
      \piso.data_r_591_sv2v_reg  <= \piso.data_li [591];
      \piso.data_r_590_sv2v_reg  <= \piso.data_li [590];
      \piso.data_r_589_sv2v_reg  <= \piso.data_li [589];
      \piso.data_r_588_sv2v_reg  <= \piso.data_li [588];
      \piso.data_r_587_sv2v_reg  <= \piso.data_li [587];
      \piso.data_r_586_sv2v_reg  <= \piso.data_li [586];
      \piso.data_r_585_sv2v_reg  <= \piso.data_li [585];
      \piso.data_r_584_sv2v_reg  <= \piso.data_li [584];
      \piso.data_r_583_sv2v_reg  <= \piso.data_li [583];
      \piso.data_r_582_sv2v_reg  <= \piso.data_li [582];
      \piso.data_r_581_sv2v_reg  <= \piso.data_li [581];
      \piso.data_r_580_sv2v_reg  <= \piso.data_li [580];
      \piso.data_r_579_sv2v_reg  <= \piso.data_li [579];
      \piso.data_r_578_sv2v_reg  <= \piso.data_li [578];
      \piso.data_r_577_sv2v_reg  <= \piso.data_li [577];
      \piso.data_r_576_sv2v_reg  <= \piso.data_li [576];
      \piso.data_r_575_sv2v_reg  <= \piso.data_li [575];
      \piso.data_r_574_sv2v_reg  <= \piso.data_li [574];
      \piso.data_r_573_sv2v_reg  <= \piso.data_li [573];
      \piso.data_r_572_sv2v_reg  <= \piso.data_li [572];
      \piso.data_r_571_sv2v_reg  <= \piso.data_li [571];
      \piso.data_r_570_sv2v_reg  <= \piso.data_li [570];
      \piso.data_r_569_sv2v_reg  <= \piso.data_li [569];
      \piso.data_r_568_sv2v_reg  <= \piso.data_li [568];
      \piso.data_r_567_sv2v_reg  <= \piso.data_li [567];
      \piso.data_r_566_sv2v_reg  <= \piso.data_li [566];
      \piso.data_r_565_sv2v_reg  <= \piso.data_li [565];
      \piso.data_r_564_sv2v_reg  <= \piso.data_li [564];
      \piso.data_r_563_sv2v_reg  <= \piso.data_li [563];
      \piso.data_r_562_sv2v_reg  <= \piso.data_li [562];
      \piso.data_r_561_sv2v_reg  <= \piso.data_li [561];
      \piso.data_r_560_sv2v_reg  <= \piso.data_li [560];
      \piso.data_r_559_sv2v_reg  <= \piso.data_li [559];
      \piso.data_r_558_sv2v_reg  <= \piso.data_li [558];
      \piso.data_r_557_sv2v_reg  <= \piso.data_li [557];
      \piso.data_r_556_sv2v_reg  <= \piso.data_li [556];
      \piso.data_r_555_sv2v_reg  <= \piso.data_li [555];
      \piso.data_r_554_sv2v_reg  <= \piso.data_li [554];
      \piso.data_r_553_sv2v_reg  <= \piso.data_li [553];
      \piso.data_r_552_sv2v_reg  <= \piso.data_li [552];
      \piso.data_r_551_sv2v_reg  <= \piso.data_li [551];
      \piso.data_r_550_sv2v_reg  <= \piso.data_li [550];
      \piso.data_r_549_sv2v_reg  <= \piso.data_li [549];
      \piso.data_r_548_sv2v_reg  <= \piso.data_li [548];
      \piso.data_r_547_sv2v_reg  <= \piso.data_li [547];
      \piso.data_r_546_sv2v_reg  <= \piso.data_li [546];
      \piso.data_r_545_sv2v_reg  <= \piso.data_li [545];
      \piso.data_r_544_sv2v_reg  <= \piso.data_li [544];
      \piso.data_r_543_sv2v_reg  <= \piso.data_li [543];
      \piso.data_r_542_sv2v_reg  <= \piso.data_li [542];
      \piso.data_r_541_sv2v_reg  <= \piso.data_li [541];
      \piso.data_r_540_sv2v_reg  <= \piso.data_li [540];
      \piso.data_r_539_sv2v_reg  <= \piso.data_li [539];
      \piso.data_r_538_sv2v_reg  <= \piso.data_li [538];
      \piso.data_r_537_sv2v_reg  <= \piso.data_li [537];
      \piso.data_r_536_sv2v_reg  <= \piso.data_li [536];
      \piso.data_r_535_sv2v_reg  <= \piso.data_li [535];
      \piso.data_r_534_sv2v_reg  <= \piso.data_li [534];
      \piso.data_r_533_sv2v_reg  <= \piso.data_li [533];
      \piso.data_r_532_sv2v_reg  <= \piso.data_li [532];
      \piso.data_r_531_sv2v_reg  <= \piso.data_li [531];
      \piso.data_r_530_sv2v_reg  <= \piso.data_li [530];
      \piso.data_r_529_sv2v_reg  <= \piso.data_li [529];
      \piso.data_r_528_sv2v_reg  <= \piso.data_li [528];
      \piso.data_r_527_sv2v_reg  <= \piso.data_li [527];
      \piso.data_r_526_sv2v_reg  <= \piso.data_li [526];
      \piso.data_r_525_sv2v_reg  <= \piso.data_li [525];
      \piso.data_r_524_sv2v_reg  <= \piso.data_li [524];
      \piso.data_r_523_sv2v_reg  <= \piso.data_li [523];
      \piso.data_r_522_sv2v_reg  <= \piso.data_li [522];
      \piso.data_r_521_sv2v_reg  <= \piso.data_li [521];
      \piso.data_r_520_sv2v_reg  <= \piso.data_li [520];
      \piso.data_r_519_sv2v_reg  <= \piso.data_li [519];
      \piso.data_r_518_sv2v_reg  <= \piso.data_li [518];
      \piso.data_r_517_sv2v_reg  <= \piso.data_li [517];
      \piso.data_r_516_sv2v_reg  <= \piso.data_li [516];
      \piso.data_r_515_sv2v_reg  <= \piso.data_li [515];
      \piso.data_r_514_sv2v_reg  <= \piso.data_li [514];
      \piso.data_r_513_sv2v_reg  <= \piso.data_li [513];
      \piso.data_r_512_sv2v_reg  <= \piso.data_li [512];
      \piso.data_r_511_sv2v_reg  <= \piso.data_li [511];
      \piso.data_r_510_sv2v_reg  <= \piso.data_li [510];
      \piso.data_r_509_sv2v_reg  <= \piso.data_li [509];
      \piso.data_r_508_sv2v_reg  <= \piso.data_li [508];
      \piso.data_r_507_sv2v_reg  <= \piso.data_li [507];
      \piso.data_r_506_sv2v_reg  <= \piso.data_li [506];
      \piso.data_r_505_sv2v_reg  <= \piso.data_li [505];
      \piso.data_r_504_sv2v_reg  <= \piso.data_li [504];
      \piso.data_r_503_sv2v_reg  <= \piso.data_li [503];
      \piso.data_r_502_sv2v_reg  <= \piso.data_li [502];
      \piso.data_r_501_sv2v_reg  <= \piso.data_li [501];
      \piso.data_r_500_sv2v_reg  <= \piso.data_li [500];
      \piso.data_r_499_sv2v_reg  <= \piso.data_li [499];
      \piso.data_r_498_sv2v_reg  <= \piso.data_li [498];
      \piso.data_r_497_sv2v_reg  <= \piso.data_li [497];
      \piso.data_r_496_sv2v_reg  <= \piso.data_li [496];
      \piso.data_r_495_sv2v_reg  <= \piso.data_li [495];
      \piso.data_r_494_sv2v_reg  <= \piso.data_li [494];
      \piso.data_r_493_sv2v_reg  <= \piso.data_li [493];
      \piso.data_r_492_sv2v_reg  <= \piso.data_li [492];
      \piso.data_r_491_sv2v_reg  <= \piso.data_li [491];
      \piso.data_r_490_sv2v_reg  <= \piso.data_li [490];
      \piso.data_r_489_sv2v_reg  <= \piso.data_li [489];
      \piso.data_r_488_sv2v_reg  <= \piso.data_li [488];
      \piso.data_r_487_sv2v_reg  <= \piso.data_li [487];
      \piso.data_r_486_sv2v_reg  <= \piso.data_li [486];
      \piso.data_r_485_sv2v_reg  <= \piso.data_li [485];
      \piso.data_r_484_sv2v_reg  <= \piso.data_li [484];
      \piso.data_r_483_sv2v_reg  <= \piso.data_li [483];
      \piso.data_r_482_sv2v_reg  <= \piso.data_li [482];
      \piso.data_r_481_sv2v_reg  <= \piso.data_li [481];
      \piso.data_r_480_sv2v_reg  <= \piso.data_li [480];
      \piso.data_r_479_sv2v_reg  <= \piso.data_li [479];
      \piso.data_r_478_sv2v_reg  <= \piso.data_li [478];
      \piso.data_r_477_sv2v_reg  <= \piso.data_li [477];
      \piso.data_r_476_sv2v_reg  <= \piso.data_li [476];
      \piso.data_r_475_sv2v_reg  <= \piso.data_li [475];
      \piso.data_r_474_sv2v_reg  <= \piso.data_li [474];
      \piso.data_r_473_sv2v_reg  <= \piso.data_li [473];
      \piso.data_r_472_sv2v_reg  <= \piso.data_li [472];
      \piso.data_r_471_sv2v_reg  <= \piso.data_li [471];
      \piso.data_r_470_sv2v_reg  <= \piso.data_li [470];
      \piso.data_r_469_sv2v_reg  <= \piso.data_li [469];
      \piso.data_r_468_sv2v_reg  <= \piso.data_li [468];
      \piso.data_r_467_sv2v_reg  <= \piso.data_li [467];
      \piso.data_r_466_sv2v_reg  <= \piso.data_li [466];
      \piso.data_r_465_sv2v_reg  <= \piso.data_li [465];
      \piso.data_r_464_sv2v_reg  <= \piso.data_li [464];
      \piso.data_r_463_sv2v_reg  <= \piso.data_li [463];
      \piso.data_r_462_sv2v_reg  <= \piso.data_li [462];
      \piso.data_r_461_sv2v_reg  <= \piso.data_li [461];
      \piso.data_r_460_sv2v_reg  <= \piso.data_li [460];
      \piso.data_r_459_sv2v_reg  <= \piso.data_li [459];
      \piso.data_r_458_sv2v_reg  <= \piso.data_li [458];
      \piso.data_r_457_sv2v_reg  <= \piso.data_li [457];
      \piso.data_r_456_sv2v_reg  <= \piso.data_li [456];
      \piso.data_r_455_sv2v_reg  <= \piso.data_li [455];
      \piso.data_r_454_sv2v_reg  <= \piso.data_li [454];
      \piso.data_r_453_sv2v_reg  <= \piso.data_li [453];
      \piso.data_r_452_sv2v_reg  <= \piso.data_li [452];
      \piso.data_r_451_sv2v_reg  <= \piso.data_li [451];
      \piso.data_r_450_sv2v_reg  <= \piso.data_li [450];
      \piso.data_r_449_sv2v_reg  <= \piso.data_li [449];
      \piso.data_r_448_sv2v_reg  <= \piso.data_li [448];
      \piso.data_r_447_sv2v_reg  <= \piso.data_li [447];
      \piso.data_r_446_sv2v_reg  <= \piso.data_li [446];
      \piso.data_r_445_sv2v_reg  <= \piso.data_li [445];
      \piso.data_r_444_sv2v_reg  <= \piso.data_li [444];
      \piso.data_r_443_sv2v_reg  <= \piso.data_li [443];
      \piso.data_r_442_sv2v_reg  <= \piso.data_li [442];
      \piso.data_r_441_sv2v_reg  <= \piso.data_li [441];
      \piso.data_r_440_sv2v_reg  <= \piso.data_li [440];
      \piso.data_r_439_sv2v_reg  <= \piso.data_li [439];
      \piso.data_r_438_sv2v_reg  <= \piso.data_li [438];
      \piso.data_r_437_sv2v_reg  <= \piso.data_li [437];
      \piso.data_r_436_sv2v_reg  <= \piso.data_li [436];
      \piso.data_r_435_sv2v_reg  <= \piso.data_li [435];
      \piso.data_r_434_sv2v_reg  <= \piso.data_li [434];
      \piso.data_r_433_sv2v_reg  <= \piso.data_li [433];
      \piso.data_r_432_sv2v_reg  <= \piso.data_li [432];
      \piso.data_r_431_sv2v_reg  <= \piso.data_li [431];
      \piso.data_r_430_sv2v_reg  <= \piso.data_li [430];
      \piso.data_r_429_sv2v_reg  <= \piso.data_li [429];
      \piso.data_r_428_sv2v_reg  <= \piso.data_li [428];
      \piso.data_r_427_sv2v_reg  <= \piso.data_li [427];
      \piso.data_r_426_sv2v_reg  <= \piso.data_li [426];
      \piso.data_r_425_sv2v_reg  <= \piso.data_li [425];
      \piso.data_r_424_sv2v_reg  <= \piso.data_li [424];
      \piso.data_r_423_sv2v_reg  <= \piso.data_li [423];
      \piso.data_r_422_sv2v_reg  <= \piso.data_li [422];
      \piso.data_r_421_sv2v_reg  <= \piso.data_li [421];
      \piso.data_r_420_sv2v_reg  <= \piso.data_li [420];
      \piso.data_r_419_sv2v_reg  <= \piso.data_li [419];
      \piso.data_r_418_sv2v_reg  <= \piso.data_li [418];
      \piso.data_r_417_sv2v_reg  <= \piso.data_li [417];
      \piso.data_r_416_sv2v_reg  <= \piso.data_li [416];
      \piso.data_r_415_sv2v_reg  <= \piso.data_li [415];
      \piso.data_r_414_sv2v_reg  <= \piso.data_li [414];
      \piso.data_r_413_sv2v_reg  <= \piso.data_li [413];
      \piso.data_r_412_sv2v_reg  <= \piso.data_li [412];
      \piso.data_r_411_sv2v_reg  <= \piso.data_li [411];
      \piso.data_r_410_sv2v_reg  <= \piso.data_li [410];
      \piso.data_r_409_sv2v_reg  <= \piso.data_li [409];
      \piso.data_r_408_sv2v_reg  <= \piso.data_li [408];
      \piso.data_r_407_sv2v_reg  <= \piso.data_li [407];
      \piso.data_r_406_sv2v_reg  <= \piso.data_li [406];
      \piso.data_r_405_sv2v_reg  <= \piso.data_li [405];
      \piso.data_r_404_sv2v_reg  <= \piso.data_li [404];
      \piso.data_r_403_sv2v_reg  <= \piso.data_li [403];
      \piso.data_r_402_sv2v_reg  <= \piso.data_li [402];
      \piso.data_r_401_sv2v_reg  <= \piso.data_li [401];
      \piso.data_r_400_sv2v_reg  <= \piso.data_li [400];
      \piso.data_r_399_sv2v_reg  <= \piso.data_li [399];
      \piso.data_r_398_sv2v_reg  <= \piso.data_li [398];
      \piso.data_r_397_sv2v_reg  <= \piso.data_li [397];
      \piso.data_r_396_sv2v_reg  <= \piso.data_li [396];
      \piso.data_r_395_sv2v_reg  <= \piso.data_li [395];
      \piso.data_r_394_sv2v_reg  <= \piso.data_li [394];
      \piso.data_r_393_sv2v_reg  <= \piso.data_li [393];
      \piso.data_r_392_sv2v_reg  <= \piso.data_li [392];
      \piso.data_r_391_sv2v_reg  <= \piso.data_li [391];
      \piso.data_r_390_sv2v_reg  <= \piso.data_li [390];
      \piso.data_r_389_sv2v_reg  <= \piso.data_li [389];
      \piso.data_r_388_sv2v_reg  <= \piso.data_li [388];
      \piso.data_r_387_sv2v_reg  <= \piso.data_li [387];
      \piso.data_r_386_sv2v_reg  <= \piso.data_li [386];
      \piso.data_r_385_sv2v_reg  <= \piso.data_li [385];
      \piso.data_r_384_sv2v_reg  <= \piso.data_li [384];
      \piso.data_r_383_sv2v_reg  <= \piso.data_li [383];
      \piso.data_r_382_sv2v_reg  <= \piso.data_li [382];
      \piso.data_r_381_sv2v_reg  <= \piso.data_li [381];
      \piso.data_r_380_sv2v_reg  <= \piso.data_li [380];
      \piso.data_r_379_sv2v_reg  <= \piso.data_li [379];
      \piso.data_r_378_sv2v_reg  <= \piso.data_li [378];
      \piso.data_r_377_sv2v_reg  <= \piso.data_li [377];
      \piso.data_r_376_sv2v_reg  <= \piso.data_li [376];
      \piso.data_r_375_sv2v_reg  <= \piso.data_li [375];
      \piso.data_r_374_sv2v_reg  <= \piso.data_li [374];
      \piso.data_r_373_sv2v_reg  <= \piso.data_li [373];
      \piso.data_r_372_sv2v_reg  <= \piso.data_li [372];
      \piso.data_r_371_sv2v_reg  <= \piso.data_li [371];
      \piso.data_r_370_sv2v_reg  <= \piso.data_li [370];
      \piso.data_r_369_sv2v_reg  <= \piso.data_li [369];
      \piso.data_r_368_sv2v_reg  <= \piso.data_li [368];
      \piso.data_r_367_sv2v_reg  <= \piso.data_li [367];
      \piso.data_r_366_sv2v_reg  <= \piso.data_li [366];
      \piso.data_r_365_sv2v_reg  <= \piso.data_li [365];
      \piso.data_r_364_sv2v_reg  <= \piso.data_li [364];
      \piso.data_r_363_sv2v_reg  <= \piso.data_li [363];
      \piso.data_r_362_sv2v_reg  <= \piso.data_li [362];
      \piso.data_r_361_sv2v_reg  <= \piso.data_li [361];
      \piso.data_r_360_sv2v_reg  <= \piso.data_li [360];
      \piso.data_r_359_sv2v_reg  <= \piso.data_li [359];
      \piso.data_r_358_sv2v_reg  <= \piso.data_li [358];
      \piso.data_r_357_sv2v_reg  <= \piso.data_li [357];
      \piso.data_r_356_sv2v_reg  <= \piso.data_li [356];
      \piso.data_r_355_sv2v_reg  <= \piso.data_li [355];
      \piso.data_r_354_sv2v_reg  <= \piso.data_li [354];
      \piso.data_r_353_sv2v_reg  <= \piso.data_li [353];
      \piso.data_r_352_sv2v_reg  <= \piso.data_li [352];
      \piso.data_r_351_sv2v_reg  <= \piso.data_li [351];
      \piso.data_r_350_sv2v_reg  <= \piso.data_li [350];
      \piso.data_r_349_sv2v_reg  <= \piso.data_li [349];
      \piso.data_r_348_sv2v_reg  <= \piso.data_li [348];
      \piso.data_r_347_sv2v_reg  <= \piso.data_li [347];
      \piso.data_r_346_sv2v_reg  <= \piso.data_li [346];
      \piso.data_r_345_sv2v_reg  <= \piso.data_li [345];
      \piso.data_r_344_sv2v_reg  <= \piso.data_li [344];
      \piso.data_r_343_sv2v_reg  <= \piso.data_li [343];
      \piso.data_r_342_sv2v_reg  <= \piso.data_li [342];
      \piso.data_r_341_sv2v_reg  <= \piso.data_li [341];
      \piso.data_r_340_sv2v_reg  <= \piso.data_li [340];
      \piso.data_r_339_sv2v_reg  <= \piso.data_li [339];
      \piso.data_r_338_sv2v_reg  <= \piso.data_li [338];
      \piso.data_r_337_sv2v_reg  <= \piso.data_li [337];
      \piso.data_r_336_sv2v_reg  <= \piso.data_li [336];
      \piso.data_r_335_sv2v_reg  <= \piso.data_li [335];
      \piso.data_r_334_sv2v_reg  <= \piso.data_li [334];
      \piso.data_r_333_sv2v_reg  <= \piso.data_li [333];
      \piso.data_r_332_sv2v_reg  <= \piso.data_li [332];
      \piso.data_r_331_sv2v_reg  <= \piso.data_li [331];
      \piso.data_r_330_sv2v_reg  <= \piso.data_li [330];
      \piso.data_r_329_sv2v_reg  <= \piso.data_li [329];
      \piso.data_r_328_sv2v_reg  <= \piso.data_li [328];
      \piso.data_r_327_sv2v_reg  <= \piso.data_li [327];
      \piso.data_r_326_sv2v_reg  <= \piso.data_li [326];
      \piso.data_r_325_sv2v_reg  <= \piso.data_li [325];
      \piso.data_r_324_sv2v_reg  <= \piso.data_li [324];
      \piso.data_r_323_sv2v_reg  <= \piso.data_li [323];
      \piso.data_r_322_sv2v_reg  <= \piso.data_li [322];
      \piso.data_r_321_sv2v_reg  <= \piso.data_li [321];
      \piso.data_r_320_sv2v_reg  <= \piso.data_li [320];
      \piso.data_r_319_sv2v_reg  <= \piso.data_li [319];
      \piso.data_r_318_sv2v_reg  <= \piso.data_li [318];
      \piso.data_r_317_sv2v_reg  <= \piso.data_li [317];
      \piso.data_r_316_sv2v_reg  <= \piso.data_li [316];
      \piso.data_r_315_sv2v_reg  <= \piso.data_li [315];
      \piso.data_r_314_sv2v_reg  <= \piso.data_li [314];
      \piso.data_r_313_sv2v_reg  <= \piso.data_li [313];
      \piso.data_r_312_sv2v_reg  <= \piso.data_li [312];
      \piso.data_r_311_sv2v_reg  <= \piso.data_li [311];
      \piso.data_r_310_sv2v_reg  <= \piso.data_li [310];
      \piso.data_r_309_sv2v_reg  <= \piso.data_li [309];
      \piso.data_r_308_sv2v_reg  <= \piso.data_li [308];
      \piso.data_r_307_sv2v_reg  <= \piso.data_li [307];
      \piso.data_r_306_sv2v_reg  <= \piso.data_li [306];
      \piso.data_r_305_sv2v_reg  <= \piso.data_li [305];
      \piso.data_r_304_sv2v_reg  <= \piso.data_li [304];
      \piso.data_r_303_sv2v_reg  <= \piso.data_li [303];
      \piso.data_r_302_sv2v_reg  <= \piso.data_li [302];
      \piso.data_r_301_sv2v_reg  <= \piso.data_li [301];
      \piso.data_r_300_sv2v_reg  <= \piso.data_li [300];
      \piso.data_r_299_sv2v_reg  <= \piso.data_li [299];
      \piso.data_r_298_sv2v_reg  <= \piso.data_li [298];
      \piso.data_r_297_sv2v_reg  <= \piso.data_li [297];
      \piso.data_r_296_sv2v_reg  <= \piso.data_li [296];
      \piso.data_r_295_sv2v_reg  <= \piso.data_li [295];
      \piso.data_r_294_sv2v_reg  <= \piso.data_li [294];
      \piso.data_r_293_sv2v_reg  <= \piso.data_li [293];
      \piso.data_r_292_sv2v_reg  <= \piso.data_li [292];
      \piso.data_r_291_sv2v_reg  <= \piso.data_li [291];
      \piso.data_r_290_sv2v_reg  <= \piso.data_li [290];
      \piso.data_r_289_sv2v_reg  <= \piso.data_li [289];
      \piso.data_r_288_sv2v_reg  <= \piso.data_li [288];
      \piso.data_r_287_sv2v_reg  <= \piso.data_li [287];
      \piso.data_r_286_sv2v_reg  <= \piso.data_li [286];
      \piso.data_r_285_sv2v_reg  <= \piso.data_li [285];
      \piso.data_r_284_sv2v_reg  <= \piso.data_li [284];
      \piso.data_r_283_sv2v_reg  <= \piso.data_li [283];
      \piso.data_r_282_sv2v_reg  <= \piso.data_li [282];
      \piso.data_r_281_sv2v_reg  <= \piso.data_li [281];
      \piso.data_r_280_sv2v_reg  <= \piso.data_li [280];
      \piso.data_r_279_sv2v_reg  <= \piso.data_li [279];
      \piso.data_r_278_sv2v_reg  <= \piso.data_li [278];
      \piso.data_r_277_sv2v_reg  <= \piso.data_li [277];
      \piso.data_r_276_sv2v_reg  <= \piso.data_li [276];
      \piso.data_r_275_sv2v_reg  <= \piso.data_li [275];
      \piso.data_r_274_sv2v_reg  <= \piso.data_li [274];
      \piso.data_r_273_sv2v_reg  <= \piso.data_li [273];
      \piso.data_r_272_sv2v_reg  <= \piso.data_li [272];
      \piso.data_r_271_sv2v_reg  <= \piso.data_li [271];
      \piso.data_r_270_sv2v_reg  <= \piso.data_li [270];
      \piso.data_r_269_sv2v_reg  <= \piso.data_li [269];
      \piso.data_r_268_sv2v_reg  <= \piso.data_li [268];
      \piso.data_r_267_sv2v_reg  <= \piso.data_li [267];
      \piso.data_r_266_sv2v_reg  <= \piso.data_li [266];
      \piso.data_r_265_sv2v_reg  <= \piso.data_li [265];
      \piso.data_r_264_sv2v_reg  <= \piso.data_li [264];
      \piso.data_r_263_sv2v_reg  <= \piso.data_li [263];
      \piso.data_r_262_sv2v_reg  <= \piso.data_li [262];
      \piso.data_r_261_sv2v_reg  <= \piso.data_li [261];
      \piso.data_r_260_sv2v_reg  <= \piso.data_li [260];
      \piso.data_r_259_sv2v_reg  <= \piso.data_li [259];
      \piso.data_r_258_sv2v_reg  <= \piso.data_li [258];
      \piso.data_r_257_sv2v_reg  <= \piso.data_li [257];
      \piso.data_r_256_sv2v_reg  <= \piso.data_li [256];
      \piso.data_r_255_sv2v_reg  <= \piso.data_li [255];
      \piso.data_r_254_sv2v_reg  <= \piso.data_li [254];
      \piso.data_r_253_sv2v_reg  <= \piso.data_li [253];
      \piso.data_r_252_sv2v_reg  <= \piso.data_li [252];
      \piso.data_r_251_sv2v_reg  <= \piso.data_li [251];
      \piso.data_r_250_sv2v_reg  <= \piso.data_li [250];
      \piso.data_r_249_sv2v_reg  <= \piso.data_li [249];
      \piso.data_r_248_sv2v_reg  <= \piso.data_li [248];
      \piso.data_r_247_sv2v_reg  <= \piso.data_li [247];
      \piso.data_r_246_sv2v_reg  <= \piso.data_li [246];
      \piso.data_r_245_sv2v_reg  <= \piso.data_li [245];
      \piso.data_r_244_sv2v_reg  <= \piso.data_li [244];
      \piso.data_r_243_sv2v_reg  <= \piso.data_li [243];
      \piso.data_r_242_sv2v_reg  <= \piso.data_li [242];
      \piso.data_r_241_sv2v_reg  <= \piso.data_li [241];
      \piso.data_r_240_sv2v_reg  <= \piso.data_li [240];
      \piso.data_r_239_sv2v_reg  <= \piso.data_li [239];
      \piso.data_r_238_sv2v_reg  <= \piso.data_li [238];
      \piso.data_r_237_sv2v_reg  <= \piso.data_li [237];
      \piso.data_r_236_sv2v_reg  <= \piso.data_li [236];
      \piso.data_r_235_sv2v_reg  <= \piso.data_li [235];
      \piso.data_r_234_sv2v_reg  <= \piso.data_li [234];
      \piso.data_r_233_sv2v_reg  <= \piso.data_li [233];
      \piso.data_r_232_sv2v_reg  <= \piso.data_li [232];
      \piso.data_r_231_sv2v_reg  <= \piso.data_li [231];
      \piso.data_r_230_sv2v_reg  <= \piso.data_li [230];
      \piso.data_r_229_sv2v_reg  <= \piso.data_li [229];
      \piso.data_r_228_sv2v_reg  <= \piso.data_li [228];
      \piso.data_r_227_sv2v_reg  <= \piso.data_li [227];
      \piso.data_r_226_sv2v_reg  <= \piso.data_li [226];
      \piso.data_r_225_sv2v_reg  <= \piso.data_li [225];
      \piso.data_r_224_sv2v_reg  <= \piso.data_li [224];
      \piso.data_r_223_sv2v_reg  <= \piso.data_li [223];
      \piso.data_r_222_sv2v_reg  <= \piso.data_li [222];
      \piso.data_r_221_sv2v_reg  <= \piso.data_li [221];
      \piso.data_r_220_sv2v_reg  <= \piso.data_li [220];
      \piso.data_r_219_sv2v_reg  <= \piso.data_li [219];
      \piso.data_r_218_sv2v_reg  <= \piso.data_li [218];
      \piso.data_r_217_sv2v_reg  <= \piso.data_li [217];
      \piso.data_r_216_sv2v_reg  <= \piso.data_li [216];
      \piso.data_r_215_sv2v_reg  <= \piso.data_li [215];
      \piso.data_r_214_sv2v_reg  <= \piso.data_li [214];
      \piso.data_r_213_sv2v_reg  <= \piso.data_li [213];
      \piso.data_r_212_sv2v_reg  <= \piso.data_li [212];
      \piso.data_r_211_sv2v_reg  <= \piso.data_li [211];
      \piso.data_r_210_sv2v_reg  <= \piso.data_li [210];
      \piso.data_r_209_sv2v_reg  <= \piso.data_li [209];
      \piso.data_r_208_sv2v_reg  <= \piso.data_li [208];
      \piso.data_r_207_sv2v_reg  <= \piso.data_li [207];
      \piso.data_r_206_sv2v_reg  <= \piso.data_li [206];
      \piso.data_r_205_sv2v_reg  <= \piso.data_li [205];
      \piso.data_r_204_sv2v_reg  <= \piso.data_li [204];
      \piso.data_r_203_sv2v_reg  <= \piso.data_li [203];
      \piso.data_r_202_sv2v_reg  <= \piso.data_li [202];
      \piso.data_r_201_sv2v_reg  <= \piso.data_li [201];
      \piso.data_r_200_sv2v_reg  <= \piso.data_li [200];
      \piso.data_r_199_sv2v_reg  <= \piso.data_li [199];
      \piso.data_r_198_sv2v_reg  <= \piso.data_li [198];
      \piso.data_r_197_sv2v_reg  <= \piso.data_li [197];
      \piso.data_r_196_sv2v_reg  <= \piso.data_li [196];
      \piso.data_r_195_sv2v_reg  <= \piso.data_li [195];
      \piso.data_r_194_sv2v_reg  <= \piso.data_li [194];
      \piso.data_r_193_sv2v_reg  <= \piso.data_li [193];
      \piso.data_r_192_sv2v_reg  <= \piso.data_li [192];
      \piso.data_r_191_sv2v_reg  <= \piso.data_li [191];
      \piso.data_r_190_sv2v_reg  <= \piso.data_li [190];
      \piso.data_r_189_sv2v_reg  <= \piso.data_li [189];
      \piso.data_r_188_sv2v_reg  <= \piso.data_li [188];
      \piso.data_r_187_sv2v_reg  <= \piso.data_li [187];
      \piso.data_r_186_sv2v_reg  <= \piso.data_li [186];
      \piso.data_r_185_sv2v_reg  <= \piso.data_li [185];
      \piso.data_r_184_sv2v_reg  <= \piso.data_li [184];
      \piso.data_r_183_sv2v_reg  <= \piso.data_li [183];
      \piso.data_r_182_sv2v_reg  <= \piso.data_li [182];
      \piso.data_r_181_sv2v_reg  <= \piso.data_li [181];
      \piso.data_r_180_sv2v_reg  <= \piso.data_li [180];
      \piso.data_r_179_sv2v_reg  <= \piso.data_li [179];
      \piso.data_r_178_sv2v_reg  <= \piso.data_li [178];
      \piso.data_r_177_sv2v_reg  <= \piso.data_li [177];
      \piso.data_r_176_sv2v_reg  <= \piso.data_li [176];
      \piso.data_r_175_sv2v_reg  <= \piso.data_li [175];
      \piso.data_r_174_sv2v_reg  <= \piso.data_li [174];
      \piso.data_r_173_sv2v_reg  <= \piso.data_li [173];
      \piso.data_r_172_sv2v_reg  <= \piso.data_li [172];
      \piso.data_r_171_sv2v_reg  <= \piso.data_li [171];
      \piso.data_r_170_sv2v_reg  <= \piso.data_li [170];
      \piso.data_r_169_sv2v_reg  <= \piso.data_li [169];
      \piso.data_r_168_sv2v_reg  <= \piso.data_li [168];
      \piso.data_r_167_sv2v_reg  <= \piso.data_li [167];
      \piso.data_r_166_sv2v_reg  <= \piso.data_li [166];
      \piso.data_r_165_sv2v_reg  <= \piso.data_li [165];
      \piso.data_r_164_sv2v_reg  <= \piso.data_li [164];
      \piso.data_r_163_sv2v_reg  <= \piso.data_li [163];
      \piso.data_r_162_sv2v_reg  <= \piso.data_li [162];
      \piso.data_r_161_sv2v_reg  <= \piso.data_li [161];
      \piso.data_r_160_sv2v_reg  <= \piso.data_li [160];
      \piso.data_r_159_sv2v_reg  <= \piso.data_li [159];
      \piso.data_r_158_sv2v_reg  <= \piso.data_li [158];
      \piso.data_r_157_sv2v_reg  <= \piso.data_li [157];
      \piso.data_r_156_sv2v_reg  <= \piso.data_li [156];
      \piso.data_r_155_sv2v_reg  <= \piso.data_li [155];
      \piso.data_r_154_sv2v_reg  <= \piso.data_li [154];
      \piso.data_r_153_sv2v_reg  <= \piso.data_li [153];
      \piso.data_r_152_sv2v_reg  <= \piso.data_li [152];
      \piso.data_r_151_sv2v_reg  <= \piso.data_li [151];
      \piso.data_r_150_sv2v_reg  <= \piso.data_li [150];
      \piso.data_r_149_sv2v_reg  <= \piso.data_li [149];
      \piso.data_r_148_sv2v_reg  <= \piso.data_li [148];
      \piso.data_r_147_sv2v_reg  <= \piso.data_li [147];
      \piso.data_r_146_sv2v_reg  <= \piso.data_li [146];
      \piso.data_r_145_sv2v_reg  <= \piso.data_li [145];
      \piso.data_r_144_sv2v_reg  <= \piso.data_li [144];
      \piso.data_r_143_sv2v_reg  <= \piso.data_li [143];
      \piso.data_r_142_sv2v_reg  <= \piso.data_li [142];
      \piso.data_r_141_sv2v_reg  <= \piso.data_li [141];
      \piso.data_r_140_sv2v_reg  <= \piso.data_li [140];
      \piso.data_r_139_sv2v_reg  <= \piso.data_li [139];
      \piso.data_r_138_sv2v_reg  <= \piso.data_li [138];
      \piso.data_r_137_sv2v_reg  <= \piso.data_li [137];
      \piso.data_r_136_sv2v_reg  <= \piso.data_li [136];
      \piso.data_r_135_sv2v_reg  <= \piso.data_li [135];
      \piso.data_r_134_sv2v_reg  <= \piso.data_li [134];
      \piso.data_r_133_sv2v_reg  <= \piso.data_li [133];
      \piso.data_r_132_sv2v_reg  <= \piso.data_li [132];
      \piso.data_r_131_sv2v_reg  <= \piso.data_li [131];
      \piso.data_r_130_sv2v_reg  <= \piso.data_li [130];
      \piso.data_r_129_sv2v_reg  <= \piso.data_li [129];
      \piso.data_r_128_sv2v_reg  <= \piso.data_li [128];
      \piso.data_r_127_sv2v_reg  <= \piso.data_li [127];
      \piso.data_r_126_sv2v_reg  <= \piso.data_li [126];
      \piso.data_r_125_sv2v_reg  <= \piso.data_li [125];
      \piso.data_r_124_sv2v_reg  <= \piso.data_li [124];
      \piso.data_r_123_sv2v_reg  <= \piso.data_li [123];
      \piso.data_r_122_sv2v_reg  <= \piso.data_li [122];
      \piso.data_r_121_sv2v_reg  <= \piso.data_li [121];
      \piso.data_r_120_sv2v_reg  <= \piso.data_li [120];
      \piso.data_r_119_sv2v_reg  <= \piso.data_li [119];
      \piso.data_r_118_sv2v_reg  <= \piso.data_li [118];
      \piso.data_r_117_sv2v_reg  <= \piso.data_li [117];
      \piso.data_r_116_sv2v_reg  <= \piso.data_li [116];
      \piso.data_r_115_sv2v_reg  <= \piso.data_li [115];
      \piso.data_r_114_sv2v_reg  <= \piso.data_li [114];
      \piso.data_r_113_sv2v_reg  <= \piso.data_li [113];
      \piso.data_r_112_sv2v_reg  <= \piso.data_li [112];
      \piso.data_r_111_sv2v_reg  <= \piso.data_li [111];
      \piso.data_r_110_sv2v_reg  <= \piso.data_li [110];
      \piso.data_r_109_sv2v_reg  <= \piso.data_li [109];
      \piso.data_r_108_sv2v_reg  <= \piso.data_li [108];
      \piso.data_r_107_sv2v_reg  <= \piso.data_li [107];
      \piso.data_r_106_sv2v_reg  <= \piso.data_li [106];
      \piso.data_r_105_sv2v_reg  <= \piso.data_li [105];
      \piso.data_r_104_sv2v_reg  <= \piso.data_li [104];
      \piso.data_r_103_sv2v_reg  <= \piso.data_li [103];
      \piso.data_r_102_sv2v_reg  <= \piso.data_li [102];
      \piso.data_r_101_sv2v_reg  <= \piso.data_li [101];
      \piso.data_r_100_sv2v_reg  <= \piso.data_li [100];
      \piso.data_r_99_sv2v_reg  <= \piso.data_li [99];
      \piso.data_r_98_sv2v_reg  <= \piso.data_li [98];
      \piso.data_r_97_sv2v_reg  <= \piso.data_li [97];
      \piso.data_r_96_sv2v_reg  <= \piso.data_li [96];
      \piso.data_r_95_sv2v_reg  <= \piso.data_li [95];
      \piso.data_r_94_sv2v_reg  <= \piso.data_li [94];
      \piso.data_r_93_sv2v_reg  <= \piso.data_li [93];
      \piso.data_r_92_sv2v_reg  <= \piso.data_li [92];
      \piso.data_r_91_sv2v_reg  <= \piso.data_li [91];
      \piso.data_r_90_sv2v_reg  <= \piso.data_li [90];
      \piso.data_r_89_sv2v_reg  <= \piso.data_li [89];
      \piso.data_r_88_sv2v_reg  <= \piso.data_li [88];
      \piso.data_r_87_sv2v_reg  <= \piso.data_li [87];
      \piso.data_r_86_sv2v_reg  <= \piso.data_li [86];
      \piso.data_r_85_sv2v_reg  <= \piso.data_li [85];
      \piso.data_r_84_sv2v_reg  <= \piso.data_li [84];
      \piso.data_r_83_sv2v_reg  <= \piso.data_li [83];
      \piso.data_r_82_sv2v_reg  <= \piso.data_li [82];
      \piso.data_r_81_sv2v_reg  <= \piso.data_li [81];
      \piso.data_r_80_sv2v_reg  <= \piso.data_li [80];
      \piso.data_r_79_sv2v_reg  <= \piso.data_li [79];
      \piso.data_r_78_sv2v_reg  <= \piso.data_li [78];
      \piso.data_r_77_sv2v_reg  <= \piso.data_li [77];
      \piso.data_r_76_sv2v_reg  <= \piso.data_li [76];
      \piso.data_r_75_sv2v_reg  <= \piso.data_li [75];
      \piso.data_r_74_sv2v_reg  <= \piso.data_li [74];
      \piso.data_r_73_sv2v_reg  <= \piso.data_li [73];
      \piso.data_r_72_sv2v_reg  <= \piso.data_li [72];
      \piso.data_r_71_sv2v_reg  <= \piso.data_li [71];
      \piso.data_r_70_sv2v_reg  <= \piso.data_li [70];
      \piso.data_r_69_sv2v_reg  <= \piso.data_li [69];
      \piso.data_r_68_sv2v_reg  <= \piso.data_li [68];
      \piso.data_r_67_sv2v_reg  <= \piso.data_li [67];
      \piso.data_r_66_sv2v_reg  <= \piso.data_li [66];
      \piso.data_r_65_sv2v_reg  <= \piso.data_li [65];
      \piso.data_r_64_sv2v_reg  <= \piso.data_li [64];
      \piso.data_r_63_sv2v_reg  <= \piso.data_li [63];
      \piso.data_r_62_sv2v_reg  <= \piso.data_li [62];
      \piso.data_r_61_sv2v_reg  <= \piso.data_li [61];
      \piso.data_r_60_sv2v_reg  <= \piso.data_li [60];
      \piso.data_r_59_sv2v_reg  <= \piso.data_li [59];
      \piso.data_r_58_sv2v_reg  <= \piso.data_li [58];
      \piso.data_r_57_sv2v_reg  <= \piso.data_li [57];
      \piso.data_r_56_sv2v_reg  <= \piso.data_li [56];
      \piso.data_r_55_sv2v_reg  <= \piso.data_li [55];
      \piso.data_r_54_sv2v_reg  <= \piso.data_li [54];
      \piso.data_r_53_sv2v_reg  <= \piso.data_li [53];
      \piso.data_r_52_sv2v_reg  <= \piso.data_li [52];
      \piso.data_r_51_sv2v_reg  <= \piso.data_li [51];
      \piso.data_r_50_sv2v_reg  <= \piso.data_li [50];
      \piso.data_r_49_sv2v_reg  <= \piso.data_li [49];
      \piso.data_r_48_sv2v_reg  <= \piso.data_li [48];
      \piso.data_r_47_sv2v_reg  <= \piso.data_li [47];
      \piso.data_r_46_sv2v_reg  <= \piso.data_li [46];
      \piso.data_r_45_sv2v_reg  <= \piso.data_li [45];
      \piso.data_r_44_sv2v_reg  <= \piso.data_li [44];
      \piso.data_r_43_sv2v_reg  <= \piso.data_li [43];
      \piso.data_r_42_sv2v_reg  <= \piso.data_li [42];
      \piso.data_r_41_sv2v_reg  <= \piso.data_li [41];
      \piso.data_r_40_sv2v_reg  <= \piso.data_li [40];
      \piso.data_r_39_sv2v_reg  <= \piso.data_li [39];
      \piso.data_r_38_sv2v_reg  <= \piso.data_li [38];
      \piso.data_r_37_sv2v_reg  <= \piso.data_li [37];
      \piso.data_r_36_sv2v_reg  <= \piso.data_li [36];
      \piso.data_r_35_sv2v_reg  <= \piso.data_li [35];
      \piso.data_r_34_sv2v_reg  <= \piso.data_li [34];
      \piso.data_r_33_sv2v_reg  <= \piso.data_li [33];
      \piso.data_r_32_sv2v_reg  <= \piso.data_li [32];
      \piso.data_r_31_sv2v_reg  <= \piso.data_li [31];
      \piso.data_r_30_sv2v_reg  <= \piso.data_li [30];
      \piso.data_r_29_sv2v_reg  <= \piso.data_li [29];
      \piso.data_r_28_sv2v_reg  <= \piso.data_li [28];
      \piso.data_r_27_sv2v_reg  <= \piso.data_li [27];
      \piso.data_r_26_sv2v_reg  <= \piso.data_li [26];
      \piso.data_r_25_sv2v_reg  <= \piso.data_li [25];
      \piso.data_r_24_sv2v_reg  <= \piso.data_li [24];
      \piso.data_r_23_sv2v_reg  <= \piso.data_li [23];
      \piso.data_r_22_sv2v_reg  <= \piso.data_li [22];
      \piso.data_r_21_sv2v_reg  <= \piso.data_li [21];
      \piso.data_r_20_sv2v_reg  <= \piso.data_li [20];
      \piso.data_r_19_sv2v_reg  <= \piso.data_li [19];
      \piso.data_r_18_sv2v_reg  <= \piso.data_li [18];
      \piso.data_r_17_sv2v_reg  <= \piso.data_li [17];
      \piso.data_r_16_sv2v_reg  <= \piso.data_li [16];
      \piso.data_r_15_sv2v_reg  <= \piso.data_li [15];
      \piso.data_r_14_sv2v_reg  <= \piso.data_li [14];
      \piso.data_r_13_sv2v_reg  <= \piso.data_li [13];
      \piso.data_r_12_sv2v_reg  <= \piso.data_li [12];
      \piso.data_r_11_sv2v_reg  <= \piso.data_li [11];
      \piso.data_r_10_sv2v_reg  <= \piso.data_li [10];
      \piso.data_r_9_sv2v_reg  <= \piso.data_li [9];
      \piso.data_r_8_sv2v_reg  <= \piso.data_li [8];
      \piso.data_r_7_sv2v_reg  <= \piso.data_li [7];
      \piso.data_r_6_sv2v_reg  <= \piso.data_li [6];
      \piso.data_r_5_sv2v_reg  <= \piso.data_li [5];
      \piso.data_r_4_sv2v_reg  <= \piso.data_li [4];
      \piso.data_r_3_sv2v_reg  <= \piso.data_li [3];
      \piso.data_r_2_sv2v_reg  <= \piso.data_li [2];
      \piso.data_r_1_sv2v_reg  <= \piso.data_li [1];
      \piso.data_r_0_sv2v_reg  <= \piso.data_li [0];
    end 
    if(reset_i) begin
      \piso.shift_ctr_r_6_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_5_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_4_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_3_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_2_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_1_sv2v_reg  <= 1'b0;
      \piso.shift_ctr_r_0_sv2v_reg  <= 1'b0;
    end else if(N285) begin
      \piso.shift_ctr_r_6_sv2v_reg  <= N15;
      \piso.shift_ctr_r_5_sv2v_reg  <= N14;
      \piso.shift_ctr_r_4_sv2v_reg  <= N13;
      \piso.shift_ctr_r_3_sv2v_reg  <= N12;
      \piso.shift_ctr_r_2_sv2v_reg  <= N11;
      \piso.shift_ctr_r_1_sv2v_reg  <= N10;
      \piso.shift_ctr_r_0_sv2v_reg  <= N9;
    end 
  end


endmodule

