

module top
(
  clk_i,
  reset_i,
  en_i,
  v_i,
  a_i,
  b_i,
  sub_i,
  ready_o,
  v_o,
  z_o,
  unimplemented_o,
  invalid_o,
  overflow_o,
  underflow_o,
  yumi_i
);

  input [127:0] a_i;
  input [127:0] b_i;
  output [127:0] z_o;
  input clk_i;
  input reset_i;
  input en_i;
  input v_i;
  input sub_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output unimplemented_o;
  output invalid_o;
  output overflow_o;
  output underflow_o;

  bsg_fpu_add_sub
  wrapper
  (
    .a_i(a_i),
    .b_i(b_i),
    .z_o(z_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(en_i),
    .v_i(v_i),
    .sub_i(sub_i),
    .yumi_i(yumi_i),
    .ready_o(ready_o),
    .v_o(v_o),
    .unimplemented_o(unimplemented_o),
    .invalid_o(invalid_o),
    .overflow_o(overflow_o),
    .underflow_o(underflow_o)
  );


endmodule



module bsg_fpu_preprocess_e_p15_m_p112
(
  a_i,
  zero_o,
  nan_o,
  sig_nan_o,
  infty_o,
  exp_zero_o,
  man_zero_o,
  denormal_o,
  sign_o,
  exp_o,
  man_o
);

  input [127:0] a_i;
  output [14:0] exp_o;
  output [111:0] man_o;
  output zero_o;
  output nan_o;
  output sig_nan_o;
  output infty_o;
  output exp_zero_o;
  output man_zero_o;
  output denormal_o;
  output sign_o;
  wire [14:0] exp_o;
  wire [111:0] man_o;
  wire zero_o,nan_o,sig_nan_o,infty_o,exp_zero_o,man_zero_o,denormal_o,sign_o,N0,N1,N2,
  N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,
  N136,N137,N138,N139,N141;
  assign man_o[111] = a_i[111];
  assign man_o[110] = a_i[110];
  assign man_o[109] = a_i[109];
  assign man_o[108] = a_i[108];
  assign man_o[107] = a_i[107];
  assign man_o[106] = a_i[106];
  assign man_o[105] = a_i[105];
  assign man_o[104] = a_i[104];
  assign man_o[103] = a_i[103];
  assign man_o[102] = a_i[102];
  assign man_o[101] = a_i[101];
  assign man_o[100] = a_i[100];
  assign man_o[99] = a_i[99];
  assign man_o[98] = a_i[98];
  assign man_o[97] = a_i[97];
  assign man_o[96] = a_i[96];
  assign man_o[95] = a_i[95];
  assign man_o[94] = a_i[94];
  assign man_o[93] = a_i[93];
  assign man_o[92] = a_i[92];
  assign man_o[91] = a_i[91];
  assign man_o[90] = a_i[90];
  assign man_o[89] = a_i[89];
  assign man_o[88] = a_i[88];
  assign man_o[87] = a_i[87];
  assign man_o[86] = a_i[86];
  assign man_o[85] = a_i[85];
  assign man_o[84] = a_i[84];
  assign man_o[83] = a_i[83];
  assign man_o[82] = a_i[82];
  assign man_o[81] = a_i[81];
  assign man_o[80] = a_i[80];
  assign man_o[79] = a_i[79];
  assign man_o[78] = a_i[78];
  assign man_o[77] = a_i[77];
  assign man_o[76] = a_i[76];
  assign man_o[75] = a_i[75];
  assign man_o[74] = a_i[74];
  assign man_o[73] = a_i[73];
  assign man_o[72] = a_i[72];
  assign man_o[71] = a_i[71];
  assign man_o[70] = a_i[70];
  assign man_o[69] = a_i[69];
  assign man_o[68] = a_i[68];
  assign man_o[67] = a_i[67];
  assign man_o[66] = a_i[66];
  assign man_o[65] = a_i[65];
  assign man_o[64] = a_i[64];
  assign man_o[63] = a_i[63];
  assign man_o[62] = a_i[62];
  assign man_o[61] = a_i[61];
  assign man_o[60] = a_i[60];
  assign man_o[59] = a_i[59];
  assign man_o[58] = a_i[58];
  assign man_o[57] = a_i[57];
  assign man_o[56] = a_i[56];
  assign man_o[55] = a_i[55];
  assign man_o[54] = a_i[54];
  assign man_o[53] = a_i[53];
  assign man_o[52] = a_i[52];
  assign man_o[51] = a_i[51];
  assign man_o[50] = a_i[50];
  assign man_o[49] = a_i[49];
  assign man_o[48] = a_i[48];
  assign man_o[47] = a_i[47];
  assign man_o[46] = a_i[46];
  assign man_o[45] = a_i[45];
  assign man_o[44] = a_i[44];
  assign man_o[43] = a_i[43];
  assign man_o[42] = a_i[42];
  assign man_o[41] = a_i[41];
  assign man_o[40] = a_i[40];
  assign man_o[39] = a_i[39];
  assign man_o[38] = a_i[38];
  assign man_o[37] = a_i[37];
  assign man_o[36] = a_i[36];
  assign man_o[35] = a_i[35];
  assign man_o[34] = a_i[34];
  assign man_o[33] = a_i[33];
  assign man_o[32] = a_i[32];
  assign man_o[31] = a_i[31];
  assign man_o[30] = a_i[30];
  assign man_o[29] = a_i[29];
  assign man_o[28] = a_i[28];
  assign man_o[27] = a_i[27];
  assign man_o[26] = a_i[26];
  assign man_o[25] = a_i[25];
  assign man_o[24] = a_i[24];
  assign man_o[23] = a_i[23];
  assign man_o[22] = a_i[22];
  assign man_o[21] = a_i[21];
  assign man_o[20] = a_i[20];
  assign man_o[19] = a_i[19];
  assign man_o[18] = a_i[18];
  assign man_o[17] = a_i[17];
  assign man_o[16] = a_i[16];
  assign man_o[15] = a_i[15];
  assign man_o[14] = a_i[14];
  assign man_o[13] = a_i[13];
  assign man_o[12] = a_i[12];
  assign man_o[11] = a_i[11];
  assign man_o[10] = a_i[10];
  assign man_o[9] = a_i[9];
  assign man_o[8] = a_i[8];
  assign man_o[7] = a_i[7];
  assign man_o[6] = a_i[6];
  assign man_o[5] = a_i[5];
  assign man_o[4] = a_i[4];
  assign man_o[3] = a_i[3];
  assign man_o[2] = a_i[2];
  assign man_o[1] = a_i[1];
  assign man_o[0] = a_i[0];
  assign exp_o[14] = a_i[126];
  assign exp_o[13] = a_i[125];
  assign exp_o[12] = a_i[124];
  assign exp_o[11] = a_i[123];
  assign exp_o[10] = a_i[122];
  assign exp_o[9] = a_i[121];
  assign exp_o[8] = a_i[120];
  assign exp_o[7] = a_i[119];
  assign exp_o[6] = a_i[118];
  assign exp_o[5] = a_i[117];
  assign exp_o[4] = a_i[116];
  assign exp_o[3] = a_i[115];
  assign exp_o[2] = a_i[114];
  assign exp_o[1] = a_i[113];
  assign exp_o[0] = a_i[112];
  assign sign_o = a_i[127];
  assign N0 = a_i[125] | a_i[126];
  assign N1 = a_i[124] | N0;
  assign N2 = a_i[123] | N1;
  assign N3 = a_i[122] | N2;
  assign N4 = a_i[121] | N3;
  assign N5 = a_i[120] | N4;
  assign N6 = a_i[119] | N5;
  assign N7 = a_i[118] | N6;
  assign N8 = a_i[117] | N7;
  assign N9 = a_i[116] | N8;
  assign N10 = a_i[115] | N9;
  assign N11 = a_i[114] | N10;
  assign N12 = a_i[113] | N11;
  assign N13 = a_i[112] | N12;
  assign exp_zero_o = ~N13;
  assign N15 = a_i[125] & a_i[126];
  assign N16 = a_i[124] & N15;
  assign N17 = a_i[123] & N16;
  assign N18 = a_i[122] & N17;
  assign N19 = a_i[121] & N18;
  assign N20 = a_i[120] & N19;
  assign N21 = a_i[119] & N20;
  assign N22 = a_i[118] & N21;
  assign N23 = a_i[117] & N22;
  assign N24 = a_i[116] & N23;
  assign N25 = a_i[115] & N24;
  assign N26 = a_i[114] & N25;
  assign N27 = a_i[113] & N26;
  assign N28 = a_i[112] & N27;
  assign N29 = a_i[110] | a_i[111];
  assign N30 = a_i[109] | N29;
  assign N31 = a_i[108] | N30;
  assign N32 = a_i[107] | N31;
  assign N33 = a_i[106] | N32;
  assign N34 = a_i[105] | N33;
  assign N35 = a_i[104] | N34;
  assign N36 = a_i[103] | N35;
  assign N37 = a_i[102] | N36;
  assign N38 = a_i[101] | N37;
  assign N39 = a_i[100] | N38;
  assign N40 = a_i[99] | N39;
  assign N41 = a_i[98] | N40;
  assign N42 = a_i[97] | N41;
  assign N43 = a_i[96] | N42;
  assign N44 = a_i[95] | N43;
  assign N45 = a_i[94] | N44;
  assign N46 = a_i[93] | N45;
  assign N47 = a_i[92] | N46;
  assign N48 = a_i[91] | N47;
  assign N49 = a_i[90] | N48;
  assign N50 = a_i[89] | N49;
  assign N51 = a_i[88] | N50;
  assign N52 = a_i[87] | N51;
  assign N53 = a_i[86] | N52;
  assign N54 = a_i[85] | N53;
  assign N55 = a_i[84] | N54;
  assign N56 = a_i[83] | N55;
  assign N57 = a_i[82] | N56;
  assign N58 = a_i[81] | N57;
  assign N59 = a_i[80] | N58;
  assign N60 = a_i[79] | N59;
  assign N61 = a_i[78] | N60;
  assign N62 = a_i[77] | N61;
  assign N63 = a_i[76] | N62;
  assign N64 = a_i[75] | N63;
  assign N65 = a_i[74] | N64;
  assign N66 = a_i[73] | N65;
  assign N67 = a_i[72] | N66;
  assign N68 = a_i[71] | N67;
  assign N69 = a_i[70] | N68;
  assign N70 = a_i[69] | N69;
  assign N71 = a_i[68] | N70;
  assign N72 = a_i[67] | N71;
  assign N73 = a_i[66] | N72;
  assign N74 = a_i[65] | N73;
  assign N75 = a_i[64] | N74;
  assign N76 = a_i[63] | N75;
  assign N77 = a_i[62] | N76;
  assign N78 = a_i[61] | N77;
  assign N79 = a_i[60] | N78;
  assign N80 = a_i[59] | N79;
  assign N81 = a_i[58] | N80;
  assign N82 = a_i[57] | N81;
  assign N83 = a_i[56] | N82;
  assign N84 = a_i[55] | N83;
  assign N85 = a_i[54] | N84;
  assign N86 = a_i[53] | N85;
  assign N87 = a_i[52] | N86;
  assign N88 = a_i[51] | N87;
  assign N89 = a_i[50] | N88;
  assign N90 = a_i[49] | N89;
  assign N91 = a_i[48] | N90;
  assign N92 = a_i[47] | N91;
  assign N93 = a_i[46] | N92;
  assign N94 = a_i[45] | N93;
  assign N95 = a_i[44] | N94;
  assign N96 = a_i[43] | N95;
  assign N97 = a_i[42] | N96;
  assign N98 = a_i[41] | N97;
  assign N99 = a_i[40] | N98;
  assign N100 = a_i[39] | N99;
  assign N101 = a_i[38] | N100;
  assign N102 = a_i[37] | N101;
  assign N103 = a_i[36] | N102;
  assign N104 = a_i[35] | N103;
  assign N105 = a_i[34] | N104;
  assign N106 = a_i[33] | N105;
  assign N107 = a_i[32] | N106;
  assign N108 = a_i[31] | N107;
  assign N109 = a_i[30] | N108;
  assign N110 = a_i[29] | N109;
  assign N111 = a_i[28] | N110;
  assign N112 = a_i[27] | N111;
  assign N113 = a_i[26] | N112;
  assign N114 = a_i[25] | N113;
  assign N115 = a_i[24] | N114;
  assign N116 = a_i[23] | N115;
  assign N117 = a_i[22] | N116;
  assign N118 = a_i[21] | N117;
  assign N119 = a_i[20] | N118;
  assign N120 = a_i[19] | N119;
  assign N121 = a_i[18] | N120;
  assign N122 = a_i[17] | N121;
  assign N123 = a_i[16] | N122;
  assign N124 = a_i[15] | N123;
  assign N125 = a_i[14] | N124;
  assign N126 = a_i[13] | N125;
  assign N127 = a_i[12] | N126;
  assign N128 = a_i[11] | N127;
  assign N129 = a_i[10] | N128;
  assign N130 = a_i[9] | N129;
  assign N131 = a_i[8] | N130;
  assign N132 = a_i[7] | N131;
  assign N133 = a_i[6] | N132;
  assign N134 = a_i[5] | N133;
  assign N135 = a_i[4] | N134;
  assign N136 = a_i[3] | N135;
  assign N137 = a_i[2] | N136;
  assign N138 = a_i[1] | N137;
  assign N139 = a_i[0] | N138;
  assign man_zero_o = ~N139;
  assign zero_o = exp_zero_o & man_zero_o;
  assign nan_o = N28 & N139;
  assign sig_nan_o = nan_o & N141;
  assign N141 = ~a_i[111];
  assign infty_o = N28 & man_zero_o;
  assign denormal_o = exp_zero_o & N139;

endmodule



module bsg_less_than_width_p15
(
  a_i,
  b_i,
  o
);

  input [14:0] a_i;
  input [14:0] b_i;
  output o;
  wire o;
  assign o = a_i < b_i;

endmodule



module bsg_scan_width_p115_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [114:0] i;
  output [114:0] o;
  wire [114:0] o;
  wire t_6__114_,t_6__113_,t_6__112_,t_6__111_,t_6__110_,t_6__109_,t_6__108_,t_6__107_,
  t_6__106_,t_6__105_,t_6__104_,t_6__103_,t_6__102_,t_6__101_,t_6__100_,t_6__99_,
  t_6__98_,t_6__97_,t_6__96_,t_6__95_,t_6__94_,t_6__93_,t_6__92_,t_6__91_,t_6__90_,
  t_6__89_,t_6__88_,t_6__87_,t_6__86_,t_6__85_,t_6__84_,t_6__83_,t_6__82_,
  t_6__81_,t_6__80_,t_6__79_,t_6__78_,t_6__77_,t_6__76_,t_6__75_,t_6__74_,t_6__73_,
  t_6__72_,t_6__71_,t_6__70_,t_6__69_,t_6__68_,t_6__67_,t_6__66_,t_6__65_,t_6__64_,
  t_6__63_,t_6__62_,t_6__61_,t_6__60_,t_6__59_,t_6__58_,t_6__57_,t_6__56_,t_6__55_,
  t_6__54_,t_6__53_,t_6__52_,t_6__51_,t_6__50_,t_6__49_,t_6__48_,t_6__47_,t_6__46_,
  t_6__45_,t_6__44_,t_6__43_,t_6__42_,t_6__41_,t_6__40_,t_6__39_,t_6__38_,t_6__37_,
  t_6__36_,t_6__35_,t_6__34_,t_6__33_,t_6__32_,t_6__31_,t_6__30_,t_6__29_,t_6__28_,
  t_6__27_,t_6__26_,t_6__25_,t_6__24_,t_6__23_,t_6__22_,t_6__21_,t_6__20_,t_6__19_,
  t_6__18_,t_6__17_,t_6__16_,t_6__15_,t_6__14_,t_6__13_,t_6__12_,t_6__11_,t_6__10_,
  t_6__9_,t_6__8_,t_6__7_,t_6__6_,t_6__5_,t_6__4_,t_6__3_,t_6__2_,t_6__1_,t_6__0_,
  t_5__114_,t_5__113_,t_5__112_,t_5__111_,t_5__110_,t_5__109_,t_5__108_,t_5__107_,
  t_5__106_,t_5__105_,t_5__104_,t_5__103_,t_5__102_,t_5__101_,t_5__100_,t_5__99_,
  t_5__98_,t_5__97_,t_5__96_,t_5__95_,t_5__94_,t_5__93_,t_5__92_,t_5__91_,t_5__90_,
  t_5__89_,t_5__88_,t_5__87_,t_5__86_,t_5__85_,t_5__84_,t_5__83_,t_5__82_,
  t_5__81_,t_5__80_,t_5__79_,t_5__78_,t_5__77_,t_5__76_,t_5__75_,t_5__74_,t_5__73_,
  t_5__72_,t_5__71_,t_5__70_,t_5__69_,t_5__68_,t_5__67_,t_5__66_,t_5__65_,t_5__64_,
  t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,t_5__55_,
  t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,t_5__46_,
  t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,t_5__37_,
  t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,t_5__28_,
  t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,t_5__19_,
  t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,t_5__11_,t_5__10_,
  t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,t_5__1_,t_5__0_,
  t_4__114_,t_4__113_,t_4__112_,t_4__111_,t_4__110_,t_4__109_,t_4__108_,t_4__107_,
  t_4__106_,t_4__105_,t_4__104_,t_4__103_,t_4__102_,t_4__101_,t_4__100_,t_4__99_,
  t_4__98_,t_4__97_,t_4__96_,t_4__95_,t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,
  t_4__89_,t_4__88_,t_4__87_,t_4__86_,t_4__85_,t_4__84_,t_4__83_,t_4__82_,
  t_4__81_,t_4__80_,t_4__79_,t_4__78_,t_4__77_,t_4__76_,t_4__75_,t_4__74_,t_4__73_,
  t_4__72_,t_4__71_,t_4__70_,t_4__69_,t_4__68_,t_4__67_,t_4__66_,t_4__65_,t_4__64_,
  t_4__63_,t_4__62_,t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,
  t_4__54_,t_4__53_,t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,
  t_4__45_,t_4__44_,t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,
  t_4__36_,t_4__35_,t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,
  t_4__27_,t_4__26_,t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,
  t_4__18_,t_4__17_,t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,
  t_4__9_,t_4__8_,t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_,
  t_3__114_,t_3__113_,t_3__112_,t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,
  t_3__106_,t_3__105_,t_3__104_,t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,
  t_3__98_,t_3__97_,t_3__96_,t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,
  t_3__89_,t_3__88_,t_3__87_,t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,
  t_3__81_,t_3__80_,t_3__79_,t_3__78_,t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,
  t_3__72_,t_3__71_,t_3__70_,t_3__69_,t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,
  t_3__63_,t_3__62_,t_3__61_,t_3__60_,t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,
  t_3__54_,t_3__53_,t_3__52_,t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,
  t_3__45_,t_3__44_,t_3__43_,t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,
  t_3__36_,t_3__35_,t_3__34_,t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,
  t_3__27_,t_3__26_,t_3__25_,t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,
  t_3__18_,t_3__17_,t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,
  t_3__9_,t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,
  t_2__114_,t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,t_2__108_,t_2__107_,
  t_2__106_,t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,t_2__100_,t_2__99_,
  t_2__98_,t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,t_2__92_,t_2__91_,t_2__90_,
  t_2__89_,t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,t_2__83_,t_2__82_,
  t_2__81_,t_2__80_,t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,t_2__74_,t_2__73_,
  t_2__72_,t_2__71_,t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,t_2__65_,t_2__64_,
  t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,t_2__56_,t_2__55_,
  t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,t_2__47_,t_2__46_,
  t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,t_2__38_,t_2__37_,
  t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,t_2__29_,t_2__28_,
  t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,t_2__21_,t_2__20_,t_2__19_,
  t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,t_2__12_,t_2__11_,t_2__10_,
  t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,
  t_1__114_,t_1__113_,t_1__112_,t_1__111_,t_1__110_,t_1__109_,t_1__108_,t_1__107_,
  t_1__106_,t_1__105_,t_1__104_,t_1__103_,t_1__102_,t_1__101_,t_1__100_,t_1__99_,
  t_1__98_,t_1__97_,t_1__96_,t_1__95_,t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,
  t_1__89_,t_1__88_,t_1__87_,t_1__86_,t_1__85_,t_1__84_,t_1__83_,t_1__82_,
  t_1__81_,t_1__80_,t_1__79_,t_1__78_,t_1__77_,t_1__76_,t_1__75_,t_1__74_,t_1__73_,
  t_1__72_,t_1__71_,t_1__70_,t_1__69_,t_1__68_,t_1__67_,t_1__66_,t_1__65_,t_1__64_,
  t_1__63_,t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,t_1__57_,t_1__56_,t_1__55_,
  t_1__54_,t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,
  t_1__45_,t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,
  t_1__36_,t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,
  t_1__27_,t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,
  t_1__18_,t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,
  t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__114_ = i[0] | 1'b0;
  assign t_1__113_ = i[1] | i[0];
  assign t_1__112_ = i[2] | i[1];
  assign t_1__111_ = i[3] | i[2];
  assign t_1__110_ = i[4] | i[3];
  assign t_1__109_ = i[5] | i[4];
  assign t_1__108_ = i[6] | i[5];
  assign t_1__107_ = i[7] | i[6];
  assign t_1__106_ = i[8] | i[7];
  assign t_1__105_ = i[9] | i[8];
  assign t_1__104_ = i[10] | i[9];
  assign t_1__103_ = i[11] | i[10];
  assign t_1__102_ = i[12] | i[11];
  assign t_1__101_ = i[13] | i[12];
  assign t_1__100_ = i[14] | i[13];
  assign t_1__99_ = i[15] | i[14];
  assign t_1__98_ = i[16] | i[15];
  assign t_1__97_ = i[17] | i[16];
  assign t_1__96_ = i[18] | i[17];
  assign t_1__95_ = i[19] | i[18];
  assign t_1__94_ = i[20] | i[19];
  assign t_1__93_ = i[21] | i[20];
  assign t_1__92_ = i[22] | i[21];
  assign t_1__91_ = i[23] | i[22];
  assign t_1__90_ = i[24] | i[23];
  assign t_1__89_ = i[25] | i[24];
  assign t_1__88_ = i[26] | i[25];
  assign t_1__87_ = i[27] | i[26];
  assign t_1__86_ = i[28] | i[27];
  assign t_1__85_ = i[29] | i[28];
  assign t_1__84_ = i[30] | i[29];
  assign t_1__83_ = i[31] | i[30];
  assign t_1__82_ = i[32] | i[31];
  assign t_1__81_ = i[33] | i[32];
  assign t_1__80_ = i[34] | i[33];
  assign t_1__79_ = i[35] | i[34];
  assign t_1__78_ = i[36] | i[35];
  assign t_1__77_ = i[37] | i[36];
  assign t_1__76_ = i[38] | i[37];
  assign t_1__75_ = i[39] | i[38];
  assign t_1__74_ = i[40] | i[39];
  assign t_1__73_ = i[41] | i[40];
  assign t_1__72_ = i[42] | i[41];
  assign t_1__71_ = i[43] | i[42];
  assign t_1__70_ = i[44] | i[43];
  assign t_1__69_ = i[45] | i[44];
  assign t_1__68_ = i[46] | i[45];
  assign t_1__67_ = i[47] | i[46];
  assign t_1__66_ = i[48] | i[47];
  assign t_1__65_ = i[49] | i[48];
  assign t_1__64_ = i[50] | i[49];
  assign t_1__63_ = i[51] | i[50];
  assign t_1__62_ = i[52] | i[51];
  assign t_1__61_ = i[53] | i[52];
  assign t_1__60_ = i[54] | i[53];
  assign t_1__59_ = i[55] | i[54];
  assign t_1__58_ = i[56] | i[55];
  assign t_1__57_ = i[57] | i[56];
  assign t_1__56_ = i[58] | i[57];
  assign t_1__55_ = i[59] | i[58];
  assign t_1__54_ = i[60] | i[59];
  assign t_1__53_ = i[61] | i[60];
  assign t_1__52_ = i[62] | i[61];
  assign t_1__51_ = i[63] | i[62];
  assign t_1__50_ = i[64] | i[63];
  assign t_1__49_ = i[65] | i[64];
  assign t_1__48_ = i[66] | i[65];
  assign t_1__47_ = i[67] | i[66];
  assign t_1__46_ = i[68] | i[67];
  assign t_1__45_ = i[69] | i[68];
  assign t_1__44_ = i[70] | i[69];
  assign t_1__43_ = i[71] | i[70];
  assign t_1__42_ = i[72] | i[71];
  assign t_1__41_ = i[73] | i[72];
  assign t_1__40_ = i[74] | i[73];
  assign t_1__39_ = i[75] | i[74];
  assign t_1__38_ = i[76] | i[75];
  assign t_1__37_ = i[77] | i[76];
  assign t_1__36_ = i[78] | i[77];
  assign t_1__35_ = i[79] | i[78];
  assign t_1__34_ = i[80] | i[79];
  assign t_1__33_ = i[81] | i[80];
  assign t_1__32_ = i[82] | i[81];
  assign t_1__31_ = i[83] | i[82];
  assign t_1__30_ = i[84] | i[83];
  assign t_1__29_ = i[85] | i[84];
  assign t_1__28_ = i[86] | i[85];
  assign t_1__27_ = i[87] | i[86];
  assign t_1__26_ = i[88] | i[87];
  assign t_1__25_ = i[89] | i[88];
  assign t_1__24_ = i[90] | i[89];
  assign t_1__23_ = i[91] | i[90];
  assign t_1__22_ = i[92] | i[91];
  assign t_1__21_ = i[93] | i[92];
  assign t_1__20_ = i[94] | i[93];
  assign t_1__19_ = i[95] | i[94];
  assign t_1__18_ = i[96] | i[95];
  assign t_1__17_ = i[97] | i[96];
  assign t_1__16_ = i[98] | i[97];
  assign t_1__15_ = i[99] | i[98];
  assign t_1__14_ = i[100] | i[99];
  assign t_1__13_ = i[101] | i[100];
  assign t_1__12_ = i[102] | i[101];
  assign t_1__11_ = i[103] | i[102];
  assign t_1__10_ = i[104] | i[103];
  assign t_1__9_ = i[105] | i[104];
  assign t_1__8_ = i[106] | i[105];
  assign t_1__7_ = i[107] | i[106];
  assign t_1__6_ = i[108] | i[107];
  assign t_1__5_ = i[109] | i[108];
  assign t_1__4_ = i[110] | i[109];
  assign t_1__3_ = i[111] | i[110];
  assign t_1__2_ = i[112] | i[111];
  assign t_1__1_ = i[113] | i[112];
  assign t_1__0_ = i[114] | i[113];
  assign t_2__114_ = t_1__114_ | 1'b0;
  assign t_2__113_ = t_1__113_ | 1'b0;
  assign t_2__112_ = t_1__112_ | t_1__114_;
  assign t_2__111_ = t_1__111_ | t_1__113_;
  assign t_2__110_ = t_1__110_ | t_1__112_;
  assign t_2__109_ = t_1__109_ | t_1__111_;
  assign t_2__108_ = t_1__108_ | t_1__110_;
  assign t_2__107_ = t_1__107_ | t_1__109_;
  assign t_2__106_ = t_1__106_ | t_1__108_;
  assign t_2__105_ = t_1__105_ | t_1__107_;
  assign t_2__104_ = t_1__104_ | t_1__106_;
  assign t_2__103_ = t_1__103_ | t_1__105_;
  assign t_2__102_ = t_1__102_ | t_1__104_;
  assign t_2__101_ = t_1__101_ | t_1__103_;
  assign t_2__100_ = t_1__100_ | t_1__102_;
  assign t_2__99_ = t_1__99_ | t_1__101_;
  assign t_2__98_ = t_1__98_ | t_1__100_;
  assign t_2__97_ = t_1__97_ | t_1__99_;
  assign t_2__96_ = t_1__96_ | t_1__98_;
  assign t_2__95_ = t_1__95_ | t_1__97_;
  assign t_2__94_ = t_1__94_ | t_1__96_;
  assign t_2__93_ = t_1__93_ | t_1__95_;
  assign t_2__92_ = t_1__92_ | t_1__94_;
  assign t_2__91_ = t_1__91_ | t_1__93_;
  assign t_2__90_ = t_1__90_ | t_1__92_;
  assign t_2__89_ = t_1__89_ | t_1__91_;
  assign t_2__88_ = t_1__88_ | t_1__90_;
  assign t_2__87_ = t_1__87_ | t_1__89_;
  assign t_2__86_ = t_1__86_ | t_1__88_;
  assign t_2__85_ = t_1__85_ | t_1__87_;
  assign t_2__84_ = t_1__84_ | t_1__86_;
  assign t_2__83_ = t_1__83_ | t_1__85_;
  assign t_2__82_ = t_1__82_ | t_1__84_;
  assign t_2__81_ = t_1__81_ | t_1__83_;
  assign t_2__80_ = t_1__80_ | t_1__82_;
  assign t_2__79_ = t_1__79_ | t_1__81_;
  assign t_2__78_ = t_1__78_ | t_1__80_;
  assign t_2__77_ = t_1__77_ | t_1__79_;
  assign t_2__76_ = t_1__76_ | t_1__78_;
  assign t_2__75_ = t_1__75_ | t_1__77_;
  assign t_2__74_ = t_1__74_ | t_1__76_;
  assign t_2__73_ = t_1__73_ | t_1__75_;
  assign t_2__72_ = t_1__72_ | t_1__74_;
  assign t_2__71_ = t_1__71_ | t_1__73_;
  assign t_2__70_ = t_1__70_ | t_1__72_;
  assign t_2__69_ = t_1__69_ | t_1__71_;
  assign t_2__68_ = t_1__68_ | t_1__70_;
  assign t_2__67_ = t_1__67_ | t_1__69_;
  assign t_2__66_ = t_1__66_ | t_1__68_;
  assign t_2__65_ = t_1__65_ | t_1__67_;
  assign t_2__64_ = t_1__64_ | t_1__66_;
  assign t_2__63_ = t_1__63_ | t_1__65_;
  assign t_2__62_ = t_1__62_ | t_1__64_;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__114_ = t_2__114_ | 1'b0;
  assign t_3__113_ = t_2__113_ | 1'b0;
  assign t_3__112_ = t_2__112_ | 1'b0;
  assign t_3__111_ = t_2__111_ | 1'b0;
  assign t_3__110_ = t_2__110_ | t_2__114_;
  assign t_3__109_ = t_2__109_ | t_2__113_;
  assign t_3__108_ = t_2__108_ | t_2__112_;
  assign t_3__107_ = t_2__107_ | t_2__111_;
  assign t_3__106_ = t_2__106_ | t_2__110_;
  assign t_3__105_ = t_2__105_ | t_2__109_;
  assign t_3__104_ = t_2__104_ | t_2__108_;
  assign t_3__103_ = t_2__103_ | t_2__107_;
  assign t_3__102_ = t_2__102_ | t_2__106_;
  assign t_3__101_ = t_2__101_ | t_2__105_;
  assign t_3__100_ = t_2__100_ | t_2__104_;
  assign t_3__99_ = t_2__99_ | t_2__103_;
  assign t_3__98_ = t_2__98_ | t_2__102_;
  assign t_3__97_ = t_2__97_ | t_2__101_;
  assign t_3__96_ = t_2__96_ | t_2__100_;
  assign t_3__95_ = t_2__95_ | t_2__99_;
  assign t_3__94_ = t_2__94_ | t_2__98_;
  assign t_3__93_ = t_2__93_ | t_2__97_;
  assign t_3__92_ = t_2__92_ | t_2__96_;
  assign t_3__91_ = t_2__91_ | t_2__95_;
  assign t_3__90_ = t_2__90_ | t_2__94_;
  assign t_3__89_ = t_2__89_ | t_2__93_;
  assign t_3__88_ = t_2__88_ | t_2__92_;
  assign t_3__87_ = t_2__87_ | t_2__91_;
  assign t_3__86_ = t_2__86_ | t_2__90_;
  assign t_3__85_ = t_2__85_ | t_2__89_;
  assign t_3__84_ = t_2__84_ | t_2__88_;
  assign t_3__83_ = t_2__83_ | t_2__87_;
  assign t_3__82_ = t_2__82_ | t_2__86_;
  assign t_3__81_ = t_2__81_ | t_2__85_;
  assign t_3__80_ = t_2__80_ | t_2__84_;
  assign t_3__79_ = t_2__79_ | t_2__83_;
  assign t_3__78_ = t_2__78_ | t_2__82_;
  assign t_3__77_ = t_2__77_ | t_2__81_;
  assign t_3__76_ = t_2__76_ | t_2__80_;
  assign t_3__75_ = t_2__75_ | t_2__79_;
  assign t_3__74_ = t_2__74_ | t_2__78_;
  assign t_3__73_ = t_2__73_ | t_2__77_;
  assign t_3__72_ = t_2__72_ | t_2__76_;
  assign t_3__71_ = t_2__71_ | t_2__75_;
  assign t_3__70_ = t_2__70_ | t_2__74_;
  assign t_3__69_ = t_2__69_ | t_2__73_;
  assign t_3__68_ = t_2__68_ | t_2__72_;
  assign t_3__67_ = t_2__67_ | t_2__71_;
  assign t_3__66_ = t_2__66_ | t_2__70_;
  assign t_3__65_ = t_2__65_ | t_2__69_;
  assign t_3__64_ = t_2__64_ | t_2__68_;
  assign t_3__63_ = t_2__63_ | t_2__67_;
  assign t_3__62_ = t_2__62_ | t_2__66_;
  assign t_3__61_ = t_2__61_ | t_2__65_;
  assign t_3__60_ = t_2__60_ | t_2__64_;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__114_ = t_3__114_ | 1'b0;
  assign t_4__113_ = t_3__113_ | 1'b0;
  assign t_4__112_ = t_3__112_ | 1'b0;
  assign t_4__111_ = t_3__111_ | 1'b0;
  assign t_4__110_ = t_3__110_ | 1'b0;
  assign t_4__109_ = t_3__109_ | 1'b0;
  assign t_4__108_ = t_3__108_ | 1'b0;
  assign t_4__107_ = t_3__107_ | 1'b0;
  assign t_4__106_ = t_3__106_ | t_3__114_;
  assign t_4__105_ = t_3__105_ | t_3__113_;
  assign t_4__104_ = t_3__104_ | t_3__112_;
  assign t_4__103_ = t_3__103_ | t_3__111_;
  assign t_4__102_ = t_3__102_ | t_3__110_;
  assign t_4__101_ = t_3__101_ | t_3__109_;
  assign t_4__100_ = t_3__100_ | t_3__108_;
  assign t_4__99_ = t_3__99_ | t_3__107_;
  assign t_4__98_ = t_3__98_ | t_3__106_;
  assign t_4__97_ = t_3__97_ | t_3__105_;
  assign t_4__96_ = t_3__96_ | t_3__104_;
  assign t_4__95_ = t_3__95_ | t_3__103_;
  assign t_4__94_ = t_3__94_ | t_3__102_;
  assign t_4__93_ = t_3__93_ | t_3__101_;
  assign t_4__92_ = t_3__92_ | t_3__100_;
  assign t_4__91_ = t_3__91_ | t_3__99_;
  assign t_4__90_ = t_3__90_ | t_3__98_;
  assign t_4__89_ = t_3__89_ | t_3__97_;
  assign t_4__88_ = t_3__88_ | t_3__96_;
  assign t_4__87_ = t_3__87_ | t_3__95_;
  assign t_4__86_ = t_3__86_ | t_3__94_;
  assign t_4__85_ = t_3__85_ | t_3__93_;
  assign t_4__84_ = t_3__84_ | t_3__92_;
  assign t_4__83_ = t_3__83_ | t_3__91_;
  assign t_4__82_ = t_3__82_ | t_3__90_;
  assign t_4__81_ = t_3__81_ | t_3__89_;
  assign t_4__80_ = t_3__80_ | t_3__88_;
  assign t_4__79_ = t_3__79_ | t_3__87_;
  assign t_4__78_ = t_3__78_ | t_3__86_;
  assign t_4__77_ = t_3__77_ | t_3__85_;
  assign t_4__76_ = t_3__76_ | t_3__84_;
  assign t_4__75_ = t_3__75_ | t_3__83_;
  assign t_4__74_ = t_3__74_ | t_3__82_;
  assign t_4__73_ = t_3__73_ | t_3__81_;
  assign t_4__72_ = t_3__72_ | t_3__80_;
  assign t_4__71_ = t_3__71_ | t_3__79_;
  assign t_4__70_ = t_3__70_ | t_3__78_;
  assign t_4__69_ = t_3__69_ | t_3__77_;
  assign t_4__68_ = t_3__68_ | t_3__76_;
  assign t_4__67_ = t_3__67_ | t_3__75_;
  assign t_4__66_ = t_3__66_ | t_3__74_;
  assign t_4__65_ = t_3__65_ | t_3__73_;
  assign t_4__64_ = t_3__64_ | t_3__72_;
  assign t_4__63_ = t_3__63_ | t_3__71_;
  assign t_4__62_ = t_3__62_ | t_3__70_;
  assign t_4__61_ = t_3__61_ | t_3__69_;
  assign t_4__60_ = t_3__60_ | t_3__68_;
  assign t_4__59_ = t_3__59_ | t_3__67_;
  assign t_4__58_ = t_3__58_ | t_3__66_;
  assign t_4__57_ = t_3__57_ | t_3__65_;
  assign t_4__56_ = t_3__56_ | t_3__64_;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__114_ = t_4__114_ | 1'b0;
  assign t_5__113_ = t_4__113_ | 1'b0;
  assign t_5__112_ = t_4__112_ | 1'b0;
  assign t_5__111_ = t_4__111_ | 1'b0;
  assign t_5__110_ = t_4__110_ | 1'b0;
  assign t_5__109_ = t_4__109_ | 1'b0;
  assign t_5__108_ = t_4__108_ | 1'b0;
  assign t_5__107_ = t_4__107_ | 1'b0;
  assign t_5__106_ = t_4__106_ | 1'b0;
  assign t_5__105_ = t_4__105_ | 1'b0;
  assign t_5__104_ = t_4__104_ | 1'b0;
  assign t_5__103_ = t_4__103_ | 1'b0;
  assign t_5__102_ = t_4__102_ | 1'b0;
  assign t_5__101_ = t_4__101_ | 1'b0;
  assign t_5__100_ = t_4__100_ | 1'b0;
  assign t_5__99_ = t_4__99_ | 1'b0;
  assign t_5__98_ = t_4__98_ | t_4__114_;
  assign t_5__97_ = t_4__97_ | t_4__113_;
  assign t_5__96_ = t_4__96_ | t_4__112_;
  assign t_5__95_ = t_4__95_ | t_4__111_;
  assign t_5__94_ = t_4__94_ | t_4__110_;
  assign t_5__93_ = t_4__93_ | t_4__109_;
  assign t_5__92_ = t_4__92_ | t_4__108_;
  assign t_5__91_ = t_4__91_ | t_4__107_;
  assign t_5__90_ = t_4__90_ | t_4__106_;
  assign t_5__89_ = t_4__89_ | t_4__105_;
  assign t_5__88_ = t_4__88_ | t_4__104_;
  assign t_5__87_ = t_4__87_ | t_4__103_;
  assign t_5__86_ = t_4__86_ | t_4__102_;
  assign t_5__85_ = t_4__85_ | t_4__101_;
  assign t_5__84_ = t_4__84_ | t_4__100_;
  assign t_5__83_ = t_4__83_ | t_4__99_;
  assign t_5__82_ = t_4__82_ | t_4__98_;
  assign t_5__81_ = t_4__81_ | t_4__97_;
  assign t_5__80_ = t_4__80_ | t_4__96_;
  assign t_5__79_ = t_4__79_ | t_4__95_;
  assign t_5__78_ = t_4__78_ | t_4__94_;
  assign t_5__77_ = t_4__77_ | t_4__93_;
  assign t_5__76_ = t_4__76_ | t_4__92_;
  assign t_5__75_ = t_4__75_ | t_4__91_;
  assign t_5__74_ = t_4__74_ | t_4__90_;
  assign t_5__73_ = t_4__73_ | t_4__89_;
  assign t_5__72_ = t_4__72_ | t_4__88_;
  assign t_5__71_ = t_4__71_ | t_4__87_;
  assign t_5__70_ = t_4__70_ | t_4__86_;
  assign t_5__69_ = t_4__69_ | t_4__85_;
  assign t_5__68_ = t_4__68_ | t_4__84_;
  assign t_5__67_ = t_4__67_ | t_4__83_;
  assign t_5__66_ = t_4__66_ | t_4__82_;
  assign t_5__65_ = t_4__65_ | t_4__81_;
  assign t_5__64_ = t_4__64_ | t_4__80_;
  assign t_5__63_ = t_4__63_ | t_4__79_;
  assign t_5__62_ = t_4__62_ | t_4__78_;
  assign t_5__61_ = t_4__61_ | t_4__77_;
  assign t_5__60_ = t_4__60_ | t_4__76_;
  assign t_5__59_ = t_4__59_ | t_4__75_;
  assign t_5__58_ = t_4__58_ | t_4__74_;
  assign t_5__57_ = t_4__57_ | t_4__73_;
  assign t_5__56_ = t_4__56_ | t_4__72_;
  assign t_5__55_ = t_4__55_ | t_4__71_;
  assign t_5__54_ = t_4__54_ | t_4__70_;
  assign t_5__53_ = t_4__53_ | t_4__69_;
  assign t_5__52_ = t_4__52_ | t_4__68_;
  assign t_5__51_ = t_4__51_ | t_4__67_;
  assign t_5__50_ = t_4__50_ | t_4__66_;
  assign t_5__49_ = t_4__49_ | t_4__65_;
  assign t_5__48_ = t_4__48_ | t_4__64_;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign t_6__114_ = t_5__114_ | 1'b0;
  assign t_6__113_ = t_5__113_ | 1'b0;
  assign t_6__112_ = t_5__112_ | 1'b0;
  assign t_6__111_ = t_5__111_ | 1'b0;
  assign t_6__110_ = t_5__110_ | 1'b0;
  assign t_6__109_ = t_5__109_ | 1'b0;
  assign t_6__108_ = t_5__108_ | 1'b0;
  assign t_6__107_ = t_5__107_ | 1'b0;
  assign t_6__106_ = t_5__106_ | 1'b0;
  assign t_6__105_ = t_5__105_ | 1'b0;
  assign t_6__104_ = t_5__104_ | 1'b0;
  assign t_6__103_ = t_5__103_ | 1'b0;
  assign t_6__102_ = t_5__102_ | 1'b0;
  assign t_6__101_ = t_5__101_ | 1'b0;
  assign t_6__100_ = t_5__100_ | 1'b0;
  assign t_6__99_ = t_5__99_ | 1'b0;
  assign t_6__98_ = t_5__98_ | 1'b0;
  assign t_6__97_ = t_5__97_ | 1'b0;
  assign t_6__96_ = t_5__96_ | 1'b0;
  assign t_6__95_ = t_5__95_ | 1'b0;
  assign t_6__94_ = t_5__94_ | 1'b0;
  assign t_6__93_ = t_5__93_ | 1'b0;
  assign t_6__92_ = t_5__92_ | 1'b0;
  assign t_6__91_ = t_5__91_ | 1'b0;
  assign t_6__90_ = t_5__90_ | 1'b0;
  assign t_6__89_ = t_5__89_ | 1'b0;
  assign t_6__88_ = t_5__88_ | 1'b0;
  assign t_6__87_ = t_5__87_ | 1'b0;
  assign t_6__86_ = t_5__86_ | 1'b0;
  assign t_6__85_ = t_5__85_ | 1'b0;
  assign t_6__84_ = t_5__84_ | 1'b0;
  assign t_6__83_ = t_5__83_ | 1'b0;
  assign t_6__82_ = t_5__82_ | t_5__114_;
  assign t_6__81_ = t_5__81_ | t_5__113_;
  assign t_6__80_ = t_5__80_ | t_5__112_;
  assign t_6__79_ = t_5__79_ | t_5__111_;
  assign t_6__78_ = t_5__78_ | t_5__110_;
  assign t_6__77_ = t_5__77_ | t_5__109_;
  assign t_6__76_ = t_5__76_ | t_5__108_;
  assign t_6__75_ = t_5__75_ | t_5__107_;
  assign t_6__74_ = t_5__74_ | t_5__106_;
  assign t_6__73_ = t_5__73_ | t_5__105_;
  assign t_6__72_ = t_5__72_ | t_5__104_;
  assign t_6__71_ = t_5__71_ | t_5__103_;
  assign t_6__70_ = t_5__70_ | t_5__102_;
  assign t_6__69_ = t_5__69_ | t_5__101_;
  assign t_6__68_ = t_5__68_ | t_5__100_;
  assign t_6__67_ = t_5__67_ | t_5__99_;
  assign t_6__66_ = t_5__66_ | t_5__98_;
  assign t_6__65_ = t_5__65_ | t_5__97_;
  assign t_6__64_ = t_5__64_ | t_5__96_;
  assign t_6__63_ = t_5__63_ | t_5__95_;
  assign t_6__62_ = t_5__62_ | t_5__94_;
  assign t_6__61_ = t_5__61_ | t_5__93_;
  assign t_6__60_ = t_5__60_ | t_5__92_;
  assign t_6__59_ = t_5__59_ | t_5__91_;
  assign t_6__58_ = t_5__58_ | t_5__90_;
  assign t_6__57_ = t_5__57_ | t_5__89_;
  assign t_6__56_ = t_5__56_ | t_5__88_;
  assign t_6__55_ = t_5__55_ | t_5__87_;
  assign t_6__54_ = t_5__54_ | t_5__86_;
  assign t_6__53_ = t_5__53_ | t_5__85_;
  assign t_6__52_ = t_5__52_ | t_5__84_;
  assign t_6__51_ = t_5__51_ | t_5__83_;
  assign t_6__50_ = t_5__50_ | t_5__82_;
  assign t_6__49_ = t_5__49_ | t_5__81_;
  assign t_6__48_ = t_5__48_ | t_5__80_;
  assign t_6__47_ = t_5__47_ | t_5__79_;
  assign t_6__46_ = t_5__46_ | t_5__78_;
  assign t_6__45_ = t_5__45_ | t_5__77_;
  assign t_6__44_ = t_5__44_ | t_5__76_;
  assign t_6__43_ = t_5__43_ | t_5__75_;
  assign t_6__42_ = t_5__42_ | t_5__74_;
  assign t_6__41_ = t_5__41_ | t_5__73_;
  assign t_6__40_ = t_5__40_ | t_5__72_;
  assign t_6__39_ = t_5__39_ | t_5__71_;
  assign t_6__38_ = t_5__38_ | t_5__70_;
  assign t_6__37_ = t_5__37_ | t_5__69_;
  assign t_6__36_ = t_5__36_ | t_5__68_;
  assign t_6__35_ = t_5__35_ | t_5__67_;
  assign t_6__34_ = t_5__34_ | t_5__66_;
  assign t_6__33_ = t_5__33_ | t_5__65_;
  assign t_6__32_ = t_5__32_ | t_5__64_;
  assign t_6__31_ = t_5__31_ | t_5__63_;
  assign t_6__30_ = t_5__30_ | t_5__62_;
  assign t_6__29_ = t_5__29_ | t_5__61_;
  assign t_6__28_ = t_5__28_ | t_5__60_;
  assign t_6__27_ = t_5__27_ | t_5__59_;
  assign t_6__26_ = t_5__26_ | t_5__58_;
  assign t_6__25_ = t_5__25_ | t_5__57_;
  assign t_6__24_ = t_5__24_ | t_5__56_;
  assign t_6__23_ = t_5__23_ | t_5__55_;
  assign t_6__22_ = t_5__22_ | t_5__54_;
  assign t_6__21_ = t_5__21_ | t_5__53_;
  assign t_6__20_ = t_5__20_ | t_5__52_;
  assign t_6__19_ = t_5__19_ | t_5__51_;
  assign t_6__18_ = t_5__18_ | t_5__50_;
  assign t_6__17_ = t_5__17_ | t_5__49_;
  assign t_6__16_ = t_5__16_ | t_5__48_;
  assign t_6__15_ = t_5__15_ | t_5__47_;
  assign t_6__14_ = t_5__14_ | t_5__46_;
  assign t_6__13_ = t_5__13_ | t_5__45_;
  assign t_6__12_ = t_5__12_ | t_5__44_;
  assign t_6__11_ = t_5__11_ | t_5__43_;
  assign t_6__10_ = t_5__10_ | t_5__42_;
  assign t_6__9_ = t_5__9_ | t_5__41_;
  assign t_6__8_ = t_5__8_ | t_5__40_;
  assign t_6__7_ = t_5__7_ | t_5__39_;
  assign t_6__6_ = t_5__6_ | t_5__38_;
  assign t_6__5_ = t_5__5_ | t_5__37_;
  assign t_6__4_ = t_5__4_ | t_5__36_;
  assign t_6__3_ = t_5__3_ | t_5__35_;
  assign t_6__2_ = t_5__2_ | t_5__34_;
  assign t_6__1_ = t_5__1_ | t_5__33_;
  assign t_6__0_ = t_5__0_ | t_5__32_;
  assign o[0] = t_6__114_ | 1'b0;
  assign o[1] = t_6__113_ | 1'b0;
  assign o[2] = t_6__112_ | 1'b0;
  assign o[3] = t_6__111_ | 1'b0;
  assign o[4] = t_6__110_ | 1'b0;
  assign o[5] = t_6__109_ | 1'b0;
  assign o[6] = t_6__108_ | 1'b0;
  assign o[7] = t_6__107_ | 1'b0;
  assign o[8] = t_6__106_ | 1'b0;
  assign o[9] = t_6__105_ | 1'b0;
  assign o[10] = t_6__104_ | 1'b0;
  assign o[11] = t_6__103_ | 1'b0;
  assign o[12] = t_6__102_ | 1'b0;
  assign o[13] = t_6__101_ | 1'b0;
  assign o[14] = t_6__100_ | 1'b0;
  assign o[15] = t_6__99_ | 1'b0;
  assign o[16] = t_6__98_ | 1'b0;
  assign o[17] = t_6__97_ | 1'b0;
  assign o[18] = t_6__96_ | 1'b0;
  assign o[19] = t_6__95_ | 1'b0;
  assign o[20] = t_6__94_ | 1'b0;
  assign o[21] = t_6__93_ | 1'b0;
  assign o[22] = t_6__92_ | 1'b0;
  assign o[23] = t_6__91_ | 1'b0;
  assign o[24] = t_6__90_ | 1'b0;
  assign o[25] = t_6__89_ | 1'b0;
  assign o[26] = t_6__88_ | 1'b0;
  assign o[27] = t_6__87_ | 1'b0;
  assign o[28] = t_6__86_ | 1'b0;
  assign o[29] = t_6__85_ | 1'b0;
  assign o[30] = t_6__84_ | 1'b0;
  assign o[31] = t_6__83_ | 1'b0;
  assign o[32] = t_6__82_ | 1'b0;
  assign o[33] = t_6__81_ | 1'b0;
  assign o[34] = t_6__80_ | 1'b0;
  assign o[35] = t_6__79_ | 1'b0;
  assign o[36] = t_6__78_ | 1'b0;
  assign o[37] = t_6__77_ | 1'b0;
  assign o[38] = t_6__76_ | 1'b0;
  assign o[39] = t_6__75_ | 1'b0;
  assign o[40] = t_6__74_ | 1'b0;
  assign o[41] = t_6__73_ | 1'b0;
  assign o[42] = t_6__72_ | 1'b0;
  assign o[43] = t_6__71_ | 1'b0;
  assign o[44] = t_6__70_ | 1'b0;
  assign o[45] = t_6__69_ | 1'b0;
  assign o[46] = t_6__68_ | 1'b0;
  assign o[47] = t_6__67_ | 1'b0;
  assign o[48] = t_6__66_ | 1'b0;
  assign o[49] = t_6__65_ | 1'b0;
  assign o[50] = t_6__64_ | 1'b0;
  assign o[51] = t_6__63_ | 1'b0;
  assign o[52] = t_6__62_ | 1'b0;
  assign o[53] = t_6__61_ | 1'b0;
  assign o[54] = t_6__60_ | 1'b0;
  assign o[55] = t_6__59_ | 1'b0;
  assign o[56] = t_6__58_ | 1'b0;
  assign o[57] = t_6__57_ | 1'b0;
  assign o[58] = t_6__56_ | 1'b0;
  assign o[59] = t_6__55_ | 1'b0;
  assign o[60] = t_6__54_ | 1'b0;
  assign o[61] = t_6__53_ | 1'b0;
  assign o[62] = t_6__52_ | 1'b0;
  assign o[63] = t_6__51_ | 1'b0;
  assign o[64] = t_6__50_ | t_6__114_;
  assign o[65] = t_6__49_ | t_6__113_;
  assign o[66] = t_6__48_ | t_6__112_;
  assign o[67] = t_6__47_ | t_6__111_;
  assign o[68] = t_6__46_ | t_6__110_;
  assign o[69] = t_6__45_ | t_6__109_;
  assign o[70] = t_6__44_ | t_6__108_;
  assign o[71] = t_6__43_ | t_6__107_;
  assign o[72] = t_6__42_ | t_6__106_;
  assign o[73] = t_6__41_ | t_6__105_;
  assign o[74] = t_6__40_ | t_6__104_;
  assign o[75] = t_6__39_ | t_6__103_;
  assign o[76] = t_6__38_ | t_6__102_;
  assign o[77] = t_6__37_ | t_6__101_;
  assign o[78] = t_6__36_ | t_6__100_;
  assign o[79] = t_6__35_ | t_6__99_;
  assign o[80] = t_6__34_ | t_6__98_;
  assign o[81] = t_6__33_ | t_6__97_;
  assign o[82] = t_6__32_ | t_6__96_;
  assign o[83] = t_6__31_ | t_6__95_;
  assign o[84] = t_6__30_ | t_6__94_;
  assign o[85] = t_6__29_ | t_6__93_;
  assign o[86] = t_6__28_ | t_6__92_;
  assign o[87] = t_6__27_ | t_6__91_;
  assign o[88] = t_6__26_ | t_6__90_;
  assign o[89] = t_6__25_ | t_6__89_;
  assign o[90] = t_6__24_ | t_6__88_;
  assign o[91] = t_6__23_ | t_6__87_;
  assign o[92] = t_6__22_ | t_6__86_;
  assign o[93] = t_6__21_ | t_6__85_;
  assign o[94] = t_6__20_ | t_6__84_;
  assign o[95] = t_6__19_ | t_6__83_;
  assign o[96] = t_6__18_ | t_6__82_;
  assign o[97] = t_6__17_ | t_6__81_;
  assign o[98] = t_6__16_ | t_6__80_;
  assign o[99] = t_6__15_ | t_6__79_;
  assign o[100] = t_6__14_ | t_6__78_;
  assign o[101] = t_6__13_ | t_6__77_;
  assign o[102] = t_6__12_ | t_6__76_;
  assign o[103] = t_6__11_ | t_6__75_;
  assign o[104] = t_6__10_ | t_6__74_;
  assign o[105] = t_6__9_ | t_6__73_;
  assign o[106] = t_6__8_ | t_6__72_;
  assign o[107] = t_6__7_ | t_6__71_;
  assign o[108] = t_6__6_ | t_6__70_;
  assign o[109] = t_6__5_ | t_6__69_;
  assign o[110] = t_6__4_ | t_6__68_;
  assign o[111] = t_6__3_ | t_6__67_;
  assign o[112] = t_6__2_ | t_6__66_;
  assign o[113] = t_6__1_ | t_6__65_;
  assign o[114] = t_6__0_ | t_6__64_;

endmodule



module bsg_fpu_sticky_width_p115
(
  i,
  shamt_i,
  sticky_o
);

  input [114:0] i;
  input [6:0] shamt_i;
  output sticky_o;
  wire sticky_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,
  N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
  N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,
  N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,
  N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,
  N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,
  N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,
  N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
  N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,
  N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,
  N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
  N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,
  N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,
  N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,
  N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,
  N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,
  N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,
  N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143;
  wire [114:0] scan_out;

  bsg_scan_width_p115_or_p1_lo_to_hi_p1
  scan0
  (
    .i(i),
    .o(scan_out)
  );

  assign N1025 = shamt_i > { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 };
  assign N0 = N5 & N6;
  assign N1 = N0 & N7;
  assign N2 = N1 & N8;
  assign N3 = N2 & N9;
  assign N4 = N3 & N10;
  assign N1027 = N4 & N11;
  assign N5 = ~shamt_i[6];
  assign N6 = ~shamt_i[5];
  assign N7 = ~shamt_i[4];
  assign N8 = ~shamt_i[3];
  assign N9 = ~shamt_i[2];
  assign N10 = ~shamt_i[0];
  assign N11 = ~shamt_i[1];
  assign N12 = shamt_i[6] & N17;
  assign N13 = N12 & N18;
  assign N14 = N13 & N19;
  assign N15 = N14 & N20;
  assign N16 = N15 & N21;
  assign N1028 = N16 & N22;
  assign N17 = ~shamt_i[5];
  assign N18 = ~shamt_i[4];
  assign N19 = ~shamt_i[3];
  assign N20 = ~shamt_i[2];
  assign N21 = ~shamt_i[0];
  assign N22 = ~shamt_i[1];
  assign N23 = N28 & N29;
  assign N24 = N23 & N30;
  assign N25 = N24 & N31;
  assign N26 = N25 & N32;
  assign N27 = N26 & shamt_i[0];
  assign N1029 = N27 & N33;
  assign N28 = ~shamt_i[6];
  assign N29 = ~shamt_i[5];
  assign N30 = ~shamt_i[4];
  assign N31 = ~shamt_i[3];
  assign N32 = ~shamt_i[2];
  assign N33 = ~shamt_i[1];
  assign N34 = N39 & N40;
  assign N35 = N34 & N41;
  assign N36 = N35 & N42;
  assign N37 = N36 & N43;
  assign N38 = N37 & N44;
  assign N1031 = N38 & shamt_i[1];
  assign N39 = ~shamt_i[6];
  assign N40 = ~shamt_i[5];
  assign N41 = ~shamt_i[4];
  assign N42 = ~shamt_i[3];
  assign N43 = ~shamt_i[2];
  assign N44 = ~shamt_i[0];
  assign N45 = N50 & N51;
  assign N46 = N45 & N52;
  assign N47 = N46 & N53;
  assign N48 = N47 & N54;
  assign N49 = N48 & shamt_i[0];
  assign N1033 = N49 & shamt_i[1];
  assign N50 = ~shamt_i[6];
  assign N51 = ~shamt_i[5];
  assign N52 = ~shamt_i[4];
  assign N53 = ~shamt_i[3];
  assign N54 = ~shamt_i[2];
  assign N55 = N60 & N61;
  assign N56 = N55 & N62;
  assign N57 = N56 & N63;
  assign N58 = N57 & shamt_i[2];
  assign N59 = N58 & N64;
  assign N1035 = N59 & N65;
  assign N60 = ~shamt_i[6];
  assign N61 = ~shamt_i[5];
  assign N62 = ~shamt_i[4];
  assign N63 = ~shamt_i[3];
  assign N64 = ~shamt_i[0];
  assign N65 = ~shamt_i[1];
  assign N66 = N71 & N72;
  assign N67 = N66 & N73;
  assign N68 = N67 & N74;
  assign N69 = N68 & shamt_i[2];
  assign N70 = N69 & shamt_i[0];
  assign N1037 = N70 & N75;
  assign N71 = ~shamt_i[6];
  assign N72 = ~shamt_i[5];
  assign N73 = ~shamt_i[4];
  assign N74 = ~shamt_i[3];
  assign N75 = ~shamt_i[1];
  assign N76 = N81 & N82;
  assign N77 = N76 & N83;
  assign N78 = N77 & N84;
  assign N79 = N78 & shamt_i[2];
  assign N80 = N79 & N85;
  assign N1039 = N80 & shamt_i[1];
  assign N81 = ~shamt_i[6];
  assign N82 = ~shamt_i[5];
  assign N83 = ~shamt_i[4];
  assign N84 = ~shamt_i[3];
  assign N85 = ~shamt_i[0];
  assign N86 = N91 & N92;
  assign N87 = N86 & N93;
  assign N88 = N87 & N94;
  assign N89 = N88 & shamt_i[2];
  assign N90 = N89 & shamt_i[0];
  assign N1041 = N90 & shamt_i[1];
  assign N91 = ~shamt_i[6];
  assign N92 = ~shamt_i[5];
  assign N93 = ~shamt_i[4];
  assign N94 = ~shamt_i[3];
  assign N95 = N100 & N101;
  assign N96 = N95 & N102;
  assign N97 = N96 & shamt_i[3];
  assign N98 = N97 & N103;
  assign N99 = N98 & N104;
  assign N1043 = N99 & N105;
  assign N100 = ~shamt_i[6];
  assign N101 = ~shamt_i[5];
  assign N102 = ~shamt_i[4];
  assign N103 = ~shamt_i[2];
  assign N104 = ~shamt_i[0];
  assign N105 = ~shamt_i[1];
  assign N106 = N111 & N112;
  assign N107 = N106 & N113;
  assign N108 = N107 & shamt_i[3];
  assign N109 = N108 & N114;
  assign N110 = N109 & shamt_i[0];
  assign N1045 = N110 & N115;
  assign N111 = ~shamt_i[6];
  assign N112 = ~shamt_i[5];
  assign N113 = ~shamt_i[4];
  assign N114 = ~shamt_i[2];
  assign N115 = ~shamt_i[1];
  assign N116 = N121 & N122;
  assign N117 = N116 & N123;
  assign N118 = N117 & shamt_i[3];
  assign N119 = N118 & N124;
  assign N120 = N119 & N125;
  assign N1047 = N120 & shamt_i[1];
  assign N121 = ~shamt_i[6];
  assign N122 = ~shamt_i[5];
  assign N123 = ~shamt_i[4];
  assign N124 = ~shamt_i[2];
  assign N125 = ~shamt_i[0];
  assign N126 = N131 & N132;
  assign N127 = N126 & N133;
  assign N128 = N127 & shamt_i[3];
  assign N129 = N128 & N134;
  assign N130 = N129 & shamt_i[0];
  assign N1049 = N130 & shamt_i[1];
  assign N131 = ~shamt_i[6];
  assign N132 = ~shamt_i[5];
  assign N133 = ~shamt_i[4];
  assign N134 = ~shamt_i[2];
  assign N135 = N140 & N141;
  assign N136 = N135 & N142;
  assign N137 = N136 & shamt_i[3];
  assign N138 = N137 & shamt_i[2];
  assign N139 = N138 & N143;
  assign N1051 = N139 & N144;
  assign N140 = ~shamt_i[6];
  assign N141 = ~shamt_i[5];
  assign N142 = ~shamt_i[4];
  assign N143 = ~shamt_i[0];
  assign N144 = ~shamt_i[1];
  assign N145 = N150 & N151;
  assign N146 = N145 & N152;
  assign N147 = N146 & shamt_i[3];
  assign N148 = N147 & shamt_i[2];
  assign N149 = N148 & shamt_i[0];
  assign N1053 = N149 & N153;
  assign N150 = ~shamt_i[6];
  assign N151 = ~shamt_i[5];
  assign N152 = ~shamt_i[4];
  assign N153 = ~shamt_i[1];
  assign N154 = N159 & N160;
  assign N155 = N154 & N161;
  assign N156 = N155 & shamt_i[3];
  assign N157 = N156 & shamt_i[2];
  assign N158 = N157 & N162;
  assign N1055 = N158 & shamt_i[1];
  assign N159 = ~shamt_i[6];
  assign N160 = ~shamt_i[5];
  assign N161 = ~shamt_i[4];
  assign N162 = ~shamt_i[0];
  assign N163 = N168 & N169;
  assign N164 = N163 & N170;
  assign N165 = N164 & shamt_i[3];
  assign N166 = N165 & shamt_i[2];
  assign N167 = N166 & shamt_i[0];
  assign N1057 = N167 & shamt_i[1];
  assign N168 = ~shamt_i[6];
  assign N169 = ~shamt_i[5];
  assign N170 = ~shamt_i[4];
  assign N171 = N176 & N177;
  assign N172 = N171 & shamt_i[4];
  assign N173 = N172 & N178;
  assign N174 = N173 & N179;
  assign N175 = N174 & N180;
  assign N1059 = N175 & N181;
  assign N176 = ~shamt_i[6];
  assign N177 = ~shamt_i[5];
  assign N178 = ~shamt_i[3];
  assign N179 = ~shamt_i[2];
  assign N180 = ~shamt_i[0];
  assign N181 = ~shamt_i[1];
  assign N182 = N187 & N188;
  assign N183 = N182 & shamt_i[4];
  assign N184 = N183 & N189;
  assign N185 = N184 & N190;
  assign N186 = N185 & shamt_i[0];
  assign N1061 = N186 & N191;
  assign N187 = ~shamt_i[6];
  assign N188 = ~shamt_i[5];
  assign N189 = ~shamt_i[3];
  assign N190 = ~shamt_i[2];
  assign N191 = ~shamt_i[1];
  assign N192 = N197 & N198;
  assign N193 = N192 & shamt_i[4];
  assign N194 = N193 & N199;
  assign N195 = N194 & N200;
  assign N196 = N195 & N201;
  assign N1063 = N196 & shamt_i[1];
  assign N197 = ~shamt_i[6];
  assign N198 = ~shamt_i[5];
  assign N199 = ~shamt_i[3];
  assign N200 = ~shamt_i[2];
  assign N201 = ~shamt_i[0];
  assign N202 = N207 & N208;
  assign N203 = N202 & shamt_i[4];
  assign N204 = N203 & N209;
  assign N205 = N204 & N210;
  assign N206 = N205 & shamt_i[0];
  assign N1065 = N206 & shamt_i[1];
  assign N207 = ~shamt_i[6];
  assign N208 = ~shamt_i[5];
  assign N209 = ~shamt_i[3];
  assign N210 = ~shamt_i[2];
  assign N211 = N216 & N217;
  assign N212 = N211 & shamt_i[4];
  assign N213 = N212 & N218;
  assign N214 = N213 & shamt_i[2];
  assign N215 = N214 & N219;
  assign N1067 = N215 & N220;
  assign N216 = ~shamt_i[6];
  assign N217 = ~shamt_i[5];
  assign N218 = ~shamt_i[3];
  assign N219 = ~shamt_i[0];
  assign N220 = ~shamt_i[1];
  assign N221 = N226 & N227;
  assign N222 = N221 & shamt_i[4];
  assign N223 = N222 & N228;
  assign N224 = N223 & shamt_i[2];
  assign N225 = N224 & shamt_i[0];
  assign N1069 = N225 & N229;
  assign N226 = ~shamt_i[6];
  assign N227 = ~shamt_i[5];
  assign N228 = ~shamt_i[3];
  assign N229 = ~shamt_i[1];
  assign N230 = N235 & N236;
  assign N231 = N230 & shamt_i[4];
  assign N232 = N231 & N237;
  assign N233 = N232 & shamt_i[2];
  assign N234 = N233 & N238;
  assign N1071 = N234 & shamt_i[1];
  assign N235 = ~shamt_i[6];
  assign N236 = ~shamt_i[5];
  assign N237 = ~shamt_i[3];
  assign N238 = ~shamt_i[0];
  assign N239 = N244 & N245;
  assign N240 = N239 & shamt_i[4];
  assign N241 = N240 & N246;
  assign N242 = N241 & shamt_i[2];
  assign N243 = N242 & shamt_i[0];
  assign N1073 = N243 & shamt_i[1];
  assign N244 = ~shamt_i[6];
  assign N245 = ~shamt_i[5];
  assign N246 = ~shamt_i[3];
  assign N247 = N252 & N253;
  assign N248 = N247 & shamt_i[4];
  assign N249 = N248 & shamt_i[3];
  assign N250 = N249 & N254;
  assign N251 = N250 & N255;
  assign N1075 = N251 & N256;
  assign N252 = ~shamt_i[6];
  assign N253 = ~shamt_i[5];
  assign N254 = ~shamt_i[2];
  assign N255 = ~shamt_i[0];
  assign N256 = ~shamt_i[1];
  assign N257 = N262 & N263;
  assign N258 = N257 & shamt_i[4];
  assign N259 = N258 & shamt_i[3];
  assign N260 = N259 & N264;
  assign N261 = N260 & shamt_i[0];
  assign N1077 = N261 & N265;
  assign N262 = ~shamt_i[6];
  assign N263 = ~shamt_i[5];
  assign N264 = ~shamt_i[2];
  assign N265 = ~shamt_i[1];
  assign N266 = N271 & N272;
  assign N267 = N266 & shamt_i[4];
  assign N268 = N267 & shamt_i[3];
  assign N269 = N268 & N273;
  assign N270 = N269 & N274;
  assign N1079 = N270 & shamt_i[1];
  assign N271 = ~shamt_i[6];
  assign N272 = ~shamt_i[5];
  assign N273 = ~shamt_i[2];
  assign N274 = ~shamt_i[0];
  assign N275 = N280 & N281;
  assign N276 = N275 & shamt_i[4];
  assign N277 = N276 & shamt_i[3];
  assign N278 = N277 & N282;
  assign N279 = N278 & shamt_i[0];
  assign N1081 = N279 & shamt_i[1];
  assign N280 = ~shamt_i[6];
  assign N281 = ~shamt_i[5];
  assign N282 = ~shamt_i[2];
  assign N283 = N288 & N289;
  assign N284 = N283 & shamt_i[4];
  assign N285 = N284 & shamt_i[3];
  assign N286 = N285 & shamt_i[2];
  assign N287 = N286 & N290;
  assign N1083 = N287 & N291;
  assign N288 = ~shamt_i[6];
  assign N289 = ~shamt_i[5];
  assign N290 = ~shamt_i[0];
  assign N291 = ~shamt_i[1];
  assign N292 = N297 & N298;
  assign N293 = N292 & shamt_i[4];
  assign N294 = N293 & shamt_i[3];
  assign N295 = N294 & shamt_i[2];
  assign N296 = N295 & shamt_i[0];
  assign N1085 = N296 & N299;
  assign N297 = ~shamt_i[6];
  assign N298 = ~shamt_i[5];
  assign N299 = ~shamt_i[1];
  assign N300 = N305 & N306;
  assign N301 = N300 & shamt_i[4];
  assign N302 = N301 & shamt_i[3];
  assign N303 = N302 & shamt_i[2];
  assign N304 = N303 & N307;
  assign N1087 = N304 & shamt_i[1];
  assign N305 = ~shamt_i[6];
  assign N306 = ~shamt_i[5];
  assign N307 = ~shamt_i[0];
  assign N308 = N313 & N314;
  assign N309 = N308 & shamt_i[4];
  assign N310 = N309 & shamt_i[3];
  assign N311 = N310 & shamt_i[2];
  assign N312 = N311 & shamt_i[0];
  assign N1089 = N312 & shamt_i[1];
  assign N313 = ~shamt_i[6];
  assign N314 = ~shamt_i[5];
  assign N315 = N320 & shamt_i[5];
  assign N316 = N315 & N321;
  assign N317 = N316 & N322;
  assign N318 = N317 & N323;
  assign N319 = N318 & N324;
  assign N1091 = N319 & N325;
  assign N320 = ~shamt_i[6];
  assign N321 = ~shamt_i[4];
  assign N322 = ~shamt_i[3];
  assign N323 = ~shamt_i[2];
  assign N324 = ~shamt_i[0];
  assign N325 = ~shamt_i[1];
  assign N326 = N331 & shamt_i[5];
  assign N327 = N326 & N332;
  assign N328 = N327 & N333;
  assign N329 = N328 & N334;
  assign N330 = N329 & shamt_i[0];
  assign N1093 = N330 & N335;
  assign N331 = ~shamt_i[6];
  assign N332 = ~shamt_i[4];
  assign N333 = ~shamt_i[3];
  assign N334 = ~shamt_i[2];
  assign N335 = ~shamt_i[1];
  assign N336 = N341 & shamt_i[5];
  assign N337 = N336 & N342;
  assign N338 = N337 & N343;
  assign N339 = N338 & N344;
  assign N340 = N339 & N345;
  assign N1095 = N340 & shamt_i[1];
  assign N341 = ~shamt_i[6];
  assign N342 = ~shamt_i[4];
  assign N343 = ~shamt_i[3];
  assign N344 = ~shamt_i[2];
  assign N345 = ~shamt_i[0];
  assign N346 = N351 & shamt_i[5];
  assign N347 = N346 & N352;
  assign N348 = N347 & N353;
  assign N349 = N348 & N354;
  assign N350 = N349 & shamt_i[0];
  assign N1097 = N350 & shamt_i[1];
  assign N351 = ~shamt_i[6];
  assign N352 = ~shamt_i[4];
  assign N353 = ~shamt_i[3];
  assign N354 = ~shamt_i[2];
  assign N355 = N360 & shamt_i[5];
  assign N356 = N355 & N361;
  assign N357 = N356 & N362;
  assign N358 = N357 & shamt_i[2];
  assign N359 = N358 & N363;
  assign N1099 = N359 & N364;
  assign N360 = ~shamt_i[6];
  assign N361 = ~shamt_i[4];
  assign N362 = ~shamt_i[3];
  assign N363 = ~shamt_i[0];
  assign N364 = ~shamt_i[1];
  assign N365 = N370 & shamt_i[5];
  assign N366 = N365 & N371;
  assign N367 = N366 & N372;
  assign N368 = N367 & shamt_i[2];
  assign N369 = N368 & shamt_i[0];
  assign N1101 = N369 & N373;
  assign N370 = ~shamt_i[6];
  assign N371 = ~shamt_i[4];
  assign N372 = ~shamt_i[3];
  assign N373 = ~shamt_i[1];
  assign N374 = N379 & shamt_i[5];
  assign N375 = N374 & N380;
  assign N376 = N375 & N381;
  assign N377 = N376 & shamt_i[2];
  assign N378 = N377 & N382;
  assign N1103 = N378 & shamt_i[1];
  assign N379 = ~shamt_i[6];
  assign N380 = ~shamt_i[4];
  assign N381 = ~shamt_i[3];
  assign N382 = ~shamt_i[0];
  assign N383 = N388 & shamt_i[5];
  assign N384 = N383 & N389;
  assign N385 = N384 & N390;
  assign N386 = N385 & shamt_i[2];
  assign N387 = N386 & shamt_i[0];
  assign N1105 = N387 & shamt_i[1];
  assign N388 = ~shamt_i[6];
  assign N389 = ~shamt_i[4];
  assign N390 = ~shamt_i[3];
  assign N391 = N396 & shamt_i[5];
  assign N392 = N391 & N397;
  assign N393 = N392 & shamt_i[3];
  assign N394 = N393 & N398;
  assign N395 = N394 & N399;
  assign N1107 = N395 & N400;
  assign N396 = ~shamt_i[6];
  assign N397 = ~shamt_i[4];
  assign N398 = ~shamt_i[2];
  assign N399 = ~shamt_i[0];
  assign N400 = ~shamt_i[1];
  assign N401 = N406 & shamt_i[5];
  assign N402 = N401 & N407;
  assign N403 = N402 & shamt_i[3];
  assign N404 = N403 & N408;
  assign N405 = N404 & shamt_i[0];
  assign N1109 = N405 & N409;
  assign N406 = ~shamt_i[6];
  assign N407 = ~shamt_i[4];
  assign N408 = ~shamt_i[2];
  assign N409 = ~shamt_i[1];
  assign N410 = N415 & shamt_i[5];
  assign N411 = N410 & N416;
  assign N412 = N411 & shamt_i[3];
  assign N413 = N412 & N417;
  assign N414 = N413 & N418;
  assign N1111 = N414 & shamt_i[1];
  assign N415 = ~shamt_i[6];
  assign N416 = ~shamt_i[4];
  assign N417 = ~shamt_i[2];
  assign N418 = ~shamt_i[0];
  assign N419 = N424 & shamt_i[5];
  assign N420 = N419 & N425;
  assign N421 = N420 & shamt_i[3];
  assign N422 = N421 & N426;
  assign N423 = N422 & shamt_i[0];
  assign N1113 = N423 & shamt_i[1];
  assign N424 = ~shamt_i[6];
  assign N425 = ~shamt_i[4];
  assign N426 = ~shamt_i[2];
  assign N427 = N432 & shamt_i[5];
  assign N428 = N427 & N433;
  assign N429 = N428 & shamt_i[3];
  assign N430 = N429 & shamt_i[2];
  assign N431 = N430 & N434;
  assign N1115 = N431 & N435;
  assign N432 = ~shamt_i[6];
  assign N433 = ~shamt_i[4];
  assign N434 = ~shamt_i[0];
  assign N435 = ~shamt_i[1];
  assign N436 = N441 & shamt_i[5];
  assign N437 = N436 & N442;
  assign N438 = N437 & shamt_i[3];
  assign N439 = N438 & shamt_i[2];
  assign N440 = N439 & shamt_i[0];
  assign N1117 = N440 & N443;
  assign N441 = ~shamt_i[6];
  assign N442 = ~shamt_i[4];
  assign N443 = ~shamt_i[1];
  assign N444 = N449 & shamt_i[5];
  assign N445 = N444 & N450;
  assign N446 = N445 & shamt_i[3];
  assign N447 = N446 & shamt_i[2];
  assign N448 = N447 & N451;
  assign N1119 = N448 & shamt_i[1];
  assign N449 = ~shamt_i[6];
  assign N450 = ~shamt_i[4];
  assign N451 = ~shamt_i[0];
  assign N452 = N457 & shamt_i[5];
  assign N453 = N452 & N458;
  assign N454 = N453 & shamt_i[3];
  assign N455 = N454 & shamt_i[2];
  assign N456 = N455 & shamt_i[0];
  assign N1121 = N456 & shamt_i[1];
  assign N457 = ~shamt_i[6];
  assign N458 = ~shamt_i[4];
  assign N459 = N464 & shamt_i[5];
  assign N460 = N459 & shamt_i[4];
  assign N461 = N460 & N465;
  assign N462 = N461 & N466;
  assign N463 = N462 & N467;
  assign N1123 = N463 & N468;
  assign N464 = ~shamt_i[6];
  assign N465 = ~shamt_i[3];
  assign N466 = ~shamt_i[2];
  assign N467 = ~shamt_i[0];
  assign N468 = ~shamt_i[1];
  assign N469 = N474 & shamt_i[5];
  assign N470 = N469 & shamt_i[4];
  assign N471 = N470 & N475;
  assign N472 = N471 & N476;
  assign N473 = N472 & shamt_i[0];
  assign N1125 = N473 & N477;
  assign N474 = ~shamt_i[6];
  assign N475 = ~shamt_i[3];
  assign N476 = ~shamt_i[2];
  assign N477 = ~shamt_i[1];
  assign N478 = N483 & shamt_i[5];
  assign N479 = N478 & shamt_i[4];
  assign N480 = N479 & N484;
  assign N481 = N480 & N485;
  assign N482 = N481 & N486;
  assign N1127 = N482 & shamt_i[1];
  assign N483 = ~shamt_i[6];
  assign N484 = ~shamt_i[3];
  assign N485 = ~shamt_i[2];
  assign N486 = ~shamt_i[0];
  assign N487 = N492 & shamt_i[5];
  assign N488 = N487 & shamt_i[4];
  assign N489 = N488 & N493;
  assign N490 = N489 & N494;
  assign N491 = N490 & shamt_i[0];
  assign N1129 = N491 & shamt_i[1];
  assign N492 = ~shamt_i[6];
  assign N493 = ~shamt_i[3];
  assign N494 = ~shamt_i[2];
  assign N495 = shamt_i[5] & shamt_i[4];
  assign N496 = N495 & N499;
  assign N497 = N496 & shamt_i[2];
  assign N498 = N497 & N500;
  assign N1131 = N498 & N501;
  assign N499 = ~shamt_i[3];
  assign N500 = ~shamt_i[0];
  assign N501 = ~shamt_i[1];
  assign N502 = shamt_i[5] & shamt_i[4];
  assign N503 = N502 & N506;
  assign N504 = N503 & shamt_i[2];
  assign N505 = N504 & shamt_i[0];
  assign N1132 = N505 & N507;
  assign N506 = ~shamt_i[3];
  assign N507 = ~shamt_i[1];
  assign N508 = shamt_i[5] & shamt_i[4];
  assign N509 = N508 & N512;
  assign N510 = N509 & shamt_i[2];
  assign N511 = N510 & N513;
  assign N1133 = N511 & shamt_i[1];
  assign N512 = ~shamt_i[3];
  assign N513 = ~shamt_i[0];
  assign N514 = shamt_i[5] & shamt_i[4];
  assign N515 = N514 & N518;
  assign N516 = N515 & shamt_i[2];
  assign N517 = N516 & shamt_i[0];
  assign N1134 = N517 & shamt_i[1];
  assign N518 = ~shamt_i[3];
  assign N519 = shamt_i[5] & shamt_i[4];
  assign N520 = N519 & shamt_i[3];
  assign N521 = N520 & N523;
  assign N522 = N521 & N524;
  assign N1135 = N522 & N525;
  assign N523 = ~shamt_i[2];
  assign N524 = ~shamt_i[0];
  assign N525 = ~shamt_i[1];
  assign N526 = shamt_i[5] & shamt_i[4];
  assign N527 = N526 & shamt_i[3];
  assign N528 = N527 & N530;
  assign N529 = N528 & shamt_i[0];
  assign N1136 = N529 & N531;
  assign N530 = ~shamt_i[2];
  assign N531 = ~shamt_i[1];
  assign N532 = shamt_i[5] & shamt_i[4];
  assign N533 = N532 & shamt_i[3];
  assign N534 = N533 & N536;
  assign N535 = N534 & N537;
  assign N1137 = N535 & shamt_i[1];
  assign N536 = ~shamt_i[2];
  assign N537 = ~shamt_i[0];
  assign N538 = shamt_i[5] & shamt_i[4];
  assign N539 = N538 & shamt_i[3];
  assign N540 = N539 & N542;
  assign N541 = N540 & shamt_i[0];
  assign N1138 = N541 & shamt_i[1];
  assign N542 = ~shamt_i[2];
  assign N543 = shamt_i[5] & shamt_i[4];
  assign N544 = N543 & shamt_i[3];
  assign N545 = N544 & shamt_i[2];
  assign N546 = N545 & N547;
  assign N1139 = N546 & N548;
  assign N547 = ~shamt_i[0];
  assign N548 = ~shamt_i[1];
  assign N549 = shamt_i[5] & shamt_i[4];
  assign N550 = N549 & shamt_i[3];
  assign N551 = N550 & shamt_i[2];
  assign N552 = N551 & shamt_i[0];
  assign N1140 = N552 & N553;
  assign N553 = ~shamt_i[1];
  assign N554 = shamt_i[5] & shamt_i[4];
  assign N555 = N554 & shamt_i[3];
  assign N556 = N555 & shamt_i[2];
  assign N557 = N556 & N558;
  assign N1141 = N557 & shamt_i[1];
  assign N558 = ~shamt_i[0];
  assign N559 = shamt_i[5] & shamt_i[4];
  assign N560 = N559 & shamt_i[3];
  assign N561 = N560 & shamt_i[2];
  assign N562 = N561 & shamt_i[0];
  assign N1142 = N562 & shamt_i[1];
  assign N563 = shamt_i[6] & N568;
  assign N564 = N563 & N569;
  assign N565 = N564 & N570;
  assign N566 = N565 & N571;
  assign N567 = N566 & shamt_i[0];
  assign N1030 = N567 & N572;
  assign N568 = ~shamt_i[5];
  assign N569 = ~shamt_i[4];
  assign N570 = ~shamt_i[3];
  assign N571 = ~shamt_i[2];
  assign N572 = ~shamt_i[1];
  assign N573 = shamt_i[6] & N578;
  assign N574 = N573 & N579;
  assign N575 = N574 & N580;
  assign N576 = N575 & N581;
  assign N577 = N576 & N582;
  assign N1032 = N577 & shamt_i[1];
  assign N578 = ~shamt_i[5];
  assign N579 = ~shamt_i[4];
  assign N580 = ~shamt_i[3];
  assign N581 = ~shamt_i[2];
  assign N582 = ~shamt_i[0];
  assign N583 = shamt_i[6] & N588;
  assign N584 = N583 & N589;
  assign N585 = N584 & N590;
  assign N586 = N585 & N591;
  assign N587 = N586 & shamt_i[0];
  assign N1034 = N587 & shamt_i[1];
  assign N588 = ~shamt_i[5];
  assign N589 = ~shamt_i[4];
  assign N590 = ~shamt_i[3];
  assign N591 = ~shamt_i[2];
  assign N592 = shamt_i[6] & N597;
  assign N593 = N592 & N598;
  assign N594 = N593 & N599;
  assign N595 = N594 & shamt_i[2];
  assign N596 = N595 & N600;
  assign N1036 = N596 & N601;
  assign N597 = ~shamt_i[5];
  assign N598 = ~shamt_i[4];
  assign N599 = ~shamt_i[3];
  assign N600 = ~shamt_i[0];
  assign N601 = ~shamt_i[1];
  assign N602 = shamt_i[6] & N607;
  assign N603 = N602 & N608;
  assign N604 = N603 & N609;
  assign N605 = N604 & shamt_i[2];
  assign N606 = N605 & shamt_i[0];
  assign N1038 = N606 & N610;
  assign N607 = ~shamt_i[5];
  assign N608 = ~shamt_i[4];
  assign N609 = ~shamt_i[3];
  assign N610 = ~shamt_i[1];
  assign N611 = shamt_i[6] & N616;
  assign N612 = N611 & N617;
  assign N613 = N612 & N618;
  assign N614 = N613 & shamt_i[2];
  assign N615 = N614 & N619;
  assign N1040 = N615 & shamt_i[1];
  assign N616 = ~shamt_i[5];
  assign N617 = ~shamt_i[4];
  assign N618 = ~shamt_i[3];
  assign N619 = ~shamt_i[0];
  assign N620 = shamt_i[6] & N625;
  assign N621 = N620 & N626;
  assign N622 = N621 & N627;
  assign N623 = N622 & shamt_i[2];
  assign N624 = N623 & shamt_i[0];
  assign N1042 = N624 & shamt_i[1];
  assign N625 = ~shamt_i[5];
  assign N626 = ~shamt_i[4];
  assign N627 = ~shamt_i[3];
  assign N628 = shamt_i[6] & N633;
  assign N629 = N628 & N634;
  assign N630 = N629 & shamt_i[3];
  assign N631 = N630 & N635;
  assign N632 = N631 & N636;
  assign N1044 = N632 & N637;
  assign N633 = ~shamt_i[5];
  assign N634 = ~shamt_i[4];
  assign N635 = ~shamt_i[2];
  assign N636 = ~shamt_i[0];
  assign N637 = ~shamt_i[1];
  assign N638 = shamt_i[6] & N643;
  assign N639 = N638 & N644;
  assign N640 = N639 & shamt_i[3];
  assign N641 = N640 & N645;
  assign N642 = N641 & shamt_i[0];
  assign N1046 = N642 & N646;
  assign N643 = ~shamt_i[5];
  assign N644 = ~shamt_i[4];
  assign N645 = ~shamt_i[2];
  assign N646 = ~shamt_i[1];
  assign N647 = shamt_i[6] & N652;
  assign N648 = N647 & N653;
  assign N649 = N648 & shamt_i[3];
  assign N650 = N649 & N654;
  assign N651 = N650 & N655;
  assign N1048 = N651 & shamt_i[1];
  assign N652 = ~shamt_i[5];
  assign N653 = ~shamt_i[4];
  assign N654 = ~shamt_i[2];
  assign N655 = ~shamt_i[0];
  assign N656 = shamt_i[6] & N661;
  assign N657 = N656 & N662;
  assign N658 = N657 & shamt_i[3];
  assign N659 = N658 & N663;
  assign N660 = N659 & shamt_i[0];
  assign N1050 = N660 & shamt_i[1];
  assign N661 = ~shamt_i[5];
  assign N662 = ~shamt_i[4];
  assign N663 = ~shamt_i[2];
  assign N664 = shamt_i[6] & N669;
  assign N665 = N664 & N670;
  assign N666 = N665 & shamt_i[3];
  assign N667 = N666 & shamt_i[2];
  assign N668 = N667 & N671;
  assign N1052 = N668 & N672;
  assign N669 = ~shamt_i[5];
  assign N670 = ~shamt_i[4];
  assign N671 = ~shamt_i[0];
  assign N672 = ~shamt_i[1];
  assign N673 = shamt_i[6] & N678;
  assign N674 = N673 & N679;
  assign N675 = N674 & shamt_i[3];
  assign N676 = N675 & shamt_i[2];
  assign N677 = N676 & shamt_i[0];
  assign N1054 = N677 & N680;
  assign N678 = ~shamt_i[5];
  assign N679 = ~shamt_i[4];
  assign N680 = ~shamt_i[1];
  assign N681 = shamt_i[6] & N686;
  assign N682 = N681 & N687;
  assign N683 = N682 & shamt_i[3];
  assign N684 = N683 & shamt_i[2];
  assign N685 = N684 & N688;
  assign N1056 = N685 & shamt_i[1];
  assign N686 = ~shamt_i[5];
  assign N687 = ~shamt_i[4];
  assign N688 = ~shamt_i[0];
  assign N689 = shamt_i[6] & N694;
  assign N690 = N689 & N695;
  assign N691 = N690 & shamt_i[3];
  assign N692 = N691 & shamt_i[2];
  assign N693 = N692 & shamt_i[0];
  assign N1058 = N693 & shamt_i[1];
  assign N694 = ~shamt_i[5];
  assign N695 = ~shamt_i[4];
  assign N696 = shamt_i[6] & N701;
  assign N697 = N696 & shamt_i[4];
  assign N698 = N697 & N702;
  assign N699 = N698 & N703;
  assign N700 = N699 & N704;
  assign N1060 = N700 & N705;
  assign N701 = ~shamt_i[5];
  assign N702 = ~shamt_i[3];
  assign N703 = ~shamt_i[2];
  assign N704 = ~shamt_i[0];
  assign N705 = ~shamt_i[1];
  assign N706 = shamt_i[6] & N711;
  assign N707 = N706 & shamt_i[4];
  assign N708 = N707 & N712;
  assign N709 = N708 & N713;
  assign N710 = N709 & shamt_i[0];
  assign N1062 = N710 & N714;
  assign N711 = ~shamt_i[5];
  assign N712 = ~shamt_i[3];
  assign N713 = ~shamt_i[2];
  assign N714 = ~shamt_i[1];
  assign N715 = shamt_i[6] & N720;
  assign N716 = N715 & shamt_i[4];
  assign N717 = N716 & N721;
  assign N718 = N717 & N722;
  assign N719 = N718 & N723;
  assign N1064 = N719 & shamt_i[1];
  assign N720 = ~shamt_i[5];
  assign N721 = ~shamt_i[3];
  assign N722 = ~shamt_i[2];
  assign N723 = ~shamt_i[0];
  assign N724 = shamt_i[6] & N729;
  assign N725 = N724 & shamt_i[4];
  assign N726 = N725 & N730;
  assign N727 = N726 & N731;
  assign N728 = N727 & shamt_i[0];
  assign N1066 = N728 & shamt_i[1];
  assign N729 = ~shamt_i[5];
  assign N730 = ~shamt_i[3];
  assign N731 = ~shamt_i[2];
  assign N732 = shamt_i[6] & shamt_i[4];
  assign N733 = N732 & N736;
  assign N734 = N733 & shamt_i[2];
  assign N735 = N734 & N737;
  assign N1068 = N735 & N738;
  assign N736 = ~shamt_i[3];
  assign N737 = ~shamt_i[0];
  assign N738 = ~shamt_i[1];
  assign N739 = shamt_i[6] & shamt_i[4];
  assign N740 = N739 & N743;
  assign N741 = N740 & shamt_i[2];
  assign N742 = N741 & shamt_i[0];
  assign N1070 = N742 & N744;
  assign N743 = ~shamt_i[3];
  assign N744 = ~shamt_i[1];
  assign N745 = shamt_i[6] & shamt_i[4];
  assign N746 = N745 & N749;
  assign N747 = N746 & shamt_i[2];
  assign N748 = N747 & N750;
  assign N1072 = N748 & shamt_i[1];
  assign N749 = ~shamt_i[3];
  assign N750 = ~shamt_i[0];
  assign N751 = shamt_i[6] & shamt_i[4];
  assign N752 = N751 & N755;
  assign N753 = N752 & shamt_i[2];
  assign N754 = N753 & shamt_i[0];
  assign N1074 = N754 & shamt_i[1];
  assign N755 = ~shamt_i[3];
  assign N756 = shamt_i[6] & shamt_i[4];
  assign N757 = N756 & shamt_i[3];
  assign N758 = N757 & N760;
  assign N759 = N758 & N761;
  assign N1076 = N759 & N762;
  assign N760 = ~shamt_i[2];
  assign N761 = ~shamt_i[0];
  assign N762 = ~shamt_i[1];
  assign N763 = shamt_i[6] & shamt_i[4];
  assign N764 = N763 & shamt_i[3];
  assign N765 = N764 & N767;
  assign N766 = N765 & shamt_i[0];
  assign N1078 = N766 & N768;
  assign N767 = ~shamt_i[2];
  assign N768 = ~shamt_i[1];
  assign N769 = shamt_i[6] & shamt_i[4];
  assign N770 = N769 & shamt_i[3];
  assign N771 = N770 & N773;
  assign N772 = N771 & N774;
  assign N1080 = N772 & shamt_i[1];
  assign N773 = ~shamt_i[2];
  assign N774 = ~shamt_i[0];
  assign N775 = shamt_i[6] & shamt_i[4];
  assign N776 = N775 & shamt_i[3];
  assign N777 = N776 & N779;
  assign N778 = N777 & shamt_i[0];
  assign N1082 = N778 & shamt_i[1];
  assign N779 = ~shamt_i[2];
  assign N780 = shamt_i[6] & shamt_i[4];
  assign N781 = N780 & shamt_i[3];
  assign N782 = N781 & shamt_i[2];
  assign N783 = N782 & N784;
  assign N1084 = N783 & N785;
  assign N784 = ~shamt_i[0];
  assign N785 = ~shamt_i[1];
  assign N786 = shamt_i[6] & shamt_i[4];
  assign N787 = N786 & shamt_i[3];
  assign N788 = N787 & shamt_i[2];
  assign N789 = N788 & shamt_i[0];
  assign N1086 = N789 & N790;
  assign N790 = ~shamt_i[1];
  assign N791 = shamt_i[6] & shamt_i[4];
  assign N792 = N791 & shamt_i[3];
  assign N793 = N792 & shamt_i[2];
  assign N794 = N793 & N795;
  assign N1088 = N794 & shamt_i[1];
  assign N795 = ~shamt_i[0];
  assign N796 = shamt_i[6] & shamt_i[4];
  assign N797 = N796 & shamt_i[3];
  assign N798 = N797 & shamt_i[2];
  assign N799 = N798 & shamt_i[0];
  assign N1090 = N799 & shamt_i[1];
  assign N800 = shamt_i[6] & shamt_i[5];
  assign N801 = N800 & N805;
  assign N802 = N801 & N806;
  assign N803 = N802 & N807;
  assign N804 = N803 & N808;
  assign N1092 = N804 & N809;
  assign N805 = ~shamt_i[4];
  assign N806 = ~shamt_i[3];
  assign N807 = ~shamt_i[2];
  assign N808 = ~shamt_i[0];
  assign N809 = ~shamt_i[1];
  assign N810 = shamt_i[6] & shamt_i[5];
  assign N811 = N810 & N815;
  assign N812 = N811 & N816;
  assign N813 = N812 & N817;
  assign N814 = N813 & shamt_i[0];
  assign N1094 = N814 & N818;
  assign N815 = ~shamt_i[4];
  assign N816 = ~shamt_i[3];
  assign N817 = ~shamt_i[2];
  assign N818 = ~shamt_i[1];
  assign N819 = shamt_i[6] & shamt_i[5];
  assign N820 = N819 & N824;
  assign N821 = N820 & N825;
  assign N822 = N821 & N826;
  assign N823 = N822 & N827;
  assign N1096 = N823 & shamt_i[1];
  assign N824 = ~shamt_i[4];
  assign N825 = ~shamt_i[3];
  assign N826 = ~shamt_i[2];
  assign N827 = ~shamt_i[0];
  assign N828 = shamt_i[6] & shamt_i[5];
  assign N829 = N828 & N833;
  assign N830 = N829 & N834;
  assign N831 = N830 & N835;
  assign N832 = N831 & shamt_i[0];
  assign N1098 = N832 & shamt_i[1];
  assign N833 = ~shamt_i[4];
  assign N834 = ~shamt_i[3];
  assign N835 = ~shamt_i[2];
  assign N836 = shamt_i[6] & shamt_i[5];
  assign N837 = N836 & N840;
  assign N838 = N837 & shamt_i[2];
  assign N839 = N838 & N841;
  assign N1100 = N839 & N842;
  assign N840 = ~shamt_i[3];
  assign N841 = ~shamt_i[0];
  assign N842 = ~shamt_i[1];
  assign N843 = shamt_i[6] & shamt_i[5];
  assign N844 = N843 & N847;
  assign N845 = N844 & shamt_i[2];
  assign N846 = N845 & shamt_i[0];
  assign N1102 = N846 & N848;
  assign N847 = ~shamt_i[3];
  assign N848 = ~shamt_i[1];
  assign N849 = shamt_i[6] & shamt_i[5];
  assign N850 = N849 & N853;
  assign N851 = N850 & shamt_i[2];
  assign N852 = N851 & N854;
  assign N1104 = N852 & shamt_i[1];
  assign N853 = ~shamt_i[3];
  assign N854 = ~shamt_i[0];
  assign N855 = shamt_i[6] & shamt_i[5];
  assign N856 = N855 & N859;
  assign N857 = N856 & shamt_i[2];
  assign N858 = N857 & shamt_i[0];
  assign N1106 = N858 & shamt_i[1];
  assign N859 = ~shamt_i[3];
  assign N860 = shamt_i[6] & shamt_i[5];
  assign N861 = N860 & shamt_i[3];
  assign N862 = N861 & N864;
  assign N863 = N862 & N865;
  assign N1108 = N863 & N866;
  assign N864 = ~shamt_i[2];
  assign N865 = ~shamt_i[0];
  assign N866 = ~shamt_i[1];
  assign N867 = shamt_i[6] & shamt_i[5];
  assign N868 = N867 & shamt_i[3];
  assign N869 = N868 & N871;
  assign N870 = N869 & shamt_i[0];
  assign N1110 = N870 & N872;
  assign N871 = ~shamt_i[2];
  assign N872 = ~shamt_i[1];
  assign N873 = shamt_i[6] & shamt_i[5];
  assign N874 = N873 & shamt_i[3];
  assign N875 = N874 & N877;
  assign N876 = N875 & N878;
  assign N1112 = N876 & shamt_i[1];
  assign N877 = ~shamt_i[2];
  assign N878 = ~shamt_i[0];
  assign N879 = shamt_i[6] & shamt_i[5];
  assign N880 = N879 & shamt_i[3];
  assign N881 = N880 & N883;
  assign N882 = N881 & shamt_i[0];
  assign N1114 = N882 & shamt_i[1];
  assign N883 = ~shamt_i[2];
  assign N884 = shamt_i[6] & shamt_i[5];
  assign N885 = N884 & shamt_i[3];
  assign N886 = N885 & shamt_i[2];
  assign N887 = N886 & N888;
  assign N1116 = N887 & N889;
  assign N888 = ~shamt_i[0];
  assign N889 = ~shamt_i[1];
  assign N890 = shamt_i[6] & shamt_i[5];
  assign N891 = N890 & shamt_i[3];
  assign N892 = N891 & shamt_i[2];
  assign N893 = N892 & shamt_i[0];
  assign N1118 = N893 & N894;
  assign N894 = ~shamt_i[1];
  assign N895 = shamt_i[6] & shamt_i[5];
  assign N896 = N895 & shamt_i[3];
  assign N897 = N896 & shamt_i[2];
  assign N898 = N897 & N899;
  assign N1120 = N898 & shamt_i[1];
  assign N899 = ~shamt_i[0];
  assign N900 = shamt_i[6] & shamt_i[5];
  assign N901 = N900 & shamt_i[3];
  assign N902 = N901 & shamt_i[2];
  assign N903 = N902 & shamt_i[0];
  assign N1122 = N903 & shamt_i[1];
  assign N1124 = shamt_i[6] & shamt_i[5] & (shamt_i[4] & N904) & N905;
  assign N904 = ~shamt_i[0];
  assign N905 = ~shamt_i[1];
  assign N1126 = shamt_i[6] & shamt_i[5] & (shamt_i[4] & shamt_i[0]) & N906;
  assign N906 = ~shamt_i[1];
  assign N1128 = shamt_i[6] & shamt_i[5] & (shamt_i[4] & N907) & shamt_i[1];
  assign N907 = ~shamt_i[0];
  assign N1130 = shamt_i[6] & shamt_i[5] & (shamt_i[4] & shamt_i[0]) & shamt_i[1];
  assign sticky_o = (N908)? scan_out[114] : 
                    (N1026)? N1143 : 1'b0;
  assign N908 = N1025;
  assign N1143 = (N909)? 1'b0 : 
                 (N910)? scan_out[0] : 
                 (N911)? scan_out[1] : 
                 (N912)? scan_out[2] : 
                 (N913)? scan_out[3] : 
                 (N914)? scan_out[4] : 
                 (N915)? scan_out[5] : 
                 (N916)? scan_out[6] : 
                 (N917)? scan_out[7] : 
                 (N918)? scan_out[8] : 
                 (N919)? scan_out[9] : 
                 (N920)? scan_out[10] : 
                 (N921)? scan_out[11] : 
                 (N922)? scan_out[12] : 
                 (N923)? scan_out[13] : 
                 (N924)? scan_out[14] : 
                 (N925)? scan_out[15] : 
                 (N926)? scan_out[16] : 
                 (N927)? scan_out[17] : 
                 (N928)? scan_out[18] : 
                 (N929)? scan_out[19] : 
                 (N930)? scan_out[20] : 
                 (N931)? scan_out[21] : 
                 (N932)? scan_out[22] : 
                 (N933)? scan_out[23] : 
                 (N934)? scan_out[24] : 
                 (N935)? scan_out[25] : 
                 (N936)? scan_out[26] : 
                 (N937)? scan_out[27] : 
                 (N938)? scan_out[28] : 
                 (N939)? scan_out[29] : 
                 (N940)? scan_out[30] : 
                 (N941)? scan_out[31] : 
                 (N942)? scan_out[32] : 
                 (N943)? scan_out[33] : 
                 (N944)? scan_out[34] : 
                 (N945)? scan_out[35] : 
                 (N946)? scan_out[36] : 
                 (N947)? scan_out[37] : 
                 (N948)? scan_out[38] : 
                 (N949)? scan_out[39] : 
                 (N950)? scan_out[40] : 
                 (N951)? scan_out[41] : 
                 (N952)? scan_out[42] : 
                 (N953)? scan_out[43] : 
                 (N954)? scan_out[44] : 
                 (N955)? scan_out[45] : 
                 (N956)? scan_out[46] : 
                 (N957)? scan_out[47] : 
                 (N958)? scan_out[48] : 
                 (N959)? scan_out[49] : 
                 (N960)? scan_out[50] : 
                 (N961)? scan_out[51] : 
                 (N962)? scan_out[52] : 
                 (N963)? scan_out[53] : 
                 (N964)? scan_out[54] : 
                 (N965)? scan_out[55] : 
                 (N966)? scan_out[56] : 
                 (N967)? scan_out[57] : 
                 (N968)? scan_out[58] : 
                 (N969)? scan_out[59] : 
                 (N970)? scan_out[60] : 
                 (N971)? scan_out[61] : 
                 (N972)? scan_out[62] : 
                 (N973)? scan_out[63] : 
                 (N974)? scan_out[64] : 
                 (N975)? scan_out[65] : 
                 (N976)? scan_out[66] : 
                 (N977)? scan_out[67] : 
                 (N978)? scan_out[68] : 
                 (N979)? scan_out[69] : 
                 (N980)? scan_out[70] : 
                 (N981)? scan_out[71] : 
                 (N982)? scan_out[72] : 
                 (N983)? scan_out[73] : 
                 (N984)? scan_out[74] : 
                 (N985)? scan_out[75] : 
                 (N986)? scan_out[76] : 
                 (N987)? scan_out[77] : 
                 (N988)? scan_out[78] : 
                 (N989)? scan_out[79] : 
                 (N990)? scan_out[80] : 
                 (N991)? scan_out[81] : 
                 (N992)? scan_out[82] : 
                 (N993)? scan_out[83] : 
                 (N994)? scan_out[84] : 
                 (N995)? scan_out[85] : 
                 (N996)? scan_out[86] : 
                 (N997)? scan_out[87] : 
                 (N998)? scan_out[88] : 
                 (N999)? scan_out[89] : 
                 (N1000)? scan_out[90] : 
                 (N1001)? scan_out[91] : 
                 (N1002)? scan_out[92] : 
                 (N1003)? scan_out[93] : 
                 (N1004)? scan_out[94] : 
                 (N1005)? scan_out[95] : 
                 (N1006)? scan_out[96] : 
                 (N1007)? scan_out[97] : 
                 (N1008)? scan_out[98] : 
                 (N1009)? scan_out[99] : 
                 (N1010)? scan_out[100] : 
                 (N1011)? scan_out[101] : 
                 (N1012)? scan_out[102] : 
                 (N1013)? scan_out[103] : 
                 (N1014)? scan_out[104] : 
                 (N1015)? scan_out[105] : 
                 (N1016)? scan_out[106] : 
                 (N1017)? scan_out[107] : 
                 (N1018)? scan_out[108] : 
                 (N1019)? scan_out[109] : 
                 (N1020)? scan_out[110] : 
                 (N1021)? scan_out[111] : 
                 (N1022)? scan_out[112] : 
                 (N1023)? scan_out[113] : 
                 (N1024)? scan_out[114] : 1'b0;
  assign N909 = N1027;
  assign N910 = N1029;
  assign N911 = N1031;
  assign N912 = N1033;
  assign N913 = N1035;
  assign N914 = N1037;
  assign N915 = N1039;
  assign N916 = N1041;
  assign N917 = N1043;
  assign N918 = N1045;
  assign N919 = N1047;
  assign N920 = N1049;
  assign N921 = N1051;
  assign N922 = N1053;
  assign N923 = N1055;
  assign N924 = N1057;
  assign N925 = N1059;
  assign N926 = N1061;
  assign N927 = N1063;
  assign N928 = N1065;
  assign N929 = N1067;
  assign N930 = N1069;
  assign N931 = N1071;
  assign N932 = N1073;
  assign N933 = N1075;
  assign N934 = N1077;
  assign N935 = N1079;
  assign N936 = N1081;
  assign N937 = N1083;
  assign N938 = N1085;
  assign N939 = N1087;
  assign N940 = N1089;
  assign N941 = N1091;
  assign N942 = N1093;
  assign N943 = N1095;
  assign N944 = N1097;
  assign N945 = N1099;
  assign N946 = N1101;
  assign N947 = N1103;
  assign N948 = N1105;
  assign N949 = N1107;
  assign N950 = N1109;
  assign N951 = N1111;
  assign N952 = N1113;
  assign N953 = N1115;
  assign N954 = N1117;
  assign N955 = N1119;
  assign N956 = N1121;
  assign N957 = N1123;
  assign N958 = N1125;
  assign N959 = N1127;
  assign N960 = N1129;
  assign N961 = N1131;
  assign N962 = N1132;
  assign N963 = N1133;
  assign N964 = N1134;
  assign N965 = N1135;
  assign N966 = N1136;
  assign N967 = N1137;
  assign N968 = N1138;
  assign N969 = N1139;
  assign N970 = N1140;
  assign N971 = N1141;
  assign N972 = N1142;
  assign N973 = N1028;
  assign N974 = N1030;
  assign N975 = N1032;
  assign N976 = N1034;
  assign N977 = N1036;
  assign N978 = N1038;
  assign N979 = N1040;
  assign N980 = N1042;
  assign N981 = N1044;
  assign N982 = N1046;
  assign N983 = N1048;
  assign N984 = N1050;
  assign N985 = N1052;
  assign N986 = N1054;
  assign N987 = N1056;
  assign N988 = N1058;
  assign N989 = N1060;
  assign N990 = N1062;
  assign N991 = N1064;
  assign N992 = N1066;
  assign N993 = N1068;
  assign N994 = N1070;
  assign N995 = N1072;
  assign N996 = N1074;
  assign N997 = N1076;
  assign N998 = N1078;
  assign N999 = N1080;
  assign N1000 = N1082;
  assign N1001 = N1084;
  assign N1002 = N1086;
  assign N1003 = N1088;
  assign N1004 = N1090;
  assign N1005 = N1092;
  assign N1006 = N1094;
  assign N1007 = N1096;
  assign N1008 = N1098;
  assign N1009 = N1100;
  assign N1010 = N1102;
  assign N1011 = N1104;
  assign N1012 = N1106;
  assign N1013 = N1108;
  assign N1014 = N1110;
  assign N1015 = N1112;
  assign N1016 = N1114;
  assign N1017 = N1116;
  assign N1018 = N1118;
  assign N1019 = N1120;
  assign N1020 = N1122;
  assign N1021 = N1124;
  assign N1022 = N1126;
  assign N1023 = N1128;
  assign N1024 = N1130;
  assign N1026 = ~N1025;

endmodule



module bsg_less_than_width_p127
(
  a_i,
  b_i,
  o
);

  input [126:0] a_i;
  input [126:0] b_i;
  output o;
  wire o;
  assign o = a_i < b_i;

endmodule



module bsg_less_than_width_p116
(
  a_i,
  b_i,
  o
);

  input [115:0] a_i;
  input [115:0] b_i;
  output o;
  wire o;
  assign o = a_i < b_i;

endmodule



module bsg_scan_width_p117_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [116:0] i;
  output [116:0] o;
  wire [116:0] o;
  wire t_6__116_,t_6__115_,t_6__114_,t_6__113_,t_6__112_,t_6__111_,t_6__110_,t_6__109_,
  t_6__108_,t_6__107_,t_6__106_,t_6__105_,t_6__104_,t_6__103_,t_6__102_,t_6__101_,
  t_6__100_,t_6__99_,t_6__98_,t_6__97_,t_6__96_,t_6__95_,t_6__94_,t_6__93_,
  t_6__92_,t_6__91_,t_6__90_,t_6__89_,t_6__88_,t_6__87_,t_6__86_,t_6__85_,t_6__84_,
  t_6__83_,t_6__82_,t_6__81_,t_6__80_,t_6__79_,t_6__78_,t_6__77_,t_6__76_,t_6__75_,
  t_6__74_,t_6__73_,t_6__72_,t_6__71_,t_6__70_,t_6__69_,t_6__68_,t_6__67_,t_6__66_,
  t_6__65_,t_6__64_,t_6__63_,t_6__62_,t_6__61_,t_6__60_,t_6__59_,t_6__58_,t_6__57_,
  t_6__56_,t_6__55_,t_6__54_,t_6__53_,t_6__52_,t_6__51_,t_6__50_,t_6__49_,t_6__48_,
  t_6__47_,t_6__46_,t_6__45_,t_6__44_,t_6__43_,t_6__42_,t_6__41_,t_6__40_,t_6__39_,
  t_6__38_,t_6__37_,t_6__36_,t_6__35_,t_6__34_,t_6__33_,t_6__32_,t_6__31_,t_6__30_,
  t_6__29_,t_6__28_,t_6__27_,t_6__26_,t_6__25_,t_6__24_,t_6__23_,t_6__22_,
  t_6__21_,t_6__20_,t_6__19_,t_6__18_,t_6__17_,t_6__16_,t_6__15_,t_6__14_,t_6__13_,
  t_6__12_,t_6__11_,t_6__10_,t_6__9_,t_6__8_,t_6__7_,t_6__6_,t_6__5_,t_6__4_,t_6__3_,
  t_6__2_,t_6__1_,t_6__0_,t_5__116_,t_5__115_,t_5__114_,t_5__113_,t_5__112_,t_5__111_,
  t_5__110_,t_5__109_,t_5__108_,t_5__107_,t_5__106_,t_5__105_,t_5__104_,t_5__103_,
  t_5__102_,t_5__101_,t_5__100_,t_5__99_,t_5__98_,t_5__97_,t_5__96_,t_5__95_,
  t_5__94_,t_5__93_,t_5__92_,t_5__91_,t_5__90_,t_5__89_,t_5__88_,t_5__87_,t_5__86_,
  t_5__85_,t_5__84_,t_5__83_,t_5__82_,t_5__81_,t_5__80_,t_5__79_,t_5__78_,t_5__77_,
  t_5__76_,t_5__75_,t_5__74_,t_5__73_,t_5__72_,t_5__71_,t_5__70_,t_5__69_,t_5__68_,
  t_5__67_,t_5__66_,t_5__65_,t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,
  t_5__58_,t_5__57_,t_5__56_,t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,
  t_5__49_,t_5__48_,t_5__47_,t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,
  t_5__41_,t_5__40_,t_5__39_,t_5__38_,t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,
  t_5__32_,t_5__31_,t_5__30_,t_5__29_,t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,
  t_5__23_,t_5__22_,t_5__21_,t_5__20_,t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,
  t_5__14_,t_5__13_,t_5__12_,t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,
  t_5__4_,t_5__3_,t_5__2_,t_5__1_,t_5__0_,t_4__116_,t_4__115_,t_4__114_,t_4__113_,
  t_4__112_,t_4__111_,t_4__110_,t_4__109_,t_4__108_,t_4__107_,t_4__106_,t_4__105_,
  t_4__104_,t_4__103_,t_4__102_,t_4__101_,t_4__100_,t_4__99_,t_4__98_,t_4__97_,
  t_4__96_,t_4__95_,t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,t_4__89_,t_4__88_,
  t_4__87_,t_4__86_,t_4__85_,t_4__84_,t_4__83_,t_4__82_,t_4__81_,t_4__80_,t_4__79_,
  t_4__78_,t_4__77_,t_4__76_,t_4__75_,t_4__74_,t_4__73_,t_4__72_,t_4__71_,t_4__70_,
  t_4__69_,t_4__68_,t_4__67_,t_4__66_,t_4__65_,t_4__64_,t_4__63_,t_4__62_,
  t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,
  t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,
  t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,
  t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,
  t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,
  t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,
  t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_,t_3__116_,t_3__115_,
  t_3__114_,t_3__113_,t_3__112_,t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,
  t_3__106_,t_3__105_,t_3__104_,t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,
  t_3__98_,t_3__97_,t_3__96_,t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,
  t_3__89_,t_3__88_,t_3__87_,t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,
  t_3__81_,t_3__80_,t_3__79_,t_3__78_,t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,
  t_3__72_,t_3__71_,t_3__70_,t_3__69_,t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,
  t_3__63_,t_3__62_,t_3__61_,t_3__60_,t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,
  t_3__54_,t_3__53_,t_3__52_,t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,
  t_3__45_,t_3__44_,t_3__43_,t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,
  t_3__36_,t_3__35_,t_3__34_,t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,
  t_3__27_,t_3__26_,t_3__25_,t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,
  t_3__18_,t_3__17_,t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,
  t_3__9_,t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,
  t_2__116_,t_2__115_,t_2__114_,t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,
  t_2__108_,t_2__107_,t_2__106_,t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,
  t_2__100_,t_2__99_,t_2__98_,t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,
  t_2__92_,t_2__91_,t_2__90_,t_2__89_,t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,
  t_2__83_,t_2__82_,t_2__81_,t_2__80_,t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,
  t_2__74_,t_2__73_,t_2__72_,t_2__71_,t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,
  t_2__65_,t_2__64_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,
  t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,
  t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,
  t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,
  t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_1__116_,t_1__115_,t_1__114_,t_1__113_,t_1__112_,t_1__111_,
  t_1__110_,t_1__109_,t_1__108_,t_1__107_,t_1__106_,t_1__105_,t_1__104_,t_1__103_,
  t_1__102_,t_1__101_,t_1__100_,t_1__99_,t_1__98_,t_1__97_,t_1__96_,t_1__95_,
  t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,t_1__89_,t_1__88_,t_1__87_,t_1__86_,
  t_1__85_,t_1__84_,t_1__83_,t_1__82_,t_1__81_,t_1__80_,t_1__79_,t_1__78_,t_1__77_,
  t_1__76_,t_1__75_,t_1__74_,t_1__73_,t_1__72_,t_1__71_,t_1__70_,t_1__69_,t_1__68_,
  t_1__67_,t_1__66_,t_1__65_,t_1__64_,t_1__63_,t_1__62_,t_1__61_,t_1__60_,t_1__59_,
  t_1__58_,t_1__57_,t_1__56_,t_1__55_,t_1__54_,t_1__53_,t_1__52_,t_1__51_,t_1__50_,
  t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,t_1__44_,t_1__43_,t_1__42_,
  t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,t_1__35_,t_1__34_,t_1__33_,
  t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,t_1__26_,t_1__25_,t_1__24_,
  t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,t_1__17_,t_1__16_,t_1__15_,
  t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,
  t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__116_ = i[0] | 1'b0;
  assign t_1__115_ = i[1] | i[0];
  assign t_1__114_ = i[2] | i[1];
  assign t_1__113_ = i[3] | i[2];
  assign t_1__112_ = i[4] | i[3];
  assign t_1__111_ = i[5] | i[4];
  assign t_1__110_ = i[6] | i[5];
  assign t_1__109_ = i[7] | i[6];
  assign t_1__108_ = i[8] | i[7];
  assign t_1__107_ = i[9] | i[8];
  assign t_1__106_ = i[10] | i[9];
  assign t_1__105_ = i[11] | i[10];
  assign t_1__104_ = i[12] | i[11];
  assign t_1__103_ = i[13] | i[12];
  assign t_1__102_ = i[14] | i[13];
  assign t_1__101_ = i[15] | i[14];
  assign t_1__100_ = i[16] | i[15];
  assign t_1__99_ = i[17] | i[16];
  assign t_1__98_ = i[18] | i[17];
  assign t_1__97_ = i[19] | i[18];
  assign t_1__96_ = i[20] | i[19];
  assign t_1__95_ = i[21] | i[20];
  assign t_1__94_ = i[22] | i[21];
  assign t_1__93_ = i[23] | i[22];
  assign t_1__92_ = i[24] | i[23];
  assign t_1__91_ = i[25] | i[24];
  assign t_1__90_ = i[26] | i[25];
  assign t_1__89_ = i[27] | i[26];
  assign t_1__88_ = i[28] | i[27];
  assign t_1__87_ = i[29] | i[28];
  assign t_1__86_ = i[30] | i[29];
  assign t_1__85_ = i[31] | i[30];
  assign t_1__84_ = i[32] | i[31];
  assign t_1__83_ = i[33] | i[32];
  assign t_1__82_ = i[34] | i[33];
  assign t_1__81_ = i[35] | i[34];
  assign t_1__80_ = i[36] | i[35];
  assign t_1__79_ = i[37] | i[36];
  assign t_1__78_ = i[38] | i[37];
  assign t_1__77_ = i[39] | i[38];
  assign t_1__76_ = i[40] | i[39];
  assign t_1__75_ = i[41] | i[40];
  assign t_1__74_ = i[42] | i[41];
  assign t_1__73_ = i[43] | i[42];
  assign t_1__72_ = i[44] | i[43];
  assign t_1__71_ = i[45] | i[44];
  assign t_1__70_ = i[46] | i[45];
  assign t_1__69_ = i[47] | i[46];
  assign t_1__68_ = i[48] | i[47];
  assign t_1__67_ = i[49] | i[48];
  assign t_1__66_ = i[50] | i[49];
  assign t_1__65_ = i[51] | i[50];
  assign t_1__64_ = i[52] | i[51];
  assign t_1__63_ = i[53] | i[52];
  assign t_1__62_ = i[54] | i[53];
  assign t_1__61_ = i[55] | i[54];
  assign t_1__60_ = i[56] | i[55];
  assign t_1__59_ = i[57] | i[56];
  assign t_1__58_ = i[58] | i[57];
  assign t_1__57_ = i[59] | i[58];
  assign t_1__56_ = i[60] | i[59];
  assign t_1__55_ = i[61] | i[60];
  assign t_1__54_ = i[62] | i[61];
  assign t_1__53_ = i[63] | i[62];
  assign t_1__52_ = i[64] | i[63];
  assign t_1__51_ = i[65] | i[64];
  assign t_1__50_ = i[66] | i[65];
  assign t_1__49_ = i[67] | i[66];
  assign t_1__48_ = i[68] | i[67];
  assign t_1__47_ = i[69] | i[68];
  assign t_1__46_ = i[70] | i[69];
  assign t_1__45_ = i[71] | i[70];
  assign t_1__44_ = i[72] | i[71];
  assign t_1__43_ = i[73] | i[72];
  assign t_1__42_ = i[74] | i[73];
  assign t_1__41_ = i[75] | i[74];
  assign t_1__40_ = i[76] | i[75];
  assign t_1__39_ = i[77] | i[76];
  assign t_1__38_ = i[78] | i[77];
  assign t_1__37_ = i[79] | i[78];
  assign t_1__36_ = i[80] | i[79];
  assign t_1__35_ = i[81] | i[80];
  assign t_1__34_ = i[82] | i[81];
  assign t_1__33_ = i[83] | i[82];
  assign t_1__32_ = i[84] | i[83];
  assign t_1__31_ = i[85] | i[84];
  assign t_1__30_ = i[86] | i[85];
  assign t_1__29_ = i[87] | i[86];
  assign t_1__28_ = i[88] | i[87];
  assign t_1__27_ = i[89] | i[88];
  assign t_1__26_ = i[90] | i[89];
  assign t_1__25_ = i[91] | i[90];
  assign t_1__24_ = i[92] | i[91];
  assign t_1__23_ = i[93] | i[92];
  assign t_1__22_ = i[94] | i[93];
  assign t_1__21_ = i[95] | i[94];
  assign t_1__20_ = i[96] | i[95];
  assign t_1__19_ = i[97] | i[96];
  assign t_1__18_ = i[98] | i[97];
  assign t_1__17_ = i[99] | i[98];
  assign t_1__16_ = i[100] | i[99];
  assign t_1__15_ = i[101] | i[100];
  assign t_1__14_ = i[102] | i[101];
  assign t_1__13_ = i[103] | i[102];
  assign t_1__12_ = i[104] | i[103];
  assign t_1__11_ = i[105] | i[104];
  assign t_1__10_ = i[106] | i[105];
  assign t_1__9_ = i[107] | i[106];
  assign t_1__8_ = i[108] | i[107];
  assign t_1__7_ = i[109] | i[108];
  assign t_1__6_ = i[110] | i[109];
  assign t_1__5_ = i[111] | i[110];
  assign t_1__4_ = i[112] | i[111];
  assign t_1__3_ = i[113] | i[112];
  assign t_1__2_ = i[114] | i[113];
  assign t_1__1_ = i[115] | i[114];
  assign t_1__0_ = i[116] | i[115];
  assign t_2__116_ = t_1__116_ | 1'b0;
  assign t_2__115_ = t_1__115_ | 1'b0;
  assign t_2__114_ = t_1__114_ | t_1__116_;
  assign t_2__113_ = t_1__113_ | t_1__115_;
  assign t_2__112_ = t_1__112_ | t_1__114_;
  assign t_2__111_ = t_1__111_ | t_1__113_;
  assign t_2__110_ = t_1__110_ | t_1__112_;
  assign t_2__109_ = t_1__109_ | t_1__111_;
  assign t_2__108_ = t_1__108_ | t_1__110_;
  assign t_2__107_ = t_1__107_ | t_1__109_;
  assign t_2__106_ = t_1__106_ | t_1__108_;
  assign t_2__105_ = t_1__105_ | t_1__107_;
  assign t_2__104_ = t_1__104_ | t_1__106_;
  assign t_2__103_ = t_1__103_ | t_1__105_;
  assign t_2__102_ = t_1__102_ | t_1__104_;
  assign t_2__101_ = t_1__101_ | t_1__103_;
  assign t_2__100_ = t_1__100_ | t_1__102_;
  assign t_2__99_ = t_1__99_ | t_1__101_;
  assign t_2__98_ = t_1__98_ | t_1__100_;
  assign t_2__97_ = t_1__97_ | t_1__99_;
  assign t_2__96_ = t_1__96_ | t_1__98_;
  assign t_2__95_ = t_1__95_ | t_1__97_;
  assign t_2__94_ = t_1__94_ | t_1__96_;
  assign t_2__93_ = t_1__93_ | t_1__95_;
  assign t_2__92_ = t_1__92_ | t_1__94_;
  assign t_2__91_ = t_1__91_ | t_1__93_;
  assign t_2__90_ = t_1__90_ | t_1__92_;
  assign t_2__89_ = t_1__89_ | t_1__91_;
  assign t_2__88_ = t_1__88_ | t_1__90_;
  assign t_2__87_ = t_1__87_ | t_1__89_;
  assign t_2__86_ = t_1__86_ | t_1__88_;
  assign t_2__85_ = t_1__85_ | t_1__87_;
  assign t_2__84_ = t_1__84_ | t_1__86_;
  assign t_2__83_ = t_1__83_ | t_1__85_;
  assign t_2__82_ = t_1__82_ | t_1__84_;
  assign t_2__81_ = t_1__81_ | t_1__83_;
  assign t_2__80_ = t_1__80_ | t_1__82_;
  assign t_2__79_ = t_1__79_ | t_1__81_;
  assign t_2__78_ = t_1__78_ | t_1__80_;
  assign t_2__77_ = t_1__77_ | t_1__79_;
  assign t_2__76_ = t_1__76_ | t_1__78_;
  assign t_2__75_ = t_1__75_ | t_1__77_;
  assign t_2__74_ = t_1__74_ | t_1__76_;
  assign t_2__73_ = t_1__73_ | t_1__75_;
  assign t_2__72_ = t_1__72_ | t_1__74_;
  assign t_2__71_ = t_1__71_ | t_1__73_;
  assign t_2__70_ = t_1__70_ | t_1__72_;
  assign t_2__69_ = t_1__69_ | t_1__71_;
  assign t_2__68_ = t_1__68_ | t_1__70_;
  assign t_2__67_ = t_1__67_ | t_1__69_;
  assign t_2__66_ = t_1__66_ | t_1__68_;
  assign t_2__65_ = t_1__65_ | t_1__67_;
  assign t_2__64_ = t_1__64_ | t_1__66_;
  assign t_2__63_ = t_1__63_ | t_1__65_;
  assign t_2__62_ = t_1__62_ | t_1__64_;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__116_ = t_2__116_ | 1'b0;
  assign t_3__115_ = t_2__115_ | 1'b0;
  assign t_3__114_ = t_2__114_ | 1'b0;
  assign t_3__113_ = t_2__113_ | 1'b0;
  assign t_3__112_ = t_2__112_ | t_2__116_;
  assign t_3__111_ = t_2__111_ | t_2__115_;
  assign t_3__110_ = t_2__110_ | t_2__114_;
  assign t_3__109_ = t_2__109_ | t_2__113_;
  assign t_3__108_ = t_2__108_ | t_2__112_;
  assign t_3__107_ = t_2__107_ | t_2__111_;
  assign t_3__106_ = t_2__106_ | t_2__110_;
  assign t_3__105_ = t_2__105_ | t_2__109_;
  assign t_3__104_ = t_2__104_ | t_2__108_;
  assign t_3__103_ = t_2__103_ | t_2__107_;
  assign t_3__102_ = t_2__102_ | t_2__106_;
  assign t_3__101_ = t_2__101_ | t_2__105_;
  assign t_3__100_ = t_2__100_ | t_2__104_;
  assign t_3__99_ = t_2__99_ | t_2__103_;
  assign t_3__98_ = t_2__98_ | t_2__102_;
  assign t_3__97_ = t_2__97_ | t_2__101_;
  assign t_3__96_ = t_2__96_ | t_2__100_;
  assign t_3__95_ = t_2__95_ | t_2__99_;
  assign t_3__94_ = t_2__94_ | t_2__98_;
  assign t_3__93_ = t_2__93_ | t_2__97_;
  assign t_3__92_ = t_2__92_ | t_2__96_;
  assign t_3__91_ = t_2__91_ | t_2__95_;
  assign t_3__90_ = t_2__90_ | t_2__94_;
  assign t_3__89_ = t_2__89_ | t_2__93_;
  assign t_3__88_ = t_2__88_ | t_2__92_;
  assign t_3__87_ = t_2__87_ | t_2__91_;
  assign t_3__86_ = t_2__86_ | t_2__90_;
  assign t_3__85_ = t_2__85_ | t_2__89_;
  assign t_3__84_ = t_2__84_ | t_2__88_;
  assign t_3__83_ = t_2__83_ | t_2__87_;
  assign t_3__82_ = t_2__82_ | t_2__86_;
  assign t_3__81_ = t_2__81_ | t_2__85_;
  assign t_3__80_ = t_2__80_ | t_2__84_;
  assign t_3__79_ = t_2__79_ | t_2__83_;
  assign t_3__78_ = t_2__78_ | t_2__82_;
  assign t_3__77_ = t_2__77_ | t_2__81_;
  assign t_3__76_ = t_2__76_ | t_2__80_;
  assign t_3__75_ = t_2__75_ | t_2__79_;
  assign t_3__74_ = t_2__74_ | t_2__78_;
  assign t_3__73_ = t_2__73_ | t_2__77_;
  assign t_3__72_ = t_2__72_ | t_2__76_;
  assign t_3__71_ = t_2__71_ | t_2__75_;
  assign t_3__70_ = t_2__70_ | t_2__74_;
  assign t_3__69_ = t_2__69_ | t_2__73_;
  assign t_3__68_ = t_2__68_ | t_2__72_;
  assign t_3__67_ = t_2__67_ | t_2__71_;
  assign t_3__66_ = t_2__66_ | t_2__70_;
  assign t_3__65_ = t_2__65_ | t_2__69_;
  assign t_3__64_ = t_2__64_ | t_2__68_;
  assign t_3__63_ = t_2__63_ | t_2__67_;
  assign t_3__62_ = t_2__62_ | t_2__66_;
  assign t_3__61_ = t_2__61_ | t_2__65_;
  assign t_3__60_ = t_2__60_ | t_2__64_;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__116_ = t_3__116_ | 1'b0;
  assign t_4__115_ = t_3__115_ | 1'b0;
  assign t_4__114_ = t_3__114_ | 1'b0;
  assign t_4__113_ = t_3__113_ | 1'b0;
  assign t_4__112_ = t_3__112_ | 1'b0;
  assign t_4__111_ = t_3__111_ | 1'b0;
  assign t_4__110_ = t_3__110_ | 1'b0;
  assign t_4__109_ = t_3__109_ | 1'b0;
  assign t_4__108_ = t_3__108_ | t_3__116_;
  assign t_4__107_ = t_3__107_ | t_3__115_;
  assign t_4__106_ = t_3__106_ | t_3__114_;
  assign t_4__105_ = t_3__105_ | t_3__113_;
  assign t_4__104_ = t_3__104_ | t_3__112_;
  assign t_4__103_ = t_3__103_ | t_3__111_;
  assign t_4__102_ = t_3__102_ | t_3__110_;
  assign t_4__101_ = t_3__101_ | t_3__109_;
  assign t_4__100_ = t_3__100_ | t_3__108_;
  assign t_4__99_ = t_3__99_ | t_3__107_;
  assign t_4__98_ = t_3__98_ | t_3__106_;
  assign t_4__97_ = t_3__97_ | t_3__105_;
  assign t_4__96_ = t_3__96_ | t_3__104_;
  assign t_4__95_ = t_3__95_ | t_3__103_;
  assign t_4__94_ = t_3__94_ | t_3__102_;
  assign t_4__93_ = t_3__93_ | t_3__101_;
  assign t_4__92_ = t_3__92_ | t_3__100_;
  assign t_4__91_ = t_3__91_ | t_3__99_;
  assign t_4__90_ = t_3__90_ | t_3__98_;
  assign t_4__89_ = t_3__89_ | t_3__97_;
  assign t_4__88_ = t_3__88_ | t_3__96_;
  assign t_4__87_ = t_3__87_ | t_3__95_;
  assign t_4__86_ = t_3__86_ | t_3__94_;
  assign t_4__85_ = t_3__85_ | t_3__93_;
  assign t_4__84_ = t_3__84_ | t_3__92_;
  assign t_4__83_ = t_3__83_ | t_3__91_;
  assign t_4__82_ = t_3__82_ | t_3__90_;
  assign t_4__81_ = t_3__81_ | t_3__89_;
  assign t_4__80_ = t_3__80_ | t_3__88_;
  assign t_4__79_ = t_3__79_ | t_3__87_;
  assign t_4__78_ = t_3__78_ | t_3__86_;
  assign t_4__77_ = t_3__77_ | t_3__85_;
  assign t_4__76_ = t_3__76_ | t_3__84_;
  assign t_4__75_ = t_3__75_ | t_3__83_;
  assign t_4__74_ = t_3__74_ | t_3__82_;
  assign t_4__73_ = t_3__73_ | t_3__81_;
  assign t_4__72_ = t_3__72_ | t_3__80_;
  assign t_4__71_ = t_3__71_ | t_3__79_;
  assign t_4__70_ = t_3__70_ | t_3__78_;
  assign t_4__69_ = t_3__69_ | t_3__77_;
  assign t_4__68_ = t_3__68_ | t_3__76_;
  assign t_4__67_ = t_3__67_ | t_3__75_;
  assign t_4__66_ = t_3__66_ | t_3__74_;
  assign t_4__65_ = t_3__65_ | t_3__73_;
  assign t_4__64_ = t_3__64_ | t_3__72_;
  assign t_4__63_ = t_3__63_ | t_3__71_;
  assign t_4__62_ = t_3__62_ | t_3__70_;
  assign t_4__61_ = t_3__61_ | t_3__69_;
  assign t_4__60_ = t_3__60_ | t_3__68_;
  assign t_4__59_ = t_3__59_ | t_3__67_;
  assign t_4__58_ = t_3__58_ | t_3__66_;
  assign t_4__57_ = t_3__57_ | t_3__65_;
  assign t_4__56_ = t_3__56_ | t_3__64_;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__116_ = t_4__116_ | 1'b0;
  assign t_5__115_ = t_4__115_ | 1'b0;
  assign t_5__114_ = t_4__114_ | 1'b0;
  assign t_5__113_ = t_4__113_ | 1'b0;
  assign t_5__112_ = t_4__112_ | 1'b0;
  assign t_5__111_ = t_4__111_ | 1'b0;
  assign t_5__110_ = t_4__110_ | 1'b0;
  assign t_5__109_ = t_4__109_ | 1'b0;
  assign t_5__108_ = t_4__108_ | 1'b0;
  assign t_5__107_ = t_4__107_ | 1'b0;
  assign t_5__106_ = t_4__106_ | 1'b0;
  assign t_5__105_ = t_4__105_ | 1'b0;
  assign t_5__104_ = t_4__104_ | 1'b0;
  assign t_5__103_ = t_4__103_ | 1'b0;
  assign t_5__102_ = t_4__102_ | 1'b0;
  assign t_5__101_ = t_4__101_ | 1'b0;
  assign t_5__100_ = t_4__100_ | t_4__116_;
  assign t_5__99_ = t_4__99_ | t_4__115_;
  assign t_5__98_ = t_4__98_ | t_4__114_;
  assign t_5__97_ = t_4__97_ | t_4__113_;
  assign t_5__96_ = t_4__96_ | t_4__112_;
  assign t_5__95_ = t_4__95_ | t_4__111_;
  assign t_5__94_ = t_4__94_ | t_4__110_;
  assign t_5__93_ = t_4__93_ | t_4__109_;
  assign t_5__92_ = t_4__92_ | t_4__108_;
  assign t_5__91_ = t_4__91_ | t_4__107_;
  assign t_5__90_ = t_4__90_ | t_4__106_;
  assign t_5__89_ = t_4__89_ | t_4__105_;
  assign t_5__88_ = t_4__88_ | t_4__104_;
  assign t_5__87_ = t_4__87_ | t_4__103_;
  assign t_5__86_ = t_4__86_ | t_4__102_;
  assign t_5__85_ = t_4__85_ | t_4__101_;
  assign t_5__84_ = t_4__84_ | t_4__100_;
  assign t_5__83_ = t_4__83_ | t_4__99_;
  assign t_5__82_ = t_4__82_ | t_4__98_;
  assign t_5__81_ = t_4__81_ | t_4__97_;
  assign t_5__80_ = t_4__80_ | t_4__96_;
  assign t_5__79_ = t_4__79_ | t_4__95_;
  assign t_5__78_ = t_4__78_ | t_4__94_;
  assign t_5__77_ = t_4__77_ | t_4__93_;
  assign t_5__76_ = t_4__76_ | t_4__92_;
  assign t_5__75_ = t_4__75_ | t_4__91_;
  assign t_5__74_ = t_4__74_ | t_4__90_;
  assign t_5__73_ = t_4__73_ | t_4__89_;
  assign t_5__72_ = t_4__72_ | t_4__88_;
  assign t_5__71_ = t_4__71_ | t_4__87_;
  assign t_5__70_ = t_4__70_ | t_4__86_;
  assign t_5__69_ = t_4__69_ | t_4__85_;
  assign t_5__68_ = t_4__68_ | t_4__84_;
  assign t_5__67_ = t_4__67_ | t_4__83_;
  assign t_5__66_ = t_4__66_ | t_4__82_;
  assign t_5__65_ = t_4__65_ | t_4__81_;
  assign t_5__64_ = t_4__64_ | t_4__80_;
  assign t_5__63_ = t_4__63_ | t_4__79_;
  assign t_5__62_ = t_4__62_ | t_4__78_;
  assign t_5__61_ = t_4__61_ | t_4__77_;
  assign t_5__60_ = t_4__60_ | t_4__76_;
  assign t_5__59_ = t_4__59_ | t_4__75_;
  assign t_5__58_ = t_4__58_ | t_4__74_;
  assign t_5__57_ = t_4__57_ | t_4__73_;
  assign t_5__56_ = t_4__56_ | t_4__72_;
  assign t_5__55_ = t_4__55_ | t_4__71_;
  assign t_5__54_ = t_4__54_ | t_4__70_;
  assign t_5__53_ = t_4__53_ | t_4__69_;
  assign t_5__52_ = t_4__52_ | t_4__68_;
  assign t_5__51_ = t_4__51_ | t_4__67_;
  assign t_5__50_ = t_4__50_ | t_4__66_;
  assign t_5__49_ = t_4__49_ | t_4__65_;
  assign t_5__48_ = t_4__48_ | t_4__64_;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign t_6__116_ = t_5__116_ | 1'b0;
  assign t_6__115_ = t_5__115_ | 1'b0;
  assign t_6__114_ = t_5__114_ | 1'b0;
  assign t_6__113_ = t_5__113_ | 1'b0;
  assign t_6__112_ = t_5__112_ | 1'b0;
  assign t_6__111_ = t_5__111_ | 1'b0;
  assign t_6__110_ = t_5__110_ | 1'b0;
  assign t_6__109_ = t_5__109_ | 1'b0;
  assign t_6__108_ = t_5__108_ | 1'b0;
  assign t_6__107_ = t_5__107_ | 1'b0;
  assign t_6__106_ = t_5__106_ | 1'b0;
  assign t_6__105_ = t_5__105_ | 1'b0;
  assign t_6__104_ = t_5__104_ | 1'b0;
  assign t_6__103_ = t_5__103_ | 1'b0;
  assign t_6__102_ = t_5__102_ | 1'b0;
  assign t_6__101_ = t_5__101_ | 1'b0;
  assign t_6__100_ = t_5__100_ | 1'b0;
  assign t_6__99_ = t_5__99_ | 1'b0;
  assign t_6__98_ = t_5__98_ | 1'b0;
  assign t_6__97_ = t_5__97_ | 1'b0;
  assign t_6__96_ = t_5__96_ | 1'b0;
  assign t_6__95_ = t_5__95_ | 1'b0;
  assign t_6__94_ = t_5__94_ | 1'b0;
  assign t_6__93_ = t_5__93_ | 1'b0;
  assign t_6__92_ = t_5__92_ | 1'b0;
  assign t_6__91_ = t_5__91_ | 1'b0;
  assign t_6__90_ = t_5__90_ | 1'b0;
  assign t_6__89_ = t_5__89_ | 1'b0;
  assign t_6__88_ = t_5__88_ | 1'b0;
  assign t_6__87_ = t_5__87_ | 1'b0;
  assign t_6__86_ = t_5__86_ | 1'b0;
  assign t_6__85_ = t_5__85_ | 1'b0;
  assign t_6__84_ = t_5__84_ | t_5__116_;
  assign t_6__83_ = t_5__83_ | t_5__115_;
  assign t_6__82_ = t_5__82_ | t_5__114_;
  assign t_6__81_ = t_5__81_ | t_5__113_;
  assign t_6__80_ = t_5__80_ | t_5__112_;
  assign t_6__79_ = t_5__79_ | t_5__111_;
  assign t_6__78_ = t_5__78_ | t_5__110_;
  assign t_6__77_ = t_5__77_ | t_5__109_;
  assign t_6__76_ = t_5__76_ | t_5__108_;
  assign t_6__75_ = t_5__75_ | t_5__107_;
  assign t_6__74_ = t_5__74_ | t_5__106_;
  assign t_6__73_ = t_5__73_ | t_5__105_;
  assign t_6__72_ = t_5__72_ | t_5__104_;
  assign t_6__71_ = t_5__71_ | t_5__103_;
  assign t_6__70_ = t_5__70_ | t_5__102_;
  assign t_6__69_ = t_5__69_ | t_5__101_;
  assign t_6__68_ = t_5__68_ | t_5__100_;
  assign t_6__67_ = t_5__67_ | t_5__99_;
  assign t_6__66_ = t_5__66_ | t_5__98_;
  assign t_6__65_ = t_5__65_ | t_5__97_;
  assign t_6__64_ = t_5__64_ | t_5__96_;
  assign t_6__63_ = t_5__63_ | t_5__95_;
  assign t_6__62_ = t_5__62_ | t_5__94_;
  assign t_6__61_ = t_5__61_ | t_5__93_;
  assign t_6__60_ = t_5__60_ | t_5__92_;
  assign t_6__59_ = t_5__59_ | t_5__91_;
  assign t_6__58_ = t_5__58_ | t_5__90_;
  assign t_6__57_ = t_5__57_ | t_5__89_;
  assign t_6__56_ = t_5__56_ | t_5__88_;
  assign t_6__55_ = t_5__55_ | t_5__87_;
  assign t_6__54_ = t_5__54_ | t_5__86_;
  assign t_6__53_ = t_5__53_ | t_5__85_;
  assign t_6__52_ = t_5__52_ | t_5__84_;
  assign t_6__51_ = t_5__51_ | t_5__83_;
  assign t_6__50_ = t_5__50_ | t_5__82_;
  assign t_6__49_ = t_5__49_ | t_5__81_;
  assign t_6__48_ = t_5__48_ | t_5__80_;
  assign t_6__47_ = t_5__47_ | t_5__79_;
  assign t_6__46_ = t_5__46_ | t_5__78_;
  assign t_6__45_ = t_5__45_ | t_5__77_;
  assign t_6__44_ = t_5__44_ | t_5__76_;
  assign t_6__43_ = t_5__43_ | t_5__75_;
  assign t_6__42_ = t_5__42_ | t_5__74_;
  assign t_6__41_ = t_5__41_ | t_5__73_;
  assign t_6__40_ = t_5__40_ | t_5__72_;
  assign t_6__39_ = t_5__39_ | t_5__71_;
  assign t_6__38_ = t_5__38_ | t_5__70_;
  assign t_6__37_ = t_5__37_ | t_5__69_;
  assign t_6__36_ = t_5__36_ | t_5__68_;
  assign t_6__35_ = t_5__35_ | t_5__67_;
  assign t_6__34_ = t_5__34_ | t_5__66_;
  assign t_6__33_ = t_5__33_ | t_5__65_;
  assign t_6__32_ = t_5__32_ | t_5__64_;
  assign t_6__31_ = t_5__31_ | t_5__63_;
  assign t_6__30_ = t_5__30_ | t_5__62_;
  assign t_6__29_ = t_5__29_ | t_5__61_;
  assign t_6__28_ = t_5__28_ | t_5__60_;
  assign t_6__27_ = t_5__27_ | t_5__59_;
  assign t_6__26_ = t_5__26_ | t_5__58_;
  assign t_6__25_ = t_5__25_ | t_5__57_;
  assign t_6__24_ = t_5__24_ | t_5__56_;
  assign t_6__23_ = t_5__23_ | t_5__55_;
  assign t_6__22_ = t_5__22_ | t_5__54_;
  assign t_6__21_ = t_5__21_ | t_5__53_;
  assign t_6__20_ = t_5__20_ | t_5__52_;
  assign t_6__19_ = t_5__19_ | t_5__51_;
  assign t_6__18_ = t_5__18_ | t_5__50_;
  assign t_6__17_ = t_5__17_ | t_5__49_;
  assign t_6__16_ = t_5__16_ | t_5__48_;
  assign t_6__15_ = t_5__15_ | t_5__47_;
  assign t_6__14_ = t_5__14_ | t_5__46_;
  assign t_6__13_ = t_5__13_ | t_5__45_;
  assign t_6__12_ = t_5__12_ | t_5__44_;
  assign t_6__11_ = t_5__11_ | t_5__43_;
  assign t_6__10_ = t_5__10_ | t_5__42_;
  assign t_6__9_ = t_5__9_ | t_5__41_;
  assign t_6__8_ = t_5__8_ | t_5__40_;
  assign t_6__7_ = t_5__7_ | t_5__39_;
  assign t_6__6_ = t_5__6_ | t_5__38_;
  assign t_6__5_ = t_5__5_ | t_5__37_;
  assign t_6__4_ = t_5__4_ | t_5__36_;
  assign t_6__3_ = t_5__3_ | t_5__35_;
  assign t_6__2_ = t_5__2_ | t_5__34_;
  assign t_6__1_ = t_5__1_ | t_5__33_;
  assign t_6__0_ = t_5__0_ | t_5__32_;
  assign o[0] = t_6__116_ | 1'b0;
  assign o[1] = t_6__115_ | 1'b0;
  assign o[2] = t_6__114_ | 1'b0;
  assign o[3] = t_6__113_ | 1'b0;
  assign o[4] = t_6__112_ | 1'b0;
  assign o[5] = t_6__111_ | 1'b0;
  assign o[6] = t_6__110_ | 1'b0;
  assign o[7] = t_6__109_ | 1'b0;
  assign o[8] = t_6__108_ | 1'b0;
  assign o[9] = t_6__107_ | 1'b0;
  assign o[10] = t_6__106_ | 1'b0;
  assign o[11] = t_6__105_ | 1'b0;
  assign o[12] = t_6__104_ | 1'b0;
  assign o[13] = t_6__103_ | 1'b0;
  assign o[14] = t_6__102_ | 1'b0;
  assign o[15] = t_6__101_ | 1'b0;
  assign o[16] = t_6__100_ | 1'b0;
  assign o[17] = t_6__99_ | 1'b0;
  assign o[18] = t_6__98_ | 1'b0;
  assign o[19] = t_6__97_ | 1'b0;
  assign o[20] = t_6__96_ | 1'b0;
  assign o[21] = t_6__95_ | 1'b0;
  assign o[22] = t_6__94_ | 1'b0;
  assign o[23] = t_6__93_ | 1'b0;
  assign o[24] = t_6__92_ | 1'b0;
  assign o[25] = t_6__91_ | 1'b0;
  assign o[26] = t_6__90_ | 1'b0;
  assign o[27] = t_6__89_ | 1'b0;
  assign o[28] = t_6__88_ | 1'b0;
  assign o[29] = t_6__87_ | 1'b0;
  assign o[30] = t_6__86_ | 1'b0;
  assign o[31] = t_6__85_ | 1'b0;
  assign o[32] = t_6__84_ | 1'b0;
  assign o[33] = t_6__83_ | 1'b0;
  assign o[34] = t_6__82_ | 1'b0;
  assign o[35] = t_6__81_ | 1'b0;
  assign o[36] = t_6__80_ | 1'b0;
  assign o[37] = t_6__79_ | 1'b0;
  assign o[38] = t_6__78_ | 1'b0;
  assign o[39] = t_6__77_ | 1'b0;
  assign o[40] = t_6__76_ | 1'b0;
  assign o[41] = t_6__75_ | 1'b0;
  assign o[42] = t_6__74_ | 1'b0;
  assign o[43] = t_6__73_ | 1'b0;
  assign o[44] = t_6__72_ | 1'b0;
  assign o[45] = t_6__71_ | 1'b0;
  assign o[46] = t_6__70_ | 1'b0;
  assign o[47] = t_6__69_ | 1'b0;
  assign o[48] = t_6__68_ | 1'b0;
  assign o[49] = t_6__67_ | 1'b0;
  assign o[50] = t_6__66_ | 1'b0;
  assign o[51] = t_6__65_ | 1'b0;
  assign o[52] = t_6__64_ | 1'b0;
  assign o[53] = t_6__63_ | 1'b0;
  assign o[54] = t_6__62_ | 1'b0;
  assign o[55] = t_6__61_ | 1'b0;
  assign o[56] = t_6__60_ | 1'b0;
  assign o[57] = t_6__59_ | 1'b0;
  assign o[58] = t_6__58_ | 1'b0;
  assign o[59] = t_6__57_ | 1'b0;
  assign o[60] = t_6__56_ | 1'b0;
  assign o[61] = t_6__55_ | 1'b0;
  assign o[62] = t_6__54_ | 1'b0;
  assign o[63] = t_6__53_ | 1'b0;
  assign o[64] = t_6__52_ | t_6__116_;
  assign o[65] = t_6__51_ | t_6__115_;
  assign o[66] = t_6__50_ | t_6__114_;
  assign o[67] = t_6__49_ | t_6__113_;
  assign o[68] = t_6__48_ | t_6__112_;
  assign o[69] = t_6__47_ | t_6__111_;
  assign o[70] = t_6__46_ | t_6__110_;
  assign o[71] = t_6__45_ | t_6__109_;
  assign o[72] = t_6__44_ | t_6__108_;
  assign o[73] = t_6__43_ | t_6__107_;
  assign o[74] = t_6__42_ | t_6__106_;
  assign o[75] = t_6__41_ | t_6__105_;
  assign o[76] = t_6__40_ | t_6__104_;
  assign o[77] = t_6__39_ | t_6__103_;
  assign o[78] = t_6__38_ | t_6__102_;
  assign o[79] = t_6__37_ | t_6__101_;
  assign o[80] = t_6__36_ | t_6__100_;
  assign o[81] = t_6__35_ | t_6__99_;
  assign o[82] = t_6__34_ | t_6__98_;
  assign o[83] = t_6__33_ | t_6__97_;
  assign o[84] = t_6__32_ | t_6__96_;
  assign o[85] = t_6__31_ | t_6__95_;
  assign o[86] = t_6__30_ | t_6__94_;
  assign o[87] = t_6__29_ | t_6__93_;
  assign o[88] = t_6__28_ | t_6__92_;
  assign o[89] = t_6__27_ | t_6__91_;
  assign o[90] = t_6__26_ | t_6__90_;
  assign o[91] = t_6__25_ | t_6__89_;
  assign o[92] = t_6__24_ | t_6__88_;
  assign o[93] = t_6__23_ | t_6__87_;
  assign o[94] = t_6__22_ | t_6__86_;
  assign o[95] = t_6__21_ | t_6__85_;
  assign o[96] = t_6__20_ | t_6__84_;
  assign o[97] = t_6__19_ | t_6__83_;
  assign o[98] = t_6__18_ | t_6__82_;
  assign o[99] = t_6__17_ | t_6__81_;
  assign o[100] = t_6__16_ | t_6__80_;
  assign o[101] = t_6__15_ | t_6__79_;
  assign o[102] = t_6__14_ | t_6__78_;
  assign o[103] = t_6__13_ | t_6__77_;
  assign o[104] = t_6__12_ | t_6__76_;
  assign o[105] = t_6__11_ | t_6__75_;
  assign o[106] = t_6__10_ | t_6__74_;
  assign o[107] = t_6__9_ | t_6__73_;
  assign o[108] = t_6__8_ | t_6__72_;
  assign o[109] = t_6__7_ | t_6__71_;
  assign o[110] = t_6__6_ | t_6__70_;
  assign o[111] = t_6__5_ | t_6__69_;
  assign o[112] = t_6__4_ | t_6__68_;
  assign o[113] = t_6__3_ | t_6__67_;
  assign o[114] = t_6__2_ | t_6__66_;
  assign o[115] = t_6__1_ | t_6__65_;
  assign o[116] = t_6__0_ | t_6__64_;

endmodule



module bsg_priority_encode_one_hot_out_width_p117_lo_to_hi_p1
(
  i,
  o
);

  input [116:0] i;
  output [116:0] o;
  wire [116:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115;
  wire [116:1] scan_lo;

  bsg_scan_width_p117_or_p1_lo_to_hi_p1
  genblk1_scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[116] = scan_lo[116] & N0;
  assign N0 = ~scan_lo[115];
  assign o[115] = scan_lo[115] & N1;
  assign N1 = ~scan_lo[114];
  assign o[114] = scan_lo[114] & N2;
  assign N2 = ~scan_lo[113];
  assign o[113] = scan_lo[113] & N3;
  assign N3 = ~scan_lo[112];
  assign o[112] = scan_lo[112] & N4;
  assign N4 = ~scan_lo[111];
  assign o[111] = scan_lo[111] & N5;
  assign N5 = ~scan_lo[110];
  assign o[110] = scan_lo[110] & N6;
  assign N6 = ~scan_lo[109];
  assign o[109] = scan_lo[109] & N7;
  assign N7 = ~scan_lo[108];
  assign o[108] = scan_lo[108] & N8;
  assign N8 = ~scan_lo[107];
  assign o[107] = scan_lo[107] & N9;
  assign N9 = ~scan_lo[106];
  assign o[106] = scan_lo[106] & N10;
  assign N10 = ~scan_lo[105];
  assign o[105] = scan_lo[105] & N11;
  assign N11 = ~scan_lo[104];
  assign o[104] = scan_lo[104] & N12;
  assign N12 = ~scan_lo[103];
  assign o[103] = scan_lo[103] & N13;
  assign N13 = ~scan_lo[102];
  assign o[102] = scan_lo[102] & N14;
  assign N14 = ~scan_lo[101];
  assign o[101] = scan_lo[101] & N15;
  assign N15 = ~scan_lo[100];
  assign o[100] = scan_lo[100] & N16;
  assign N16 = ~scan_lo[99];
  assign o[99] = scan_lo[99] & N17;
  assign N17 = ~scan_lo[98];
  assign o[98] = scan_lo[98] & N18;
  assign N18 = ~scan_lo[97];
  assign o[97] = scan_lo[97] & N19;
  assign N19 = ~scan_lo[96];
  assign o[96] = scan_lo[96] & N20;
  assign N20 = ~scan_lo[95];
  assign o[95] = scan_lo[95] & N21;
  assign N21 = ~scan_lo[94];
  assign o[94] = scan_lo[94] & N22;
  assign N22 = ~scan_lo[93];
  assign o[93] = scan_lo[93] & N23;
  assign N23 = ~scan_lo[92];
  assign o[92] = scan_lo[92] & N24;
  assign N24 = ~scan_lo[91];
  assign o[91] = scan_lo[91] & N25;
  assign N25 = ~scan_lo[90];
  assign o[90] = scan_lo[90] & N26;
  assign N26 = ~scan_lo[89];
  assign o[89] = scan_lo[89] & N27;
  assign N27 = ~scan_lo[88];
  assign o[88] = scan_lo[88] & N28;
  assign N28 = ~scan_lo[87];
  assign o[87] = scan_lo[87] & N29;
  assign N29 = ~scan_lo[86];
  assign o[86] = scan_lo[86] & N30;
  assign N30 = ~scan_lo[85];
  assign o[85] = scan_lo[85] & N31;
  assign N31 = ~scan_lo[84];
  assign o[84] = scan_lo[84] & N32;
  assign N32 = ~scan_lo[83];
  assign o[83] = scan_lo[83] & N33;
  assign N33 = ~scan_lo[82];
  assign o[82] = scan_lo[82] & N34;
  assign N34 = ~scan_lo[81];
  assign o[81] = scan_lo[81] & N35;
  assign N35 = ~scan_lo[80];
  assign o[80] = scan_lo[80] & N36;
  assign N36 = ~scan_lo[79];
  assign o[79] = scan_lo[79] & N37;
  assign N37 = ~scan_lo[78];
  assign o[78] = scan_lo[78] & N38;
  assign N38 = ~scan_lo[77];
  assign o[77] = scan_lo[77] & N39;
  assign N39 = ~scan_lo[76];
  assign o[76] = scan_lo[76] & N40;
  assign N40 = ~scan_lo[75];
  assign o[75] = scan_lo[75] & N41;
  assign N41 = ~scan_lo[74];
  assign o[74] = scan_lo[74] & N42;
  assign N42 = ~scan_lo[73];
  assign o[73] = scan_lo[73] & N43;
  assign N43 = ~scan_lo[72];
  assign o[72] = scan_lo[72] & N44;
  assign N44 = ~scan_lo[71];
  assign o[71] = scan_lo[71] & N45;
  assign N45 = ~scan_lo[70];
  assign o[70] = scan_lo[70] & N46;
  assign N46 = ~scan_lo[69];
  assign o[69] = scan_lo[69] & N47;
  assign N47 = ~scan_lo[68];
  assign o[68] = scan_lo[68] & N48;
  assign N48 = ~scan_lo[67];
  assign o[67] = scan_lo[67] & N49;
  assign N49 = ~scan_lo[66];
  assign o[66] = scan_lo[66] & N50;
  assign N50 = ~scan_lo[65];
  assign o[65] = scan_lo[65] & N51;
  assign N51 = ~scan_lo[64];
  assign o[64] = scan_lo[64] & N52;
  assign N52 = ~scan_lo[63];
  assign o[63] = scan_lo[63] & N53;
  assign N53 = ~scan_lo[62];
  assign o[62] = scan_lo[62] & N54;
  assign N54 = ~scan_lo[61];
  assign o[61] = scan_lo[61] & N55;
  assign N55 = ~scan_lo[60];
  assign o[60] = scan_lo[60] & N56;
  assign N56 = ~scan_lo[59];
  assign o[59] = scan_lo[59] & N57;
  assign N57 = ~scan_lo[58];
  assign o[58] = scan_lo[58] & N58;
  assign N58 = ~scan_lo[57];
  assign o[57] = scan_lo[57] & N59;
  assign N59 = ~scan_lo[56];
  assign o[56] = scan_lo[56] & N60;
  assign N60 = ~scan_lo[55];
  assign o[55] = scan_lo[55] & N61;
  assign N61 = ~scan_lo[54];
  assign o[54] = scan_lo[54] & N62;
  assign N62 = ~scan_lo[53];
  assign o[53] = scan_lo[53] & N63;
  assign N63 = ~scan_lo[52];
  assign o[52] = scan_lo[52] & N64;
  assign N64 = ~scan_lo[51];
  assign o[51] = scan_lo[51] & N65;
  assign N65 = ~scan_lo[50];
  assign o[50] = scan_lo[50] & N66;
  assign N66 = ~scan_lo[49];
  assign o[49] = scan_lo[49] & N67;
  assign N67 = ~scan_lo[48];
  assign o[48] = scan_lo[48] & N68;
  assign N68 = ~scan_lo[47];
  assign o[47] = scan_lo[47] & N69;
  assign N69 = ~scan_lo[46];
  assign o[46] = scan_lo[46] & N70;
  assign N70 = ~scan_lo[45];
  assign o[45] = scan_lo[45] & N71;
  assign N71 = ~scan_lo[44];
  assign o[44] = scan_lo[44] & N72;
  assign N72 = ~scan_lo[43];
  assign o[43] = scan_lo[43] & N73;
  assign N73 = ~scan_lo[42];
  assign o[42] = scan_lo[42] & N74;
  assign N74 = ~scan_lo[41];
  assign o[41] = scan_lo[41] & N75;
  assign N75 = ~scan_lo[40];
  assign o[40] = scan_lo[40] & N76;
  assign N76 = ~scan_lo[39];
  assign o[39] = scan_lo[39] & N77;
  assign N77 = ~scan_lo[38];
  assign o[38] = scan_lo[38] & N78;
  assign N78 = ~scan_lo[37];
  assign o[37] = scan_lo[37] & N79;
  assign N79 = ~scan_lo[36];
  assign o[36] = scan_lo[36] & N80;
  assign N80 = ~scan_lo[35];
  assign o[35] = scan_lo[35] & N81;
  assign N81 = ~scan_lo[34];
  assign o[34] = scan_lo[34] & N82;
  assign N82 = ~scan_lo[33];
  assign o[33] = scan_lo[33] & N83;
  assign N83 = ~scan_lo[32];
  assign o[32] = scan_lo[32] & N84;
  assign N84 = ~scan_lo[31];
  assign o[31] = scan_lo[31] & N85;
  assign N85 = ~scan_lo[30];
  assign o[30] = scan_lo[30] & N86;
  assign N86 = ~scan_lo[29];
  assign o[29] = scan_lo[29] & N87;
  assign N87 = ~scan_lo[28];
  assign o[28] = scan_lo[28] & N88;
  assign N88 = ~scan_lo[27];
  assign o[27] = scan_lo[27] & N89;
  assign N89 = ~scan_lo[26];
  assign o[26] = scan_lo[26] & N90;
  assign N90 = ~scan_lo[25];
  assign o[25] = scan_lo[25] & N91;
  assign N91 = ~scan_lo[24];
  assign o[24] = scan_lo[24] & N92;
  assign N92 = ~scan_lo[23];
  assign o[23] = scan_lo[23] & N93;
  assign N93 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N94;
  assign N94 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N95;
  assign N95 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N96;
  assign N96 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N97;
  assign N97 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N98;
  assign N98 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N99;
  assign N99 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N100;
  assign N100 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N101;
  assign N101 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N102;
  assign N102 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N103;
  assign N103 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N104;
  assign N104 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N105;
  assign N105 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N106;
  assign N106 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N107;
  assign N107 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N108;
  assign N108 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N109;
  assign N109 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N110;
  assign N110 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N111;
  assign N111 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N112;
  assign N112 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N113;
  assign N113 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N114;
  assign N114 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N115;
  assign N115 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_encode_one_hot_width_p16
(
  i,
  addr_o,
  v_o
);

  input [15:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;
  wire [5:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p8
  aligned_left
  (
    .i(i[7:0]),
    .addr_o(aligned_addrs[2:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p8
  aligned_right
  (
    .i(i[15:8]),
    .addr_o(aligned_addrs[5:3]),
    .v_o(addr_o[3])
  );

  assign v_o = addr_o[3] | aligned_vs[0];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[5];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[4];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[3];

endmodule



module bsg_encode_one_hot_width_p32
(
  i,
  addr_o,
  v_o
);

  input [31:0] i;
  output [4:0] addr_o;
  output v_o;
  wire [4:0] addr_o;
  wire v_o;
  wire [7:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p16
  aligned_left
  (
    .i(i[15:0]),
    .addr_o(aligned_addrs[3:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p16
  aligned_right
  (
    .i(i[31:16]),
    .addr_o(aligned_addrs[7:4]),
    .v_o(addr_o[4])
  );

  assign v_o = addr_o[4] | aligned_vs[0];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[7];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[6];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[5];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[4];

endmodule



module bsg_encode_one_hot_width_p64
(
  i,
  addr_o,
  v_o
);

  input [63:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o;
  wire [9:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p32
  aligned_left
  (
    .i(i[31:0]),
    .addr_o(aligned_addrs[4:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p32
  aligned_right
  (
    .i(i[63:32]),
    .addr_o(aligned_addrs[9:5]),
    .v_o(addr_o[5])
  );

  assign v_o = addr_o[5] | aligned_vs[0];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[9];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[8];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[7];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[6];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[5];

endmodule



module bsg_encode_one_hot_width_p128
(
  i,
  addr_o,
  v_o
);

  input [127:0] i;
  output [6:0] addr_o;
  output v_o;
  wire [6:0] addr_o;
  wire v_o;
  wire [11:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p64
  aligned_left
  (
    .i(i[63:0]),
    .addr_o(aligned_addrs[5:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p64
  aligned_right
  (
    .i(i[127:64]),
    .addr_o(aligned_addrs[11:6]),
    .v_o(addr_o[6])
  );

  assign v_o = addr_o[6] | aligned_vs[0];
  assign addr_o[5] = aligned_addrs[5] | aligned_addrs[11];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[10];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[9];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[8];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[7];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[6];

endmodule



module bsg_encode_one_hot_width_p117_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [116:0] i;
  output [6:0] addr_o;
  output v_o;
  wire [6:0] addr_o;
  wire v_o;

  bsg_encode_one_hot_width_p128
  unaligned_align
  (
    .i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, i }),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_priority_encode_width_p117_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [116:0] i;
  output [6:0] addr_o;
  output v_o;
  wire [6:0] addr_o;
  wire v_o;
  wire [116:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p117_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p117_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_fpu_clz_width_p117
(
  i,
  num_zero_o
);

  input [116:0] i;
  output [6:0] num_zero_o;
  wire [6:0] num_zero_o;

  bsg_priority_encode_width_p117_lo_to_hi_p1
  pe0
  (
    .i({ i[0:0], i[1:1], i[2:2], i[3:3], i[4:4], i[5:5], i[6:6], i[7:7], i[8:8], i[9:9], i[10:10], i[11:11], i[12:12], i[13:13], i[14:14], i[15:15], i[16:16], i[17:17], i[18:18], i[19:19], i[20:20], i[21:21], i[22:22], i[23:23], i[24:24], i[25:25], i[26:26], i[27:27], i[28:28], i[29:29], i[30:30], i[31:31], i[32:32], i[33:33], i[34:34], i[35:35], i[36:36], i[37:37], i[38:38], i[39:39], i[40:40], i[41:41], i[42:42], i[43:43], i[44:44], i[45:45], i[46:46], i[47:47], i[48:48], i[49:49], i[50:50], i[51:51], i[52:52], i[53:53], i[54:54], i[55:55], i[56:56], i[57:57], i[58:58], i[59:59], i[60:60], i[61:61], i[62:62], i[63:63], i[64:64], i[65:65], i[66:66], i[67:67], i[68:68], i[69:69], i[70:70], i[71:71], i[72:72], i[73:73], i[74:74], i[75:75], i[76:76], i[77:77], i[78:78], i[79:79], i[80:80], i[81:81], i[82:82], i[83:83], i[84:84], i[85:85], i[86:86], i[87:87], i[88:88], i[89:89], i[90:90], i[91:91], i[92:92], i[93:93], i[94:94], i[95:95], i[96:96], i[97:97], i[98:98], i[99:99], i[100:100], i[101:101], i[102:102], i[103:103], i[104:104], i[105:105], i[106:106], i[107:107], i[108:108], i[109:109], i[110:110], i[111:111], i[112:112], i[113:113], i[114:114], i[115:115], i[116:116] }),
    .addr_o(num_zero_o)
  );


endmodule



module bsg_fpu_add_sub
(
  clk_i,
  reset_i,
  en_i,
  v_i,
  a_i,
  b_i,
  sub_i,
  ready_o,
  v_o,
  z_o,
  unimplemented_o,
  invalid_o,
  overflow_o,
  underflow_o,
  yumi_i
);

  input [127:0] a_i;
  input [127:0] b_i;
  output [127:0] z_o;
  input clk_i;
  input reset_i;
  input en_i;
  input v_i;
  input sub_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output unimplemented_o;
  output invalid_o;
  output overflow_o;
  output underflow_o;
  wire [127:0] z_o;
  wire ready_o,unimplemented_o,invalid_o,overflow_o,underflow_o,N0,N1,N2,N3,N4,N5,N6,
  N7,N8,N9,stall,a_zero,a_nan,a_sig_nan,a_infty,exp_a_zero,a_denormal,sign_a,b_zero,
  b_nan,b_sig_nan,b_infty,exp_b_zero,b_denormal,sign_b,exp_a_less,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,mag_a_less,final_sign,do_sub,
  N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,larger_exp_man_less,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,
  N277,reduce_o,all_zero,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,adjusted_exp_cout,round_up,N395,
  N396,N397,N398,N399,N400,N401,N402,carry_into_exp,N403,N404,N405,N406,N407,N408,
  N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,
  N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,
  N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,
  N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,
  N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,
  N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,
  N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,
  N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,
  N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,
  N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,
  N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,
  N601,N602,N603,N604,N605,N606,N607;
  wire [14:0] exp_a,exp_b,larger_exp,diff_ab,diff_ba,exp_diff,adjusted_exp;
  wire [111:0] man_a,man_b,larger_exp_man,smaller_exp_man;
  wire [115:0] smaller_exp_man_shifted,larger_mag_man,smaller_mag_man,shifted_adder_output;
  wire [116:0] adder_output;
  wire [6:0] num_zero;
  wire [126:0] rounded;
  reg a_denormal_1_r,v_1_r,b_denormal_1_r,final_sign_1_r,do_sub_1_r,a_sig_nan_1_r,
  b_sig_nan_1_r,a_nan_1_r,b_nan_1_r,a_infty_1_r,b_infty_1_r,a_denormal_2_r,v_2_r,
  b_denormal_2_r,final_sign_2_r,do_sub_2_r,a_sig_nan_2_r,b_sig_nan_2_r,a_nan_2_r,
  b_nan_2_r,a_infty_2_r,b_infty_2_r,adjusted_exp_cout_3_r,v_o,final_sign_3_r,
  round_up_3_r,all_zero_3_r,a_sig_nan_3_r,b_sig_nan_3_r,a_nan_3_r,b_nan_3_r,a_infty_3_r,
  b_infty_3_r,do_sub_3_r,a_denormal_3_r,b_denormal_3_r;
  reg [14:0] larger_exp_1_r,larger_exp_2_r;
  reg [115:0] smaller_exp_man_shifted_1_r,larger_exp_man_padded_1_r;
  reg [116:0] adder_output_2_r;
  reg [126:0] pre_roundup_3_r;

  bsg_fpu_preprocess_e_p15_m_p112
  a_preprocess
  (
    .a_i(a_i),
    .zero_o(a_zero),
    .nan_o(a_nan),
    .sig_nan_o(a_sig_nan),
    .infty_o(a_infty),
    .exp_zero_o(exp_a_zero),
    .denormal_o(a_denormal),
    .sign_o(sign_a),
    .exp_o(exp_a),
    .man_o(man_a)
  );


  bsg_fpu_preprocess_e_p15_m_p112
  b_preprocess
  (
    .a_i(b_i),
    .zero_o(b_zero),
    .nan_o(b_nan),
    .sig_nan_o(b_sig_nan),
    .infty_o(b_infty),
    .exp_zero_o(exp_b_zero),
    .denormal_o(b_denormal),
    .sign_o(sign_b),
    .exp_o(exp_b),
    .man_o(man_b)
  );


  bsg_less_than_width_p15
  lt_exp
  (
    .a_i(exp_a),
    .b_i(exp_b),
    .o(exp_a_less)
  );


  bsg_fpu_sticky_width_p115
  sticky0
  (
    .i({ 1'b1, smaller_exp_man, 1'b0, 1'b0 }),
    .shamt_i(exp_diff[6:0]),
    .sticky_o(smaller_exp_man_shifted[0])
  );


  bsg_less_than_width_p127
  lt_mag
  (
    .a_i(a_i[126:0]),
    .b_i(b_i[126:0]),
    .o(mag_a_less)
  );

  assign smaller_exp_man_shifted[115:1] = { 1'b1, smaller_exp_man, 1'b0, 1'b0 } >> exp_diff;

  bsg_less_than_width_p116
  lt_man_norm
  (
    .a_i(larger_exp_man_padded_1_r),
    .b_i(smaller_exp_man_shifted_1_r),
    .o(larger_exp_man_less)
  );


  bsg_fpu_clz_width_p117
  clz
  (
    .i(adder_output_2_r),
    .num_zero_o(num_zero)
  );


  bsg_reduce
  reduce0
  (
    .i(adder_output_2_r),
    .o(reduce_o)
  );

  assign N449 = pre_roundup_3_r[125] | pre_roundup_3_r[126];
  assign N450 = pre_roundup_3_r[124] | N449;
  assign N451 = pre_roundup_3_r[123] | N450;
  assign N452 = pre_roundup_3_r[122] | N451;
  assign N453 = pre_roundup_3_r[121] | N452;
  assign N454 = pre_roundup_3_r[120] | N453;
  assign N455 = pre_roundup_3_r[119] | N454;
  assign N456 = pre_roundup_3_r[118] | N455;
  assign N457 = pre_roundup_3_r[117] | N456;
  assign N458 = pre_roundup_3_r[116] | N457;
  assign N459 = pre_roundup_3_r[115] | N458;
  assign N460 = pre_roundup_3_r[114] | N459;
  assign N461 = pre_roundup_3_r[113] | N460;
  assign N462 = pre_roundup_3_r[112] | N461;
  assign N463 = ~N462;
  assign { N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279 } = adder_output_2_r[115:0] << num_zero;
  assign N464 = pre_roundup_3_r[125] & pre_roundup_3_r[126];
  assign N465 = pre_roundup_3_r[124] & N464;
  assign N466 = pre_roundup_3_r[123] & N465;
  assign N467 = pre_roundup_3_r[122] & N466;
  assign N468 = pre_roundup_3_r[121] & N467;
  assign N469 = pre_roundup_3_r[120] & N468;
  assign N470 = pre_roundup_3_r[119] & N469;
  assign N471 = pre_roundup_3_r[118] & N470;
  assign N472 = pre_roundup_3_r[117] & N471;
  assign N473 = pre_roundup_3_r[116] & N472;
  assign N474 = pre_roundup_3_r[115] & N473;
  assign N475 = pre_roundup_3_r[114] & N474;
  assign N476 = pre_roundup_3_r[113] & N475;
  assign N477 = pre_roundup_3_r[112] & N476;
  assign rounded = pre_roundup_3_r + round_up_3_r;
  assign { adjusted_exp_cout, adjusted_exp } = larger_exp_2_r - num_zero;
  assign diff_ba = exp_b - exp_a;
  assign diff_ab = exp_a - exp_b;
  assign larger_exp = { N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11 } + 1'b1;
  assign { N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153 } = larger_mag_man + { do_sub_1_r, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152 };
  assign adder_output = { N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153 } + do_sub_1_r;
  assign { N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11 } = (N0)? exp_b : 
                                                                                         (N1)? exp_a : 1'b0;
  assign N0 = exp_a_less;
  assign N1 = N10;
  assign exp_diff = (N0)? diff_ba : 
                    (N1)? diff_ab : 1'b0;
  assign larger_exp_man = (N0)? man_b : 
                          (N1)? man_a : 1'b0;
  assign smaller_exp_man = (N0)? man_a : 
                           (N1)? man_b : 1'b0;
  assign N29 = (N2)? 1'b1 : 
               (N35)? 1'b1 : 
               (N28)? 1'b0 : 1'b0;
  assign N2 = reset_i;
  assign N30 = (N2)? 1'b0 : 
               (N35)? v_i : 1'b0;
  assign N31 = (N2)? 1'b0 : 
               (N35)? v_i : 
               (N28)? 1'b0 : 1'b0;
  assign N32 = (N2)? 1'b0 : 
               (N35)? v_i : 
               (N28)? 1'b0 : 1'b0;
  assign N33 = (N2)? 1'b0 : 
               (N35)? v_i : 
               (N28)? 1'b0 : 1'b0;
  assign larger_mag_man = (N3)? smaller_exp_man_shifted_1_r : 
                          (N4)? larger_exp_man_padded_1_r : 1'b0;
  assign N3 = larger_exp_man_less;
  assign N4 = N36;
  assign smaller_mag_man = (N3)? larger_exp_man_padded_1_r : 
                           (N4)? smaller_exp_man_shifted_1_r : 1'b0;
  assign N273 = (N2)? 1'b1 : 
                (N277)? 1'b1 : 
                (N272)? 1'b0 : 1'b0;
  assign N274 = (N2)? 1'b0 : 
                (N277)? v_1_r : 1'b0;
  assign N275 = (N2)? 1'b0 : 
                (N277)? v_1_r : 
                (N272)? 1'b0 : 1'b0;
  assign N276 = (N2)? 1'b0 : 
                (N277)? v_1_r : 
                (N272)? 1'b0 : 1'b0;
  assign shifted_adder_output = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N6)? { N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279 } : 1'b0;
  assign N5 = all_zero;
  assign N6 = N278;
  assign N398 = (N2)? 1'b1 : 
                (N402)? 1'b1 : 
                (N397)? 1'b0 : 1'b0;
  assign N399 = (N2)? 1'b0 : 
                (N402)? v_2_r : 1'b0;
  assign N400 = (N2)? 1'b0 : 
                (N402)? v_2_r : 
                (N397)? 1'b0 : 1'b0;
  assign N401 = (N2)? 1'b0 : 
                (N402)? v_2_r : 
                (N397)? 1'b0 : 1'b0;
  assign N422 = (N7)? 1'b0 : 
                (N8)? final_sign_3_r : 1'b0;
  assign N7 = do_sub_3_r;
  assign N8 = N421;
  assign unimplemented_o = (N9)? 1'b0 : 
                           (N424)? 1'b0 : 
                           (N427)? 1'b0 : 
                           (N430)? 1'b0 : 
                           (N433)? 1'b0 : 
                           (N436)? 1'b1 : 
                           (N439)? 1'b0 : 
                           (N442)? 1'b0 : 
                           (N445)? 1'b0 : 
                           (N448)? 1'b0 : 
                           (N420)? 1'b0 : 1'b0;
  assign N9 = N403;
  assign invalid_o = (N9)? 1'b1 : 
                     (N424)? 1'b0 : 
                     (N427)? do_sub_3_r : 
                     (N430)? 1'b0 : 
                     (N433)? 1'b0 : 
                     (N436)? 1'b0 : 
                     (N439)? 1'b0 : 
                     (N442)? 1'b0 : 
                     (N445)? 1'b0 : 
                     (N448)? 1'b0 : 
                     (N420)? 1'b0 : 1'b0;
  assign overflow_o = (N9)? 1'b0 : 
                      (N424)? 1'b0 : 
                      (N427)? 1'b0 : 
                      (N430)? 1'b0 : 
                      (N433)? 1'b0 : 
                      (N436)? 1'b0 : 
                      (N439)? 1'b0 : 
                      (N442)? 1'b0 : 
                      (N445)? 1'b1 : 
                      (N448)? 1'b0 : 
                      (N420)? 1'b0 : 1'b0;
  assign underflow_o = (N9)? 1'b0 : 
                       (N424)? 1'b0 : 
                       (N427)? 1'b0 : 
                       (N430)? 1'b0 : 
                       (N433)? 1'b0 : 
                       (N436)? 1'b0 : 
                       (N439)? 1'b0 : 
                       (N442)? 1'b1 : 
                       (N445)? 1'b0 : 
                       (N448)? 1'b1 : 
                       (N420)? 1'b0 : 1'b0;
  assign z_o = (N9)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
               (N424)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N427)? { N422, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, do_sub_3_r, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N430)? { final_sign_3_r, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N433)? { final_sign_3_r, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N436)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N439)? { final_sign_3_r, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N442)? { final_sign_3_r, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N445)? { final_sign_3_r, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N448)? { final_sign_3_r, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
               (N420)? { final_sign_3_r, rounded } : 1'b0;
  assign stall = v_o & N478;
  assign N478 = ~yumi_i;
  assign ready_o = N479 & en_i;
  assign N479 = ~stall;
  assign N10 = ~exp_a_less;
  assign final_sign = N485 | N488;
  assign N485 = N481 | N484;
  assign N481 = sign_a & N480;
  assign N480 = ~mag_a_less;
  assign N484 = N483 & sub_i;
  assign N483 = N482 & mag_a_less;
  assign N482 = ~sign_b;
  assign N488 = N486 & N487;
  assign N486 = sign_b & mag_a_less;
  assign N487 = ~sub_i;
  assign do_sub = N489 ^ sign_b;
  assign N489 = sub_i ^ sign_a;
  assign N26 = N479 & en_i;
  assign N27 = N26 | reset_i;
  assign N28 = ~N27;
  assign N34 = ~reset_i;
  assign N35 = N26 & N34;
  assign N36 = ~larger_exp_man_less;
  assign N37 = do_sub_1_r ^ smaller_mag_man[115];
  assign N38 = do_sub_1_r ^ smaller_mag_man[114];
  assign N39 = do_sub_1_r ^ smaller_mag_man[113];
  assign N40 = do_sub_1_r ^ smaller_mag_man[112];
  assign N41 = do_sub_1_r ^ smaller_mag_man[111];
  assign N42 = do_sub_1_r ^ smaller_mag_man[110];
  assign N43 = do_sub_1_r ^ smaller_mag_man[109];
  assign N44 = do_sub_1_r ^ smaller_mag_man[108];
  assign N45 = do_sub_1_r ^ smaller_mag_man[107];
  assign N46 = do_sub_1_r ^ smaller_mag_man[106];
  assign N47 = do_sub_1_r ^ smaller_mag_man[105];
  assign N48 = do_sub_1_r ^ smaller_mag_man[104];
  assign N49 = do_sub_1_r ^ smaller_mag_man[103];
  assign N50 = do_sub_1_r ^ smaller_mag_man[102];
  assign N51 = do_sub_1_r ^ smaller_mag_man[101];
  assign N52 = do_sub_1_r ^ smaller_mag_man[100];
  assign N53 = do_sub_1_r ^ smaller_mag_man[99];
  assign N54 = do_sub_1_r ^ smaller_mag_man[98];
  assign N55 = do_sub_1_r ^ smaller_mag_man[97];
  assign N56 = do_sub_1_r ^ smaller_mag_man[96];
  assign N57 = do_sub_1_r ^ smaller_mag_man[95];
  assign N58 = do_sub_1_r ^ smaller_mag_man[94];
  assign N59 = do_sub_1_r ^ smaller_mag_man[93];
  assign N60 = do_sub_1_r ^ smaller_mag_man[92];
  assign N61 = do_sub_1_r ^ smaller_mag_man[91];
  assign N62 = do_sub_1_r ^ smaller_mag_man[90];
  assign N63 = do_sub_1_r ^ smaller_mag_man[89];
  assign N64 = do_sub_1_r ^ smaller_mag_man[88];
  assign N65 = do_sub_1_r ^ smaller_mag_man[87];
  assign N66 = do_sub_1_r ^ smaller_mag_man[86];
  assign N67 = do_sub_1_r ^ smaller_mag_man[85];
  assign N68 = do_sub_1_r ^ smaller_mag_man[84];
  assign N69 = do_sub_1_r ^ smaller_mag_man[83];
  assign N70 = do_sub_1_r ^ smaller_mag_man[82];
  assign N71 = do_sub_1_r ^ smaller_mag_man[81];
  assign N72 = do_sub_1_r ^ smaller_mag_man[80];
  assign N73 = do_sub_1_r ^ smaller_mag_man[79];
  assign N74 = do_sub_1_r ^ smaller_mag_man[78];
  assign N75 = do_sub_1_r ^ smaller_mag_man[77];
  assign N76 = do_sub_1_r ^ smaller_mag_man[76];
  assign N77 = do_sub_1_r ^ smaller_mag_man[75];
  assign N78 = do_sub_1_r ^ smaller_mag_man[74];
  assign N79 = do_sub_1_r ^ smaller_mag_man[73];
  assign N80 = do_sub_1_r ^ smaller_mag_man[72];
  assign N81 = do_sub_1_r ^ smaller_mag_man[71];
  assign N82 = do_sub_1_r ^ smaller_mag_man[70];
  assign N83 = do_sub_1_r ^ smaller_mag_man[69];
  assign N84 = do_sub_1_r ^ smaller_mag_man[68];
  assign N85 = do_sub_1_r ^ smaller_mag_man[67];
  assign N86 = do_sub_1_r ^ smaller_mag_man[66];
  assign N87 = do_sub_1_r ^ smaller_mag_man[65];
  assign N88 = do_sub_1_r ^ smaller_mag_man[64];
  assign N89 = do_sub_1_r ^ smaller_mag_man[63];
  assign N90 = do_sub_1_r ^ smaller_mag_man[62];
  assign N91 = do_sub_1_r ^ smaller_mag_man[61];
  assign N92 = do_sub_1_r ^ smaller_mag_man[60];
  assign N93 = do_sub_1_r ^ smaller_mag_man[59];
  assign N94 = do_sub_1_r ^ smaller_mag_man[58];
  assign N95 = do_sub_1_r ^ smaller_mag_man[57];
  assign N96 = do_sub_1_r ^ smaller_mag_man[56];
  assign N97 = do_sub_1_r ^ smaller_mag_man[55];
  assign N98 = do_sub_1_r ^ smaller_mag_man[54];
  assign N99 = do_sub_1_r ^ smaller_mag_man[53];
  assign N100 = do_sub_1_r ^ smaller_mag_man[52];
  assign N101 = do_sub_1_r ^ smaller_mag_man[51];
  assign N102 = do_sub_1_r ^ smaller_mag_man[50];
  assign N103 = do_sub_1_r ^ smaller_mag_man[49];
  assign N104 = do_sub_1_r ^ smaller_mag_man[48];
  assign N105 = do_sub_1_r ^ smaller_mag_man[47];
  assign N106 = do_sub_1_r ^ smaller_mag_man[46];
  assign N107 = do_sub_1_r ^ smaller_mag_man[45];
  assign N108 = do_sub_1_r ^ smaller_mag_man[44];
  assign N109 = do_sub_1_r ^ smaller_mag_man[43];
  assign N110 = do_sub_1_r ^ smaller_mag_man[42];
  assign N111 = do_sub_1_r ^ smaller_mag_man[41];
  assign N112 = do_sub_1_r ^ smaller_mag_man[40];
  assign N113 = do_sub_1_r ^ smaller_mag_man[39];
  assign N114 = do_sub_1_r ^ smaller_mag_man[38];
  assign N115 = do_sub_1_r ^ smaller_mag_man[37];
  assign N116 = do_sub_1_r ^ smaller_mag_man[36];
  assign N117 = do_sub_1_r ^ smaller_mag_man[35];
  assign N118 = do_sub_1_r ^ smaller_mag_man[34];
  assign N119 = do_sub_1_r ^ smaller_mag_man[33];
  assign N120 = do_sub_1_r ^ smaller_mag_man[32];
  assign N121 = do_sub_1_r ^ smaller_mag_man[31];
  assign N122 = do_sub_1_r ^ smaller_mag_man[30];
  assign N123 = do_sub_1_r ^ smaller_mag_man[29];
  assign N124 = do_sub_1_r ^ smaller_mag_man[28];
  assign N125 = do_sub_1_r ^ smaller_mag_man[27];
  assign N126 = do_sub_1_r ^ smaller_mag_man[26];
  assign N127 = do_sub_1_r ^ smaller_mag_man[25];
  assign N128 = do_sub_1_r ^ smaller_mag_man[24];
  assign N129 = do_sub_1_r ^ smaller_mag_man[23];
  assign N130 = do_sub_1_r ^ smaller_mag_man[22];
  assign N131 = do_sub_1_r ^ smaller_mag_man[21];
  assign N132 = do_sub_1_r ^ smaller_mag_man[20];
  assign N133 = do_sub_1_r ^ smaller_mag_man[19];
  assign N134 = do_sub_1_r ^ smaller_mag_man[18];
  assign N135 = do_sub_1_r ^ smaller_mag_man[17];
  assign N136 = do_sub_1_r ^ smaller_mag_man[16];
  assign N137 = do_sub_1_r ^ smaller_mag_man[15];
  assign N138 = do_sub_1_r ^ smaller_mag_man[14];
  assign N139 = do_sub_1_r ^ smaller_mag_man[13];
  assign N140 = do_sub_1_r ^ smaller_mag_man[12];
  assign N141 = do_sub_1_r ^ smaller_mag_man[11];
  assign N142 = do_sub_1_r ^ smaller_mag_man[10];
  assign N143 = do_sub_1_r ^ smaller_mag_man[9];
  assign N144 = do_sub_1_r ^ smaller_mag_man[8];
  assign N145 = do_sub_1_r ^ smaller_mag_man[7];
  assign N146 = do_sub_1_r ^ smaller_mag_man[6];
  assign N147 = do_sub_1_r ^ smaller_mag_man[5];
  assign N148 = do_sub_1_r ^ smaller_mag_man[4];
  assign N149 = do_sub_1_r ^ smaller_mag_man[3];
  assign N150 = do_sub_1_r ^ smaller_mag_man[2];
  assign N151 = do_sub_1_r ^ smaller_mag_man[1];
  assign N152 = do_sub_1_r ^ smaller_mag_man[0];
  assign N270 = N479 & en_i;
  assign N271 = N270 | reset_i;
  assign N272 = ~N271;
  assign N277 = N270 & N34;
  assign all_zero = ~reduce_o;
  assign N278 = ~all_zero;
  assign round_up = shifted_adder_output[3] & N492;
  assign N492 = N491 | shifted_adder_output[4];
  assign N491 = N490 | shifted_adder_output[0];
  assign N490 = shifted_adder_output[2] | shifted_adder_output[1];
  assign N395 = N479 & en_i;
  assign N396 = N395 | reset_i;
  assign N397 = ~N396;
  assign N402 = N395 & N34;
  assign carry_into_exp = N603 & pre_roundup_3_r[0];
  assign N603 = N602 & pre_roundup_3_r[1];
  assign N602 = N601 & pre_roundup_3_r[2];
  assign N601 = N600 & pre_roundup_3_r[3];
  assign N600 = N599 & pre_roundup_3_r[4];
  assign N599 = N598 & pre_roundup_3_r[5];
  assign N598 = N597 & pre_roundup_3_r[6];
  assign N597 = N596 & pre_roundup_3_r[7];
  assign N596 = N595 & pre_roundup_3_r[8];
  assign N595 = N594 & pre_roundup_3_r[9];
  assign N594 = N593 & pre_roundup_3_r[10];
  assign N593 = N592 & pre_roundup_3_r[11];
  assign N592 = N591 & pre_roundup_3_r[12];
  assign N591 = N590 & pre_roundup_3_r[13];
  assign N590 = N589 & pre_roundup_3_r[14];
  assign N589 = N588 & pre_roundup_3_r[15];
  assign N588 = N587 & pre_roundup_3_r[16];
  assign N587 = N586 & pre_roundup_3_r[17];
  assign N586 = N585 & pre_roundup_3_r[18];
  assign N585 = N584 & pre_roundup_3_r[19];
  assign N584 = N583 & pre_roundup_3_r[20];
  assign N583 = N582 & pre_roundup_3_r[21];
  assign N582 = N581 & pre_roundup_3_r[22];
  assign N581 = N580 & pre_roundup_3_r[23];
  assign N580 = N579 & pre_roundup_3_r[24];
  assign N579 = N578 & pre_roundup_3_r[25];
  assign N578 = N577 & pre_roundup_3_r[26];
  assign N577 = N576 & pre_roundup_3_r[27];
  assign N576 = N575 & pre_roundup_3_r[28];
  assign N575 = N574 & pre_roundup_3_r[29];
  assign N574 = N573 & pre_roundup_3_r[30];
  assign N573 = N572 & pre_roundup_3_r[31];
  assign N572 = N571 & pre_roundup_3_r[32];
  assign N571 = N570 & pre_roundup_3_r[33];
  assign N570 = N569 & pre_roundup_3_r[34];
  assign N569 = N568 & pre_roundup_3_r[35];
  assign N568 = N567 & pre_roundup_3_r[36];
  assign N567 = N566 & pre_roundup_3_r[37];
  assign N566 = N565 & pre_roundup_3_r[38];
  assign N565 = N564 & pre_roundup_3_r[39];
  assign N564 = N563 & pre_roundup_3_r[40];
  assign N563 = N562 & pre_roundup_3_r[41];
  assign N562 = N561 & pre_roundup_3_r[42];
  assign N561 = N560 & pre_roundup_3_r[43];
  assign N560 = N559 & pre_roundup_3_r[44];
  assign N559 = N558 & pre_roundup_3_r[45];
  assign N558 = N557 & pre_roundup_3_r[46];
  assign N557 = N556 & pre_roundup_3_r[47];
  assign N556 = N555 & pre_roundup_3_r[48];
  assign N555 = N554 & pre_roundup_3_r[49];
  assign N554 = N553 & pre_roundup_3_r[50];
  assign N553 = N552 & pre_roundup_3_r[51];
  assign N552 = N551 & pre_roundup_3_r[52];
  assign N551 = N550 & pre_roundup_3_r[53];
  assign N550 = N549 & pre_roundup_3_r[54];
  assign N549 = N548 & pre_roundup_3_r[55];
  assign N548 = N547 & pre_roundup_3_r[56];
  assign N547 = N546 & pre_roundup_3_r[57];
  assign N546 = N545 & pre_roundup_3_r[58];
  assign N545 = N544 & pre_roundup_3_r[59];
  assign N544 = N543 & pre_roundup_3_r[60];
  assign N543 = N542 & pre_roundup_3_r[61];
  assign N542 = N541 & pre_roundup_3_r[62];
  assign N541 = N540 & pre_roundup_3_r[63];
  assign N540 = N539 & pre_roundup_3_r[64];
  assign N539 = N538 & pre_roundup_3_r[65];
  assign N538 = N537 & pre_roundup_3_r[66];
  assign N537 = N536 & pre_roundup_3_r[67];
  assign N536 = N535 & pre_roundup_3_r[68];
  assign N535 = N534 & pre_roundup_3_r[69];
  assign N534 = N533 & pre_roundup_3_r[70];
  assign N533 = N532 & pre_roundup_3_r[71];
  assign N532 = N531 & pre_roundup_3_r[72];
  assign N531 = N530 & pre_roundup_3_r[73];
  assign N530 = N529 & pre_roundup_3_r[74];
  assign N529 = N528 & pre_roundup_3_r[75];
  assign N528 = N527 & pre_roundup_3_r[76];
  assign N527 = N526 & pre_roundup_3_r[77];
  assign N526 = N525 & pre_roundup_3_r[78];
  assign N525 = N524 & pre_roundup_3_r[79];
  assign N524 = N523 & pre_roundup_3_r[80];
  assign N523 = N522 & pre_roundup_3_r[81];
  assign N522 = N521 & pre_roundup_3_r[82];
  assign N521 = N520 & pre_roundup_3_r[83];
  assign N520 = N519 & pre_roundup_3_r[84];
  assign N519 = N518 & pre_roundup_3_r[85];
  assign N518 = N517 & pre_roundup_3_r[86];
  assign N517 = N516 & pre_roundup_3_r[87];
  assign N516 = N515 & pre_roundup_3_r[88];
  assign N515 = N514 & pre_roundup_3_r[89];
  assign N514 = N513 & pre_roundup_3_r[90];
  assign N513 = N512 & pre_roundup_3_r[91];
  assign N512 = N511 & pre_roundup_3_r[92];
  assign N511 = N510 & pre_roundup_3_r[93];
  assign N510 = N509 & pre_roundup_3_r[94];
  assign N509 = N508 & pre_roundup_3_r[95];
  assign N508 = N507 & pre_roundup_3_r[96];
  assign N507 = N506 & pre_roundup_3_r[97];
  assign N506 = N505 & pre_roundup_3_r[98];
  assign N505 = N504 & pre_roundup_3_r[99];
  assign N504 = N503 & pre_roundup_3_r[100];
  assign N503 = N502 & pre_roundup_3_r[101];
  assign N502 = N501 & pre_roundup_3_r[102];
  assign N501 = N500 & pre_roundup_3_r[103];
  assign N500 = N499 & pre_roundup_3_r[104];
  assign N499 = N498 & pre_roundup_3_r[105];
  assign N498 = N497 & pre_roundup_3_r[106];
  assign N497 = N496 & pre_roundup_3_r[107];
  assign N496 = N495 & pre_roundup_3_r[108];
  assign N495 = N494 & pre_roundup_3_r[109];
  assign N494 = N493 & pre_roundup_3_r[110];
  assign N493 = round_up_3_r & pre_roundup_3_r[111];
  assign N403 = a_sig_nan_3_r | b_sig_nan_3_r;
  assign N404 = a_nan_3_r | b_nan_3_r;
  assign N405 = a_infty_3_r & b_infty_3_r;
  assign N406 = a_infty_3_r & N604;
  assign N604 = ~b_infty_3_r;
  assign N407 = N605 & b_infty_3_r;
  assign N605 = ~a_infty_3_r;
  assign N408 = a_denormal_3_r | b_denormal_3_r;
  assign N409 = N477 & N606;
  assign N606 = pre_roundup_3_r[112] | carry_into_exp;
  assign N410 = N463 & N607;
  assign N607 = ~carry_into_exp;
  assign N411 = N404 | N403;
  assign N412 = N405 | N411;
  assign N413 = N406 | N412;
  assign N414 = N407 | N413;
  assign N415 = N408 | N414;
  assign N416 = all_zero_3_r | N415;
  assign N417 = adjusted_exp_cout_3_r | N416;
  assign N418 = N409 | N417;
  assign N419 = N410 | N418;
  assign N420 = ~N419;
  assign N421 = ~do_sub_3_r;
  assign N423 = ~N403;
  assign N424 = N404 & N423;
  assign N425 = ~N404;
  assign N426 = N423 & N425;
  assign N427 = N405 & N426;
  assign N428 = ~N405;
  assign N429 = N426 & N428;
  assign N430 = N406 & N429;
  assign N431 = ~N406;
  assign N432 = N429 & N431;
  assign N433 = N407 & N432;
  assign N434 = ~N407;
  assign N435 = N432 & N434;
  assign N436 = N408 & N435;
  assign N437 = ~N408;
  assign N438 = N435 & N437;
  assign N439 = all_zero_3_r & N438;
  assign N440 = ~all_zero_3_r;
  assign N441 = N438 & N440;
  assign N442 = adjusted_exp_cout_3_r & N441;
  assign N443 = ~adjusted_exp_cout_3_r;
  assign N444 = N441 & N443;
  assign N445 = N409 & N444;
  assign N446 = ~N409;
  assign N447 = N444 & N446;
  assign N448 = N410 & N447;

  always @(posedge clk_i) begin
    if(N31) begin
      a_denormal_1_r <= a_denormal;
      b_denormal_1_r <= b_denormal;
      final_sign_1_r <= final_sign;
      { larger_exp_man_padded_1_r[115:25] } <= { 1'b1, larger_exp_man[111:22] };
      a_sig_nan_1_r <= a_sig_nan;
      b_sig_nan_1_r <= b_sig_nan;
      a_nan_1_r <= a_nan;
      b_nan_1_r <= b_nan;
      a_infty_1_r <= a_infty;
      b_infty_1_r <= b_infty;
    end 
    if(N29) begin
      v_1_r <= N30;
    end 
    if(N32) begin
      do_sub_1_r <= do_sub;
      { smaller_exp_man_shifted_1_r[115:42] } <= { smaller_exp_man_shifted[115:42] };
      { larger_exp_man_padded_1_r[24:0] } <= { larger_exp_man[21:0], 1'b0, 1'b0, 1'b0 };
    end 
    if(N33) begin
      { larger_exp_1_r[14:0] } <= { larger_exp[14:0] };
      { smaller_exp_man_shifted_1_r[41:0] } <= { smaller_exp_man_shifted[41:0] };
    end 
    if(N275) begin
      a_denormal_2_r <= a_denormal_1_r;
      b_denormal_2_r <= b_denormal_1_r;
      { larger_exp_2_r[0:0] } <= { larger_exp_1_r[0:0] };
      { adder_output_2_r[116:28] } <= { adder_output[116:28] };
      final_sign_2_r <= final_sign_1_r;
      do_sub_2_r <= do_sub_1_r;
      a_sig_nan_2_r <= a_sig_nan_1_r;
      b_sig_nan_2_r <= b_sig_nan_1_r;
      a_nan_2_r <= a_nan_1_r;
      b_nan_2_r <= b_nan_1_r;
      a_infty_2_r <= a_infty_1_r;
      b_infty_2_r <= b_infty_1_r;
    end 
    if(N273) begin
      v_2_r <= N274;
    end 
    if(N276) begin
      { larger_exp_2_r[14:1] } <= { larger_exp_1_r[14:1] };
      { adder_output_2_r[27:0] } <= { adder_output[27:0] };
    end 
    if(N400) begin
      adjusted_exp_cout_3_r <= adjusted_exp_cout;
      final_sign_3_r <= final_sign_2_r;
      { pre_roundup_3_r[126:41], pre_roundup_3_r[0:0] } <= { adjusted_exp[14:0], shifted_adder_output[115:45], shifted_adder_output[4:4] };
      round_up_3_r <= round_up;
      all_zero_3_r <= all_zero;
      a_sig_nan_3_r <= a_sig_nan_2_r;
      b_sig_nan_3_r <= b_sig_nan_2_r;
      a_nan_3_r <= a_nan_2_r;
      b_nan_3_r <= b_nan_2_r;
      a_infty_3_r <= a_infty_2_r;
      b_infty_3_r <= b_infty_2_r;
      do_sub_3_r <= do_sub_2_r;
      a_denormal_3_r <= a_denormal_2_r;
      b_denormal_3_r <= b_denormal_2_r;
    end 
    if(N398) begin
      v_o <= N399;
    end 
    if(N401) begin
      { pre_roundup_3_r[40:1] } <= { shifted_adder_output[44:5] };
    end 
  end


endmodule

