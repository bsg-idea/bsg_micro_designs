

module top
(
  clk_i,
  reset_i,
  ready_o,
  v_i,
  data_i,
  v_o,
  data_o,
  ready_i
);

  input [31:0] data_i;
  output [49:0] v_o;
  output [1599:0] data_o;
  input [49:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output ready_o;

  bsg_front_side_bus_hop_in
  wrapper
  (
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .ready_i(ready_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [63:0] mem;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[62] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[61] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[60] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[59] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[58] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[57] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[56] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[55] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[45] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[44] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[43] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[42] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[41] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[40] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[39] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[38] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[37] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[36] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[35] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[34] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[33] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[63:32] } <= { w_data_i[31:0] };
    end 
    if(N7) begin
      { mem[31:0] } <= { w_data_i[31:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bsg_front_side_bus_hop_in
(
  clk_i,
  reset_i,
  ready_o,
  v_i,
  data_i,
  v_o,
  data_o,
  ready_i
);

  input [31:0] data_i;
  output [49:0] v_o;
  output [1599:0] data_o;
  input [49:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output ready_o;
  wire [49:0] v_o,sent_n;
  wire [1599:0] data_o;
  wire ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,fifo_v,fifo_yumi,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597;
  reg [49:0] sent_r;
  assign data_o[63] = data_o[31];
  assign data_o[95] = data_o[31];
  assign data_o[127] = data_o[31];
  assign data_o[159] = data_o[31];
  assign data_o[191] = data_o[31];
  assign data_o[223] = data_o[31];
  assign data_o[255] = data_o[31];
  assign data_o[287] = data_o[31];
  assign data_o[319] = data_o[31];
  assign data_o[351] = data_o[31];
  assign data_o[383] = data_o[31];
  assign data_o[415] = data_o[31];
  assign data_o[447] = data_o[31];
  assign data_o[479] = data_o[31];
  assign data_o[511] = data_o[31];
  assign data_o[543] = data_o[31];
  assign data_o[575] = data_o[31];
  assign data_o[607] = data_o[31];
  assign data_o[639] = data_o[31];
  assign data_o[671] = data_o[31];
  assign data_o[703] = data_o[31];
  assign data_o[735] = data_o[31];
  assign data_o[767] = data_o[31];
  assign data_o[799] = data_o[31];
  assign data_o[831] = data_o[31];
  assign data_o[863] = data_o[31];
  assign data_o[895] = data_o[31];
  assign data_o[927] = data_o[31];
  assign data_o[959] = data_o[31];
  assign data_o[991] = data_o[31];
  assign data_o[1023] = data_o[31];
  assign data_o[1055] = data_o[31];
  assign data_o[1087] = data_o[31];
  assign data_o[1119] = data_o[31];
  assign data_o[1151] = data_o[31];
  assign data_o[1183] = data_o[31];
  assign data_o[1215] = data_o[31];
  assign data_o[1247] = data_o[31];
  assign data_o[1279] = data_o[31];
  assign data_o[1311] = data_o[31];
  assign data_o[1343] = data_o[31];
  assign data_o[1375] = data_o[31];
  assign data_o[1407] = data_o[31];
  assign data_o[1439] = data_o[31];
  assign data_o[1471] = data_o[31];
  assign data_o[1503] = data_o[31];
  assign data_o[1535] = data_o[31];
  assign data_o[1567] = data_o[31];
  assign data_o[1599] = data_o[31];
  assign data_o[62] = data_o[30];
  assign data_o[94] = data_o[30];
  assign data_o[126] = data_o[30];
  assign data_o[158] = data_o[30];
  assign data_o[190] = data_o[30];
  assign data_o[222] = data_o[30];
  assign data_o[254] = data_o[30];
  assign data_o[286] = data_o[30];
  assign data_o[318] = data_o[30];
  assign data_o[350] = data_o[30];
  assign data_o[382] = data_o[30];
  assign data_o[414] = data_o[30];
  assign data_o[446] = data_o[30];
  assign data_o[478] = data_o[30];
  assign data_o[510] = data_o[30];
  assign data_o[542] = data_o[30];
  assign data_o[574] = data_o[30];
  assign data_o[606] = data_o[30];
  assign data_o[638] = data_o[30];
  assign data_o[670] = data_o[30];
  assign data_o[702] = data_o[30];
  assign data_o[734] = data_o[30];
  assign data_o[766] = data_o[30];
  assign data_o[798] = data_o[30];
  assign data_o[830] = data_o[30];
  assign data_o[862] = data_o[30];
  assign data_o[894] = data_o[30];
  assign data_o[926] = data_o[30];
  assign data_o[958] = data_o[30];
  assign data_o[990] = data_o[30];
  assign data_o[1022] = data_o[30];
  assign data_o[1054] = data_o[30];
  assign data_o[1086] = data_o[30];
  assign data_o[1118] = data_o[30];
  assign data_o[1150] = data_o[30];
  assign data_o[1182] = data_o[30];
  assign data_o[1214] = data_o[30];
  assign data_o[1246] = data_o[30];
  assign data_o[1278] = data_o[30];
  assign data_o[1310] = data_o[30];
  assign data_o[1342] = data_o[30];
  assign data_o[1374] = data_o[30];
  assign data_o[1406] = data_o[30];
  assign data_o[1438] = data_o[30];
  assign data_o[1470] = data_o[30];
  assign data_o[1502] = data_o[30];
  assign data_o[1534] = data_o[30];
  assign data_o[1566] = data_o[30];
  assign data_o[1598] = data_o[30];
  assign data_o[61] = data_o[29];
  assign data_o[93] = data_o[29];
  assign data_o[125] = data_o[29];
  assign data_o[157] = data_o[29];
  assign data_o[189] = data_o[29];
  assign data_o[221] = data_o[29];
  assign data_o[253] = data_o[29];
  assign data_o[285] = data_o[29];
  assign data_o[317] = data_o[29];
  assign data_o[349] = data_o[29];
  assign data_o[381] = data_o[29];
  assign data_o[413] = data_o[29];
  assign data_o[445] = data_o[29];
  assign data_o[477] = data_o[29];
  assign data_o[509] = data_o[29];
  assign data_o[541] = data_o[29];
  assign data_o[573] = data_o[29];
  assign data_o[605] = data_o[29];
  assign data_o[637] = data_o[29];
  assign data_o[669] = data_o[29];
  assign data_o[701] = data_o[29];
  assign data_o[733] = data_o[29];
  assign data_o[765] = data_o[29];
  assign data_o[797] = data_o[29];
  assign data_o[829] = data_o[29];
  assign data_o[861] = data_o[29];
  assign data_o[893] = data_o[29];
  assign data_o[925] = data_o[29];
  assign data_o[957] = data_o[29];
  assign data_o[989] = data_o[29];
  assign data_o[1021] = data_o[29];
  assign data_o[1053] = data_o[29];
  assign data_o[1085] = data_o[29];
  assign data_o[1117] = data_o[29];
  assign data_o[1149] = data_o[29];
  assign data_o[1181] = data_o[29];
  assign data_o[1213] = data_o[29];
  assign data_o[1245] = data_o[29];
  assign data_o[1277] = data_o[29];
  assign data_o[1309] = data_o[29];
  assign data_o[1341] = data_o[29];
  assign data_o[1373] = data_o[29];
  assign data_o[1405] = data_o[29];
  assign data_o[1437] = data_o[29];
  assign data_o[1469] = data_o[29];
  assign data_o[1501] = data_o[29];
  assign data_o[1533] = data_o[29];
  assign data_o[1565] = data_o[29];
  assign data_o[1597] = data_o[29];
  assign data_o[60] = data_o[28];
  assign data_o[92] = data_o[28];
  assign data_o[124] = data_o[28];
  assign data_o[156] = data_o[28];
  assign data_o[188] = data_o[28];
  assign data_o[220] = data_o[28];
  assign data_o[252] = data_o[28];
  assign data_o[284] = data_o[28];
  assign data_o[316] = data_o[28];
  assign data_o[348] = data_o[28];
  assign data_o[380] = data_o[28];
  assign data_o[412] = data_o[28];
  assign data_o[444] = data_o[28];
  assign data_o[476] = data_o[28];
  assign data_o[508] = data_o[28];
  assign data_o[540] = data_o[28];
  assign data_o[572] = data_o[28];
  assign data_o[604] = data_o[28];
  assign data_o[636] = data_o[28];
  assign data_o[668] = data_o[28];
  assign data_o[700] = data_o[28];
  assign data_o[732] = data_o[28];
  assign data_o[764] = data_o[28];
  assign data_o[796] = data_o[28];
  assign data_o[828] = data_o[28];
  assign data_o[860] = data_o[28];
  assign data_o[892] = data_o[28];
  assign data_o[924] = data_o[28];
  assign data_o[956] = data_o[28];
  assign data_o[988] = data_o[28];
  assign data_o[1020] = data_o[28];
  assign data_o[1052] = data_o[28];
  assign data_o[1084] = data_o[28];
  assign data_o[1116] = data_o[28];
  assign data_o[1148] = data_o[28];
  assign data_o[1180] = data_o[28];
  assign data_o[1212] = data_o[28];
  assign data_o[1244] = data_o[28];
  assign data_o[1276] = data_o[28];
  assign data_o[1308] = data_o[28];
  assign data_o[1340] = data_o[28];
  assign data_o[1372] = data_o[28];
  assign data_o[1404] = data_o[28];
  assign data_o[1436] = data_o[28];
  assign data_o[1468] = data_o[28];
  assign data_o[1500] = data_o[28];
  assign data_o[1532] = data_o[28];
  assign data_o[1564] = data_o[28];
  assign data_o[1596] = data_o[28];
  assign data_o[59] = data_o[27];
  assign data_o[91] = data_o[27];
  assign data_o[123] = data_o[27];
  assign data_o[155] = data_o[27];
  assign data_o[187] = data_o[27];
  assign data_o[219] = data_o[27];
  assign data_o[251] = data_o[27];
  assign data_o[283] = data_o[27];
  assign data_o[315] = data_o[27];
  assign data_o[347] = data_o[27];
  assign data_o[379] = data_o[27];
  assign data_o[411] = data_o[27];
  assign data_o[443] = data_o[27];
  assign data_o[475] = data_o[27];
  assign data_o[507] = data_o[27];
  assign data_o[539] = data_o[27];
  assign data_o[571] = data_o[27];
  assign data_o[603] = data_o[27];
  assign data_o[635] = data_o[27];
  assign data_o[667] = data_o[27];
  assign data_o[699] = data_o[27];
  assign data_o[731] = data_o[27];
  assign data_o[763] = data_o[27];
  assign data_o[795] = data_o[27];
  assign data_o[827] = data_o[27];
  assign data_o[859] = data_o[27];
  assign data_o[891] = data_o[27];
  assign data_o[923] = data_o[27];
  assign data_o[955] = data_o[27];
  assign data_o[987] = data_o[27];
  assign data_o[1019] = data_o[27];
  assign data_o[1051] = data_o[27];
  assign data_o[1083] = data_o[27];
  assign data_o[1115] = data_o[27];
  assign data_o[1147] = data_o[27];
  assign data_o[1179] = data_o[27];
  assign data_o[1211] = data_o[27];
  assign data_o[1243] = data_o[27];
  assign data_o[1275] = data_o[27];
  assign data_o[1307] = data_o[27];
  assign data_o[1339] = data_o[27];
  assign data_o[1371] = data_o[27];
  assign data_o[1403] = data_o[27];
  assign data_o[1435] = data_o[27];
  assign data_o[1467] = data_o[27];
  assign data_o[1499] = data_o[27];
  assign data_o[1531] = data_o[27];
  assign data_o[1563] = data_o[27];
  assign data_o[1595] = data_o[27];
  assign data_o[58] = data_o[26];
  assign data_o[90] = data_o[26];
  assign data_o[122] = data_o[26];
  assign data_o[154] = data_o[26];
  assign data_o[186] = data_o[26];
  assign data_o[218] = data_o[26];
  assign data_o[250] = data_o[26];
  assign data_o[282] = data_o[26];
  assign data_o[314] = data_o[26];
  assign data_o[346] = data_o[26];
  assign data_o[378] = data_o[26];
  assign data_o[410] = data_o[26];
  assign data_o[442] = data_o[26];
  assign data_o[474] = data_o[26];
  assign data_o[506] = data_o[26];
  assign data_o[538] = data_o[26];
  assign data_o[570] = data_o[26];
  assign data_o[602] = data_o[26];
  assign data_o[634] = data_o[26];
  assign data_o[666] = data_o[26];
  assign data_o[698] = data_o[26];
  assign data_o[730] = data_o[26];
  assign data_o[762] = data_o[26];
  assign data_o[794] = data_o[26];
  assign data_o[826] = data_o[26];
  assign data_o[858] = data_o[26];
  assign data_o[890] = data_o[26];
  assign data_o[922] = data_o[26];
  assign data_o[954] = data_o[26];
  assign data_o[986] = data_o[26];
  assign data_o[1018] = data_o[26];
  assign data_o[1050] = data_o[26];
  assign data_o[1082] = data_o[26];
  assign data_o[1114] = data_o[26];
  assign data_o[1146] = data_o[26];
  assign data_o[1178] = data_o[26];
  assign data_o[1210] = data_o[26];
  assign data_o[1242] = data_o[26];
  assign data_o[1274] = data_o[26];
  assign data_o[1306] = data_o[26];
  assign data_o[1338] = data_o[26];
  assign data_o[1370] = data_o[26];
  assign data_o[1402] = data_o[26];
  assign data_o[1434] = data_o[26];
  assign data_o[1466] = data_o[26];
  assign data_o[1498] = data_o[26];
  assign data_o[1530] = data_o[26];
  assign data_o[1562] = data_o[26];
  assign data_o[1594] = data_o[26];
  assign data_o[57] = data_o[25];
  assign data_o[89] = data_o[25];
  assign data_o[121] = data_o[25];
  assign data_o[153] = data_o[25];
  assign data_o[185] = data_o[25];
  assign data_o[217] = data_o[25];
  assign data_o[249] = data_o[25];
  assign data_o[281] = data_o[25];
  assign data_o[313] = data_o[25];
  assign data_o[345] = data_o[25];
  assign data_o[377] = data_o[25];
  assign data_o[409] = data_o[25];
  assign data_o[441] = data_o[25];
  assign data_o[473] = data_o[25];
  assign data_o[505] = data_o[25];
  assign data_o[537] = data_o[25];
  assign data_o[569] = data_o[25];
  assign data_o[601] = data_o[25];
  assign data_o[633] = data_o[25];
  assign data_o[665] = data_o[25];
  assign data_o[697] = data_o[25];
  assign data_o[729] = data_o[25];
  assign data_o[761] = data_o[25];
  assign data_o[793] = data_o[25];
  assign data_o[825] = data_o[25];
  assign data_o[857] = data_o[25];
  assign data_o[889] = data_o[25];
  assign data_o[921] = data_o[25];
  assign data_o[953] = data_o[25];
  assign data_o[985] = data_o[25];
  assign data_o[1017] = data_o[25];
  assign data_o[1049] = data_o[25];
  assign data_o[1081] = data_o[25];
  assign data_o[1113] = data_o[25];
  assign data_o[1145] = data_o[25];
  assign data_o[1177] = data_o[25];
  assign data_o[1209] = data_o[25];
  assign data_o[1241] = data_o[25];
  assign data_o[1273] = data_o[25];
  assign data_o[1305] = data_o[25];
  assign data_o[1337] = data_o[25];
  assign data_o[1369] = data_o[25];
  assign data_o[1401] = data_o[25];
  assign data_o[1433] = data_o[25];
  assign data_o[1465] = data_o[25];
  assign data_o[1497] = data_o[25];
  assign data_o[1529] = data_o[25];
  assign data_o[1561] = data_o[25];
  assign data_o[1593] = data_o[25];
  assign data_o[56] = data_o[24];
  assign data_o[88] = data_o[24];
  assign data_o[120] = data_o[24];
  assign data_o[152] = data_o[24];
  assign data_o[184] = data_o[24];
  assign data_o[216] = data_o[24];
  assign data_o[248] = data_o[24];
  assign data_o[280] = data_o[24];
  assign data_o[312] = data_o[24];
  assign data_o[344] = data_o[24];
  assign data_o[376] = data_o[24];
  assign data_o[408] = data_o[24];
  assign data_o[440] = data_o[24];
  assign data_o[472] = data_o[24];
  assign data_o[504] = data_o[24];
  assign data_o[536] = data_o[24];
  assign data_o[568] = data_o[24];
  assign data_o[600] = data_o[24];
  assign data_o[632] = data_o[24];
  assign data_o[664] = data_o[24];
  assign data_o[696] = data_o[24];
  assign data_o[728] = data_o[24];
  assign data_o[760] = data_o[24];
  assign data_o[792] = data_o[24];
  assign data_o[824] = data_o[24];
  assign data_o[856] = data_o[24];
  assign data_o[888] = data_o[24];
  assign data_o[920] = data_o[24];
  assign data_o[952] = data_o[24];
  assign data_o[984] = data_o[24];
  assign data_o[1016] = data_o[24];
  assign data_o[1048] = data_o[24];
  assign data_o[1080] = data_o[24];
  assign data_o[1112] = data_o[24];
  assign data_o[1144] = data_o[24];
  assign data_o[1176] = data_o[24];
  assign data_o[1208] = data_o[24];
  assign data_o[1240] = data_o[24];
  assign data_o[1272] = data_o[24];
  assign data_o[1304] = data_o[24];
  assign data_o[1336] = data_o[24];
  assign data_o[1368] = data_o[24];
  assign data_o[1400] = data_o[24];
  assign data_o[1432] = data_o[24];
  assign data_o[1464] = data_o[24];
  assign data_o[1496] = data_o[24];
  assign data_o[1528] = data_o[24];
  assign data_o[1560] = data_o[24];
  assign data_o[1592] = data_o[24];
  assign data_o[55] = data_o[23];
  assign data_o[87] = data_o[23];
  assign data_o[119] = data_o[23];
  assign data_o[151] = data_o[23];
  assign data_o[183] = data_o[23];
  assign data_o[215] = data_o[23];
  assign data_o[247] = data_o[23];
  assign data_o[279] = data_o[23];
  assign data_o[311] = data_o[23];
  assign data_o[343] = data_o[23];
  assign data_o[375] = data_o[23];
  assign data_o[407] = data_o[23];
  assign data_o[439] = data_o[23];
  assign data_o[471] = data_o[23];
  assign data_o[503] = data_o[23];
  assign data_o[535] = data_o[23];
  assign data_o[567] = data_o[23];
  assign data_o[599] = data_o[23];
  assign data_o[631] = data_o[23];
  assign data_o[663] = data_o[23];
  assign data_o[695] = data_o[23];
  assign data_o[727] = data_o[23];
  assign data_o[759] = data_o[23];
  assign data_o[791] = data_o[23];
  assign data_o[823] = data_o[23];
  assign data_o[855] = data_o[23];
  assign data_o[887] = data_o[23];
  assign data_o[919] = data_o[23];
  assign data_o[951] = data_o[23];
  assign data_o[983] = data_o[23];
  assign data_o[1015] = data_o[23];
  assign data_o[1047] = data_o[23];
  assign data_o[1079] = data_o[23];
  assign data_o[1111] = data_o[23];
  assign data_o[1143] = data_o[23];
  assign data_o[1175] = data_o[23];
  assign data_o[1207] = data_o[23];
  assign data_o[1239] = data_o[23];
  assign data_o[1271] = data_o[23];
  assign data_o[1303] = data_o[23];
  assign data_o[1335] = data_o[23];
  assign data_o[1367] = data_o[23];
  assign data_o[1399] = data_o[23];
  assign data_o[1431] = data_o[23];
  assign data_o[1463] = data_o[23];
  assign data_o[1495] = data_o[23];
  assign data_o[1527] = data_o[23];
  assign data_o[1559] = data_o[23];
  assign data_o[1591] = data_o[23];
  assign data_o[54] = data_o[22];
  assign data_o[86] = data_o[22];
  assign data_o[118] = data_o[22];
  assign data_o[150] = data_o[22];
  assign data_o[182] = data_o[22];
  assign data_o[214] = data_o[22];
  assign data_o[246] = data_o[22];
  assign data_o[278] = data_o[22];
  assign data_o[310] = data_o[22];
  assign data_o[342] = data_o[22];
  assign data_o[374] = data_o[22];
  assign data_o[406] = data_o[22];
  assign data_o[438] = data_o[22];
  assign data_o[470] = data_o[22];
  assign data_o[502] = data_o[22];
  assign data_o[534] = data_o[22];
  assign data_o[566] = data_o[22];
  assign data_o[598] = data_o[22];
  assign data_o[630] = data_o[22];
  assign data_o[662] = data_o[22];
  assign data_o[694] = data_o[22];
  assign data_o[726] = data_o[22];
  assign data_o[758] = data_o[22];
  assign data_o[790] = data_o[22];
  assign data_o[822] = data_o[22];
  assign data_o[854] = data_o[22];
  assign data_o[886] = data_o[22];
  assign data_o[918] = data_o[22];
  assign data_o[950] = data_o[22];
  assign data_o[982] = data_o[22];
  assign data_o[1014] = data_o[22];
  assign data_o[1046] = data_o[22];
  assign data_o[1078] = data_o[22];
  assign data_o[1110] = data_o[22];
  assign data_o[1142] = data_o[22];
  assign data_o[1174] = data_o[22];
  assign data_o[1206] = data_o[22];
  assign data_o[1238] = data_o[22];
  assign data_o[1270] = data_o[22];
  assign data_o[1302] = data_o[22];
  assign data_o[1334] = data_o[22];
  assign data_o[1366] = data_o[22];
  assign data_o[1398] = data_o[22];
  assign data_o[1430] = data_o[22];
  assign data_o[1462] = data_o[22];
  assign data_o[1494] = data_o[22];
  assign data_o[1526] = data_o[22];
  assign data_o[1558] = data_o[22];
  assign data_o[1590] = data_o[22];
  assign data_o[53] = data_o[21];
  assign data_o[85] = data_o[21];
  assign data_o[117] = data_o[21];
  assign data_o[149] = data_o[21];
  assign data_o[181] = data_o[21];
  assign data_o[213] = data_o[21];
  assign data_o[245] = data_o[21];
  assign data_o[277] = data_o[21];
  assign data_o[309] = data_o[21];
  assign data_o[341] = data_o[21];
  assign data_o[373] = data_o[21];
  assign data_o[405] = data_o[21];
  assign data_o[437] = data_o[21];
  assign data_o[469] = data_o[21];
  assign data_o[501] = data_o[21];
  assign data_o[533] = data_o[21];
  assign data_o[565] = data_o[21];
  assign data_o[597] = data_o[21];
  assign data_o[629] = data_o[21];
  assign data_o[661] = data_o[21];
  assign data_o[693] = data_o[21];
  assign data_o[725] = data_o[21];
  assign data_o[757] = data_o[21];
  assign data_o[789] = data_o[21];
  assign data_o[821] = data_o[21];
  assign data_o[853] = data_o[21];
  assign data_o[885] = data_o[21];
  assign data_o[917] = data_o[21];
  assign data_o[949] = data_o[21];
  assign data_o[981] = data_o[21];
  assign data_o[1013] = data_o[21];
  assign data_o[1045] = data_o[21];
  assign data_o[1077] = data_o[21];
  assign data_o[1109] = data_o[21];
  assign data_o[1141] = data_o[21];
  assign data_o[1173] = data_o[21];
  assign data_o[1205] = data_o[21];
  assign data_o[1237] = data_o[21];
  assign data_o[1269] = data_o[21];
  assign data_o[1301] = data_o[21];
  assign data_o[1333] = data_o[21];
  assign data_o[1365] = data_o[21];
  assign data_o[1397] = data_o[21];
  assign data_o[1429] = data_o[21];
  assign data_o[1461] = data_o[21];
  assign data_o[1493] = data_o[21];
  assign data_o[1525] = data_o[21];
  assign data_o[1557] = data_o[21];
  assign data_o[1589] = data_o[21];
  assign data_o[52] = data_o[20];
  assign data_o[84] = data_o[20];
  assign data_o[116] = data_o[20];
  assign data_o[148] = data_o[20];
  assign data_o[180] = data_o[20];
  assign data_o[212] = data_o[20];
  assign data_o[244] = data_o[20];
  assign data_o[276] = data_o[20];
  assign data_o[308] = data_o[20];
  assign data_o[340] = data_o[20];
  assign data_o[372] = data_o[20];
  assign data_o[404] = data_o[20];
  assign data_o[436] = data_o[20];
  assign data_o[468] = data_o[20];
  assign data_o[500] = data_o[20];
  assign data_o[532] = data_o[20];
  assign data_o[564] = data_o[20];
  assign data_o[596] = data_o[20];
  assign data_o[628] = data_o[20];
  assign data_o[660] = data_o[20];
  assign data_o[692] = data_o[20];
  assign data_o[724] = data_o[20];
  assign data_o[756] = data_o[20];
  assign data_o[788] = data_o[20];
  assign data_o[820] = data_o[20];
  assign data_o[852] = data_o[20];
  assign data_o[884] = data_o[20];
  assign data_o[916] = data_o[20];
  assign data_o[948] = data_o[20];
  assign data_o[980] = data_o[20];
  assign data_o[1012] = data_o[20];
  assign data_o[1044] = data_o[20];
  assign data_o[1076] = data_o[20];
  assign data_o[1108] = data_o[20];
  assign data_o[1140] = data_o[20];
  assign data_o[1172] = data_o[20];
  assign data_o[1204] = data_o[20];
  assign data_o[1236] = data_o[20];
  assign data_o[1268] = data_o[20];
  assign data_o[1300] = data_o[20];
  assign data_o[1332] = data_o[20];
  assign data_o[1364] = data_o[20];
  assign data_o[1396] = data_o[20];
  assign data_o[1428] = data_o[20];
  assign data_o[1460] = data_o[20];
  assign data_o[1492] = data_o[20];
  assign data_o[1524] = data_o[20];
  assign data_o[1556] = data_o[20];
  assign data_o[1588] = data_o[20];
  assign data_o[51] = data_o[19];
  assign data_o[83] = data_o[19];
  assign data_o[115] = data_o[19];
  assign data_o[147] = data_o[19];
  assign data_o[179] = data_o[19];
  assign data_o[211] = data_o[19];
  assign data_o[243] = data_o[19];
  assign data_o[275] = data_o[19];
  assign data_o[307] = data_o[19];
  assign data_o[339] = data_o[19];
  assign data_o[371] = data_o[19];
  assign data_o[403] = data_o[19];
  assign data_o[435] = data_o[19];
  assign data_o[467] = data_o[19];
  assign data_o[499] = data_o[19];
  assign data_o[531] = data_o[19];
  assign data_o[563] = data_o[19];
  assign data_o[595] = data_o[19];
  assign data_o[627] = data_o[19];
  assign data_o[659] = data_o[19];
  assign data_o[691] = data_o[19];
  assign data_o[723] = data_o[19];
  assign data_o[755] = data_o[19];
  assign data_o[787] = data_o[19];
  assign data_o[819] = data_o[19];
  assign data_o[851] = data_o[19];
  assign data_o[883] = data_o[19];
  assign data_o[915] = data_o[19];
  assign data_o[947] = data_o[19];
  assign data_o[979] = data_o[19];
  assign data_o[1011] = data_o[19];
  assign data_o[1043] = data_o[19];
  assign data_o[1075] = data_o[19];
  assign data_o[1107] = data_o[19];
  assign data_o[1139] = data_o[19];
  assign data_o[1171] = data_o[19];
  assign data_o[1203] = data_o[19];
  assign data_o[1235] = data_o[19];
  assign data_o[1267] = data_o[19];
  assign data_o[1299] = data_o[19];
  assign data_o[1331] = data_o[19];
  assign data_o[1363] = data_o[19];
  assign data_o[1395] = data_o[19];
  assign data_o[1427] = data_o[19];
  assign data_o[1459] = data_o[19];
  assign data_o[1491] = data_o[19];
  assign data_o[1523] = data_o[19];
  assign data_o[1555] = data_o[19];
  assign data_o[1587] = data_o[19];
  assign data_o[50] = data_o[18];
  assign data_o[82] = data_o[18];
  assign data_o[114] = data_o[18];
  assign data_o[146] = data_o[18];
  assign data_o[178] = data_o[18];
  assign data_o[210] = data_o[18];
  assign data_o[242] = data_o[18];
  assign data_o[274] = data_o[18];
  assign data_o[306] = data_o[18];
  assign data_o[338] = data_o[18];
  assign data_o[370] = data_o[18];
  assign data_o[402] = data_o[18];
  assign data_o[434] = data_o[18];
  assign data_o[466] = data_o[18];
  assign data_o[498] = data_o[18];
  assign data_o[530] = data_o[18];
  assign data_o[562] = data_o[18];
  assign data_o[594] = data_o[18];
  assign data_o[626] = data_o[18];
  assign data_o[658] = data_o[18];
  assign data_o[690] = data_o[18];
  assign data_o[722] = data_o[18];
  assign data_o[754] = data_o[18];
  assign data_o[786] = data_o[18];
  assign data_o[818] = data_o[18];
  assign data_o[850] = data_o[18];
  assign data_o[882] = data_o[18];
  assign data_o[914] = data_o[18];
  assign data_o[946] = data_o[18];
  assign data_o[978] = data_o[18];
  assign data_o[1010] = data_o[18];
  assign data_o[1042] = data_o[18];
  assign data_o[1074] = data_o[18];
  assign data_o[1106] = data_o[18];
  assign data_o[1138] = data_o[18];
  assign data_o[1170] = data_o[18];
  assign data_o[1202] = data_o[18];
  assign data_o[1234] = data_o[18];
  assign data_o[1266] = data_o[18];
  assign data_o[1298] = data_o[18];
  assign data_o[1330] = data_o[18];
  assign data_o[1362] = data_o[18];
  assign data_o[1394] = data_o[18];
  assign data_o[1426] = data_o[18];
  assign data_o[1458] = data_o[18];
  assign data_o[1490] = data_o[18];
  assign data_o[1522] = data_o[18];
  assign data_o[1554] = data_o[18];
  assign data_o[1586] = data_o[18];
  assign data_o[49] = data_o[17];
  assign data_o[81] = data_o[17];
  assign data_o[113] = data_o[17];
  assign data_o[145] = data_o[17];
  assign data_o[177] = data_o[17];
  assign data_o[209] = data_o[17];
  assign data_o[241] = data_o[17];
  assign data_o[273] = data_o[17];
  assign data_o[305] = data_o[17];
  assign data_o[337] = data_o[17];
  assign data_o[369] = data_o[17];
  assign data_o[401] = data_o[17];
  assign data_o[433] = data_o[17];
  assign data_o[465] = data_o[17];
  assign data_o[497] = data_o[17];
  assign data_o[529] = data_o[17];
  assign data_o[561] = data_o[17];
  assign data_o[593] = data_o[17];
  assign data_o[625] = data_o[17];
  assign data_o[657] = data_o[17];
  assign data_o[689] = data_o[17];
  assign data_o[721] = data_o[17];
  assign data_o[753] = data_o[17];
  assign data_o[785] = data_o[17];
  assign data_o[817] = data_o[17];
  assign data_o[849] = data_o[17];
  assign data_o[881] = data_o[17];
  assign data_o[913] = data_o[17];
  assign data_o[945] = data_o[17];
  assign data_o[977] = data_o[17];
  assign data_o[1009] = data_o[17];
  assign data_o[1041] = data_o[17];
  assign data_o[1073] = data_o[17];
  assign data_o[1105] = data_o[17];
  assign data_o[1137] = data_o[17];
  assign data_o[1169] = data_o[17];
  assign data_o[1201] = data_o[17];
  assign data_o[1233] = data_o[17];
  assign data_o[1265] = data_o[17];
  assign data_o[1297] = data_o[17];
  assign data_o[1329] = data_o[17];
  assign data_o[1361] = data_o[17];
  assign data_o[1393] = data_o[17];
  assign data_o[1425] = data_o[17];
  assign data_o[1457] = data_o[17];
  assign data_o[1489] = data_o[17];
  assign data_o[1521] = data_o[17];
  assign data_o[1553] = data_o[17];
  assign data_o[1585] = data_o[17];
  assign data_o[48] = data_o[16];
  assign data_o[80] = data_o[16];
  assign data_o[112] = data_o[16];
  assign data_o[144] = data_o[16];
  assign data_o[176] = data_o[16];
  assign data_o[208] = data_o[16];
  assign data_o[240] = data_o[16];
  assign data_o[272] = data_o[16];
  assign data_o[304] = data_o[16];
  assign data_o[336] = data_o[16];
  assign data_o[368] = data_o[16];
  assign data_o[400] = data_o[16];
  assign data_o[432] = data_o[16];
  assign data_o[464] = data_o[16];
  assign data_o[496] = data_o[16];
  assign data_o[528] = data_o[16];
  assign data_o[560] = data_o[16];
  assign data_o[592] = data_o[16];
  assign data_o[624] = data_o[16];
  assign data_o[656] = data_o[16];
  assign data_o[688] = data_o[16];
  assign data_o[720] = data_o[16];
  assign data_o[752] = data_o[16];
  assign data_o[784] = data_o[16];
  assign data_o[816] = data_o[16];
  assign data_o[848] = data_o[16];
  assign data_o[880] = data_o[16];
  assign data_o[912] = data_o[16];
  assign data_o[944] = data_o[16];
  assign data_o[976] = data_o[16];
  assign data_o[1008] = data_o[16];
  assign data_o[1040] = data_o[16];
  assign data_o[1072] = data_o[16];
  assign data_o[1104] = data_o[16];
  assign data_o[1136] = data_o[16];
  assign data_o[1168] = data_o[16];
  assign data_o[1200] = data_o[16];
  assign data_o[1232] = data_o[16];
  assign data_o[1264] = data_o[16];
  assign data_o[1296] = data_o[16];
  assign data_o[1328] = data_o[16];
  assign data_o[1360] = data_o[16];
  assign data_o[1392] = data_o[16];
  assign data_o[1424] = data_o[16];
  assign data_o[1456] = data_o[16];
  assign data_o[1488] = data_o[16];
  assign data_o[1520] = data_o[16];
  assign data_o[1552] = data_o[16];
  assign data_o[1584] = data_o[16];
  assign data_o[47] = data_o[15];
  assign data_o[79] = data_o[15];
  assign data_o[111] = data_o[15];
  assign data_o[143] = data_o[15];
  assign data_o[175] = data_o[15];
  assign data_o[207] = data_o[15];
  assign data_o[239] = data_o[15];
  assign data_o[271] = data_o[15];
  assign data_o[303] = data_o[15];
  assign data_o[335] = data_o[15];
  assign data_o[367] = data_o[15];
  assign data_o[399] = data_o[15];
  assign data_o[431] = data_o[15];
  assign data_o[463] = data_o[15];
  assign data_o[495] = data_o[15];
  assign data_o[527] = data_o[15];
  assign data_o[559] = data_o[15];
  assign data_o[591] = data_o[15];
  assign data_o[623] = data_o[15];
  assign data_o[655] = data_o[15];
  assign data_o[687] = data_o[15];
  assign data_o[719] = data_o[15];
  assign data_o[751] = data_o[15];
  assign data_o[783] = data_o[15];
  assign data_o[815] = data_o[15];
  assign data_o[847] = data_o[15];
  assign data_o[879] = data_o[15];
  assign data_o[911] = data_o[15];
  assign data_o[943] = data_o[15];
  assign data_o[975] = data_o[15];
  assign data_o[1007] = data_o[15];
  assign data_o[1039] = data_o[15];
  assign data_o[1071] = data_o[15];
  assign data_o[1103] = data_o[15];
  assign data_o[1135] = data_o[15];
  assign data_o[1167] = data_o[15];
  assign data_o[1199] = data_o[15];
  assign data_o[1231] = data_o[15];
  assign data_o[1263] = data_o[15];
  assign data_o[1295] = data_o[15];
  assign data_o[1327] = data_o[15];
  assign data_o[1359] = data_o[15];
  assign data_o[1391] = data_o[15];
  assign data_o[1423] = data_o[15];
  assign data_o[1455] = data_o[15];
  assign data_o[1487] = data_o[15];
  assign data_o[1519] = data_o[15];
  assign data_o[1551] = data_o[15];
  assign data_o[1583] = data_o[15];
  assign data_o[46] = data_o[14];
  assign data_o[78] = data_o[14];
  assign data_o[110] = data_o[14];
  assign data_o[142] = data_o[14];
  assign data_o[174] = data_o[14];
  assign data_o[206] = data_o[14];
  assign data_o[238] = data_o[14];
  assign data_o[270] = data_o[14];
  assign data_o[302] = data_o[14];
  assign data_o[334] = data_o[14];
  assign data_o[366] = data_o[14];
  assign data_o[398] = data_o[14];
  assign data_o[430] = data_o[14];
  assign data_o[462] = data_o[14];
  assign data_o[494] = data_o[14];
  assign data_o[526] = data_o[14];
  assign data_o[558] = data_o[14];
  assign data_o[590] = data_o[14];
  assign data_o[622] = data_o[14];
  assign data_o[654] = data_o[14];
  assign data_o[686] = data_o[14];
  assign data_o[718] = data_o[14];
  assign data_o[750] = data_o[14];
  assign data_o[782] = data_o[14];
  assign data_o[814] = data_o[14];
  assign data_o[846] = data_o[14];
  assign data_o[878] = data_o[14];
  assign data_o[910] = data_o[14];
  assign data_o[942] = data_o[14];
  assign data_o[974] = data_o[14];
  assign data_o[1006] = data_o[14];
  assign data_o[1038] = data_o[14];
  assign data_o[1070] = data_o[14];
  assign data_o[1102] = data_o[14];
  assign data_o[1134] = data_o[14];
  assign data_o[1166] = data_o[14];
  assign data_o[1198] = data_o[14];
  assign data_o[1230] = data_o[14];
  assign data_o[1262] = data_o[14];
  assign data_o[1294] = data_o[14];
  assign data_o[1326] = data_o[14];
  assign data_o[1358] = data_o[14];
  assign data_o[1390] = data_o[14];
  assign data_o[1422] = data_o[14];
  assign data_o[1454] = data_o[14];
  assign data_o[1486] = data_o[14];
  assign data_o[1518] = data_o[14];
  assign data_o[1550] = data_o[14];
  assign data_o[1582] = data_o[14];
  assign data_o[45] = data_o[13];
  assign data_o[77] = data_o[13];
  assign data_o[109] = data_o[13];
  assign data_o[141] = data_o[13];
  assign data_o[173] = data_o[13];
  assign data_o[205] = data_o[13];
  assign data_o[237] = data_o[13];
  assign data_o[269] = data_o[13];
  assign data_o[301] = data_o[13];
  assign data_o[333] = data_o[13];
  assign data_o[365] = data_o[13];
  assign data_o[397] = data_o[13];
  assign data_o[429] = data_o[13];
  assign data_o[461] = data_o[13];
  assign data_o[493] = data_o[13];
  assign data_o[525] = data_o[13];
  assign data_o[557] = data_o[13];
  assign data_o[589] = data_o[13];
  assign data_o[621] = data_o[13];
  assign data_o[653] = data_o[13];
  assign data_o[685] = data_o[13];
  assign data_o[717] = data_o[13];
  assign data_o[749] = data_o[13];
  assign data_o[781] = data_o[13];
  assign data_o[813] = data_o[13];
  assign data_o[845] = data_o[13];
  assign data_o[877] = data_o[13];
  assign data_o[909] = data_o[13];
  assign data_o[941] = data_o[13];
  assign data_o[973] = data_o[13];
  assign data_o[1005] = data_o[13];
  assign data_o[1037] = data_o[13];
  assign data_o[1069] = data_o[13];
  assign data_o[1101] = data_o[13];
  assign data_o[1133] = data_o[13];
  assign data_o[1165] = data_o[13];
  assign data_o[1197] = data_o[13];
  assign data_o[1229] = data_o[13];
  assign data_o[1261] = data_o[13];
  assign data_o[1293] = data_o[13];
  assign data_o[1325] = data_o[13];
  assign data_o[1357] = data_o[13];
  assign data_o[1389] = data_o[13];
  assign data_o[1421] = data_o[13];
  assign data_o[1453] = data_o[13];
  assign data_o[1485] = data_o[13];
  assign data_o[1517] = data_o[13];
  assign data_o[1549] = data_o[13];
  assign data_o[1581] = data_o[13];
  assign data_o[44] = data_o[12];
  assign data_o[76] = data_o[12];
  assign data_o[108] = data_o[12];
  assign data_o[140] = data_o[12];
  assign data_o[172] = data_o[12];
  assign data_o[204] = data_o[12];
  assign data_o[236] = data_o[12];
  assign data_o[268] = data_o[12];
  assign data_o[300] = data_o[12];
  assign data_o[332] = data_o[12];
  assign data_o[364] = data_o[12];
  assign data_o[396] = data_o[12];
  assign data_o[428] = data_o[12];
  assign data_o[460] = data_o[12];
  assign data_o[492] = data_o[12];
  assign data_o[524] = data_o[12];
  assign data_o[556] = data_o[12];
  assign data_o[588] = data_o[12];
  assign data_o[620] = data_o[12];
  assign data_o[652] = data_o[12];
  assign data_o[684] = data_o[12];
  assign data_o[716] = data_o[12];
  assign data_o[748] = data_o[12];
  assign data_o[780] = data_o[12];
  assign data_o[812] = data_o[12];
  assign data_o[844] = data_o[12];
  assign data_o[876] = data_o[12];
  assign data_o[908] = data_o[12];
  assign data_o[940] = data_o[12];
  assign data_o[972] = data_o[12];
  assign data_o[1004] = data_o[12];
  assign data_o[1036] = data_o[12];
  assign data_o[1068] = data_o[12];
  assign data_o[1100] = data_o[12];
  assign data_o[1132] = data_o[12];
  assign data_o[1164] = data_o[12];
  assign data_o[1196] = data_o[12];
  assign data_o[1228] = data_o[12];
  assign data_o[1260] = data_o[12];
  assign data_o[1292] = data_o[12];
  assign data_o[1324] = data_o[12];
  assign data_o[1356] = data_o[12];
  assign data_o[1388] = data_o[12];
  assign data_o[1420] = data_o[12];
  assign data_o[1452] = data_o[12];
  assign data_o[1484] = data_o[12];
  assign data_o[1516] = data_o[12];
  assign data_o[1548] = data_o[12];
  assign data_o[1580] = data_o[12];
  assign data_o[43] = data_o[11];
  assign data_o[75] = data_o[11];
  assign data_o[107] = data_o[11];
  assign data_o[139] = data_o[11];
  assign data_o[171] = data_o[11];
  assign data_o[203] = data_o[11];
  assign data_o[235] = data_o[11];
  assign data_o[267] = data_o[11];
  assign data_o[299] = data_o[11];
  assign data_o[331] = data_o[11];
  assign data_o[363] = data_o[11];
  assign data_o[395] = data_o[11];
  assign data_o[427] = data_o[11];
  assign data_o[459] = data_o[11];
  assign data_o[491] = data_o[11];
  assign data_o[523] = data_o[11];
  assign data_o[555] = data_o[11];
  assign data_o[587] = data_o[11];
  assign data_o[619] = data_o[11];
  assign data_o[651] = data_o[11];
  assign data_o[683] = data_o[11];
  assign data_o[715] = data_o[11];
  assign data_o[747] = data_o[11];
  assign data_o[779] = data_o[11];
  assign data_o[811] = data_o[11];
  assign data_o[843] = data_o[11];
  assign data_o[875] = data_o[11];
  assign data_o[907] = data_o[11];
  assign data_o[939] = data_o[11];
  assign data_o[971] = data_o[11];
  assign data_o[1003] = data_o[11];
  assign data_o[1035] = data_o[11];
  assign data_o[1067] = data_o[11];
  assign data_o[1099] = data_o[11];
  assign data_o[1131] = data_o[11];
  assign data_o[1163] = data_o[11];
  assign data_o[1195] = data_o[11];
  assign data_o[1227] = data_o[11];
  assign data_o[1259] = data_o[11];
  assign data_o[1291] = data_o[11];
  assign data_o[1323] = data_o[11];
  assign data_o[1355] = data_o[11];
  assign data_o[1387] = data_o[11];
  assign data_o[1419] = data_o[11];
  assign data_o[1451] = data_o[11];
  assign data_o[1483] = data_o[11];
  assign data_o[1515] = data_o[11];
  assign data_o[1547] = data_o[11];
  assign data_o[1579] = data_o[11];
  assign data_o[42] = data_o[10];
  assign data_o[74] = data_o[10];
  assign data_o[106] = data_o[10];
  assign data_o[138] = data_o[10];
  assign data_o[170] = data_o[10];
  assign data_o[202] = data_o[10];
  assign data_o[234] = data_o[10];
  assign data_o[266] = data_o[10];
  assign data_o[298] = data_o[10];
  assign data_o[330] = data_o[10];
  assign data_o[362] = data_o[10];
  assign data_o[394] = data_o[10];
  assign data_o[426] = data_o[10];
  assign data_o[458] = data_o[10];
  assign data_o[490] = data_o[10];
  assign data_o[522] = data_o[10];
  assign data_o[554] = data_o[10];
  assign data_o[586] = data_o[10];
  assign data_o[618] = data_o[10];
  assign data_o[650] = data_o[10];
  assign data_o[682] = data_o[10];
  assign data_o[714] = data_o[10];
  assign data_o[746] = data_o[10];
  assign data_o[778] = data_o[10];
  assign data_o[810] = data_o[10];
  assign data_o[842] = data_o[10];
  assign data_o[874] = data_o[10];
  assign data_o[906] = data_o[10];
  assign data_o[938] = data_o[10];
  assign data_o[970] = data_o[10];
  assign data_o[1002] = data_o[10];
  assign data_o[1034] = data_o[10];
  assign data_o[1066] = data_o[10];
  assign data_o[1098] = data_o[10];
  assign data_o[1130] = data_o[10];
  assign data_o[1162] = data_o[10];
  assign data_o[1194] = data_o[10];
  assign data_o[1226] = data_o[10];
  assign data_o[1258] = data_o[10];
  assign data_o[1290] = data_o[10];
  assign data_o[1322] = data_o[10];
  assign data_o[1354] = data_o[10];
  assign data_o[1386] = data_o[10];
  assign data_o[1418] = data_o[10];
  assign data_o[1450] = data_o[10];
  assign data_o[1482] = data_o[10];
  assign data_o[1514] = data_o[10];
  assign data_o[1546] = data_o[10];
  assign data_o[1578] = data_o[10];
  assign data_o[41] = data_o[9];
  assign data_o[73] = data_o[9];
  assign data_o[105] = data_o[9];
  assign data_o[137] = data_o[9];
  assign data_o[169] = data_o[9];
  assign data_o[201] = data_o[9];
  assign data_o[233] = data_o[9];
  assign data_o[265] = data_o[9];
  assign data_o[297] = data_o[9];
  assign data_o[329] = data_o[9];
  assign data_o[361] = data_o[9];
  assign data_o[393] = data_o[9];
  assign data_o[425] = data_o[9];
  assign data_o[457] = data_o[9];
  assign data_o[489] = data_o[9];
  assign data_o[521] = data_o[9];
  assign data_o[553] = data_o[9];
  assign data_o[585] = data_o[9];
  assign data_o[617] = data_o[9];
  assign data_o[649] = data_o[9];
  assign data_o[681] = data_o[9];
  assign data_o[713] = data_o[9];
  assign data_o[745] = data_o[9];
  assign data_o[777] = data_o[9];
  assign data_o[809] = data_o[9];
  assign data_o[841] = data_o[9];
  assign data_o[873] = data_o[9];
  assign data_o[905] = data_o[9];
  assign data_o[937] = data_o[9];
  assign data_o[969] = data_o[9];
  assign data_o[1001] = data_o[9];
  assign data_o[1033] = data_o[9];
  assign data_o[1065] = data_o[9];
  assign data_o[1097] = data_o[9];
  assign data_o[1129] = data_o[9];
  assign data_o[1161] = data_o[9];
  assign data_o[1193] = data_o[9];
  assign data_o[1225] = data_o[9];
  assign data_o[1257] = data_o[9];
  assign data_o[1289] = data_o[9];
  assign data_o[1321] = data_o[9];
  assign data_o[1353] = data_o[9];
  assign data_o[1385] = data_o[9];
  assign data_o[1417] = data_o[9];
  assign data_o[1449] = data_o[9];
  assign data_o[1481] = data_o[9];
  assign data_o[1513] = data_o[9];
  assign data_o[1545] = data_o[9];
  assign data_o[1577] = data_o[9];
  assign data_o[40] = data_o[8];
  assign data_o[72] = data_o[8];
  assign data_o[104] = data_o[8];
  assign data_o[136] = data_o[8];
  assign data_o[168] = data_o[8];
  assign data_o[200] = data_o[8];
  assign data_o[232] = data_o[8];
  assign data_o[264] = data_o[8];
  assign data_o[296] = data_o[8];
  assign data_o[328] = data_o[8];
  assign data_o[360] = data_o[8];
  assign data_o[392] = data_o[8];
  assign data_o[424] = data_o[8];
  assign data_o[456] = data_o[8];
  assign data_o[488] = data_o[8];
  assign data_o[520] = data_o[8];
  assign data_o[552] = data_o[8];
  assign data_o[584] = data_o[8];
  assign data_o[616] = data_o[8];
  assign data_o[648] = data_o[8];
  assign data_o[680] = data_o[8];
  assign data_o[712] = data_o[8];
  assign data_o[744] = data_o[8];
  assign data_o[776] = data_o[8];
  assign data_o[808] = data_o[8];
  assign data_o[840] = data_o[8];
  assign data_o[872] = data_o[8];
  assign data_o[904] = data_o[8];
  assign data_o[936] = data_o[8];
  assign data_o[968] = data_o[8];
  assign data_o[1000] = data_o[8];
  assign data_o[1032] = data_o[8];
  assign data_o[1064] = data_o[8];
  assign data_o[1096] = data_o[8];
  assign data_o[1128] = data_o[8];
  assign data_o[1160] = data_o[8];
  assign data_o[1192] = data_o[8];
  assign data_o[1224] = data_o[8];
  assign data_o[1256] = data_o[8];
  assign data_o[1288] = data_o[8];
  assign data_o[1320] = data_o[8];
  assign data_o[1352] = data_o[8];
  assign data_o[1384] = data_o[8];
  assign data_o[1416] = data_o[8];
  assign data_o[1448] = data_o[8];
  assign data_o[1480] = data_o[8];
  assign data_o[1512] = data_o[8];
  assign data_o[1544] = data_o[8];
  assign data_o[1576] = data_o[8];
  assign data_o[39] = data_o[7];
  assign data_o[71] = data_o[7];
  assign data_o[103] = data_o[7];
  assign data_o[135] = data_o[7];
  assign data_o[167] = data_o[7];
  assign data_o[199] = data_o[7];
  assign data_o[231] = data_o[7];
  assign data_o[263] = data_o[7];
  assign data_o[295] = data_o[7];
  assign data_o[327] = data_o[7];
  assign data_o[359] = data_o[7];
  assign data_o[391] = data_o[7];
  assign data_o[423] = data_o[7];
  assign data_o[455] = data_o[7];
  assign data_o[487] = data_o[7];
  assign data_o[519] = data_o[7];
  assign data_o[551] = data_o[7];
  assign data_o[583] = data_o[7];
  assign data_o[615] = data_o[7];
  assign data_o[647] = data_o[7];
  assign data_o[679] = data_o[7];
  assign data_o[711] = data_o[7];
  assign data_o[743] = data_o[7];
  assign data_o[775] = data_o[7];
  assign data_o[807] = data_o[7];
  assign data_o[839] = data_o[7];
  assign data_o[871] = data_o[7];
  assign data_o[903] = data_o[7];
  assign data_o[935] = data_o[7];
  assign data_o[967] = data_o[7];
  assign data_o[999] = data_o[7];
  assign data_o[1031] = data_o[7];
  assign data_o[1063] = data_o[7];
  assign data_o[1095] = data_o[7];
  assign data_o[1127] = data_o[7];
  assign data_o[1159] = data_o[7];
  assign data_o[1191] = data_o[7];
  assign data_o[1223] = data_o[7];
  assign data_o[1255] = data_o[7];
  assign data_o[1287] = data_o[7];
  assign data_o[1319] = data_o[7];
  assign data_o[1351] = data_o[7];
  assign data_o[1383] = data_o[7];
  assign data_o[1415] = data_o[7];
  assign data_o[1447] = data_o[7];
  assign data_o[1479] = data_o[7];
  assign data_o[1511] = data_o[7];
  assign data_o[1543] = data_o[7];
  assign data_o[1575] = data_o[7];
  assign data_o[38] = data_o[6];
  assign data_o[70] = data_o[6];
  assign data_o[102] = data_o[6];
  assign data_o[134] = data_o[6];
  assign data_o[166] = data_o[6];
  assign data_o[198] = data_o[6];
  assign data_o[230] = data_o[6];
  assign data_o[262] = data_o[6];
  assign data_o[294] = data_o[6];
  assign data_o[326] = data_o[6];
  assign data_o[358] = data_o[6];
  assign data_o[390] = data_o[6];
  assign data_o[422] = data_o[6];
  assign data_o[454] = data_o[6];
  assign data_o[486] = data_o[6];
  assign data_o[518] = data_o[6];
  assign data_o[550] = data_o[6];
  assign data_o[582] = data_o[6];
  assign data_o[614] = data_o[6];
  assign data_o[646] = data_o[6];
  assign data_o[678] = data_o[6];
  assign data_o[710] = data_o[6];
  assign data_o[742] = data_o[6];
  assign data_o[774] = data_o[6];
  assign data_o[806] = data_o[6];
  assign data_o[838] = data_o[6];
  assign data_o[870] = data_o[6];
  assign data_o[902] = data_o[6];
  assign data_o[934] = data_o[6];
  assign data_o[966] = data_o[6];
  assign data_o[998] = data_o[6];
  assign data_o[1030] = data_o[6];
  assign data_o[1062] = data_o[6];
  assign data_o[1094] = data_o[6];
  assign data_o[1126] = data_o[6];
  assign data_o[1158] = data_o[6];
  assign data_o[1190] = data_o[6];
  assign data_o[1222] = data_o[6];
  assign data_o[1254] = data_o[6];
  assign data_o[1286] = data_o[6];
  assign data_o[1318] = data_o[6];
  assign data_o[1350] = data_o[6];
  assign data_o[1382] = data_o[6];
  assign data_o[1414] = data_o[6];
  assign data_o[1446] = data_o[6];
  assign data_o[1478] = data_o[6];
  assign data_o[1510] = data_o[6];
  assign data_o[1542] = data_o[6];
  assign data_o[1574] = data_o[6];
  assign data_o[37] = data_o[5];
  assign data_o[69] = data_o[5];
  assign data_o[101] = data_o[5];
  assign data_o[133] = data_o[5];
  assign data_o[165] = data_o[5];
  assign data_o[197] = data_o[5];
  assign data_o[229] = data_o[5];
  assign data_o[261] = data_o[5];
  assign data_o[293] = data_o[5];
  assign data_o[325] = data_o[5];
  assign data_o[357] = data_o[5];
  assign data_o[389] = data_o[5];
  assign data_o[421] = data_o[5];
  assign data_o[453] = data_o[5];
  assign data_o[485] = data_o[5];
  assign data_o[517] = data_o[5];
  assign data_o[549] = data_o[5];
  assign data_o[581] = data_o[5];
  assign data_o[613] = data_o[5];
  assign data_o[645] = data_o[5];
  assign data_o[677] = data_o[5];
  assign data_o[709] = data_o[5];
  assign data_o[741] = data_o[5];
  assign data_o[773] = data_o[5];
  assign data_o[805] = data_o[5];
  assign data_o[837] = data_o[5];
  assign data_o[869] = data_o[5];
  assign data_o[901] = data_o[5];
  assign data_o[933] = data_o[5];
  assign data_o[965] = data_o[5];
  assign data_o[997] = data_o[5];
  assign data_o[1029] = data_o[5];
  assign data_o[1061] = data_o[5];
  assign data_o[1093] = data_o[5];
  assign data_o[1125] = data_o[5];
  assign data_o[1157] = data_o[5];
  assign data_o[1189] = data_o[5];
  assign data_o[1221] = data_o[5];
  assign data_o[1253] = data_o[5];
  assign data_o[1285] = data_o[5];
  assign data_o[1317] = data_o[5];
  assign data_o[1349] = data_o[5];
  assign data_o[1381] = data_o[5];
  assign data_o[1413] = data_o[5];
  assign data_o[1445] = data_o[5];
  assign data_o[1477] = data_o[5];
  assign data_o[1509] = data_o[5];
  assign data_o[1541] = data_o[5];
  assign data_o[1573] = data_o[5];
  assign data_o[36] = data_o[4];
  assign data_o[68] = data_o[4];
  assign data_o[100] = data_o[4];
  assign data_o[132] = data_o[4];
  assign data_o[164] = data_o[4];
  assign data_o[196] = data_o[4];
  assign data_o[228] = data_o[4];
  assign data_o[260] = data_o[4];
  assign data_o[292] = data_o[4];
  assign data_o[324] = data_o[4];
  assign data_o[356] = data_o[4];
  assign data_o[388] = data_o[4];
  assign data_o[420] = data_o[4];
  assign data_o[452] = data_o[4];
  assign data_o[484] = data_o[4];
  assign data_o[516] = data_o[4];
  assign data_o[548] = data_o[4];
  assign data_o[580] = data_o[4];
  assign data_o[612] = data_o[4];
  assign data_o[644] = data_o[4];
  assign data_o[676] = data_o[4];
  assign data_o[708] = data_o[4];
  assign data_o[740] = data_o[4];
  assign data_o[772] = data_o[4];
  assign data_o[804] = data_o[4];
  assign data_o[836] = data_o[4];
  assign data_o[868] = data_o[4];
  assign data_o[900] = data_o[4];
  assign data_o[932] = data_o[4];
  assign data_o[964] = data_o[4];
  assign data_o[996] = data_o[4];
  assign data_o[1028] = data_o[4];
  assign data_o[1060] = data_o[4];
  assign data_o[1092] = data_o[4];
  assign data_o[1124] = data_o[4];
  assign data_o[1156] = data_o[4];
  assign data_o[1188] = data_o[4];
  assign data_o[1220] = data_o[4];
  assign data_o[1252] = data_o[4];
  assign data_o[1284] = data_o[4];
  assign data_o[1316] = data_o[4];
  assign data_o[1348] = data_o[4];
  assign data_o[1380] = data_o[4];
  assign data_o[1412] = data_o[4];
  assign data_o[1444] = data_o[4];
  assign data_o[1476] = data_o[4];
  assign data_o[1508] = data_o[4];
  assign data_o[1540] = data_o[4];
  assign data_o[1572] = data_o[4];
  assign data_o[35] = data_o[3];
  assign data_o[67] = data_o[3];
  assign data_o[99] = data_o[3];
  assign data_o[131] = data_o[3];
  assign data_o[163] = data_o[3];
  assign data_o[195] = data_o[3];
  assign data_o[227] = data_o[3];
  assign data_o[259] = data_o[3];
  assign data_o[291] = data_o[3];
  assign data_o[323] = data_o[3];
  assign data_o[355] = data_o[3];
  assign data_o[387] = data_o[3];
  assign data_o[419] = data_o[3];
  assign data_o[451] = data_o[3];
  assign data_o[483] = data_o[3];
  assign data_o[515] = data_o[3];
  assign data_o[547] = data_o[3];
  assign data_o[579] = data_o[3];
  assign data_o[611] = data_o[3];
  assign data_o[643] = data_o[3];
  assign data_o[675] = data_o[3];
  assign data_o[707] = data_o[3];
  assign data_o[739] = data_o[3];
  assign data_o[771] = data_o[3];
  assign data_o[803] = data_o[3];
  assign data_o[835] = data_o[3];
  assign data_o[867] = data_o[3];
  assign data_o[899] = data_o[3];
  assign data_o[931] = data_o[3];
  assign data_o[963] = data_o[3];
  assign data_o[995] = data_o[3];
  assign data_o[1027] = data_o[3];
  assign data_o[1059] = data_o[3];
  assign data_o[1091] = data_o[3];
  assign data_o[1123] = data_o[3];
  assign data_o[1155] = data_o[3];
  assign data_o[1187] = data_o[3];
  assign data_o[1219] = data_o[3];
  assign data_o[1251] = data_o[3];
  assign data_o[1283] = data_o[3];
  assign data_o[1315] = data_o[3];
  assign data_o[1347] = data_o[3];
  assign data_o[1379] = data_o[3];
  assign data_o[1411] = data_o[3];
  assign data_o[1443] = data_o[3];
  assign data_o[1475] = data_o[3];
  assign data_o[1507] = data_o[3];
  assign data_o[1539] = data_o[3];
  assign data_o[1571] = data_o[3];
  assign data_o[34] = data_o[2];
  assign data_o[66] = data_o[2];
  assign data_o[98] = data_o[2];
  assign data_o[130] = data_o[2];
  assign data_o[162] = data_o[2];
  assign data_o[194] = data_o[2];
  assign data_o[226] = data_o[2];
  assign data_o[258] = data_o[2];
  assign data_o[290] = data_o[2];
  assign data_o[322] = data_o[2];
  assign data_o[354] = data_o[2];
  assign data_o[386] = data_o[2];
  assign data_o[418] = data_o[2];
  assign data_o[450] = data_o[2];
  assign data_o[482] = data_o[2];
  assign data_o[514] = data_o[2];
  assign data_o[546] = data_o[2];
  assign data_o[578] = data_o[2];
  assign data_o[610] = data_o[2];
  assign data_o[642] = data_o[2];
  assign data_o[674] = data_o[2];
  assign data_o[706] = data_o[2];
  assign data_o[738] = data_o[2];
  assign data_o[770] = data_o[2];
  assign data_o[802] = data_o[2];
  assign data_o[834] = data_o[2];
  assign data_o[866] = data_o[2];
  assign data_o[898] = data_o[2];
  assign data_o[930] = data_o[2];
  assign data_o[962] = data_o[2];
  assign data_o[994] = data_o[2];
  assign data_o[1026] = data_o[2];
  assign data_o[1058] = data_o[2];
  assign data_o[1090] = data_o[2];
  assign data_o[1122] = data_o[2];
  assign data_o[1154] = data_o[2];
  assign data_o[1186] = data_o[2];
  assign data_o[1218] = data_o[2];
  assign data_o[1250] = data_o[2];
  assign data_o[1282] = data_o[2];
  assign data_o[1314] = data_o[2];
  assign data_o[1346] = data_o[2];
  assign data_o[1378] = data_o[2];
  assign data_o[1410] = data_o[2];
  assign data_o[1442] = data_o[2];
  assign data_o[1474] = data_o[2];
  assign data_o[1506] = data_o[2];
  assign data_o[1538] = data_o[2];
  assign data_o[1570] = data_o[2];
  assign data_o[33] = data_o[1];
  assign data_o[65] = data_o[1];
  assign data_o[97] = data_o[1];
  assign data_o[129] = data_o[1];
  assign data_o[161] = data_o[1];
  assign data_o[193] = data_o[1];
  assign data_o[225] = data_o[1];
  assign data_o[257] = data_o[1];
  assign data_o[289] = data_o[1];
  assign data_o[321] = data_o[1];
  assign data_o[353] = data_o[1];
  assign data_o[385] = data_o[1];
  assign data_o[417] = data_o[1];
  assign data_o[449] = data_o[1];
  assign data_o[481] = data_o[1];
  assign data_o[513] = data_o[1];
  assign data_o[545] = data_o[1];
  assign data_o[577] = data_o[1];
  assign data_o[609] = data_o[1];
  assign data_o[641] = data_o[1];
  assign data_o[673] = data_o[1];
  assign data_o[705] = data_o[1];
  assign data_o[737] = data_o[1];
  assign data_o[769] = data_o[1];
  assign data_o[801] = data_o[1];
  assign data_o[833] = data_o[1];
  assign data_o[865] = data_o[1];
  assign data_o[897] = data_o[1];
  assign data_o[929] = data_o[1];
  assign data_o[961] = data_o[1];
  assign data_o[993] = data_o[1];
  assign data_o[1025] = data_o[1];
  assign data_o[1057] = data_o[1];
  assign data_o[1089] = data_o[1];
  assign data_o[1121] = data_o[1];
  assign data_o[1153] = data_o[1];
  assign data_o[1185] = data_o[1];
  assign data_o[1217] = data_o[1];
  assign data_o[1249] = data_o[1];
  assign data_o[1281] = data_o[1];
  assign data_o[1313] = data_o[1];
  assign data_o[1345] = data_o[1];
  assign data_o[1377] = data_o[1];
  assign data_o[1409] = data_o[1];
  assign data_o[1441] = data_o[1];
  assign data_o[1473] = data_o[1];
  assign data_o[1505] = data_o[1];
  assign data_o[1537] = data_o[1];
  assign data_o[1569] = data_o[1];
  assign data_o[32] = data_o[0];
  assign data_o[64] = data_o[0];
  assign data_o[96] = data_o[0];
  assign data_o[128] = data_o[0];
  assign data_o[160] = data_o[0];
  assign data_o[192] = data_o[0];
  assign data_o[224] = data_o[0];
  assign data_o[256] = data_o[0];
  assign data_o[288] = data_o[0];
  assign data_o[320] = data_o[0];
  assign data_o[352] = data_o[0];
  assign data_o[384] = data_o[0];
  assign data_o[416] = data_o[0];
  assign data_o[448] = data_o[0];
  assign data_o[480] = data_o[0];
  assign data_o[512] = data_o[0];
  assign data_o[544] = data_o[0];
  assign data_o[576] = data_o[0];
  assign data_o[608] = data_o[0];
  assign data_o[640] = data_o[0];
  assign data_o[672] = data_o[0];
  assign data_o[704] = data_o[0];
  assign data_o[736] = data_o[0];
  assign data_o[768] = data_o[0];
  assign data_o[800] = data_o[0];
  assign data_o[832] = data_o[0];
  assign data_o[864] = data_o[0];
  assign data_o[896] = data_o[0];
  assign data_o[928] = data_o[0];
  assign data_o[960] = data_o[0];
  assign data_o[992] = data_o[0];
  assign data_o[1024] = data_o[0];
  assign data_o[1056] = data_o[0];
  assign data_o[1088] = data_o[0];
  assign data_o[1120] = data_o[0];
  assign data_o[1152] = data_o[0];
  assign data_o[1184] = data_o[0];
  assign data_o[1216] = data_o[0];
  assign data_o[1248] = data_o[0];
  assign data_o[1280] = data_o[0];
  assign data_o[1312] = data_o[0];
  assign data_o[1344] = data_o[0];
  assign data_o[1376] = data_o[0];
  assign data_o[1408] = data_o[0];
  assign data_o[1440] = data_o[0];
  assign data_o[1472] = data_o[0];
  assign data_o[1504] = data_o[0];
  assign data_o[1536] = data_o[0];
  assign data_o[1568] = data_o[0];

  bsg_two_fifo_width_p32
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_i(v_i),
    .v_o(fifo_v),
    .data_o(data_o[31:0]),
    .yumi_i(fifo_yumi)
  );

  assign N153 = (N0)? 1'b0 : 
                (N1)? N152 : 1'b0;
  assign N0 = N151;
  assign N1 = N150;
  assign sent_n[0] = (N2)? 1'b1 : 
                     (N155)? sent_r[0] : 1'b0;
  assign N2 = N154;
  assign N159 = (N3)? 1'b0 : 
                (N4)? N158 : 1'b0;
  assign N3 = N157;
  assign N4 = N156;
  assign sent_n[1] = (N5)? 1'b1 : 
                     (N161)? sent_r[1] : 1'b0;
  assign N5 = N160;
  assign N165 = (N6)? 1'b0 : 
                (N7)? N164 : 1'b0;
  assign N6 = N163;
  assign N7 = N162;
  assign sent_n[2] = (N8)? 1'b1 : 
                     (N167)? sent_r[2] : 1'b0;
  assign N8 = N166;
  assign N171 = (N9)? 1'b0 : 
                (N10)? N170 : 1'b0;
  assign N9 = N169;
  assign N10 = N168;
  assign sent_n[3] = (N11)? 1'b1 : 
                     (N173)? sent_r[3] : 1'b0;
  assign N11 = N172;
  assign N177 = (N12)? 1'b0 : 
                (N13)? N176 : 1'b0;
  assign N12 = N175;
  assign N13 = N174;
  assign sent_n[4] = (N14)? 1'b1 : 
                     (N179)? sent_r[4] : 1'b0;
  assign N14 = N178;
  assign N183 = (N15)? 1'b0 : 
                (N16)? N182 : 1'b0;
  assign N15 = N181;
  assign N16 = N180;
  assign sent_n[5] = (N17)? 1'b1 : 
                     (N185)? sent_r[5] : 1'b0;
  assign N17 = N184;
  assign N189 = (N18)? 1'b0 : 
                (N19)? N188 : 1'b0;
  assign N18 = N187;
  assign N19 = N186;
  assign sent_n[6] = (N20)? 1'b1 : 
                     (N191)? sent_r[6] : 1'b0;
  assign N20 = N190;
  assign N195 = (N21)? 1'b0 : 
                (N22)? N194 : 1'b0;
  assign N21 = N193;
  assign N22 = N192;
  assign sent_n[7] = (N23)? 1'b1 : 
                     (N197)? sent_r[7] : 1'b0;
  assign N23 = N196;
  assign N201 = (N24)? 1'b0 : 
                (N25)? N200 : 1'b0;
  assign N24 = N199;
  assign N25 = N198;
  assign sent_n[8] = (N26)? 1'b1 : 
                     (N203)? sent_r[8] : 1'b0;
  assign N26 = N202;
  assign N207 = (N27)? 1'b0 : 
                (N28)? N206 : 1'b0;
  assign N27 = N205;
  assign N28 = N204;
  assign sent_n[9] = (N29)? 1'b1 : 
                     (N209)? sent_r[9] : 1'b0;
  assign N29 = N208;
  assign N213 = (N30)? 1'b0 : 
                (N31)? N212 : 1'b0;
  assign N30 = N211;
  assign N31 = N210;
  assign sent_n[10] = (N32)? 1'b1 : 
                      (N215)? sent_r[10] : 1'b0;
  assign N32 = N214;
  assign N219 = (N33)? 1'b0 : 
                (N34)? N218 : 1'b0;
  assign N33 = N217;
  assign N34 = N216;
  assign sent_n[11] = (N35)? 1'b1 : 
                      (N221)? sent_r[11] : 1'b0;
  assign N35 = N220;
  assign N225 = (N36)? 1'b0 : 
                (N37)? N224 : 1'b0;
  assign N36 = N223;
  assign N37 = N222;
  assign sent_n[12] = (N38)? 1'b1 : 
                      (N227)? sent_r[12] : 1'b0;
  assign N38 = N226;
  assign N231 = (N39)? 1'b0 : 
                (N40)? N230 : 1'b0;
  assign N39 = N229;
  assign N40 = N228;
  assign sent_n[13] = (N41)? 1'b1 : 
                      (N233)? sent_r[13] : 1'b0;
  assign N41 = N232;
  assign N237 = (N42)? 1'b0 : 
                (N43)? N236 : 1'b0;
  assign N42 = N235;
  assign N43 = N234;
  assign sent_n[14] = (N44)? 1'b1 : 
                      (N239)? sent_r[14] : 1'b0;
  assign N44 = N238;
  assign N243 = (N45)? 1'b0 : 
                (N46)? N242 : 1'b0;
  assign N45 = N241;
  assign N46 = N240;
  assign sent_n[15] = (N47)? 1'b1 : 
                      (N245)? sent_r[15] : 1'b0;
  assign N47 = N244;
  assign N249 = (N48)? 1'b0 : 
                (N49)? N248 : 1'b0;
  assign N48 = N247;
  assign N49 = N246;
  assign sent_n[16] = (N50)? 1'b1 : 
                      (N251)? sent_r[16] : 1'b0;
  assign N50 = N250;
  assign N255 = (N51)? 1'b0 : 
                (N52)? N254 : 1'b0;
  assign N51 = N253;
  assign N52 = N252;
  assign sent_n[17] = (N53)? 1'b1 : 
                      (N257)? sent_r[17] : 1'b0;
  assign N53 = N256;
  assign N261 = (N54)? 1'b0 : 
                (N55)? N260 : 1'b0;
  assign N54 = N259;
  assign N55 = N258;
  assign sent_n[18] = (N56)? 1'b1 : 
                      (N263)? sent_r[18] : 1'b0;
  assign N56 = N262;
  assign N267 = (N57)? 1'b0 : 
                (N58)? N266 : 1'b0;
  assign N57 = N265;
  assign N58 = N264;
  assign sent_n[19] = (N59)? 1'b1 : 
                      (N269)? sent_r[19] : 1'b0;
  assign N59 = N268;
  assign N273 = (N60)? 1'b0 : 
                (N61)? N272 : 1'b0;
  assign N60 = N271;
  assign N61 = N270;
  assign sent_n[20] = (N62)? 1'b1 : 
                      (N275)? sent_r[20] : 1'b0;
  assign N62 = N274;
  assign N279 = (N63)? 1'b0 : 
                (N64)? N278 : 1'b0;
  assign N63 = N277;
  assign N64 = N276;
  assign sent_n[21] = (N65)? 1'b1 : 
                      (N281)? sent_r[21] : 1'b0;
  assign N65 = N280;
  assign N285 = (N66)? 1'b0 : 
                (N67)? N284 : 1'b0;
  assign N66 = N283;
  assign N67 = N282;
  assign sent_n[22] = (N68)? 1'b1 : 
                      (N287)? sent_r[22] : 1'b0;
  assign N68 = N286;
  assign N291 = (N69)? 1'b0 : 
                (N70)? N290 : 1'b0;
  assign N69 = N289;
  assign N70 = N288;
  assign sent_n[23] = (N71)? 1'b1 : 
                      (N293)? sent_r[23] : 1'b0;
  assign N71 = N292;
  assign N297 = (N72)? 1'b0 : 
                (N73)? N296 : 1'b0;
  assign N72 = N295;
  assign N73 = N294;
  assign sent_n[24] = (N74)? 1'b1 : 
                      (N299)? sent_r[24] : 1'b0;
  assign N74 = N298;
  assign N303 = (N75)? 1'b0 : 
                (N76)? N302 : 1'b0;
  assign N75 = N301;
  assign N76 = N300;
  assign sent_n[25] = (N77)? 1'b1 : 
                      (N305)? sent_r[25] : 1'b0;
  assign N77 = N304;
  assign N309 = (N78)? 1'b0 : 
                (N79)? N308 : 1'b0;
  assign N78 = N307;
  assign N79 = N306;
  assign sent_n[26] = (N80)? 1'b1 : 
                      (N311)? sent_r[26] : 1'b0;
  assign N80 = N310;
  assign N315 = (N81)? 1'b0 : 
                (N82)? N314 : 1'b0;
  assign N81 = N313;
  assign N82 = N312;
  assign sent_n[27] = (N83)? 1'b1 : 
                      (N317)? sent_r[27] : 1'b0;
  assign N83 = N316;
  assign N321 = (N84)? 1'b0 : 
                (N85)? N320 : 1'b0;
  assign N84 = N319;
  assign N85 = N318;
  assign sent_n[28] = (N86)? 1'b1 : 
                      (N323)? sent_r[28] : 1'b0;
  assign N86 = N322;
  assign N327 = (N87)? 1'b0 : 
                (N88)? N326 : 1'b0;
  assign N87 = N325;
  assign N88 = N324;
  assign sent_n[29] = (N89)? 1'b1 : 
                      (N329)? sent_r[29] : 1'b0;
  assign N89 = N328;
  assign N333 = (N90)? 1'b0 : 
                (N91)? N332 : 1'b0;
  assign N90 = N331;
  assign N91 = N330;
  assign sent_n[30] = (N92)? 1'b1 : 
                      (N335)? sent_r[30] : 1'b0;
  assign N92 = N334;
  assign N339 = (N93)? 1'b0 : 
                (N94)? N338 : 1'b0;
  assign N93 = N337;
  assign N94 = N336;
  assign sent_n[31] = (N95)? 1'b1 : 
                      (N341)? sent_r[31] : 1'b0;
  assign N95 = N340;
  assign N345 = (N96)? 1'b0 : 
                (N97)? N344 : 1'b0;
  assign N96 = N343;
  assign N97 = N342;
  assign sent_n[32] = (N98)? 1'b1 : 
                      (N347)? sent_r[32] : 1'b0;
  assign N98 = N346;
  assign N351 = (N99)? 1'b0 : 
                (N100)? N350 : 1'b0;
  assign N99 = N349;
  assign N100 = N348;
  assign sent_n[33] = (N101)? 1'b1 : 
                      (N353)? sent_r[33] : 1'b0;
  assign N101 = N352;
  assign N357 = (N102)? 1'b0 : 
                (N103)? N356 : 1'b0;
  assign N102 = N355;
  assign N103 = N354;
  assign sent_n[34] = (N104)? 1'b1 : 
                      (N359)? sent_r[34] : 1'b0;
  assign N104 = N358;
  assign N363 = (N105)? 1'b0 : 
                (N106)? N362 : 1'b0;
  assign N105 = N361;
  assign N106 = N360;
  assign sent_n[35] = (N107)? 1'b1 : 
                      (N365)? sent_r[35] : 1'b0;
  assign N107 = N364;
  assign N369 = (N108)? 1'b0 : 
                (N109)? N368 : 1'b0;
  assign N108 = N367;
  assign N109 = N366;
  assign sent_n[36] = (N110)? 1'b1 : 
                      (N371)? sent_r[36] : 1'b0;
  assign N110 = N370;
  assign N375 = (N111)? 1'b0 : 
                (N112)? N374 : 1'b0;
  assign N111 = N373;
  assign N112 = N372;
  assign sent_n[37] = (N113)? 1'b1 : 
                      (N377)? sent_r[37] : 1'b0;
  assign N113 = N376;
  assign N381 = (N114)? 1'b0 : 
                (N115)? N380 : 1'b0;
  assign N114 = N379;
  assign N115 = N378;
  assign sent_n[38] = (N116)? 1'b1 : 
                      (N383)? sent_r[38] : 1'b0;
  assign N116 = N382;
  assign N387 = (N117)? 1'b0 : 
                (N118)? N386 : 1'b0;
  assign N117 = N385;
  assign N118 = N384;
  assign sent_n[39] = (N119)? 1'b1 : 
                      (N389)? sent_r[39] : 1'b0;
  assign N119 = N388;
  assign N393 = (N120)? 1'b0 : 
                (N121)? N392 : 1'b0;
  assign N120 = N391;
  assign N121 = N390;
  assign sent_n[40] = (N122)? 1'b1 : 
                      (N395)? sent_r[40] : 1'b0;
  assign N122 = N394;
  assign N399 = (N123)? 1'b0 : 
                (N124)? N398 : 1'b0;
  assign N123 = N397;
  assign N124 = N396;
  assign sent_n[41] = (N125)? 1'b1 : 
                      (N401)? sent_r[41] : 1'b0;
  assign N125 = N400;
  assign N405 = (N126)? 1'b0 : 
                (N127)? N404 : 1'b0;
  assign N126 = N403;
  assign N127 = N402;
  assign sent_n[42] = (N128)? 1'b1 : 
                      (N407)? sent_r[42] : 1'b0;
  assign N128 = N406;
  assign N411 = (N129)? 1'b0 : 
                (N130)? N410 : 1'b0;
  assign N129 = N409;
  assign N130 = N408;
  assign sent_n[43] = (N131)? 1'b1 : 
                      (N413)? sent_r[43] : 1'b0;
  assign N131 = N412;
  assign N417 = (N132)? 1'b0 : 
                (N133)? N416 : 1'b0;
  assign N132 = N415;
  assign N133 = N414;
  assign sent_n[44] = (N134)? 1'b1 : 
                      (N419)? sent_r[44] : 1'b0;
  assign N134 = N418;
  assign N423 = (N135)? 1'b0 : 
                (N136)? N422 : 1'b0;
  assign N135 = N421;
  assign N136 = N420;
  assign sent_n[45] = (N137)? 1'b1 : 
                      (N425)? sent_r[45] : 1'b0;
  assign N137 = N424;
  assign N429 = (N138)? 1'b0 : 
                (N139)? N428 : 1'b0;
  assign N138 = N427;
  assign N139 = N426;
  assign sent_n[46] = (N140)? 1'b1 : 
                      (N431)? sent_r[46] : 1'b0;
  assign N140 = N430;
  assign N435 = (N141)? 1'b0 : 
                (N142)? N434 : 1'b0;
  assign N141 = N433;
  assign N142 = N432;
  assign sent_n[47] = (N143)? 1'b1 : 
                      (N437)? sent_r[47] : 1'b0;
  assign N143 = N436;
  assign N441 = (N144)? 1'b0 : 
                (N145)? N440 : 1'b0;
  assign N144 = N439;
  assign N145 = N438;
  assign sent_n[48] = (N146)? 1'b1 : 
                      (N443)? sent_r[48] : 1'b0;
  assign N146 = N442;
  assign N447 = (N147)? 1'b0 : 
                (N148)? N446 : 1'b0;
  assign N147 = N445;
  assign N148 = N444;
  assign sent_n[49] = (N149)? 1'b1 : 
                      (N449)? sent_r[49] : 1'b0;
  assign N149 = N448;
  assign v_o[0] = fifo_v & N450;
  assign N450 = ~sent_r[0];
  assign N150 = ~reset_i;
  assign N151 = reset_i;
  assign N152 = sent_n[0] & N451;
  assign N451 = ~fifo_yumi;
  assign N154 = v_o[0] & ready_i[0];
  assign N155 = ~N154;
  assign v_o[1] = fifo_v & N452;
  assign N452 = ~sent_r[1];
  assign N156 = ~reset_i;
  assign N157 = reset_i;
  assign N158 = sent_n[1] & N453;
  assign N453 = ~fifo_yumi;
  assign N160 = v_o[1] & ready_i[1];
  assign N161 = ~N160;
  assign v_o[2] = fifo_v & N454;
  assign N454 = ~sent_r[2];
  assign N162 = ~reset_i;
  assign N163 = reset_i;
  assign N164 = sent_n[2] & N455;
  assign N455 = ~fifo_yumi;
  assign N166 = v_o[2] & ready_i[2];
  assign N167 = ~N166;
  assign v_o[3] = fifo_v & N456;
  assign N456 = ~sent_r[3];
  assign N168 = ~reset_i;
  assign N169 = reset_i;
  assign N170 = sent_n[3] & N457;
  assign N457 = ~fifo_yumi;
  assign N172 = v_o[3] & ready_i[3];
  assign N173 = ~N172;
  assign v_o[4] = fifo_v & N458;
  assign N458 = ~sent_r[4];
  assign N174 = ~reset_i;
  assign N175 = reset_i;
  assign N176 = sent_n[4] & N459;
  assign N459 = ~fifo_yumi;
  assign N178 = v_o[4] & ready_i[4];
  assign N179 = ~N178;
  assign v_o[5] = fifo_v & N460;
  assign N460 = ~sent_r[5];
  assign N180 = ~reset_i;
  assign N181 = reset_i;
  assign N182 = sent_n[5] & N461;
  assign N461 = ~fifo_yumi;
  assign N184 = v_o[5] & ready_i[5];
  assign N185 = ~N184;
  assign v_o[6] = fifo_v & N462;
  assign N462 = ~sent_r[6];
  assign N186 = ~reset_i;
  assign N187 = reset_i;
  assign N188 = sent_n[6] & N463;
  assign N463 = ~fifo_yumi;
  assign N190 = v_o[6] & ready_i[6];
  assign N191 = ~N190;
  assign v_o[7] = fifo_v & N464;
  assign N464 = ~sent_r[7];
  assign N192 = ~reset_i;
  assign N193 = reset_i;
  assign N194 = sent_n[7] & N465;
  assign N465 = ~fifo_yumi;
  assign N196 = v_o[7] & ready_i[7];
  assign N197 = ~N196;
  assign v_o[8] = fifo_v & N466;
  assign N466 = ~sent_r[8];
  assign N198 = ~reset_i;
  assign N199 = reset_i;
  assign N200 = sent_n[8] & N467;
  assign N467 = ~fifo_yumi;
  assign N202 = v_o[8] & ready_i[8];
  assign N203 = ~N202;
  assign v_o[9] = fifo_v & N468;
  assign N468 = ~sent_r[9];
  assign N204 = ~reset_i;
  assign N205 = reset_i;
  assign N206 = sent_n[9] & N469;
  assign N469 = ~fifo_yumi;
  assign N208 = v_o[9] & ready_i[9];
  assign N209 = ~N208;
  assign v_o[10] = fifo_v & N470;
  assign N470 = ~sent_r[10];
  assign N210 = ~reset_i;
  assign N211 = reset_i;
  assign N212 = sent_n[10] & N471;
  assign N471 = ~fifo_yumi;
  assign N214 = v_o[10] & ready_i[10];
  assign N215 = ~N214;
  assign v_o[11] = fifo_v & N472;
  assign N472 = ~sent_r[11];
  assign N216 = ~reset_i;
  assign N217 = reset_i;
  assign N218 = sent_n[11] & N473;
  assign N473 = ~fifo_yumi;
  assign N220 = v_o[11] & ready_i[11];
  assign N221 = ~N220;
  assign v_o[12] = fifo_v & N474;
  assign N474 = ~sent_r[12];
  assign N222 = ~reset_i;
  assign N223 = reset_i;
  assign N224 = sent_n[12] & N475;
  assign N475 = ~fifo_yumi;
  assign N226 = v_o[12] & ready_i[12];
  assign N227 = ~N226;
  assign v_o[13] = fifo_v & N476;
  assign N476 = ~sent_r[13];
  assign N228 = ~reset_i;
  assign N229 = reset_i;
  assign N230 = sent_n[13] & N477;
  assign N477 = ~fifo_yumi;
  assign N232 = v_o[13] & ready_i[13];
  assign N233 = ~N232;
  assign v_o[14] = fifo_v & N478;
  assign N478 = ~sent_r[14];
  assign N234 = ~reset_i;
  assign N235 = reset_i;
  assign N236 = sent_n[14] & N479;
  assign N479 = ~fifo_yumi;
  assign N238 = v_o[14] & ready_i[14];
  assign N239 = ~N238;
  assign v_o[15] = fifo_v & N480;
  assign N480 = ~sent_r[15];
  assign N240 = ~reset_i;
  assign N241 = reset_i;
  assign N242 = sent_n[15] & N481;
  assign N481 = ~fifo_yumi;
  assign N244 = v_o[15] & ready_i[15];
  assign N245 = ~N244;
  assign v_o[16] = fifo_v & N482;
  assign N482 = ~sent_r[16];
  assign N246 = ~reset_i;
  assign N247 = reset_i;
  assign N248 = sent_n[16] & N483;
  assign N483 = ~fifo_yumi;
  assign N250 = v_o[16] & ready_i[16];
  assign N251 = ~N250;
  assign v_o[17] = fifo_v & N484;
  assign N484 = ~sent_r[17];
  assign N252 = ~reset_i;
  assign N253 = reset_i;
  assign N254 = sent_n[17] & N485;
  assign N485 = ~fifo_yumi;
  assign N256 = v_o[17] & ready_i[17];
  assign N257 = ~N256;
  assign v_o[18] = fifo_v & N486;
  assign N486 = ~sent_r[18];
  assign N258 = ~reset_i;
  assign N259 = reset_i;
  assign N260 = sent_n[18] & N487;
  assign N487 = ~fifo_yumi;
  assign N262 = v_o[18] & ready_i[18];
  assign N263 = ~N262;
  assign v_o[19] = fifo_v & N488;
  assign N488 = ~sent_r[19];
  assign N264 = ~reset_i;
  assign N265 = reset_i;
  assign N266 = sent_n[19] & N489;
  assign N489 = ~fifo_yumi;
  assign N268 = v_o[19] & ready_i[19];
  assign N269 = ~N268;
  assign v_o[20] = fifo_v & N490;
  assign N490 = ~sent_r[20];
  assign N270 = ~reset_i;
  assign N271 = reset_i;
  assign N272 = sent_n[20] & N491;
  assign N491 = ~fifo_yumi;
  assign N274 = v_o[20] & ready_i[20];
  assign N275 = ~N274;
  assign v_o[21] = fifo_v & N492;
  assign N492 = ~sent_r[21];
  assign N276 = ~reset_i;
  assign N277 = reset_i;
  assign N278 = sent_n[21] & N493;
  assign N493 = ~fifo_yumi;
  assign N280 = v_o[21] & ready_i[21];
  assign N281 = ~N280;
  assign v_o[22] = fifo_v & N494;
  assign N494 = ~sent_r[22];
  assign N282 = ~reset_i;
  assign N283 = reset_i;
  assign N284 = sent_n[22] & N495;
  assign N495 = ~fifo_yumi;
  assign N286 = v_o[22] & ready_i[22];
  assign N287 = ~N286;
  assign v_o[23] = fifo_v & N496;
  assign N496 = ~sent_r[23];
  assign N288 = ~reset_i;
  assign N289 = reset_i;
  assign N290 = sent_n[23] & N497;
  assign N497 = ~fifo_yumi;
  assign N292 = v_o[23] & ready_i[23];
  assign N293 = ~N292;
  assign v_o[24] = fifo_v & N498;
  assign N498 = ~sent_r[24];
  assign N294 = ~reset_i;
  assign N295 = reset_i;
  assign N296 = sent_n[24] & N499;
  assign N499 = ~fifo_yumi;
  assign N298 = v_o[24] & ready_i[24];
  assign N299 = ~N298;
  assign v_o[25] = fifo_v & N500;
  assign N500 = ~sent_r[25];
  assign N300 = ~reset_i;
  assign N301 = reset_i;
  assign N302 = sent_n[25] & N501;
  assign N501 = ~fifo_yumi;
  assign N304 = v_o[25] & ready_i[25];
  assign N305 = ~N304;
  assign v_o[26] = fifo_v & N502;
  assign N502 = ~sent_r[26];
  assign N306 = ~reset_i;
  assign N307 = reset_i;
  assign N308 = sent_n[26] & N503;
  assign N503 = ~fifo_yumi;
  assign N310 = v_o[26] & ready_i[26];
  assign N311 = ~N310;
  assign v_o[27] = fifo_v & N504;
  assign N504 = ~sent_r[27];
  assign N312 = ~reset_i;
  assign N313 = reset_i;
  assign N314 = sent_n[27] & N505;
  assign N505 = ~fifo_yumi;
  assign N316 = v_o[27] & ready_i[27];
  assign N317 = ~N316;
  assign v_o[28] = fifo_v & N506;
  assign N506 = ~sent_r[28];
  assign N318 = ~reset_i;
  assign N319 = reset_i;
  assign N320 = sent_n[28] & N507;
  assign N507 = ~fifo_yumi;
  assign N322 = v_o[28] & ready_i[28];
  assign N323 = ~N322;
  assign v_o[29] = fifo_v & N508;
  assign N508 = ~sent_r[29];
  assign N324 = ~reset_i;
  assign N325 = reset_i;
  assign N326 = sent_n[29] & N509;
  assign N509 = ~fifo_yumi;
  assign N328 = v_o[29] & ready_i[29];
  assign N329 = ~N328;
  assign v_o[30] = fifo_v & N510;
  assign N510 = ~sent_r[30];
  assign N330 = ~reset_i;
  assign N331 = reset_i;
  assign N332 = sent_n[30] & N511;
  assign N511 = ~fifo_yumi;
  assign N334 = v_o[30] & ready_i[30];
  assign N335 = ~N334;
  assign v_o[31] = fifo_v & N512;
  assign N512 = ~sent_r[31];
  assign N336 = ~reset_i;
  assign N337 = reset_i;
  assign N338 = sent_n[31] & N513;
  assign N513 = ~fifo_yumi;
  assign N340 = v_o[31] & ready_i[31];
  assign N341 = ~N340;
  assign v_o[32] = fifo_v & N514;
  assign N514 = ~sent_r[32];
  assign N342 = ~reset_i;
  assign N343 = reset_i;
  assign N344 = sent_n[32] & N515;
  assign N515 = ~fifo_yumi;
  assign N346 = v_o[32] & ready_i[32];
  assign N347 = ~N346;
  assign v_o[33] = fifo_v & N516;
  assign N516 = ~sent_r[33];
  assign N348 = ~reset_i;
  assign N349 = reset_i;
  assign N350 = sent_n[33] & N517;
  assign N517 = ~fifo_yumi;
  assign N352 = v_o[33] & ready_i[33];
  assign N353 = ~N352;
  assign v_o[34] = fifo_v & N518;
  assign N518 = ~sent_r[34];
  assign N354 = ~reset_i;
  assign N355 = reset_i;
  assign N356 = sent_n[34] & N519;
  assign N519 = ~fifo_yumi;
  assign N358 = v_o[34] & ready_i[34];
  assign N359 = ~N358;
  assign v_o[35] = fifo_v & N520;
  assign N520 = ~sent_r[35];
  assign N360 = ~reset_i;
  assign N361 = reset_i;
  assign N362 = sent_n[35] & N521;
  assign N521 = ~fifo_yumi;
  assign N364 = v_o[35] & ready_i[35];
  assign N365 = ~N364;
  assign v_o[36] = fifo_v & N522;
  assign N522 = ~sent_r[36];
  assign N366 = ~reset_i;
  assign N367 = reset_i;
  assign N368 = sent_n[36] & N523;
  assign N523 = ~fifo_yumi;
  assign N370 = v_o[36] & ready_i[36];
  assign N371 = ~N370;
  assign v_o[37] = fifo_v & N524;
  assign N524 = ~sent_r[37];
  assign N372 = ~reset_i;
  assign N373 = reset_i;
  assign N374 = sent_n[37] & N525;
  assign N525 = ~fifo_yumi;
  assign N376 = v_o[37] & ready_i[37];
  assign N377 = ~N376;
  assign v_o[38] = fifo_v & N526;
  assign N526 = ~sent_r[38];
  assign N378 = ~reset_i;
  assign N379 = reset_i;
  assign N380 = sent_n[38] & N527;
  assign N527 = ~fifo_yumi;
  assign N382 = v_o[38] & ready_i[38];
  assign N383 = ~N382;
  assign v_o[39] = fifo_v & N528;
  assign N528 = ~sent_r[39];
  assign N384 = ~reset_i;
  assign N385 = reset_i;
  assign N386 = sent_n[39] & N529;
  assign N529 = ~fifo_yumi;
  assign N388 = v_o[39] & ready_i[39];
  assign N389 = ~N388;
  assign v_o[40] = fifo_v & N530;
  assign N530 = ~sent_r[40];
  assign N390 = ~reset_i;
  assign N391 = reset_i;
  assign N392 = sent_n[40] & N531;
  assign N531 = ~fifo_yumi;
  assign N394 = v_o[40] & ready_i[40];
  assign N395 = ~N394;
  assign v_o[41] = fifo_v & N532;
  assign N532 = ~sent_r[41];
  assign N396 = ~reset_i;
  assign N397 = reset_i;
  assign N398 = sent_n[41] & N533;
  assign N533 = ~fifo_yumi;
  assign N400 = v_o[41] & ready_i[41];
  assign N401 = ~N400;
  assign v_o[42] = fifo_v & N534;
  assign N534 = ~sent_r[42];
  assign N402 = ~reset_i;
  assign N403 = reset_i;
  assign N404 = sent_n[42] & N535;
  assign N535 = ~fifo_yumi;
  assign N406 = v_o[42] & ready_i[42];
  assign N407 = ~N406;
  assign v_o[43] = fifo_v & N536;
  assign N536 = ~sent_r[43];
  assign N408 = ~reset_i;
  assign N409 = reset_i;
  assign N410 = sent_n[43] & N537;
  assign N537 = ~fifo_yumi;
  assign N412 = v_o[43] & ready_i[43];
  assign N413 = ~N412;
  assign v_o[44] = fifo_v & N538;
  assign N538 = ~sent_r[44];
  assign N414 = ~reset_i;
  assign N415 = reset_i;
  assign N416 = sent_n[44] & N539;
  assign N539 = ~fifo_yumi;
  assign N418 = v_o[44] & ready_i[44];
  assign N419 = ~N418;
  assign v_o[45] = fifo_v & N540;
  assign N540 = ~sent_r[45];
  assign N420 = ~reset_i;
  assign N421 = reset_i;
  assign N422 = sent_n[45] & N541;
  assign N541 = ~fifo_yumi;
  assign N424 = v_o[45] & ready_i[45];
  assign N425 = ~N424;
  assign v_o[46] = fifo_v & N542;
  assign N542 = ~sent_r[46];
  assign N426 = ~reset_i;
  assign N427 = reset_i;
  assign N428 = sent_n[46] & N543;
  assign N543 = ~fifo_yumi;
  assign N430 = v_o[46] & ready_i[46];
  assign N431 = ~N430;
  assign v_o[47] = fifo_v & N544;
  assign N544 = ~sent_r[47];
  assign N432 = ~reset_i;
  assign N433 = reset_i;
  assign N434 = sent_n[47] & N545;
  assign N545 = ~fifo_yumi;
  assign N436 = v_o[47] & ready_i[47];
  assign N437 = ~N436;
  assign v_o[48] = fifo_v & N546;
  assign N546 = ~sent_r[48];
  assign N438 = ~reset_i;
  assign N439 = reset_i;
  assign N440 = sent_n[48] & N547;
  assign N547 = ~fifo_yumi;
  assign N442 = v_o[48] & ready_i[48];
  assign N443 = ~N442;
  assign v_o[49] = fifo_v & N548;
  assign N548 = ~sent_r[49];
  assign N444 = ~reset_i;
  assign N445 = reset_i;
  assign N446 = sent_n[49] & N549;
  assign N549 = ~fifo_yumi;
  assign N448 = v_o[49] & ready_i[49];
  assign N449 = ~N448;
  assign fifo_yumi = N597 & sent_n[0];
  assign N597 = N596 & sent_n[1];
  assign N596 = N595 & sent_n[2];
  assign N595 = N594 & sent_n[3];
  assign N594 = N593 & sent_n[4];
  assign N593 = N592 & sent_n[5];
  assign N592 = N591 & sent_n[6];
  assign N591 = N590 & sent_n[7];
  assign N590 = N589 & sent_n[8];
  assign N589 = N588 & sent_n[9];
  assign N588 = N587 & sent_n[10];
  assign N587 = N586 & sent_n[11];
  assign N586 = N585 & sent_n[12];
  assign N585 = N584 & sent_n[13];
  assign N584 = N583 & sent_n[14];
  assign N583 = N582 & sent_n[15];
  assign N582 = N581 & sent_n[16];
  assign N581 = N580 & sent_n[17];
  assign N580 = N579 & sent_n[18];
  assign N579 = N578 & sent_n[19];
  assign N578 = N577 & sent_n[20];
  assign N577 = N576 & sent_n[21];
  assign N576 = N575 & sent_n[22];
  assign N575 = N574 & sent_n[23];
  assign N574 = N573 & sent_n[24];
  assign N573 = N572 & sent_n[25];
  assign N572 = N571 & sent_n[26];
  assign N571 = N570 & sent_n[27];
  assign N570 = N569 & sent_n[28];
  assign N569 = N568 & sent_n[29];
  assign N568 = N567 & sent_n[30];
  assign N567 = N566 & sent_n[31];
  assign N566 = N565 & sent_n[32];
  assign N565 = N564 & sent_n[33];
  assign N564 = N563 & sent_n[34];
  assign N563 = N562 & sent_n[35];
  assign N562 = N561 & sent_n[36];
  assign N561 = N560 & sent_n[37];
  assign N560 = N559 & sent_n[38];
  assign N559 = N558 & sent_n[39];
  assign N558 = N557 & sent_n[40];
  assign N557 = N556 & sent_n[41];
  assign N556 = N555 & sent_n[42];
  assign N555 = N554 & sent_n[43];
  assign N554 = N553 & sent_n[44];
  assign N553 = N552 & sent_n[45];
  assign N552 = N551 & sent_n[46];
  assign N551 = N550 & sent_n[47];
  assign N550 = sent_n[49] & sent_n[48];

  always @(posedge clk_i) begin
    if(1'b1) begin
      { sent_r[49:0] } <= { N447, N441, N435, N429, N423, N417, N411, N405, N399, N393, N387, N381, N375, N369, N363, N357, N351, N345, N339, N333, N327, N321, N315, N309, N303, N297, N291, N285, N279, N273, N267, N261, N255, N249, N243, N237, N231, N225, N219, N213, N207, N201, N195, N189, N183, N177, N171, N165, N159, N153 };
    end 
  end


endmodule

